module heichips25_example_large (clk,
    ena,
    rst_n,
    ui_in,
    uio_in,
    uio_oe,
    uio_out,
    uo_out);
 input clk;
 input ena;
 input rst_n;
 input [7:0] ui_in;
 input [7:0] uio_in;
 output [7:0] uio_oe;
 output [7:0] uio_out;
 output [7:0] uo_out;

 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire _09_;
 wire _10_;
 wire _11_;
 wire _12_;
 wire _13_;
 wire _14_;
 wire _15_;
 wire _16_;
 wire _17_;
 wire _18_;
 wire _19_;
 wire _20_;
 wire _21_;
 wire _22_;
 wire _23_;
 wire _24_;
 wire _25_;
 wire _26_;
 wire _27_;
 wire _28_;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net40;
 wire net17;
 wire net18;
 wire net19;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net1;
 wire net2;
 wire net3;
 wire net4;
 wire net5;
 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net25;

 sg13g2_and2_1 _29_ (.A(net1),
    .B(net9),
    .X(_00_));
 sg13g2_and2_1 _30_ (.A(net2),
    .B(net10),
    .X(_01_));
 sg13g2_xor2_1 _31_ (.B(net10),
    .A(net2),
    .X(_02_));
 sg13g2_xor2_1 _32_ (.B(_02_),
    .A(_00_),
    .X(net18));
 sg13g2_a21oi_2 _33_ (.B1(_01_),
    .Y(_03_),
    .A2(_02_),
    .A1(_00_));
 sg13g2_and2_1 _34_ (.A(net3),
    .B(net11),
    .X(_04_));
 sg13g2_xnor2_1 _35_ (.Y(_05_),
    .A(net3),
    .B(net11));
 sg13g2_nor2_1 _36_ (.A(_03_),
    .B(_05_),
    .Y(_06_));
 sg13g2_xor2_1 _37_ (.B(_05_),
    .A(_03_),
    .X(net19));
 sg13g2_or2_1 _38_ (.X(_07_),
    .B(net12),
    .A(net4));
 sg13g2_and2_1 _39_ (.A(net4),
    .B(net12),
    .X(_08_));
 sg13g2_xor2_1 _40_ (.B(net12),
    .A(net4),
    .X(_09_));
 sg13g2_nor2_1 _41_ (.A(_04_),
    .B(_06_),
    .Y(_10_));
 sg13g2_xnor2_1 _42_ (.Y(net20),
    .A(_09_),
    .B(_10_));
 sg13g2_nand2b_1 _43_ (.Y(_11_),
    .B(_09_),
    .A_N(_05_));
 sg13g2_a21oi_1 _44_ (.A1(_04_),
    .A2(_07_),
    .Y(_12_),
    .B1(_08_));
 sg13g2_o21ai_1 _45_ (.B1(_12_),
    .Y(_13_),
    .A1(_03_),
    .A2(_11_));
 sg13g2_nand2_1 _46_ (.Y(_14_),
    .A(net5),
    .B(net13));
 sg13g2_xor2_1 _47_ (.B(net13),
    .A(net5),
    .X(_15_));
 sg13g2_inv_1 _48_ (.Y(_16_),
    .A(_15_));
 sg13g2_nand2_1 _49_ (.Y(_17_),
    .A(_13_),
    .B(_15_));
 sg13g2_xnor2_1 _50_ (.Y(net21),
    .A(_13_),
    .B(_16_));
 sg13g2_nor2_1 _51_ (.A(net6),
    .B(net14),
    .Y(_18_));
 sg13g2_xnor2_1 _52_ (.Y(_19_),
    .A(net6),
    .B(net14));
 sg13g2_nand2_1 _53_ (.Y(_20_),
    .A(_14_),
    .B(_17_));
 sg13g2_xnor2_1 _54_ (.Y(net22),
    .A(_19_),
    .B(_20_));
 sg13g2_nor2_1 _55_ (.A(_16_),
    .B(_19_),
    .Y(_21_));
 sg13g2_nor2_1 _56_ (.A(_14_),
    .B(_18_),
    .Y(_22_));
 sg13g2_a221oi_1 _57_ (.B2(_21_),
    .C1(_22_),
    .B1(_13_),
    .A1(net6),
    .Y(_23_),
    .A2(net14));
 sg13g2_nand2_1 _58_ (.Y(_24_),
    .A(net7),
    .B(net15));
 sg13g2_nor2_1 _59_ (.A(net7),
    .B(net15),
    .Y(_25_));
 sg13g2_xor2_1 _60_ (.B(net15),
    .A(net7),
    .X(_26_));
 sg13g2_xnor2_1 _61_ (.Y(net23),
    .A(_23_),
    .B(_26_));
 sg13g2_o21ai_1 _62_ (.B1(_24_),
    .Y(_27_),
    .A1(_23_),
    .A2(_25_));
 sg13g2_xnor2_1 _63_ (.Y(_28_),
    .A(net8),
    .B(net16));
 sg13g2_xnor2_1 _64_ (.Y(net24),
    .A(_27_),
    .B(_28_));
 sg13g2_xor2_1 _65_ (.B(net9),
    .A(net1),
    .X(net17));
 sg13g2_tielo heichips25_example_large_26 (.L_LO(net26));
 sg13g2_tielo heichips25_example_large_27 (.L_LO(net27));
 sg13g2_tielo heichips25_example_large_28 (.L_LO(net28));
 sg13g2_tielo heichips25_example_large_29 (.L_LO(net29));
 sg13g2_tielo heichips25_example_large_30 (.L_LO(net30));
 sg13g2_tielo heichips25_example_large_31 (.L_LO(net31));
 sg13g2_tielo heichips25_example_large_32 (.L_LO(net32));
 sg13g2_tielo heichips25_example_large_33 (.L_LO(net33));
 sg13g2_tielo heichips25_example_large_34 (.L_LO(net34));
 sg13g2_tielo heichips25_example_large_35 (.L_LO(net35));
 sg13g2_tielo heichips25_example_large_36 (.L_LO(net36));
 sg13g2_tielo heichips25_example_large_37 (.L_LO(net37));
 sg13g2_tielo heichips25_example_large_38 (.L_LO(net38));
 sg13g2_tielo heichips25_example_large_39 (.L_LO(net39));
 sg13g2_tielo heichips25_example_large_40 (.L_LO(net40));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_buf_1 input1 (.A(ui_in[0]),
    .X(net1));
 sg13g2_buf_1 input2 (.A(ui_in[1]),
    .X(net2));
 sg13g2_buf_1 input3 (.A(ui_in[2]),
    .X(net3));
 sg13g2_buf_1 input4 (.A(ui_in[3]),
    .X(net4));
 sg13g2_buf_1 input5 (.A(ui_in[4]),
    .X(net5));
 sg13g2_buf_1 input6 (.A(ui_in[5]),
    .X(net6));
 sg13g2_buf_1 input7 (.A(ui_in[6]),
    .X(net7));
 sg13g2_buf_1 input8 (.A(ui_in[7]),
    .X(net8));
 sg13g2_buf_1 input9 (.A(uio_in[0]),
    .X(net9));
 sg13g2_buf_1 input10 (.A(uio_in[1]),
    .X(net10));
 sg13g2_buf_1 input11 (.A(uio_in[2]),
    .X(net11));
 sg13g2_buf_1 input12 (.A(uio_in[3]),
    .X(net12));
 sg13g2_buf_1 input13 (.A(uio_in[4]),
    .X(net13));
 sg13g2_buf_2 input14 (.A(uio_in[5]),
    .X(net14));
 sg13g2_buf_1 input15 (.A(uio_in[6]),
    .X(net15));
 sg13g2_buf_1 input16 (.A(uio_in[7]),
    .X(net16));
 sg13g2_buf_1 output17 (.A(net17),
    .X(uo_out[0]));
 sg13g2_buf_1 output18 (.A(net18),
    .X(uo_out[1]));
 sg13g2_buf_1 output19 (.A(net19),
    .X(uo_out[2]));
 sg13g2_buf_1 output20 (.A(net20),
    .X(uo_out[3]));
 sg13g2_buf_1 output21 (.A(net21),
    .X(uo_out[4]));
 sg13g2_buf_1 output22 (.A(net22),
    .X(uo_out[5]));
 sg13g2_buf_1 output23 (.A(net23),
    .X(uo_out[6]));
 sg13g2_buf_1 output24 (.A(net24),
    .X(uo_out[7]));
 sg13g2_tielo heichips25_example_large_25 (.L_LO(net25));
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_168 ();
 sg13g2_decap_8 FILLER_0_175 ();
 sg13g2_decap_8 FILLER_0_182 ();
 sg13g2_decap_8 FILLER_0_189 ();
 sg13g2_decap_8 FILLER_0_196 ();
 sg13g2_decap_8 FILLER_0_203 ();
 sg13g2_decap_8 FILLER_0_210 ();
 sg13g2_decap_8 FILLER_0_217 ();
 sg13g2_decap_8 FILLER_0_224 ();
 sg13g2_decap_8 FILLER_0_231 ();
 sg13g2_decap_8 FILLER_0_238 ();
 sg13g2_decap_8 FILLER_0_245 ();
 sg13g2_decap_8 FILLER_0_252 ();
 sg13g2_decap_8 FILLER_0_259 ();
 sg13g2_decap_8 FILLER_0_266 ();
 sg13g2_decap_8 FILLER_0_273 ();
 sg13g2_decap_8 FILLER_0_280 ();
 sg13g2_decap_8 FILLER_0_287 ();
 sg13g2_decap_8 FILLER_0_294 ();
 sg13g2_decap_8 FILLER_0_301 ();
 sg13g2_decap_8 FILLER_0_308 ();
 sg13g2_decap_8 FILLER_0_315 ();
 sg13g2_decap_8 FILLER_0_322 ();
 sg13g2_decap_8 FILLER_0_329 ();
 sg13g2_decap_8 FILLER_0_336 ();
 sg13g2_decap_8 FILLER_0_343 ();
 sg13g2_decap_8 FILLER_0_350 ();
 sg13g2_decap_8 FILLER_0_357 ();
 sg13g2_decap_8 FILLER_0_364 ();
 sg13g2_decap_8 FILLER_0_371 ();
 sg13g2_decap_8 FILLER_0_378 ();
 sg13g2_decap_8 FILLER_0_385 ();
 sg13g2_decap_8 FILLER_0_392 ();
 sg13g2_decap_8 FILLER_0_399 ();
 sg13g2_decap_8 FILLER_0_406 ();
 sg13g2_decap_8 FILLER_0_413 ();
 sg13g2_decap_8 FILLER_0_420 ();
 sg13g2_decap_8 FILLER_0_427 ();
 sg13g2_decap_8 FILLER_0_434 ();
 sg13g2_decap_8 FILLER_0_441 ();
 sg13g2_decap_8 FILLER_0_448 ();
 sg13g2_decap_8 FILLER_0_455 ();
 sg13g2_decap_8 FILLER_0_462 ();
 sg13g2_decap_8 FILLER_0_469 ();
 sg13g2_decap_8 FILLER_0_476 ();
 sg13g2_decap_8 FILLER_0_483 ();
 sg13g2_decap_8 FILLER_0_490 ();
 sg13g2_decap_8 FILLER_0_497 ();
 sg13g2_decap_8 FILLER_0_504 ();
 sg13g2_decap_8 FILLER_0_511 ();
 sg13g2_decap_8 FILLER_0_518 ();
 sg13g2_decap_8 FILLER_0_525 ();
 sg13g2_decap_8 FILLER_0_532 ();
 sg13g2_decap_8 FILLER_0_539 ();
 sg13g2_decap_8 FILLER_0_546 ();
 sg13g2_decap_8 FILLER_0_553 ();
 sg13g2_decap_8 FILLER_0_560 ();
 sg13g2_decap_8 FILLER_0_567 ();
 sg13g2_decap_8 FILLER_0_574 ();
 sg13g2_decap_8 FILLER_0_581 ();
 sg13g2_decap_8 FILLER_0_588 ();
 sg13g2_decap_8 FILLER_0_595 ();
 sg13g2_decap_8 FILLER_0_602 ();
 sg13g2_decap_8 FILLER_0_609 ();
 sg13g2_decap_8 FILLER_0_616 ();
 sg13g2_decap_8 FILLER_0_623 ();
 sg13g2_decap_8 FILLER_0_630 ();
 sg13g2_decap_8 FILLER_0_637 ();
 sg13g2_decap_8 FILLER_0_644 ();
 sg13g2_decap_8 FILLER_0_651 ();
 sg13g2_decap_8 FILLER_0_658 ();
 sg13g2_decap_8 FILLER_0_665 ();
 sg13g2_decap_8 FILLER_0_672 ();
 sg13g2_decap_8 FILLER_0_679 ();
 sg13g2_decap_8 FILLER_0_686 ();
 sg13g2_decap_8 FILLER_0_693 ();
 sg13g2_decap_8 FILLER_0_700 ();
 sg13g2_decap_8 FILLER_0_707 ();
 sg13g2_decap_8 FILLER_0_714 ();
 sg13g2_decap_8 FILLER_0_721 ();
 sg13g2_decap_8 FILLER_0_728 ();
 sg13g2_decap_8 FILLER_0_735 ();
 sg13g2_decap_8 FILLER_0_742 ();
 sg13g2_decap_8 FILLER_0_749 ();
 sg13g2_decap_8 FILLER_0_756 ();
 sg13g2_decap_8 FILLER_0_763 ();
 sg13g2_decap_8 FILLER_0_770 ();
 sg13g2_decap_8 FILLER_0_777 ();
 sg13g2_decap_8 FILLER_0_784 ();
 sg13g2_decap_8 FILLER_0_791 ();
 sg13g2_decap_8 FILLER_0_798 ();
 sg13g2_decap_8 FILLER_0_805 ();
 sg13g2_decap_8 FILLER_0_812 ();
 sg13g2_decap_8 FILLER_0_819 ();
 sg13g2_decap_8 FILLER_0_826 ();
 sg13g2_decap_8 FILLER_0_833 ();
 sg13g2_decap_8 FILLER_0_840 ();
 sg13g2_decap_8 FILLER_0_847 ();
 sg13g2_decap_8 FILLER_0_854 ();
 sg13g2_decap_8 FILLER_0_861 ();
 sg13g2_decap_8 FILLER_0_868 ();
 sg13g2_decap_8 FILLER_0_875 ();
 sg13g2_decap_8 FILLER_0_882 ();
 sg13g2_decap_8 FILLER_0_889 ();
 sg13g2_decap_8 FILLER_0_896 ();
 sg13g2_decap_8 FILLER_0_903 ();
 sg13g2_decap_8 FILLER_0_910 ();
 sg13g2_decap_8 FILLER_0_917 ();
 sg13g2_decap_8 FILLER_0_924 ();
 sg13g2_decap_8 FILLER_0_931 ();
 sg13g2_decap_8 FILLER_0_938 ();
 sg13g2_decap_8 FILLER_0_945 ();
 sg13g2_decap_8 FILLER_0_952 ();
 sg13g2_decap_8 FILLER_0_959 ();
 sg13g2_decap_8 FILLER_0_966 ();
 sg13g2_decap_8 FILLER_0_973 ();
 sg13g2_decap_8 FILLER_0_980 ();
 sg13g2_decap_8 FILLER_0_987 ();
 sg13g2_decap_8 FILLER_0_994 ();
 sg13g2_decap_8 FILLER_0_1001 ();
 sg13g2_decap_8 FILLER_0_1008 ();
 sg13g2_decap_8 FILLER_0_1015 ();
 sg13g2_decap_8 FILLER_0_1022 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_7 ();
 sg13g2_decap_8 FILLER_1_14 ();
 sg13g2_decap_8 FILLER_1_21 ();
 sg13g2_decap_8 FILLER_1_28 ();
 sg13g2_decap_8 FILLER_1_35 ();
 sg13g2_decap_8 FILLER_1_42 ();
 sg13g2_decap_8 FILLER_1_49 ();
 sg13g2_decap_8 FILLER_1_56 ();
 sg13g2_decap_8 FILLER_1_63 ();
 sg13g2_decap_8 FILLER_1_70 ();
 sg13g2_decap_8 FILLER_1_77 ();
 sg13g2_decap_8 FILLER_1_84 ();
 sg13g2_decap_8 FILLER_1_91 ();
 sg13g2_decap_8 FILLER_1_98 ();
 sg13g2_decap_8 FILLER_1_105 ();
 sg13g2_decap_8 FILLER_1_112 ();
 sg13g2_decap_8 FILLER_1_119 ();
 sg13g2_decap_8 FILLER_1_126 ();
 sg13g2_decap_8 FILLER_1_133 ();
 sg13g2_decap_8 FILLER_1_140 ();
 sg13g2_decap_8 FILLER_1_147 ();
 sg13g2_decap_8 FILLER_1_154 ();
 sg13g2_decap_8 FILLER_1_161 ();
 sg13g2_decap_8 FILLER_1_168 ();
 sg13g2_decap_8 FILLER_1_175 ();
 sg13g2_decap_8 FILLER_1_182 ();
 sg13g2_decap_8 FILLER_1_189 ();
 sg13g2_decap_8 FILLER_1_196 ();
 sg13g2_decap_8 FILLER_1_203 ();
 sg13g2_decap_8 FILLER_1_210 ();
 sg13g2_decap_8 FILLER_1_217 ();
 sg13g2_decap_8 FILLER_1_224 ();
 sg13g2_decap_8 FILLER_1_231 ();
 sg13g2_decap_8 FILLER_1_238 ();
 sg13g2_decap_8 FILLER_1_245 ();
 sg13g2_decap_8 FILLER_1_252 ();
 sg13g2_decap_8 FILLER_1_259 ();
 sg13g2_decap_8 FILLER_1_266 ();
 sg13g2_decap_8 FILLER_1_273 ();
 sg13g2_decap_8 FILLER_1_280 ();
 sg13g2_decap_8 FILLER_1_287 ();
 sg13g2_decap_8 FILLER_1_294 ();
 sg13g2_decap_8 FILLER_1_301 ();
 sg13g2_decap_8 FILLER_1_308 ();
 sg13g2_decap_8 FILLER_1_315 ();
 sg13g2_decap_8 FILLER_1_322 ();
 sg13g2_decap_8 FILLER_1_329 ();
 sg13g2_decap_8 FILLER_1_336 ();
 sg13g2_decap_8 FILLER_1_343 ();
 sg13g2_decap_8 FILLER_1_350 ();
 sg13g2_decap_8 FILLER_1_357 ();
 sg13g2_decap_8 FILLER_1_364 ();
 sg13g2_decap_8 FILLER_1_371 ();
 sg13g2_decap_8 FILLER_1_378 ();
 sg13g2_decap_8 FILLER_1_385 ();
 sg13g2_decap_8 FILLER_1_392 ();
 sg13g2_decap_8 FILLER_1_399 ();
 sg13g2_decap_8 FILLER_1_406 ();
 sg13g2_decap_8 FILLER_1_413 ();
 sg13g2_decap_8 FILLER_1_420 ();
 sg13g2_decap_8 FILLER_1_427 ();
 sg13g2_decap_8 FILLER_1_434 ();
 sg13g2_decap_8 FILLER_1_441 ();
 sg13g2_decap_8 FILLER_1_448 ();
 sg13g2_decap_8 FILLER_1_455 ();
 sg13g2_decap_8 FILLER_1_462 ();
 sg13g2_decap_8 FILLER_1_469 ();
 sg13g2_decap_8 FILLER_1_476 ();
 sg13g2_decap_8 FILLER_1_483 ();
 sg13g2_decap_8 FILLER_1_490 ();
 sg13g2_decap_8 FILLER_1_497 ();
 sg13g2_decap_8 FILLER_1_504 ();
 sg13g2_decap_8 FILLER_1_511 ();
 sg13g2_decap_8 FILLER_1_518 ();
 sg13g2_decap_8 FILLER_1_525 ();
 sg13g2_decap_8 FILLER_1_532 ();
 sg13g2_decap_8 FILLER_1_539 ();
 sg13g2_decap_8 FILLER_1_546 ();
 sg13g2_decap_8 FILLER_1_553 ();
 sg13g2_decap_8 FILLER_1_560 ();
 sg13g2_decap_8 FILLER_1_567 ();
 sg13g2_decap_8 FILLER_1_574 ();
 sg13g2_decap_8 FILLER_1_581 ();
 sg13g2_decap_8 FILLER_1_588 ();
 sg13g2_decap_8 FILLER_1_595 ();
 sg13g2_decap_8 FILLER_1_602 ();
 sg13g2_decap_8 FILLER_1_609 ();
 sg13g2_decap_8 FILLER_1_616 ();
 sg13g2_decap_8 FILLER_1_623 ();
 sg13g2_decap_8 FILLER_1_630 ();
 sg13g2_decap_8 FILLER_1_637 ();
 sg13g2_decap_8 FILLER_1_644 ();
 sg13g2_decap_8 FILLER_1_651 ();
 sg13g2_decap_8 FILLER_1_658 ();
 sg13g2_decap_8 FILLER_1_665 ();
 sg13g2_decap_8 FILLER_1_672 ();
 sg13g2_decap_8 FILLER_1_679 ();
 sg13g2_decap_8 FILLER_1_686 ();
 sg13g2_decap_8 FILLER_1_693 ();
 sg13g2_decap_8 FILLER_1_700 ();
 sg13g2_decap_8 FILLER_1_707 ();
 sg13g2_decap_8 FILLER_1_714 ();
 sg13g2_decap_8 FILLER_1_721 ();
 sg13g2_decap_8 FILLER_1_728 ();
 sg13g2_decap_8 FILLER_1_735 ();
 sg13g2_decap_8 FILLER_1_742 ();
 sg13g2_decap_8 FILLER_1_749 ();
 sg13g2_decap_8 FILLER_1_756 ();
 sg13g2_decap_8 FILLER_1_763 ();
 sg13g2_decap_8 FILLER_1_770 ();
 sg13g2_decap_8 FILLER_1_777 ();
 sg13g2_decap_8 FILLER_1_784 ();
 sg13g2_decap_8 FILLER_1_791 ();
 sg13g2_decap_8 FILLER_1_798 ();
 sg13g2_decap_8 FILLER_1_805 ();
 sg13g2_decap_8 FILLER_1_812 ();
 sg13g2_decap_8 FILLER_1_819 ();
 sg13g2_decap_8 FILLER_1_826 ();
 sg13g2_decap_8 FILLER_1_833 ();
 sg13g2_decap_8 FILLER_1_840 ();
 sg13g2_decap_8 FILLER_1_847 ();
 sg13g2_decap_8 FILLER_1_854 ();
 sg13g2_decap_8 FILLER_1_861 ();
 sg13g2_decap_8 FILLER_1_868 ();
 sg13g2_decap_8 FILLER_1_875 ();
 sg13g2_decap_8 FILLER_1_882 ();
 sg13g2_decap_8 FILLER_1_889 ();
 sg13g2_decap_8 FILLER_1_896 ();
 sg13g2_decap_8 FILLER_1_903 ();
 sg13g2_decap_8 FILLER_1_910 ();
 sg13g2_decap_8 FILLER_1_917 ();
 sg13g2_decap_8 FILLER_1_924 ();
 sg13g2_decap_8 FILLER_1_931 ();
 sg13g2_decap_8 FILLER_1_938 ();
 sg13g2_decap_8 FILLER_1_945 ();
 sg13g2_decap_8 FILLER_1_952 ();
 sg13g2_decap_8 FILLER_1_959 ();
 sg13g2_decap_8 FILLER_1_966 ();
 sg13g2_decap_8 FILLER_1_973 ();
 sg13g2_decap_8 FILLER_1_980 ();
 sg13g2_decap_8 FILLER_1_987 ();
 sg13g2_decap_8 FILLER_1_994 ();
 sg13g2_decap_8 FILLER_1_1001 ();
 sg13g2_decap_8 FILLER_1_1008 ();
 sg13g2_decap_8 FILLER_1_1015 ();
 sg13g2_decap_8 FILLER_1_1022 ();
 sg13g2_decap_8 FILLER_2_4 ();
 sg13g2_decap_8 FILLER_2_11 ();
 sg13g2_decap_8 FILLER_2_18 ();
 sg13g2_decap_8 FILLER_2_25 ();
 sg13g2_decap_8 FILLER_2_32 ();
 sg13g2_decap_8 FILLER_2_39 ();
 sg13g2_decap_8 FILLER_2_46 ();
 sg13g2_decap_8 FILLER_2_53 ();
 sg13g2_decap_8 FILLER_2_60 ();
 sg13g2_decap_8 FILLER_2_67 ();
 sg13g2_decap_8 FILLER_2_74 ();
 sg13g2_decap_8 FILLER_2_81 ();
 sg13g2_decap_8 FILLER_2_88 ();
 sg13g2_decap_8 FILLER_2_95 ();
 sg13g2_decap_8 FILLER_2_102 ();
 sg13g2_decap_8 FILLER_2_109 ();
 sg13g2_decap_8 FILLER_2_116 ();
 sg13g2_decap_8 FILLER_2_123 ();
 sg13g2_decap_8 FILLER_2_130 ();
 sg13g2_decap_8 FILLER_2_137 ();
 sg13g2_decap_8 FILLER_2_144 ();
 sg13g2_decap_8 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_158 ();
 sg13g2_decap_8 FILLER_2_165 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_2_200 ();
 sg13g2_decap_8 FILLER_2_207 ();
 sg13g2_decap_8 FILLER_2_214 ();
 sg13g2_decap_8 FILLER_2_221 ();
 sg13g2_decap_8 FILLER_2_228 ();
 sg13g2_decap_8 FILLER_2_235 ();
 sg13g2_decap_8 FILLER_2_242 ();
 sg13g2_decap_8 FILLER_2_249 ();
 sg13g2_decap_8 FILLER_2_256 ();
 sg13g2_decap_8 FILLER_2_263 ();
 sg13g2_decap_8 FILLER_2_270 ();
 sg13g2_decap_8 FILLER_2_277 ();
 sg13g2_decap_8 FILLER_2_284 ();
 sg13g2_decap_8 FILLER_2_291 ();
 sg13g2_decap_8 FILLER_2_298 ();
 sg13g2_decap_8 FILLER_2_305 ();
 sg13g2_decap_8 FILLER_2_312 ();
 sg13g2_decap_8 FILLER_2_319 ();
 sg13g2_decap_8 FILLER_2_326 ();
 sg13g2_decap_8 FILLER_2_333 ();
 sg13g2_decap_8 FILLER_2_340 ();
 sg13g2_decap_8 FILLER_2_347 ();
 sg13g2_decap_8 FILLER_2_354 ();
 sg13g2_decap_8 FILLER_2_361 ();
 sg13g2_decap_8 FILLER_2_368 ();
 sg13g2_decap_8 FILLER_2_375 ();
 sg13g2_decap_8 FILLER_2_382 ();
 sg13g2_decap_8 FILLER_2_389 ();
 sg13g2_decap_8 FILLER_2_396 ();
 sg13g2_decap_8 FILLER_2_403 ();
 sg13g2_decap_8 FILLER_2_410 ();
 sg13g2_decap_8 FILLER_2_417 ();
 sg13g2_decap_8 FILLER_2_424 ();
 sg13g2_decap_8 FILLER_2_431 ();
 sg13g2_decap_8 FILLER_2_438 ();
 sg13g2_decap_8 FILLER_2_445 ();
 sg13g2_decap_8 FILLER_2_452 ();
 sg13g2_decap_8 FILLER_2_459 ();
 sg13g2_decap_8 FILLER_2_466 ();
 sg13g2_decap_8 FILLER_2_473 ();
 sg13g2_decap_8 FILLER_2_480 ();
 sg13g2_decap_8 FILLER_2_487 ();
 sg13g2_decap_8 FILLER_2_494 ();
 sg13g2_decap_8 FILLER_2_501 ();
 sg13g2_decap_8 FILLER_2_508 ();
 sg13g2_decap_8 FILLER_2_515 ();
 sg13g2_decap_8 FILLER_2_522 ();
 sg13g2_decap_8 FILLER_2_529 ();
 sg13g2_decap_8 FILLER_2_536 ();
 sg13g2_decap_8 FILLER_2_543 ();
 sg13g2_decap_8 FILLER_2_550 ();
 sg13g2_decap_8 FILLER_2_557 ();
 sg13g2_decap_8 FILLER_2_564 ();
 sg13g2_decap_8 FILLER_2_571 ();
 sg13g2_decap_8 FILLER_2_578 ();
 sg13g2_decap_8 FILLER_2_585 ();
 sg13g2_decap_8 FILLER_2_592 ();
 sg13g2_decap_8 FILLER_2_599 ();
 sg13g2_decap_8 FILLER_2_606 ();
 sg13g2_decap_8 FILLER_2_613 ();
 sg13g2_decap_8 FILLER_2_620 ();
 sg13g2_decap_8 FILLER_2_627 ();
 sg13g2_decap_8 FILLER_2_634 ();
 sg13g2_decap_8 FILLER_2_641 ();
 sg13g2_decap_8 FILLER_2_648 ();
 sg13g2_decap_8 FILLER_2_655 ();
 sg13g2_decap_8 FILLER_2_662 ();
 sg13g2_decap_8 FILLER_2_669 ();
 sg13g2_decap_8 FILLER_2_676 ();
 sg13g2_decap_8 FILLER_2_683 ();
 sg13g2_decap_8 FILLER_2_690 ();
 sg13g2_decap_8 FILLER_2_697 ();
 sg13g2_decap_8 FILLER_2_704 ();
 sg13g2_decap_8 FILLER_2_711 ();
 sg13g2_decap_8 FILLER_2_718 ();
 sg13g2_decap_8 FILLER_2_725 ();
 sg13g2_decap_8 FILLER_2_732 ();
 sg13g2_decap_8 FILLER_2_739 ();
 sg13g2_decap_8 FILLER_2_746 ();
 sg13g2_decap_8 FILLER_2_753 ();
 sg13g2_decap_8 FILLER_2_760 ();
 sg13g2_decap_8 FILLER_2_767 ();
 sg13g2_decap_8 FILLER_2_774 ();
 sg13g2_decap_8 FILLER_2_781 ();
 sg13g2_decap_8 FILLER_2_788 ();
 sg13g2_decap_8 FILLER_2_795 ();
 sg13g2_decap_8 FILLER_2_802 ();
 sg13g2_decap_8 FILLER_2_809 ();
 sg13g2_decap_8 FILLER_2_816 ();
 sg13g2_decap_8 FILLER_2_823 ();
 sg13g2_decap_8 FILLER_2_830 ();
 sg13g2_decap_8 FILLER_2_837 ();
 sg13g2_decap_8 FILLER_2_844 ();
 sg13g2_decap_8 FILLER_2_851 ();
 sg13g2_decap_8 FILLER_2_858 ();
 sg13g2_decap_8 FILLER_2_865 ();
 sg13g2_decap_8 FILLER_2_872 ();
 sg13g2_decap_8 FILLER_2_879 ();
 sg13g2_decap_8 FILLER_2_886 ();
 sg13g2_decap_8 FILLER_2_893 ();
 sg13g2_decap_8 FILLER_2_900 ();
 sg13g2_decap_8 FILLER_2_907 ();
 sg13g2_decap_8 FILLER_2_914 ();
 sg13g2_decap_8 FILLER_2_921 ();
 sg13g2_decap_8 FILLER_2_928 ();
 sg13g2_decap_8 FILLER_2_935 ();
 sg13g2_decap_8 FILLER_2_942 ();
 sg13g2_decap_8 FILLER_2_949 ();
 sg13g2_decap_8 FILLER_2_956 ();
 sg13g2_decap_8 FILLER_2_963 ();
 sg13g2_decap_8 FILLER_2_970 ();
 sg13g2_decap_8 FILLER_2_977 ();
 sg13g2_decap_8 FILLER_2_984 ();
 sg13g2_decap_8 FILLER_2_991 ();
 sg13g2_decap_8 FILLER_2_998 ();
 sg13g2_decap_8 FILLER_2_1005 ();
 sg13g2_decap_8 FILLER_2_1012 ();
 sg13g2_decap_8 FILLER_2_1019 ();
 sg13g2_fill_2 FILLER_2_1026 ();
 sg13g2_fill_1 FILLER_2_1028 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_7 ();
 sg13g2_decap_8 FILLER_3_14 ();
 sg13g2_decap_8 FILLER_3_21 ();
 sg13g2_decap_8 FILLER_3_28 ();
 sg13g2_decap_8 FILLER_3_35 ();
 sg13g2_decap_8 FILLER_3_42 ();
 sg13g2_decap_8 FILLER_3_49 ();
 sg13g2_decap_8 FILLER_3_56 ();
 sg13g2_decap_8 FILLER_3_63 ();
 sg13g2_decap_8 FILLER_3_70 ();
 sg13g2_decap_8 FILLER_3_77 ();
 sg13g2_decap_8 FILLER_3_84 ();
 sg13g2_decap_8 FILLER_3_91 ();
 sg13g2_decap_8 FILLER_3_98 ();
 sg13g2_decap_8 FILLER_3_105 ();
 sg13g2_decap_8 FILLER_3_112 ();
 sg13g2_decap_8 FILLER_3_119 ();
 sg13g2_decap_8 FILLER_3_126 ();
 sg13g2_decap_8 FILLER_3_133 ();
 sg13g2_decap_8 FILLER_3_140 ();
 sg13g2_decap_8 FILLER_3_147 ();
 sg13g2_decap_8 FILLER_3_154 ();
 sg13g2_decap_8 FILLER_3_161 ();
 sg13g2_decap_8 FILLER_3_168 ();
 sg13g2_decap_8 FILLER_3_175 ();
 sg13g2_decap_8 FILLER_3_182 ();
 sg13g2_decap_8 FILLER_3_189 ();
 sg13g2_decap_8 FILLER_3_196 ();
 sg13g2_decap_8 FILLER_3_203 ();
 sg13g2_decap_8 FILLER_3_210 ();
 sg13g2_decap_8 FILLER_3_217 ();
 sg13g2_decap_8 FILLER_3_224 ();
 sg13g2_decap_8 FILLER_3_231 ();
 sg13g2_decap_8 FILLER_3_238 ();
 sg13g2_decap_8 FILLER_3_245 ();
 sg13g2_decap_8 FILLER_3_252 ();
 sg13g2_decap_8 FILLER_3_259 ();
 sg13g2_decap_8 FILLER_3_266 ();
 sg13g2_decap_8 FILLER_3_273 ();
 sg13g2_decap_8 FILLER_3_280 ();
 sg13g2_decap_8 FILLER_3_287 ();
 sg13g2_decap_8 FILLER_3_294 ();
 sg13g2_decap_8 FILLER_3_301 ();
 sg13g2_decap_8 FILLER_3_308 ();
 sg13g2_decap_8 FILLER_3_315 ();
 sg13g2_decap_8 FILLER_3_322 ();
 sg13g2_decap_8 FILLER_3_329 ();
 sg13g2_decap_8 FILLER_3_336 ();
 sg13g2_decap_8 FILLER_3_343 ();
 sg13g2_decap_8 FILLER_3_350 ();
 sg13g2_decap_8 FILLER_3_357 ();
 sg13g2_decap_8 FILLER_3_364 ();
 sg13g2_decap_8 FILLER_3_371 ();
 sg13g2_decap_8 FILLER_3_378 ();
 sg13g2_decap_8 FILLER_3_385 ();
 sg13g2_decap_8 FILLER_3_392 ();
 sg13g2_decap_8 FILLER_3_399 ();
 sg13g2_decap_8 FILLER_3_406 ();
 sg13g2_decap_8 FILLER_3_413 ();
 sg13g2_decap_8 FILLER_3_420 ();
 sg13g2_decap_8 FILLER_3_427 ();
 sg13g2_decap_8 FILLER_3_434 ();
 sg13g2_decap_8 FILLER_3_441 ();
 sg13g2_decap_8 FILLER_3_448 ();
 sg13g2_decap_8 FILLER_3_455 ();
 sg13g2_decap_8 FILLER_3_462 ();
 sg13g2_decap_8 FILLER_3_469 ();
 sg13g2_decap_8 FILLER_3_476 ();
 sg13g2_decap_8 FILLER_3_483 ();
 sg13g2_decap_8 FILLER_3_490 ();
 sg13g2_decap_8 FILLER_3_497 ();
 sg13g2_decap_8 FILLER_3_504 ();
 sg13g2_decap_8 FILLER_3_511 ();
 sg13g2_decap_8 FILLER_3_518 ();
 sg13g2_decap_8 FILLER_3_525 ();
 sg13g2_decap_8 FILLER_3_532 ();
 sg13g2_decap_8 FILLER_3_539 ();
 sg13g2_decap_8 FILLER_3_546 ();
 sg13g2_decap_8 FILLER_3_553 ();
 sg13g2_decap_8 FILLER_3_560 ();
 sg13g2_decap_8 FILLER_3_567 ();
 sg13g2_decap_8 FILLER_3_574 ();
 sg13g2_decap_8 FILLER_3_581 ();
 sg13g2_decap_8 FILLER_3_588 ();
 sg13g2_decap_8 FILLER_3_595 ();
 sg13g2_decap_8 FILLER_3_602 ();
 sg13g2_decap_8 FILLER_3_609 ();
 sg13g2_decap_8 FILLER_3_616 ();
 sg13g2_decap_8 FILLER_3_623 ();
 sg13g2_decap_8 FILLER_3_630 ();
 sg13g2_decap_8 FILLER_3_637 ();
 sg13g2_decap_8 FILLER_3_644 ();
 sg13g2_decap_8 FILLER_3_651 ();
 sg13g2_decap_8 FILLER_3_658 ();
 sg13g2_decap_8 FILLER_3_665 ();
 sg13g2_decap_8 FILLER_3_672 ();
 sg13g2_decap_8 FILLER_3_679 ();
 sg13g2_decap_8 FILLER_3_686 ();
 sg13g2_decap_8 FILLER_3_693 ();
 sg13g2_decap_8 FILLER_3_700 ();
 sg13g2_decap_8 FILLER_3_707 ();
 sg13g2_decap_8 FILLER_3_714 ();
 sg13g2_decap_8 FILLER_3_721 ();
 sg13g2_decap_8 FILLER_3_728 ();
 sg13g2_decap_8 FILLER_3_735 ();
 sg13g2_decap_8 FILLER_3_742 ();
 sg13g2_decap_8 FILLER_3_749 ();
 sg13g2_decap_8 FILLER_3_756 ();
 sg13g2_decap_8 FILLER_3_763 ();
 sg13g2_decap_8 FILLER_3_770 ();
 sg13g2_decap_8 FILLER_3_777 ();
 sg13g2_decap_8 FILLER_3_784 ();
 sg13g2_decap_8 FILLER_3_791 ();
 sg13g2_decap_8 FILLER_3_798 ();
 sg13g2_decap_8 FILLER_3_805 ();
 sg13g2_decap_8 FILLER_3_812 ();
 sg13g2_decap_8 FILLER_3_819 ();
 sg13g2_decap_8 FILLER_3_826 ();
 sg13g2_decap_8 FILLER_3_833 ();
 sg13g2_decap_8 FILLER_3_840 ();
 sg13g2_decap_8 FILLER_3_847 ();
 sg13g2_decap_8 FILLER_3_854 ();
 sg13g2_decap_8 FILLER_3_861 ();
 sg13g2_decap_8 FILLER_3_868 ();
 sg13g2_decap_8 FILLER_3_875 ();
 sg13g2_decap_8 FILLER_3_882 ();
 sg13g2_decap_8 FILLER_3_889 ();
 sg13g2_decap_8 FILLER_3_896 ();
 sg13g2_decap_8 FILLER_3_903 ();
 sg13g2_decap_8 FILLER_3_910 ();
 sg13g2_decap_8 FILLER_3_917 ();
 sg13g2_decap_8 FILLER_3_924 ();
 sg13g2_decap_8 FILLER_3_931 ();
 sg13g2_decap_8 FILLER_3_938 ();
 sg13g2_decap_8 FILLER_3_945 ();
 sg13g2_decap_8 FILLER_3_952 ();
 sg13g2_decap_8 FILLER_3_959 ();
 sg13g2_decap_8 FILLER_3_966 ();
 sg13g2_decap_8 FILLER_3_973 ();
 sg13g2_decap_8 FILLER_3_980 ();
 sg13g2_decap_8 FILLER_3_987 ();
 sg13g2_decap_8 FILLER_3_994 ();
 sg13g2_decap_8 FILLER_3_1001 ();
 sg13g2_decap_8 FILLER_3_1008 ();
 sg13g2_decap_8 FILLER_3_1015 ();
 sg13g2_decap_8 FILLER_3_1022 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_7 ();
 sg13g2_decap_8 FILLER_4_14 ();
 sg13g2_decap_8 FILLER_4_21 ();
 sg13g2_decap_8 FILLER_4_28 ();
 sg13g2_decap_8 FILLER_4_35 ();
 sg13g2_decap_8 FILLER_4_42 ();
 sg13g2_decap_8 FILLER_4_49 ();
 sg13g2_decap_8 FILLER_4_56 ();
 sg13g2_decap_8 FILLER_4_63 ();
 sg13g2_decap_8 FILLER_4_70 ();
 sg13g2_decap_8 FILLER_4_77 ();
 sg13g2_decap_8 FILLER_4_84 ();
 sg13g2_decap_8 FILLER_4_91 ();
 sg13g2_decap_8 FILLER_4_98 ();
 sg13g2_decap_8 FILLER_4_105 ();
 sg13g2_decap_8 FILLER_4_112 ();
 sg13g2_decap_8 FILLER_4_119 ();
 sg13g2_decap_8 FILLER_4_126 ();
 sg13g2_decap_8 FILLER_4_133 ();
 sg13g2_decap_8 FILLER_4_140 ();
 sg13g2_decap_8 FILLER_4_147 ();
 sg13g2_decap_8 FILLER_4_154 ();
 sg13g2_decap_8 FILLER_4_161 ();
 sg13g2_decap_8 FILLER_4_168 ();
 sg13g2_decap_8 FILLER_4_175 ();
 sg13g2_decap_8 FILLER_4_182 ();
 sg13g2_decap_8 FILLER_4_189 ();
 sg13g2_decap_8 FILLER_4_196 ();
 sg13g2_decap_8 FILLER_4_203 ();
 sg13g2_decap_8 FILLER_4_210 ();
 sg13g2_decap_8 FILLER_4_217 ();
 sg13g2_decap_8 FILLER_4_224 ();
 sg13g2_decap_8 FILLER_4_231 ();
 sg13g2_decap_8 FILLER_4_238 ();
 sg13g2_decap_8 FILLER_4_245 ();
 sg13g2_decap_8 FILLER_4_252 ();
 sg13g2_decap_8 FILLER_4_259 ();
 sg13g2_decap_8 FILLER_4_266 ();
 sg13g2_decap_8 FILLER_4_273 ();
 sg13g2_decap_8 FILLER_4_280 ();
 sg13g2_decap_8 FILLER_4_287 ();
 sg13g2_decap_8 FILLER_4_294 ();
 sg13g2_decap_8 FILLER_4_301 ();
 sg13g2_decap_8 FILLER_4_308 ();
 sg13g2_decap_8 FILLER_4_315 ();
 sg13g2_decap_8 FILLER_4_322 ();
 sg13g2_decap_8 FILLER_4_329 ();
 sg13g2_decap_8 FILLER_4_336 ();
 sg13g2_decap_8 FILLER_4_343 ();
 sg13g2_decap_8 FILLER_4_350 ();
 sg13g2_decap_8 FILLER_4_357 ();
 sg13g2_decap_8 FILLER_4_364 ();
 sg13g2_decap_8 FILLER_4_371 ();
 sg13g2_decap_8 FILLER_4_378 ();
 sg13g2_decap_8 FILLER_4_385 ();
 sg13g2_decap_8 FILLER_4_392 ();
 sg13g2_decap_8 FILLER_4_399 ();
 sg13g2_decap_8 FILLER_4_406 ();
 sg13g2_decap_8 FILLER_4_413 ();
 sg13g2_decap_8 FILLER_4_420 ();
 sg13g2_decap_8 FILLER_4_427 ();
 sg13g2_decap_8 FILLER_4_434 ();
 sg13g2_decap_8 FILLER_4_441 ();
 sg13g2_decap_8 FILLER_4_448 ();
 sg13g2_decap_8 FILLER_4_455 ();
 sg13g2_decap_8 FILLER_4_462 ();
 sg13g2_decap_8 FILLER_4_469 ();
 sg13g2_decap_8 FILLER_4_476 ();
 sg13g2_decap_8 FILLER_4_483 ();
 sg13g2_decap_8 FILLER_4_490 ();
 sg13g2_decap_8 FILLER_4_497 ();
 sg13g2_decap_8 FILLER_4_504 ();
 sg13g2_decap_8 FILLER_4_511 ();
 sg13g2_decap_8 FILLER_4_518 ();
 sg13g2_decap_8 FILLER_4_525 ();
 sg13g2_decap_8 FILLER_4_532 ();
 sg13g2_decap_8 FILLER_4_539 ();
 sg13g2_decap_8 FILLER_4_546 ();
 sg13g2_decap_8 FILLER_4_553 ();
 sg13g2_decap_8 FILLER_4_560 ();
 sg13g2_decap_8 FILLER_4_567 ();
 sg13g2_decap_8 FILLER_4_574 ();
 sg13g2_decap_8 FILLER_4_581 ();
 sg13g2_decap_8 FILLER_4_588 ();
 sg13g2_decap_8 FILLER_4_595 ();
 sg13g2_decap_8 FILLER_4_602 ();
 sg13g2_decap_8 FILLER_4_609 ();
 sg13g2_decap_8 FILLER_4_616 ();
 sg13g2_decap_8 FILLER_4_623 ();
 sg13g2_decap_8 FILLER_4_630 ();
 sg13g2_decap_8 FILLER_4_637 ();
 sg13g2_decap_8 FILLER_4_644 ();
 sg13g2_decap_8 FILLER_4_651 ();
 sg13g2_decap_8 FILLER_4_658 ();
 sg13g2_decap_8 FILLER_4_665 ();
 sg13g2_decap_8 FILLER_4_672 ();
 sg13g2_decap_8 FILLER_4_679 ();
 sg13g2_decap_8 FILLER_4_686 ();
 sg13g2_decap_8 FILLER_4_693 ();
 sg13g2_decap_8 FILLER_4_700 ();
 sg13g2_decap_8 FILLER_4_707 ();
 sg13g2_decap_8 FILLER_4_714 ();
 sg13g2_decap_8 FILLER_4_721 ();
 sg13g2_decap_8 FILLER_4_728 ();
 sg13g2_decap_8 FILLER_4_735 ();
 sg13g2_decap_8 FILLER_4_742 ();
 sg13g2_decap_8 FILLER_4_749 ();
 sg13g2_decap_8 FILLER_4_756 ();
 sg13g2_decap_8 FILLER_4_763 ();
 sg13g2_decap_8 FILLER_4_770 ();
 sg13g2_decap_8 FILLER_4_777 ();
 sg13g2_decap_8 FILLER_4_784 ();
 sg13g2_decap_8 FILLER_4_791 ();
 sg13g2_decap_8 FILLER_4_798 ();
 sg13g2_decap_8 FILLER_4_805 ();
 sg13g2_decap_8 FILLER_4_812 ();
 sg13g2_decap_8 FILLER_4_819 ();
 sg13g2_decap_8 FILLER_4_826 ();
 sg13g2_decap_8 FILLER_4_833 ();
 sg13g2_decap_8 FILLER_4_840 ();
 sg13g2_decap_8 FILLER_4_847 ();
 sg13g2_decap_8 FILLER_4_854 ();
 sg13g2_decap_8 FILLER_4_861 ();
 sg13g2_decap_8 FILLER_4_868 ();
 sg13g2_decap_8 FILLER_4_875 ();
 sg13g2_decap_8 FILLER_4_882 ();
 sg13g2_decap_8 FILLER_4_889 ();
 sg13g2_decap_8 FILLER_4_896 ();
 sg13g2_decap_8 FILLER_4_903 ();
 sg13g2_decap_8 FILLER_4_910 ();
 sg13g2_decap_8 FILLER_4_917 ();
 sg13g2_decap_8 FILLER_4_924 ();
 sg13g2_decap_8 FILLER_4_931 ();
 sg13g2_decap_8 FILLER_4_938 ();
 sg13g2_decap_8 FILLER_4_945 ();
 sg13g2_decap_8 FILLER_4_952 ();
 sg13g2_decap_8 FILLER_4_959 ();
 sg13g2_decap_8 FILLER_4_966 ();
 sg13g2_decap_8 FILLER_4_973 ();
 sg13g2_decap_8 FILLER_4_980 ();
 sg13g2_decap_8 FILLER_4_987 ();
 sg13g2_decap_8 FILLER_4_994 ();
 sg13g2_decap_8 FILLER_4_1001 ();
 sg13g2_decap_8 FILLER_4_1008 ();
 sg13g2_decap_8 FILLER_4_1015 ();
 sg13g2_decap_8 FILLER_4_1022 ();
 sg13g2_decap_8 FILLER_5_4 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_decap_8 FILLER_5_158 ();
 sg13g2_decap_8 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_172 ();
 sg13g2_decap_8 FILLER_5_179 ();
 sg13g2_decap_8 FILLER_5_186 ();
 sg13g2_decap_8 FILLER_5_193 ();
 sg13g2_decap_8 FILLER_5_200 ();
 sg13g2_decap_8 FILLER_5_207 ();
 sg13g2_decap_8 FILLER_5_214 ();
 sg13g2_decap_8 FILLER_5_221 ();
 sg13g2_decap_8 FILLER_5_228 ();
 sg13g2_decap_8 FILLER_5_235 ();
 sg13g2_decap_8 FILLER_5_242 ();
 sg13g2_decap_8 FILLER_5_249 ();
 sg13g2_decap_8 FILLER_5_256 ();
 sg13g2_decap_8 FILLER_5_263 ();
 sg13g2_decap_8 FILLER_5_270 ();
 sg13g2_decap_8 FILLER_5_277 ();
 sg13g2_decap_8 FILLER_5_284 ();
 sg13g2_decap_8 FILLER_5_291 ();
 sg13g2_decap_8 FILLER_5_298 ();
 sg13g2_decap_8 FILLER_5_305 ();
 sg13g2_decap_8 FILLER_5_312 ();
 sg13g2_decap_8 FILLER_5_319 ();
 sg13g2_decap_8 FILLER_5_326 ();
 sg13g2_decap_8 FILLER_5_333 ();
 sg13g2_decap_8 FILLER_5_340 ();
 sg13g2_decap_8 FILLER_5_347 ();
 sg13g2_decap_8 FILLER_5_354 ();
 sg13g2_decap_8 FILLER_5_361 ();
 sg13g2_decap_8 FILLER_5_368 ();
 sg13g2_decap_8 FILLER_5_375 ();
 sg13g2_decap_8 FILLER_5_382 ();
 sg13g2_decap_8 FILLER_5_389 ();
 sg13g2_decap_8 FILLER_5_396 ();
 sg13g2_decap_8 FILLER_5_403 ();
 sg13g2_decap_8 FILLER_5_410 ();
 sg13g2_decap_8 FILLER_5_417 ();
 sg13g2_decap_8 FILLER_5_424 ();
 sg13g2_decap_8 FILLER_5_431 ();
 sg13g2_decap_8 FILLER_5_438 ();
 sg13g2_decap_8 FILLER_5_445 ();
 sg13g2_decap_8 FILLER_5_452 ();
 sg13g2_decap_8 FILLER_5_459 ();
 sg13g2_decap_8 FILLER_5_466 ();
 sg13g2_decap_8 FILLER_5_473 ();
 sg13g2_decap_8 FILLER_5_480 ();
 sg13g2_decap_8 FILLER_5_487 ();
 sg13g2_decap_8 FILLER_5_494 ();
 sg13g2_decap_8 FILLER_5_501 ();
 sg13g2_decap_8 FILLER_5_508 ();
 sg13g2_decap_8 FILLER_5_515 ();
 sg13g2_decap_8 FILLER_5_522 ();
 sg13g2_decap_8 FILLER_5_529 ();
 sg13g2_decap_8 FILLER_5_536 ();
 sg13g2_decap_8 FILLER_5_543 ();
 sg13g2_decap_8 FILLER_5_550 ();
 sg13g2_decap_8 FILLER_5_557 ();
 sg13g2_decap_8 FILLER_5_564 ();
 sg13g2_decap_8 FILLER_5_571 ();
 sg13g2_decap_8 FILLER_5_578 ();
 sg13g2_decap_8 FILLER_5_585 ();
 sg13g2_decap_8 FILLER_5_592 ();
 sg13g2_decap_8 FILLER_5_599 ();
 sg13g2_decap_8 FILLER_5_606 ();
 sg13g2_decap_8 FILLER_5_613 ();
 sg13g2_decap_8 FILLER_5_620 ();
 sg13g2_decap_8 FILLER_5_627 ();
 sg13g2_decap_8 FILLER_5_634 ();
 sg13g2_decap_8 FILLER_5_641 ();
 sg13g2_decap_8 FILLER_5_648 ();
 sg13g2_decap_8 FILLER_5_655 ();
 sg13g2_decap_8 FILLER_5_662 ();
 sg13g2_decap_8 FILLER_5_669 ();
 sg13g2_decap_8 FILLER_5_676 ();
 sg13g2_decap_8 FILLER_5_683 ();
 sg13g2_decap_8 FILLER_5_690 ();
 sg13g2_decap_8 FILLER_5_697 ();
 sg13g2_decap_8 FILLER_5_704 ();
 sg13g2_decap_8 FILLER_5_711 ();
 sg13g2_decap_8 FILLER_5_718 ();
 sg13g2_decap_8 FILLER_5_725 ();
 sg13g2_decap_8 FILLER_5_732 ();
 sg13g2_decap_8 FILLER_5_739 ();
 sg13g2_decap_8 FILLER_5_746 ();
 sg13g2_decap_8 FILLER_5_753 ();
 sg13g2_decap_8 FILLER_5_760 ();
 sg13g2_decap_8 FILLER_5_767 ();
 sg13g2_decap_8 FILLER_5_774 ();
 sg13g2_decap_8 FILLER_5_781 ();
 sg13g2_decap_8 FILLER_5_788 ();
 sg13g2_decap_8 FILLER_5_795 ();
 sg13g2_decap_8 FILLER_5_802 ();
 sg13g2_decap_8 FILLER_5_809 ();
 sg13g2_decap_8 FILLER_5_816 ();
 sg13g2_decap_8 FILLER_5_823 ();
 sg13g2_decap_8 FILLER_5_830 ();
 sg13g2_decap_8 FILLER_5_837 ();
 sg13g2_decap_8 FILLER_5_844 ();
 sg13g2_decap_8 FILLER_5_851 ();
 sg13g2_decap_8 FILLER_5_858 ();
 sg13g2_decap_8 FILLER_5_865 ();
 sg13g2_decap_8 FILLER_5_872 ();
 sg13g2_decap_8 FILLER_5_879 ();
 sg13g2_decap_8 FILLER_5_886 ();
 sg13g2_decap_8 FILLER_5_893 ();
 sg13g2_decap_8 FILLER_5_900 ();
 sg13g2_decap_8 FILLER_5_907 ();
 sg13g2_decap_8 FILLER_5_914 ();
 sg13g2_decap_8 FILLER_5_921 ();
 sg13g2_decap_8 FILLER_5_928 ();
 sg13g2_decap_8 FILLER_5_935 ();
 sg13g2_decap_8 FILLER_5_942 ();
 sg13g2_decap_8 FILLER_5_949 ();
 sg13g2_decap_8 FILLER_5_956 ();
 sg13g2_decap_8 FILLER_5_963 ();
 sg13g2_decap_8 FILLER_5_970 ();
 sg13g2_decap_8 FILLER_5_977 ();
 sg13g2_decap_8 FILLER_5_984 ();
 sg13g2_decap_8 FILLER_5_991 ();
 sg13g2_decap_8 FILLER_5_998 ();
 sg13g2_decap_8 FILLER_5_1005 ();
 sg13g2_decap_8 FILLER_5_1012 ();
 sg13g2_decap_8 FILLER_5_1019 ();
 sg13g2_fill_2 FILLER_5_1026 ();
 sg13g2_fill_1 FILLER_5_1028 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_7 ();
 sg13g2_decap_8 FILLER_6_14 ();
 sg13g2_decap_8 FILLER_6_21 ();
 sg13g2_decap_8 FILLER_6_28 ();
 sg13g2_decap_8 FILLER_6_35 ();
 sg13g2_decap_8 FILLER_6_42 ();
 sg13g2_decap_8 FILLER_6_49 ();
 sg13g2_decap_8 FILLER_6_56 ();
 sg13g2_decap_8 FILLER_6_63 ();
 sg13g2_decap_8 FILLER_6_70 ();
 sg13g2_decap_8 FILLER_6_77 ();
 sg13g2_decap_8 FILLER_6_84 ();
 sg13g2_decap_8 FILLER_6_91 ();
 sg13g2_decap_8 FILLER_6_98 ();
 sg13g2_decap_8 FILLER_6_105 ();
 sg13g2_decap_8 FILLER_6_112 ();
 sg13g2_decap_8 FILLER_6_119 ();
 sg13g2_decap_8 FILLER_6_126 ();
 sg13g2_decap_8 FILLER_6_133 ();
 sg13g2_decap_8 FILLER_6_140 ();
 sg13g2_decap_8 FILLER_6_147 ();
 sg13g2_decap_8 FILLER_6_154 ();
 sg13g2_decap_8 FILLER_6_161 ();
 sg13g2_decap_8 FILLER_6_168 ();
 sg13g2_decap_8 FILLER_6_175 ();
 sg13g2_decap_8 FILLER_6_182 ();
 sg13g2_decap_8 FILLER_6_189 ();
 sg13g2_decap_8 FILLER_6_196 ();
 sg13g2_decap_8 FILLER_6_203 ();
 sg13g2_decap_8 FILLER_6_210 ();
 sg13g2_decap_8 FILLER_6_217 ();
 sg13g2_decap_8 FILLER_6_224 ();
 sg13g2_decap_8 FILLER_6_231 ();
 sg13g2_decap_8 FILLER_6_238 ();
 sg13g2_decap_8 FILLER_6_245 ();
 sg13g2_decap_8 FILLER_6_252 ();
 sg13g2_decap_8 FILLER_6_259 ();
 sg13g2_decap_8 FILLER_6_266 ();
 sg13g2_decap_8 FILLER_6_273 ();
 sg13g2_decap_8 FILLER_6_280 ();
 sg13g2_decap_8 FILLER_6_287 ();
 sg13g2_decap_8 FILLER_6_294 ();
 sg13g2_decap_8 FILLER_6_301 ();
 sg13g2_decap_8 FILLER_6_308 ();
 sg13g2_decap_8 FILLER_6_315 ();
 sg13g2_decap_8 FILLER_6_322 ();
 sg13g2_decap_8 FILLER_6_329 ();
 sg13g2_decap_8 FILLER_6_336 ();
 sg13g2_decap_8 FILLER_6_343 ();
 sg13g2_decap_8 FILLER_6_350 ();
 sg13g2_decap_8 FILLER_6_357 ();
 sg13g2_decap_8 FILLER_6_364 ();
 sg13g2_decap_8 FILLER_6_371 ();
 sg13g2_decap_8 FILLER_6_378 ();
 sg13g2_decap_8 FILLER_6_385 ();
 sg13g2_decap_8 FILLER_6_392 ();
 sg13g2_decap_8 FILLER_6_399 ();
 sg13g2_decap_8 FILLER_6_406 ();
 sg13g2_decap_8 FILLER_6_413 ();
 sg13g2_decap_8 FILLER_6_420 ();
 sg13g2_decap_8 FILLER_6_427 ();
 sg13g2_decap_8 FILLER_6_434 ();
 sg13g2_decap_8 FILLER_6_441 ();
 sg13g2_decap_8 FILLER_6_448 ();
 sg13g2_decap_8 FILLER_6_455 ();
 sg13g2_decap_8 FILLER_6_462 ();
 sg13g2_decap_8 FILLER_6_469 ();
 sg13g2_decap_8 FILLER_6_476 ();
 sg13g2_decap_8 FILLER_6_483 ();
 sg13g2_decap_8 FILLER_6_490 ();
 sg13g2_decap_8 FILLER_6_497 ();
 sg13g2_decap_8 FILLER_6_504 ();
 sg13g2_decap_8 FILLER_6_511 ();
 sg13g2_decap_8 FILLER_6_518 ();
 sg13g2_decap_8 FILLER_6_525 ();
 sg13g2_decap_8 FILLER_6_532 ();
 sg13g2_decap_8 FILLER_6_539 ();
 sg13g2_decap_8 FILLER_6_546 ();
 sg13g2_decap_8 FILLER_6_553 ();
 sg13g2_decap_8 FILLER_6_560 ();
 sg13g2_decap_8 FILLER_6_567 ();
 sg13g2_decap_8 FILLER_6_574 ();
 sg13g2_decap_8 FILLER_6_581 ();
 sg13g2_decap_8 FILLER_6_588 ();
 sg13g2_decap_8 FILLER_6_595 ();
 sg13g2_decap_8 FILLER_6_602 ();
 sg13g2_decap_8 FILLER_6_609 ();
 sg13g2_decap_8 FILLER_6_616 ();
 sg13g2_decap_8 FILLER_6_623 ();
 sg13g2_decap_8 FILLER_6_630 ();
 sg13g2_decap_8 FILLER_6_637 ();
 sg13g2_decap_8 FILLER_6_644 ();
 sg13g2_decap_8 FILLER_6_651 ();
 sg13g2_decap_8 FILLER_6_658 ();
 sg13g2_decap_8 FILLER_6_665 ();
 sg13g2_decap_8 FILLER_6_672 ();
 sg13g2_decap_8 FILLER_6_679 ();
 sg13g2_decap_8 FILLER_6_686 ();
 sg13g2_decap_8 FILLER_6_693 ();
 sg13g2_decap_8 FILLER_6_700 ();
 sg13g2_decap_8 FILLER_6_707 ();
 sg13g2_decap_8 FILLER_6_714 ();
 sg13g2_decap_8 FILLER_6_721 ();
 sg13g2_decap_8 FILLER_6_728 ();
 sg13g2_decap_8 FILLER_6_735 ();
 sg13g2_decap_8 FILLER_6_742 ();
 sg13g2_decap_8 FILLER_6_749 ();
 sg13g2_decap_8 FILLER_6_756 ();
 sg13g2_decap_8 FILLER_6_763 ();
 sg13g2_decap_8 FILLER_6_770 ();
 sg13g2_decap_8 FILLER_6_777 ();
 sg13g2_decap_8 FILLER_6_784 ();
 sg13g2_decap_8 FILLER_6_791 ();
 sg13g2_decap_8 FILLER_6_798 ();
 sg13g2_decap_8 FILLER_6_805 ();
 sg13g2_decap_8 FILLER_6_812 ();
 sg13g2_decap_8 FILLER_6_819 ();
 sg13g2_decap_8 FILLER_6_826 ();
 sg13g2_decap_8 FILLER_6_833 ();
 sg13g2_decap_8 FILLER_6_840 ();
 sg13g2_decap_8 FILLER_6_847 ();
 sg13g2_decap_8 FILLER_6_854 ();
 sg13g2_decap_8 FILLER_6_861 ();
 sg13g2_decap_8 FILLER_6_868 ();
 sg13g2_decap_8 FILLER_6_875 ();
 sg13g2_decap_8 FILLER_6_882 ();
 sg13g2_decap_8 FILLER_6_889 ();
 sg13g2_decap_8 FILLER_6_896 ();
 sg13g2_decap_8 FILLER_6_903 ();
 sg13g2_decap_8 FILLER_6_910 ();
 sg13g2_decap_8 FILLER_6_917 ();
 sg13g2_decap_8 FILLER_6_924 ();
 sg13g2_decap_8 FILLER_6_931 ();
 sg13g2_decap_8 FILLER_6_938 ();
 sg13g2_decap_8 FILLER_6_945 ();
 sg13g2_decap_8 FILLER_6_952 ();
 sg13g2_decap_8 FILLER_6_959 ();
 sg13g2_decap_8 FILLER_6_966 ();
 sg13g2_decap_8 FILLER_6_973 ();
 sg13g2_decap_8 FILLER_6_980 ();
 sg13g2_decap_8 FILLER_6_987 ();
 sg13g2_decap_8 FILLER_6_994 ();
 sg13g2_decap_8 FILLER_6_1001 ();
 sg13g2_decap_8 FILLER_6_1008 ();
 sg13g2_decap_8 FILLER_6_1015 ();
 sg13g2_decap_8 FILLER_6_1022 ();
 sg13g2_decap_8 FILLER_7_4 ();
 sg13g2_decap_8 FILLER_7_11 ();
 sg13g2_decap_8 FILLER_7_18 ();
 sg13g2_decap_8 FILLER_7_25 ();
 sg13g2_decap_8 FILLER_7_32 ();
 sg13g2_decap_8 FILLER_7_39 ();
 sg13g2_decap_8 FILLER_7_46 ();
 sg13g2_decap_8 FILLER_7_53 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_decap_8 FILLER_7_67 ();
 sg13g2_decap_8 FILLER_7_74 ();
 sg13g2_decap_8 FILLER_7_81 ();
 sg13g2_decap_8 FILLER_7_88 ();
 sg13g2_decap_8 FILLER_7_95 ();
 sg13g2_decap_8 FILLER_7_102 ();
 sg13g2_decap_8 FILLER_7_109 ();
 sg13g2_decap_8 FILLER_7_116 ();
 sg13g2_decap_8 FILLER_7_123 ();
 sg13g2_decap_8 FILLER_7_130 ();
 sg13g2_decap_8 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_151 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_decap_8 FILLER_7_172 ();
 sg13g2_decap_8 FILLER_7_179 ();
 sg13g2_decap_8 FILLER_7_186 ();
 sg13g2_decap_8 FILLER_7_193 ();
 sg13g2_decap_8 FILLER_7_200 ();
 sg13g2_decap_8 FILLER_7_207 ();
 sg13g2_decap_8 FILLER_7_214 ();
 sg13g2_decap_8 FILLER_7_221 ();
 sg13g2_decap_8 FILLER_7_228 ();
 sg13g2_decap_8 FILLER_7_235 ();
 sg13g2_decap_8 FILLER_7_242 ();
 sg13g2_decap_8 FILLER_7_249 ();
 sg13g2_decap_8 FILLER_7_256 ();
 sg13g2_decap_8 FILLER_7_263 ();
 sg13g2_decap_8 FILLER_7_270 ();
 sg13g2_decap_8 FILLER_7_277 ();
 sg13g2_decap_8 FILLER_7_284 ();
 sg13g2_decap_8 FILLER_7_291 ();
 sg13g2_decap_8 FILLER_7_298 ();
 sg13g2_decap_8 FILLER_7_305 ();
 sg13g2_decap_8 FILLER_7_312 ();
 sg13g2_decap_8 FILLER_7_319 ();
 sg13g2_decap_8 FILLER_7_326 ();
 sg13g2_decap_8 FILLER_7_333 ();
 sg13g2_decap_8 FILLER_7_340 ();
 sg13g2_decap_8 FILLER_7_347 ();
 sg13g2_decap_8 FILLER_7_354 ();
 sg13g2_decap_8 FILLER_7_361 ();
 sg13g2_decap_8 FILLER_7_368 ();
 sg13g2_decap_8 FILLER_7_375 ();
 sg13g2_decap_8 FILLER_7_382 ();
 sg13g2_decap_8 FILLER_7_389 ();
 sg13g2_decap_8 FILLER_7_396 ();
 sg13g2_decap_8 FILLER_7_403 ();
 sg13g2_decap_8 FILLER_7_410 ();
 sg13g2_decap_8 FILLER_7_417 ();
 sg13g2_decap_8 FILLER_7_424 ();
 sg13g2_decap_8 FILLER_7_431 ();
 sg13g2_decap_8 FILLER_7_438 ();
 sg13g2_decap_8 FILLER_7_445 ();
 sg13g2_decap_8 FILLER_7_452 ();
 sg13g2_decap_8 FILLER_7_459 ();
 sg13g2_decap_8 FILLER_7_466 ();
 sg13g2_decap_8 FILLER_7_473 ();
 sg13g2_decap_8 FILLER_7_480 ();
 sg13g2_decap_8 FILLER_7_487 ();
 sg13g2_decap_8 FILLER_7_494 ();
 sg13g2_decap_8 FILLER_7_501 ();
 sg13g2_decap_8 FILLER_7_508 ();
 sg13g2_decap_8 FILLER_7_515 ();
 sg13g2_decap_8 FILLER_7_522 ();
 sg13g2_decap_8 FILLER_7_529 ();
 sg13g2_decap_8 FILLER_7_536 ();
 sg13g2_decap_8 FILLER_7_543 ();
 sg13g2_decap_8 FILLER_7_550 ();
 sg13g2_decap_8 FILLER_7_557 ();
 sg13g2_decap_8 FILLER_7_564 ();
 sg13g2_decap_8 FILLER_7_571 ();
 sg13g2_decap_8 FILLER_7_578 ();
 sg13g2_decap_8 FILLER_7_585 ();
 sg13g2_decap_8 FILLER_7_592 ();
 sg13g2_decap_8 FILLER_7_599 ();
 sg13g2_decap_8 FILLER_7_606 ();
 sg13g2_decap_8 FILLER_7_613 ();
 sg13g2_decap_8 FILLER_7_620 ();
 sg13g2_decap_8 FILLER_7_627 ();
 sg13g2_decap_8 FILLER_7_634 ();
 sg13g2_decap_8 FILLER_7_641 ();
 sg13g2_decap_8 FILLER_7_648 ();
 sg13g2_decap_8 FILLER_7_655 ();
 sg13g2_decap_8 FILLER_7_662 ();
 sg13g2_decap_8 FILLER_7_669 ();
 sg13g2_decap_8 FILLER_7_676 ();
 sg13g2_decap_8 FILLER_7_683 ();
 sg13g2_decap_8 FILLER_7_690 ();
 sg13g2_decap_8 FILLER_7_697 ();
 sg13g2_decap_8 FILLER_7_704 ();
 sg13g2_decap_8 FILLER_7_711 ();
 sg13g2_decap_8 FILLER_7_718 ();
 sg13g2_decap_8 FILLER_7_725 ();
 sg13g2_decap_8 FILLER_7_732 ();
 sg13g2_decap_8 FILLER_7_739 ();
 sg13g2_decap_8 FILLER_7_746 ();
 sg13g2_decap_8 FILLER_7_753 ();
 sg13g2_decap_8 FILLER_7_760 ();
 sg13g2_decap_8 FILLER_7_767 ();
 sg13g2_decap_8 FILLER_7_774 ();
 sg13g2_decap_8 FILLER_7_781 ();
 sg13g2_decap_8 FILLER_7_788 ();
 sg13g2_decap_8 FILLER_7_795 ();
 sg13g2_decap_8 FILLER_7_802 ();
 sg13g2_decap_8 FILLER_7_809 ();
 sg13g2_decap_8 FILLER_7_816 ();
 sg13g2_decap_8 FILLER_7_823 ();
 sg13g2_decap_8 FILLER_7_830 ();
 sg13g2_decap_8 FILLER_7_837 ();
 sg13g2_decap_8 FILLER_7_844 ();
 sg13g2_decap_8 FILLER_7_851 ();
 sg13g2_decap_8 FILLER_7_858 ();
 sg13g2_decap_8 FILLER_7_865 ();
 sg13g2_decap_8 FILLER_7_872 ();
 sg13g2_decap_8 FILLER_7_879 ();
 sg13g2_decap_8 FILLER_7_886 ();
 sg13g2_decap_8 FILLER_7_893 ();
 sg13g2_decap_8 FILLER_7_900 ();
 sg13g2_decap_8 FILLER_7_907 ();
 sg13g2_decap_8 FILLER_7_914 ();
 sg13g2_decap_8 FILLER_7_921 ();
 sg13g2_decap_8 FILLER_7_928 ();
 sg13g2_decap_8 FILLER_7_935 ();
 sg13g2_decap_8 FILLER_7_942 ();
 sg13g2_decap_8 FILLER_7_949 ();
 sg13g2_decap_8 FILLER_7_956 ();
 sg13g2_decap_8 FILLER_7_963 ();
 sg13g2_decap_8 FILLER_7_970 ();
 sg13g2_decap_8 FILLER_7_977 ();
 sg13g2_decap_8 FILLER_7_984 ();
 sg13g2_decap_8 FILLER_7_991 ();
 sg13g2_decap_8 FILLER_7_998 ();
 sg13g2_decap_8 FILLER_7_1005 ();
 sg13g2_decap_8 FILLER_7_1012 ();
 sg13g2_decap_8 FILLER_7_1019 ();
 sg13g2_fill_2 FILLER_7_1026 ();
 sg13g2_fill_1 FILLER_7_1028 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_8 FILLER_8_182 ();
 sg13g2_decap_8 FILLER_8_189 ();
 sg13g2_decap_8 FILLER_8_196 ();
 sg13g2_decap_8 FILLER_8_203 ();
 sg13g2_decap_8 FILLER_8_210 ();
 sg13g2_decap_8 FILLER_8_217 ();
 sg13g2_decap_8 FILLER_8_224 ();
 sg13g2_decap_8 FILLER_8_231 ();
 sg13g2_decap_8 FILLER_8_238 ();
 sg13g2_decap_8 FILLER_8_245 ();
 sg13g2_decap_8 FILLER_8_252 ();
 sg13g2_decap_8 FILLER_8_259 ();
 sg13g2_decap_8 FILLER_8_266 ();
 sg13g2_decap_8 FILLER_8_273 ();
 sg13g2_decap_8 FILLER_8_280 ();
 sg13g2_decap_8 FILLER_8_287 ();
 sg13g2_decap_8 FILLER_8_294 ();
 sg13g2_decap_8 FILLER_8_301 ();
 sg13g2_decap_8 FILLER_8_308 ();
 sg13g2_decap_8 FILLER_8_315 ();
 sg13g2_decap_8 FILLER_8_322 ();
 sg13g2_decap_8 FILLER_8_329 ();
 sg13g2_decap_8 FILLER_8_336 ();
 sg13g2_decap_8 FILLER_8_343 ();
 sg13g2_decap_8 FILLER_8_350 ();
 sg13g2_decap_8 FILLER_8_357 ();
 sg13g2_decap_8 FILLER_8_364 ();
 sg13g2_decap_8 FILLER_8_371 ();
 sg13g2_decap_8 FILLER_8_378 ();
 sg13g2_decap_8 FILLER_8_385 ();
 sg13g2_decap_8 FILLER_8_392 ();
 sg13g2_decap_8 FILLER_8_399 ();
 sg13g2_decap_8 FILLER_8_406 ();
 sg13g2_decap_8 FILLER_8_413 ();
 sg13g2_decap_8 FILLER_8_420 ();
 sg13g2_decap_8 FILLER_8_427 ();
 sg13g2_decap_8 FILLER_8_434 ();
 sg13g2_decap_8 FILLER_8_441 ();
 sg13g2_decap_8 FILLER_8_448 ();
 sg13g2_decap_8 FILLER_8_455 ();
 sg13g2_decap_8 FILLER_8_462 ();
 sg13g2_decap_8 FILLER_8_469 ();
 sg13g2_decap_8 FILLER_8_476 ();
 sg13g2_decap_8 FILLER_8_483 ();
 sg13g2_decap_8 FILLER_8_490 ();
 sg13g2_decap_8 FILLER_8_497 ();
 sg13g2_decap_8 FILLER_8_504 ();
 sg13g2_decap_8 FILLER_8_511 ();
 sg13g2_decap_8 FILLER_8_518 ();
 sg13g2_decap_8 FILLER_8_525 ();
 sg13g2_decap_8 FILLER_8_532 ();
 sg13g2_decap_8 FILLER_8_539 ();
 sg13g2_decap_8 FILLER_8_546 ();
 sg13g2_decap_8 FILLER_8_553 ();
 sg13g2_decap_8 FILLER_8_560 ();
 sg13g2_decap_8 FILLER_8_567 ();
 sg13g2_decap_8 FILLER_8_574 ();
 sg13g2_decap_8 FILLER_8_581 ();
 sg13g2_decap_8 FILLER_8_588 ();
 sg13g2_decap_8 FILLER_8_595 ();
 sg13g2_decap_8 FILLER_8_602 ();
 sg13g2_decap_8 FILLER_8_609 ();
 sg13g2_decap_8 FILLER_8_616 ();
 sg13g2_decap_8 FILLER_8_623 ();
 sg13g2_decap_8 FILLER_8_630 ();
 sg13g2_decap_8 FILLER_8_637 ();
 sg13g2_decap_8 FILLER_8_644 ();
 sg13g2_decap_8 FILLER_8_651 ();
 sg13g2_decap_8 FILLER_8_658 ();
 sg13g2_decap_8 FILLER_8_665 ();
 sg13g2_decap_8 FILLER_8_672 ();
 sg13g2_decap_8 FILLER_8_679 ();
 sg13g2_decap_8 FILLER_8_686 ();
 sg13g2_decap_8 FILLER_8_693 ();
 sg13g2_decap_8 FILLER_8_700 ();
 sg13g2_decap_8 FILLER_8_707 ();
 sg13g2_decap_8 FILLER_8_714 ();
 sg13g2_decap_8 FILLER_8_721 ();
 sg13g2_decap_8 FILLER_8_728 ();
 sg13g2_decap_8 FILLER_8_735 ();
 sg13g2_decap_8 FILLER_8_742 ();
 sg13g2_decap_8 FILLER_8_749 ();
 sg13g2_decap_8 FILLER_8_756 ();
 sg13g2_decap_8 FILLER_8_763 ();
 sg13g2_decap_8 FILLER_8_770 ();
 sg13g2_decap_8 FILLER_8_777 ();
 sg13g2_decap_8 FILLER_8_784 ();
 sg13g2_decap_8 FILLER_8_791 ();
 sg13g2_decap_8 FILLER_8_798 ();
 sg13g2_decap_8 FILLER_8_805 ();
 sg13g2_decap_8 FILLER_8_812 ();
 sg13g2_decap_8 FILLER_8_819 ();
 sg13g2_decap_8 FILLER_8_826 ();
 sg13g2_decap_8 FILLER_8_833 ();
 sg13g2_decap_8 FILLER_8_840 ();
 sg13g2_decap_8 FILLER_8_847 ();
 sg13g2_decap_8 FILLER_8_854 ();
 sg13g2_decap_8 FILLER_8_861 ();
 sg13g2_decap_8 FILLER_8_868 ();
 sg13g2_decap_8 FILLER_8_875 ();
 sg13g2_decap_8 FILLER_8_882 ();
 sg13g2_decap_8 FILLER_8_889 ();
 sg13g2_decap_8 FILLER_8_896 ();
 sg13g2_decap_8 FILLER_8_903 ();
 sg13g2_decap_8 FILLER_8_910 ();
 sg13g2_decap_8 FILLER_8_917 ();
 sg13g2_decap_8 FILLER_8_924 ();
 sg13g2_decap_8 FILLER_8_931 ();
 sg13g2_decap_8 FILLER_8_938 ();
 sg13g2_decap_8 FILLER_8_945 ();
 sg13g2_decap_8 FILLER_8_952 ();
 sg13g2_decap_8 FILLER_8_959 ();
 sg13g2_decap_8 FILLER_8_966 ();
 sg13g2_decap_8 FILLER_8_973 ();
 sg13g2_decap_8 FILLER_8_980 ();
 sg13g2_decap_8 FILLER_8_987 ();
 sg13g2_decap_8 FILLER_8_994 ();
 sg13g2_decap_8 FILLER_8_1001 ();
 sg13g2_decap_8 FILLER_8_1008 ();
 sg13g2_decap_8 FILLER_8_1015 ();
 sg13g2_decap_8 FILLER_8_1022 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_decap_8 FILLER_9_7 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_decap_8 FILLER_9_126 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_8 FILLER_9_196 ();
 sg13g2_decap_8 FILLER_9_203 ();
 sg13g2_decap_8 FILLER_9_210 ();
 sg13g2_decap_8 FILLER_9_217 ();
 sg13g2_decap_8 FILLER_9_224 ();
 sg13g2_decap_8 FILLER_9_231 ();
 sg13g2_decap_8 FILLER_9_238 ();
 sg13g2_decap_8 FILLER_9_245 ();
 sg13g2_decap_8 FILLER_9_252 ();
 sg13g2_decap_8 FILLER_9_259 ();
 sg13g2_decap_8 FILLER_9_266 ();
 sg13g2_decap_8 FILLER_9_273 ();
 sg13g2_decap_8 FILLER_9_280 ();
 sg13g2_decap_8 FILLER_9_287 ();
 sg13g2_decap_8 FILLER_9_294 ();
 sg13g2_decap_8 FILLER_9_301 ();
 sg13g2_decap_8 FILLER_9_308 ();
 sg13g2_decap_8 FILLER_9_315 ();
 sg13g2_decap_8 FILLER_9_322 ();
 sg13g2_decap_8 FILLER_9_329 ();
 sg13g2_decap_8 FILLER_9_336 ();
 sg13g2_decap_8 FILLER_9_343 ();
 sg13g2_decap_8 FILLER_9_350 ();
 sg13g2_decap_8 FILLER_9_357 ();
 sg13g2_decap_8 FILLER_9_364 ();
 sg13g2_decap_8 FILLER_9_371 ();
 sg13g2_decap_8 FILLER_9_378 ();
 sg13g2_decap_8 FILLER_9_385 ();
 sg13g2_decap_8 FILLER_9_392 ();
 sg13g2_decap_8 FILLER_9_399 ();
 sg13g2_decap_8 FILLER_9_406 ();
 sg13g2_decap_8 FILLER_9_413 ();
 sg13g2_decap_8 FILLER_9_420 ();
 sg13g2_decap_8 FILLER_9_427 ();
 sg13g2_decap_8 FILLER_9_434 ();
 sg13g2_decap_8 FILLER_9_441 ();
 sg13g2_decap_8 FILLER_9_448 ();
 sg13g2_decap_8 FILLER_9_455 ();
 sg13g2_decap_8 FILLER_9_462 ();
 sg13g2_decap_8 FILLER_9_469 ();
 sg13g2_decap_8 FILLER_9_476 ();
 sg13g2_decap_8 FILLER_9_483 ();
 sg13g2_decap_8 FILLER_9_490 ();
 sg13g2_decap_8 FILLER_9_497 ();
 sg13g2_decap_8 FILLER_9_504 ();
 sg13g2_decap_8 FILLER_9_511 ();
 sg13g2_decap_8 FILLER_9_518 ();
 sg13g2_decap_8 FILLER_9_525 ();
 sg13g2_decap_8 FILLER_9_532 ();
 sg13g2_decap_8 FILLER_9_539 ();
 sg13g2_decap_8 FILLER_9_546 ();
 sg13g2_decap_8 FILLER_9_553 ();
 sg13g2_decap_8 FILLER_9_560 ();
 sg13g2_decap_8 FILLER_9_567 ();
 sg13g2_decap_8 FILLER_9_574 ();
 sg13g2_decap_8 FILLER_9_581 ();
 sg13g2_decap_8 FILLER_9_588 ();
 sg13g2_decap_8 FILLER_9_595 ();
 sg13g2_decap_8 FILLER_9_602 ();
 sg13g2_decap_8 FILLER_9_609 ();
 sg13g2_decap_8 FILLER_9_616 ();
 sg13g2_decap_8 FILLER_9_623 ();
 sg13g2_decap_8 FILLER_9_630 ();
 sg13g2_decap_8 FILLER_9_637 ();
 sg13g2_decap_8 FILLER_9_644 ();
 sg13g2_decap_8 FILLER_9_651 ();
 sg13g2_decap_8 FILLER_9_658 ();
 sg13g2_decap_8 FILLER_9_665 ();
 sg13g2_decap_8 FILLER_9_672 ();
 sg13g2_decap_8 FILLER_9_679 ();
 sg13g2_decap_8 FILLER_9_686 ();
 sg13g2_decap_8 FILLER_9_693 ();
 sg13g2_decap_8 FILLER_9_700 ();
 sg13g2_decap_8 FILLER_9_707 ();
 sg13g2_decap_8 FILLER_9_714 ();
 sg13g2_decap_8 FILLER_9_721 ();
 sg13g2_decap_8 FILLER_9_728 ();
 sg13g2_decap_8 FILLER_9_735 ();
 sg13g2_decap_8 FILLER_9_742 ();
 sg13g2_decap_8 FILLER_9_749 ();
 sg13g2_decap_8 FILLER_9_756 ();
 sg13g2_decap_8 FILLER_9_763 ();
 sg13g2_decap_8 FILLER_9_770 ();
 sg13g2_decap_8 FILLER_9_777 ();
 sg13g2_decap_8 FILLER_9_784 ();
 sg13g2_decap_8 FILLER_9_791 ();
 sg13g2_decap_8 FILLER_9_798 ();
 sg13g2_decap_8 FILLER_9_805 ();
 sg13g2_decap_8 FILLER_9_812 ();
 sg13g2_decap_8 FILLER_9_819 ();
 sg13g2_decap_8 FILLER_9_826 ();
 sg13g2_decap_8 FILLER_9_833 ();
 sg13g2_decap_8 FILLER_9_840 ();
 sg13g2_decap_8 FILLER_9_847 ();
 sg13g2_decap_8 FILLER_9_854 ();
 sg13g2_decap_8 FILLER_9_861 ();
 sg13g2_decap_8 FILLER_9_868 ();
 sg13g2_decap_8 FILLER_9_875 ();
 sg13g2_decap_8 FILLER_9_882 ();
 sg13g2_decap_8 FILLER_9_889 ();
 sg13g2_decap_8 FILLER_9_896 ();
 sg13g2_decap_8 FILLER_9_903 ();
 sg13g2_decap_8 FILLER_9_910 ();
 sg13g2_decap_8 FILLER_9_917 ();
 sg13g2_decap_8 FILLER_9_924 ();
 sg13g2_decap_8 FILLER_9_931 ();
 sg13g2_decap_8 FILLER_9_938 ();
 sg13g2_decap_8 FILLER_9_945 ();
 sg13g2_decap_8 FILLER_9_952 ();
 sg13g2_decap_8 FILLER_9_959 ();
 sg13g2_decap_8 FILLER_9_966 ();
 sg13g2_decap_8 FILLER_9_973 ();
 sg13g2_decap_8 FILLER_9_980 ();
 sg13g2_decap_8 FILLER_9_987 ();
 sg13g2_decap_8 FILLER_9_994 ();
 sg13g2_decap_8 FILLER_9_1001 ();
 sg13g2_decap_8 FILLER_9_1008 ();
 sg13g2_decap_8 FILLER_9_1015 ();
 sg13g2_decap_8 FILLER_9_1022 ();
 sg13g2_decap_8 FILLER_10_4 ();
 sg13g2_decap_8 FILLER_10_11 ();
 sg13g2_decap_8 FILLER_10_18 ();
 sg13g2_decap_8 FILLER_10_25 ();
 sg13g2_decap_8 FILLER_10_32 ();
 sg13g2_decap_8 FILLER_10_39 ();
 sg13g2_decap_8 FILLER_10_46 ();
 sg13g2_decap_8 FILLER_10_53 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_decap_8 FILLER_10_67 ();
 sg13g2_decap_8 FILLER_10_74 ();
 sg13g2_decap_8 FILLER_10_81 ();
 sg13g2_decap_8 FILLER_10_88 ();
 sg13g2_decap_8 FILLER_10_95 ();
 sg13g2_decap_8 FILLER_10_102 ();
 sg13g2_decap_8 FILLER_10_109 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_123 ();
 sg13g2_decap_8 FILLER_10_130 ();
 sg13g2_decap_8 FILLER_10_137 ();
 sg13g2_decap_8 FILLER_10_144 ();
 sg13g2_decap_8 FILLER_10_151 ();
 sg13g2_decap_8 FILLER_10_158 ();
 sg13g2_decap_8 FILLER_10_165 ();
 sg13g2_decap_8 FILLER_10_172 ();
 sg13g2_decap_8 FILLER_10_179 ();
 sg13g2_decap_8 FILLER_10_186 ();
 sg13g2_decap_8 FILLER_10_193 ();
 sg13g2_decap_8 FILLER_10_200 ();
 sg13g2_decap_8 FILLER_10_207 ();
 sg13g2_decap_8 FILLER_10_214 ();
 sg13g2_decap_8 FILLER_10_221 ();
 sg13g2_decap_8 FILLER_10_228 ();
 sg13g2_decap_8 FILLER_10_235 ();
 sg13g2_decap_8 FILLER_10_242 ();
 sg13g2_decap_8 FILLER_10_249 ();
 sg13g2_decap_8 FILLER_10_256 ();
 sg13g2_decap_8 FILLER_10_263 ();
 sg13g2_decap_8 FILLER_10_270 ();
 sg13g2_decap_8 FILLER_10_277 ();
 sg13g2_decap_8 FILLER_10_284 ();
 sg13g2_decap_8 FILLER_10_291 ();
 sg13g2_decap_8 FILLER_10_298 ();
 sg13g2_decap_8 FILLER_10_305 ();
 sg13g2_decap_8 FILLER_10_312 ();
 sg13g2_decap_8 FILLER_10_319 ();
 sg13g2_decap_8 FILLER_10_326 ();
 sg13g2_decap_8 FILLER_10_333 ();
 sg13g2_decap_8 FILLER_10_340 ();
 sg13g2_decap_8 FILLER_10_347 ();
 sg13g2_decap_8 FILLER_10_354 ();
 sg13g2_decap_8 FILLER_10_361 ();
 sg13g2_decap_8 FILLER_10_368 ();
 sg13g2_decap_8 FILLER_10_375 ();
 sg13g2_decap_8 FILLER_10_382 ();
 sg13g2_decap_8 FILLER_10_389 ();
 sg13g2_decap_8 FILLER_10_396 ();
 sg13g2_decap_8 FILLER_10_403 ();
 sg13g2_decap_8 FILLER_10_410 ();
 sg13g2_decap_8 FILLER_10_417 ();
 sg13g2_decap_8 FILLER_10_424 ();
 sg13g2_decap_8 FILLER_10_431 ();
 sg13g2_decap_8 FILLER_10_438 ();
 sg13g2_decap_8 FILLER_10_445 ();
 sg13g2_decap_8 FILLER_10_452 ();
 sg13g2_decap_8 FILLER_10_459 ();
 sg13g2_decap_8 FILLER_10_466 ();
 sg13g2_decap_8 FILLER_10_473 ();
 sg13g2_decap_8 FILLER_10_480 ();
 sg13g2_decap_8 FILLER_10_487 ();
 sg13g2_decap_8 FILLER_10_494 ();
 sg13g2_decap_8 FILLER_10_501 ();
 sg13g2_decap_8 FILLER_10_508 ();
 sg13g2_decap_8 FILLER_10_515 ();
 sg13g2_decap_8 FILLER_10_522 ();
 sg13g2_decap_8 FILLER_10_529 ();
 sg13g2_decap_8 FILLER_10_536 ();
 sg13g2_decap_8 FILLER_10_543 ();
 sg13g2_decap_8 FILLER_10_550 ();
 sg13g2_decap_8 FILLER_10_557 ();
 sg13g2_decap_8 FILLER_10_564 ();
 sg13g2_decap_8 FILLER_10_571 ();
 sg13g2_decap_8 FILLER_10_578 ();
 sg13g2_decap_8 FILLER_10_585 ();
 sg13g2_decap_8 FILLER_10_592 ();
 sg13g2_decap_8 FILLER_10_599 ();
 sg13g2_decap_8 FILLER_10_606 ();
 sg13g2_decap_8 FILLER_10_613 ();
 sg13g2_decap_8 FILLER_10_620 ();
 sg13g2_decap_8 FILLER_10_627 ();
 sg13g2_decap_8 FILLER_10_634 ();
 sg13g2_decap_8 FILLER_10_641 ();
 sg13g2_decap_8 FILLER_10_648 ();
 sg13g2_decap_8 FILLER_10_655 ();
 sg13g2_decap_8 FILLER_10_662 ();
 sg13g2_decap_8 FILLER_10_669 ();
 sg13g2_decap_8 FILLER_10_676 ();
 sg13g2_decap_8 FILLER_10_683 ();
 sg13g2_decap_8 FILLER_10_690 ();
 sg13g2_decap_8 FILLER_10_697 ();
 sg13g2_decap_8 FILLER_10_704 ();
 sg13g2_decap_8 FILLER_10_711 ();
 sg13g2_decap_8 FILLER_10_718 ();
 sg13g2_decap_8 FILLER_10_725 ();
 sg13g2_decap_8 FILLER_10_732 ();
 sg13g2_decap_8 FILLER_10_739 ();
 sg13g2_decap_8 FILLER_10_746 ();
 sg13g2_decap_8 FILLER_10_753 ();
 sg13g2_decap_8 FILLER_10_760 ();
 sg13g2_decap_8 FILLER_10_767 ();
 sg13g2_decap_8 FILLER_10_774 ();
 sg13g2_decap_8 FILLER_10_781 ();
 sg13g2_decap_8 FILLER_10_788 ();
 sg13g2_decap_8 FILLER_10_795 ();
 sg13g2_decap_8 FILLER_10_802 ();
 sg13g2_decap_8 FILLER_10_809 ();
 sg13g2_decap_8 FILLER_10_816 ();
 sg13g2_decap_8 FILLER_10_823 ();
 sg13g2_decap_8 FILLER_10_830 ();
 sg13g2_decap_8 FILLER_10_837 ();
 sg13g2_decap_8 FILLER_10_844 ();
 sg13g2_decap_8 FILLER_10_851 ();
 sg13g2_decap_8 FILLER_10_858 ();
 sg13g2_decap_8 FILLER_10_865 ();
 sg13g2_decap_8 FILLER_10_872 ();
 sg13g2_decap_8 FILLER_10_879 ();
 sg13g2_decap_8 FILLER_10_886 ();
 sg13g2_decap_8 FILLER_10_893 ();
 sg13g2_decap_8 FILLER_10_900 ();
 sg13g2_decap_8 FILLER_10_907 ();
 sg13g2_decap_8 FILLER_10_914 ();
 sg13g2_decap_8 FILLER_10_921 ();
 sg13g2_decap_8 FILLER_10_928 ();
 sg13g2_decap_8 FILLER_10_935 ();
 sg13g2_decap_8 FILLER_10_942 ();
 sg13g2_decap_8 FILLER_10_949 ();
 sg13g2_decap_8 FILLER_10_956 ();
 sg13g2_decap_8 FILLER_10_963 ();
 sg13g2_decap_8 FILLER_10_970 ();
 sg13g2_decap_8 FILLER_10_977 ();
 sg13g2_decap_8 FILLER_10_984 ();
 sg13g2_decap_8 FILLER_10_991 ();
 sg13g2_decap_8 FILLER_10_998 ();
 sg13g2_decap_8 FILLER_10_1005 ();
 sg13g2_decap_8 FILLER_10_1012 ();
 sg13g2_decap_8 FILLER_10_1019 ();
 sg13g2_fill_2 FILLER_10_1026 ();
 sg13g2_fill_1 FILLER_10_1028 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_8 FILLER_11_196 ();
 sg13g2_decap_8 FILLER_11_203 ();
 sg13g2_decap_8 FILLER_11_210 ();
 sg13g2_decap_8 FILLER_11_217 ();
 sg13g2_decap_8 FILLER_11_224 ();
 sg13g2_decap_8 FILLER_11_231 ();
 sg13g2_decap_8 FILLER_11_238 ();
 sg13g2_decap_8 FILLER_11_245 ();
 sg13g2_decap_8 FILLER_11_252 ();
 sg13g2_decap_8 FILLER_11_259 ();
 sg13g2_decap_8 FILLER_11_266 ();
 sg13g2_decap_8 FILLER_11_273 ();
 sg13g2_decap_8 FILLER_11_280 ();
 sg13g2_decap_8 FILLER_11_287 ();
 sg13g2_decap_8 FILLER_11_294 ();
 sg13g2_decap_8 FILLER_11_301 ();
 sg13g2_decap_8 FILLER_11_308 ();
 sg13g2_decap_8 FILLER_11_315 ();
 sg13g2_decap_8 FILLER_11_322 ();
 sg13g2_decap_8 FILLER_11_329 ();
 sg13g2_decap_8 FILLER_11_336 ();
 sg13g2_decap_8 FILLER_11_343 ();
 sg13g2_decap_8 FILLER_11_350 ();
 sg13g2_decap_8 FILLER_11_357 ();
 sg13g2_decap_8 FILLER_11_364 ();
 sg13g2_decap_8 FILLER_11_371 ();
 sg13g2_decap_8 FILLER_11_378 ();
 sg13g2_decap_8 FILLER_11_385 ();
 sg13g2_decap_8 FILLER_11_392 ();
 sg13g2_decap_8 FILLER_11_399 ();
 sg13g2_decap_8 FILLER_11_406 ();
 sg13g2_decap_8 FILLER_11_413 ();
 sg13g2_decap_8 FILLER_11_420 ();
 sg13g2_decap_8 FILLER_11_427 ();
 sg13g2_decap_8 FILLER_11_434 ();
 sg13g2_decap_8 FILLER_11_441 ();
 sg13g2_decap_8 FILLER_11_448 ();
 sg13g2_decap_8 FILLER_11_455 ();
 sg13g2_decap_8 FILLER_11_462 ();
 sg13g2_decap_8 FILLER_11_469 ();
 sg13g2_decap_8 FILLER_11_476 ();
 sg13g2_decap_8 FILLER_11_483 ();
 sg13g2_decap_8 FILLER_11_490 ();
 sg13g2_decap_8 FILLER_11_497 ();
 sg13g2_decap_8 FILLER_11_504 ();
 sg13g2_decap_8 FILLER_11_511 ();
 sg13g2_decap_8 FILLER_11_518 ();
 sg13g2_decap_8 FILLER_11_525 ();
 sg13g2_decap_8 FILLER_11_532 ();
 sg13g2_decap_8 FILLER_11_539 ();
 sg13g2_decap_8 FILLER_11_546 ();
 sg13g2_decap_8 FILLER_11_553 ();
 sg13g2_decap_8 FILLER_11_560 ();
 sg13g2_decap_8 FILLER_11_567 ();
 sg13g2_decap_8 FILLER_11_574 ();
 sg13g2_decap_8 FILLER_11_581 ();
 sg13g2_decap_8 FILLER_11_588 ();
 sg13g2_decap_8 FILLER_11_595 ();
 sg13g2_decap_8 FILLER_11_602 ();
 sg13g2_decap_8 FILLER_11_609 ();
 sg13g2_decap_8 FILLER_11_616 ();
 sg13g2_decap_8 FILLER_11_623 ();
 sg13g2_decap_8 FILLER_11_630 ();
 sg13g2_decap_8 FILLER_11_637 ();
 sg13g2_decap_8 FILLER_11_644 ();
 sg13g2_decap_8 FILLER_11_651 ();
 sg13g2_decap_8 FILLER_11_658 ();
 sg13g2_decap_8 FILLER_11_665 ();
 sg13g2_decap_8 FILLER_11_672 ();
 sg13g2_decap_8 FILLER_11_679 ();
 sg13g2_decap_8 FILLER_11_686 ();
 sg13g2_decap_8 FILLER_11_693 ();
 sg13g2_decap_8 FILLER_11_700 ();
 sg13g2_decap_8 FILLER_11_707 ();
 sg13g2_decap_8 FILLER_11_714 ();
 sg13g2_decap_8 FILLER_11_721 ();
 sg13g2_decap_8 FILLER_11_728 ();
 sg13g2_decap_8 FILLER_11_735 ();
 sg13g2_decap_8 FILLER_11_742 ();
 sg13g2_decap_8 FILLER_11_749 ();
 sg13g2_decap_8 FILLER_11_756 ();
 sg13g2_decap_8 FILLER_11_763 ();
 sg13g2_decap_8 FILLER_11_770 ();
 sg13g2_decap_8 FILLER_11_777 ();
 sg13g2_decap_8 FILLER_11_784 ();
 sg13g2_decap_8 FILLER_11_791 ();
 sg13g2_decap_8 FILLER_11_798 ();
 sg13g2_decap_8 FILLER_11_805 ();
 sg13g2_decap_8 FILLER_11_812 ();
 sg13g2_decap_8 FILLER_11_819 ();
 sg13g2_decap_8 FILLER_11_826 ();
 sg13g2_decap_8 FILLER_11_833 ();
 sg13g2_decap_8 FILLER_11_840 ();
 sg13g2_decap_8 FILLER_11_847 ();
 sg13g2_decap_8 FILLER_11_854 ();
 sg13g2_decap_8 FILLER_11_861 ();
 sg13g2_decap_8 FILLER_11_868 ();
 sg13g2_decap_8 FILLER_11_875 ();
 sg13g2_decap_8 FILLER_11_882 ();
 sg13g2_decap_8 FILLER_11_889 ();
 sg13g2_decap_8 FILLER_11_896 ();
 sg13g2_decap_8 FILLER_11_903 ();
 sg13g2_decap_8 FILLER_11_910 ();
 sg13g2_decap_8 FILLER_11_917 ();
 sg13g2_decap_8 FILLER_11_924 ();
 sg13g2_decap_8 FILLER_11_931 ();
 sg13g2_decap_8 FILLER_11_938 ();
 sg13g2_decap_8 FILLER_11_945 ();
 sg13g2_decap_8 FILLER_11_952 ();
 sg13g2_decap_8 FILLER_11_959 ();
 sg13g2_decap_8 FILLER_11_966 ();
 sg13g2_decap_8 FILLER_11_973 ();
 sg13g2_decap_8 FILLER_11_980 ();
 sg13g2_decap_8 FILLER_11_987 ();
 sg13g2_decap_8 FILLER_11_994 ();
 sg13g2_decap_8 FILLER_11_1001 ();
 sg13g2_decap_8 FILLER_11_1008 ();
 sg13g2_decap_8 FILLER_11_1015 ();
 sg13g2_decap_8 FILLER_11_1022 ();
 sg13g2_decap_8 FILLER_12_4 ();
 sg13g2_decap_8 FILLER_12_11 ();
 sg13g2_decap_8 FILLER_12_18 ();
 sg13g2_decap_8 FILLER_12_25 ();
 sg13g2_decap_8 FILLER_12_32 ();
 sg13g2_decap_8 FILLER_12_39 ();
 sg13g2_decap_8 FILLER_12_46 ();
 sg13g2_decap_8 FILLER_12_53 ();
 sg13g2_decap_8 FILLER_12_60 ();
 sg13g2_decap_8 FILLER_12_67 ();
 sg13g2_decap_8 FILLER_12_74 ();
 sg13g2_decap_8 FILLER_12_81 ();
 sg13g2_decap_8 FILLER_12_88 ();
 sg13g2_decap_8 FILLER_12_95 ();
 sg13g2_decap_8 FILLER_12_102 ();
 sg13g2_decap_8 FILLER_12_109 ();
 sg13g2_decap_8 FILLER_12_116 ();
 sg13g2_decap_8 FILLER_12_123 ();
 sg13g2_decap_8 FILLER_12_130 ();
 sg13g2_decap_8 FILLER_12_137 ();
 sg13g2_decap_8 FILLER_12_144 ();
 sg13g2_decap_8 FILLER_12_151 ();
 sg13g2_decap_8 FILLER_12_158 ();
 sg13g2_decap_8 FILLER_12_165 ();
 sg13g2_decap_8 FILLER_12_172 ();
 sg13g2_decap_8 FILLER_12_179 ();
 sg13g2_decap_8 FILLER_12_186 ();
 sg13g2_decap_8 FILLER_12_193 ();
 sg13g2_decap_8 FILLER_12_200 ();
 sg13g2_decap_8 FILLER_12_207 ();
 sg13g2_decap_8 FILLER_12_214 ();
 sg13g2_decap_8 FILLER_12_221 ();
 sg13g2_decap_8 FILLER_12_228 ();
 sg13g2_decap_8 FILLER_12_235 ();
 sg13g2_decap_8 FILLER_12_242 ();
 sg13g2_decap_8 FILLER_12_249 ();
 sg13g2_decap_8 FILLER_12_256 ();
 sg13g2_decap_8 FILLER_12_263 ();
 sg13g2_decap_8 FILLER_12_270 ();
 sg13g2_decap_8 FILLER_12_277 ();
 sg13g2_decap_8 FILLER_12_284 ();
 sg13g2_decap_8 FILLER_12_291 ();
 sg13g2_decap_8 FILLER_12_298 ();
 sg13g2_decap_8 FILLER_12_305 ();
 sg13g2_decap_8 FILLER_12_312 ();
 sg13g2_decap_8 FILLER_12_319 ();
 sg13g2_decap_8 FILLER_12_326 ();
 sg13g2_decap_8 FILLER_12_333 ();
 sg13g2_decap_8 FILLER_12_340 ();
 sg13g2_decap_8 FILLER_12_347 ();
 sg13g2_decap_8 FILLER_12_354 ();
 sg13g2_decap_8 FILLER_12_361 ();
 sg13g2_decap_8 FILLER_12_368 ();
 sg13g2_decap_8 FILLER_12_375 ();
 sg13g2_decap_8 FILLER_12_382 ();
 sg13g2_decap_8 FILLER_12_389 ();
 sg13g2_decap_8 FILLER_12_396 ();
 sg13g2_decap_8 FILLER_12_403 ();
 sg13g2_decap_8 FILLER_12_410 ();
 sg13g2_decap_8 FILLER_12_417 ();
 sg13g2_decap_8 FILLER_12_424 ();
 sg13g2_decap_8 FILLER_12_431 ();
 sg13g2_decap_8 FILLER_12_438 ();
 sg13g2_decap_8 FILLER_12_445 ();
 sg13g2_decap_8 FILLER_12_452 ();
 sg13g2_decap_8 FILLER_12_459 ();
 sg13g2_decap_8 FILLER_12_466 ();
 sg13g2_decap_8 FILLER_12_473 ();
 sg13g2_decap_8 FILLER_12_480 ();
 sg13g2_decap_8 FILLER_12_487 ();
 sg13g2_decap_8 FILLER_12_494 ();
 sg13g2_decap_8 FILLER_12_501 ();
 sg13g2_decap_8 FILLER_12_508 ();
 sg13g2_decap_8 FILLER_12_515 ();
 sg13g2_decap_8 FILLER_12_522 ();
 sg13g2_decap_8 FILLER_12_529 ();
 sg13g2_decap_8 FILLER_12_536 ();
 sg13g2_decap_8 FILLER_12_543 ();
 sg13g2_decap_8 FILLER_12_550 ();
 sg13g2_decap_8 FILLER_12_557 ();
 sg13g2_decap_8 FILLER_12_564 ();
 sg13g2_decap_8 FILLER_12_571 ();
 sg13g2_decap_8 FILLER_12_578 ();
 sg13g2_decap_8 FILLER_12_585 ();
 sg13g2_decap_8 FILLER_12_592 ();
 sg13g2_decap_8 FILLER_12_599 ();
 sg13g2_decap_8 FILLER_12_606 ();
 sg13g2_decap_8 FILLER_12_613 ();
 sg13g2_decap_8 FILLER_12_620 ();
 sg13g2_decap_8 FILLER_12_627 ();
 sg13g2_decap_8 FILLER_12_634 ();
 sg13g2_decap_8 FILLER_12_641 ();
 sg13g2_decap_8 FILLER_12_648 ();
 sg13g2_decap_8 FILLER_12_655 ();
 sg13g2_decap_8 FILLER_12_662 ();
 sg13g2_decap_8 FILLER_12_669 ();
 sg13g2_decap_8 FILLER_12_676 ();
 sg13g2_decap_8 FILLER_12_683 ();
 sg13g2_decap_8 FILLER_12_690 ();
 sg13g2_decap_8 FILLER_12_697 ();
 sg13g2_decap_8 FILLER_12_704 ();
 sg13g2_decap_8 FILLER_12_711 ();
 sg13g2_decap_8 FILLER_12_718 ();
 sg13g2_decap_8 FILLER_12_725 ();
 sg13g2_decap_8 FILLER_12_732 ();
 sg13g2_decap_8 FILLER_12_739 ();
 sg13g2_decap_8 FILLER_12_746 ();
 sg13g2_decap_8 FILLER_12_753 ();
 sg13g2_decap_8 FILLER_12_760 ();
 sg13g2_decap_8 FILLER_12_767 ();
 sg13g2_decap_8 FILLER_12_774 ();
 sg13g2_decap_8 FILLER_12_781 ();
 sg13g2_decap_8 FILLER_12_788 ();
 sg13g2_decap_8 FILLER_12_795 ();
 sg13g2_decap_8 FILLER_12_802 ();
 sg13g2_decap_8 FILLER_12_809 ();
 sg13g2_decap_8 FILLER_12_816 ();
 sg13g2_decap_8 FILLER_12_823 ();
 sg13g2_decap_8 FILLER_12_830 ();
 sg13g2_decap_8 FILLER_12_837 ();
 sg13g2_decap_8 FILLER_12_844 ();
 sg13g2_decap_8 FILLER_12_851 ();
 sg13g2_decap_8 FILLER_12_858 ();
 sg13g2_decap_8 FILLER_12_865 ();
 sg13g2_decap_8 FILLER_12_872 ();
 sg13g2_decap_8 FILLER_12_879 ();
 sg13g2_decap_8 FILLER_12_886 ();
 sg13g2_decap_8 FILLER_12_893 ();
 sg13g2_decap_8 FILLER_12_900 ();
 sg13g2_decap_8 FILLER_12_907 ();
 sg13g2_decap_8 FILLER_12_914 ();
 sg13g2_decap_8 FILLER_12_921 ();
 sg13g2_decap_8 FILLER_12_928 ();
 sg13g2_decap_8 FILLER_12_935 ();
 sg13g2_decap_8 FILLER_12_942 ();
 sg13g2_decap_8 FILLER_12_949 ();
 sg13g2_decap_8 FILLER_12_956 ();
 sg13g2_decap_8 FILLER_12_963 ();
 sg13g2_decap_8 FILLER_12_970 ();
 sg13g2_decap_8 FILLER_12_977 ();
 sg13g2_decap_8 FILLER_12_984 ();
 sg13g2_decap_8 FILLER_12_991 ();
 sg13g2_decap_8 FILLER_12_998 ();
 sg13g2_decap_8 FILLER_12_1005 ();
 sg13g2_decap_8 FILLER_12_1012 ();
 sg13g2_decap_8 FILLER_12_1019 ();
 sg13g2_fill_2 FILLER_12_1026 ();
 sg13g2_fill_1 FILLER_12_1028 ();
 sg13g2_decap_8 FILLER_13_0 ();
 sg13g2_decap_8 FILLER_13_7 ();
 sg13g2_decap_8 FILLER_13_14 ();
 sg13g2_decap_8 FILLER_13_21 ();
 sg13g2_decap_8 FILLER_13_28 ();
 sg13g2_decap_8 FILLER_13_35 ();
 sg13g2_decap_8 FILLER_13_42 ();
 sg13g2_decap_8 FILLER_13_49 ();
 sg13g2_decap_8 FILLER_13_56 ();
 sg13g2_decap_8 FILLER_13_63 ();
 sg13g2_decap_8 FILLER_13_70 ();
 sg13g2_decap_8 FILLER_13_77 ();
 sg13g2_decap_8 FILLER_13_84 ();
 sg13g2_decap_8 FILLER_13_91 ();
 sg13g2_decap_8 FILLER_13_98 ();
 sg13g2_decap_8 FILLER_13_105 ();
 sg13g2_decap_8 FILLER_13_112 ();
 sg13g2_decap_8 FILLER_13_119 ();
 sg13g2_decap_8 FILLER_13_126 ();
 sg13g2_decap_8 FILLER_13_133 ();
 sg13g2_decap_8 FILLER_13_140 ();
 sg13g2_decap_8 FILLER_13_147 ();
 sg13g2_decap_8 FILLER_13_154 ();
 sg13g2_decap_8 FILLER_13_161 ();
 sg13g2_decap_8 FILLER_13_168 ();
 sg13g2_decap_8 FILLER_13_175 ();
 sg13g2_decap_8 FILLER_13_182 ();
 sg13g2_decap_8 FILLER_13_189 ();
 sg13g2_decap_8 FILLER_13_196 ();
 sg13g2_decap_8 FILLER_13_203 ();
 sg13g2_decap_8 FILLER_13_210 ();
 sg13g2_decap_8 FILLER_13_217 ();
 sg13g2_decap_8 FILLER_13_224 ();
 sg13g2_decap_8 FILLER_13_231 ();
 sg13g2_decap_8 FILLER_13_238 ();
 sg13g2_decap_8 FILLER_13_245 ();
 sg13g2_decap_8 FILLER_13_252 ();
 sg13g2_decap_8 FILLER_13_259 ();
 sg13g2_decap_8 FILLER_13_266 ();
 sg13g2_decap_8 FILLER_13_273 ();
 sg13g2_decap_8 FILLER_13_280 ();
 sg13g2_decap_8 FILLER_13_287 ();
 sg13g2_decap_8 FILLER_13_294 ();
 sg13g2_decap_8 FILLER_13_301 ();
 sg13g2_decap_8 FILLER_13_308 ();
 sg13g2_decap_8 FILLER_13_315 ();
 sg13g2_decap_8 FILLER_13_322 ();
 sg13g2_decap_8 FILLER_13_329 ();
 sg13g2_decap_8 FILLER_13_336 ();
 sg13g2_decap_8 FILLER_13_343 ();
 sg13g2_decap_8 FILLER_13_350 ();
 sg13g2_decap_8 FILLER_13_357 ();
 sg13g2_decap_8 FILLER_13_364 ();
 sg13g2_decap_8 FILLER_13_371 ();
 sg13g2_decap_8 FILLER_13_378 ();
 sg13g2_decap_8 FILLER_13_385 ();
 sg13g2_decap_8 FILLER_13_392 ();
 sg13g2_decap_8 FILLER_13_399 ();
 sg13g2_decap_8 FILLER_13_406 ();
 sg13g2_decap_8 FILLER_13_413 ();
 sg13g2_decap_8 FILLER_13_420 ();
 sg13g2_decap_8 FILLER_13_427 ();
 sg13g2_decap_8 FILLER_13_434 ();
 sg13g2_decap_8 FILLER_13_441 ();
 sg13g2_decap_8 FILLER_13_448 ();
 sg13g2_decap_8 FILLER_13_455 ();
 sg13g2_decap_8 FILLER_13_462 ();
 sg13g2_decap_8 FILLER_13_469 ();
 sg13g2_decap_8 FILLER_13_476 ();
 sg13g2_decap_8 FILLER_13_483 ();
 sg13g2_decap_8 FILLER_13_490 ();
 sg13g2_decap_8 FILLER_13_497 ();
 sg13g2_decap_8 FILLER_13_504 ();
 sg13g2_decap_8 FILLER_13_511 ();
 sg13g2_decap_8 FILLER_13_518 ();
 sg13g2_decap_8 FILLER_13_525 ();
 sg13g2_decap_8 FILLER_13_532 ();
 sg13g2_decap_8 FILLER_13_539 ();
 sg13g2_decap_8 FILLER_13_546 ();
 sg13g2_decap_8 FILLER_13_553 ();
 sg13g2_decap_8 FILLER_13_560 ();
 sg13g2_decap_8 FILLER_13_567 ();
 sg13g2_decap_8 FILLER_13_574 ();
 sg13g2_decap_8 FILLER_13_581 ();
 sg13g2_decap_8 FILLER_13_588 ();
 sg13g2_decap_8 FILLER_13_595 ();
 sg13g2_decap_8 FILLER_13_602 ();
 sg13g2_decap_8 FILLER_13_609 ();
 sg13g2_decap_8 FILLER_13_616 ();
 sg13g2_decap_8 FILLER_13_623 ();
 sg13g2_decap_8 FILLER_13_630 ();
 sg13g2_decap_8 FILLER_13_637 ();
 sg13g2_decap_8 FILLER_13_644 ();
 sg13g2_decap_8 FILLER_13_651 ();
 sg13g2_decap_8 FILLER_13_658 ();
 sg13g2_decap_8 FILLER_13_665 ();
 sg13g2_decap_8 FILLER_13_672 ();
 sg13g2_decap_8 FILLER_13_679 ();
 sg13g2_decap_8 FILLER_13_686 ();
 sg13g2_decap_8 FILLER_13_693 ();
 sg13g2_decap_8 FILLER_13_700 ();
 sg13g2_decap_8 FILLER_13_707 ();
 sg13g2_decap_8 FILLER_13_714 ();
 sg13g2_decap_8 FILLER_13_721 ();
 sg13g2_decap_8 FILLER_13_728 ();
 sg13g2_decap_8 FILLER_13_735 ();
 sg13g2_decap_8 FILLER_13_742 ();
 sg13g2_decap_8 FILLER_13_749 ();
 sg13g2_decap_8 FILLER_13_756 ();
 sg13g2_decap_8 FILLER_13_763 ();
 sg13g2_decap_8 FILLER_13_770 ();
 sg13g2_decap_8 FILLER_13_777 ();
 sg13g2_decap_8 FILLER_13_784 ();
 sg13g2_decap_8 FILLER_13_791 ();
 sg13g2_decap_8 FILLER_13_798 ();
 sg13g2_decap_8 FILLER_13_805 ();
 sg13g2_decap_8 FILLER_13_812 ();
 sg13g2_decap_8 FILLER_13_819 ();
 sg13g2_decap_8 FILLER_13_826 ();
 sg13g2_decap_8 FILLER_13_833 ();
 sg13g2_decap_8 FILLER_13_840 ();
 sg13g2_decap_8 FILLER_13_847 ();
 sg13g2_decap_8 FILLER_13_854 ();
 sg13g2_decap_8 FILLER_13_861 ();
 sg13g2_decap_8 FILLER_13_868 ();
 sg13g2_decap_8 FILLER_13_875 ();
 sg13g2_decap_8 FILLER_13_882 ();
 sg13g2_decap_8 FILLER_13_889 ();
 sg13g2_decap_8 FILLER_13_896 ();
 sg13g2_decap_8 FILLER_13_903 ();
 sg13g2_decap_8 FILLER_13_910 ();
 sg13g2_decap_8 FILLER_13_917 ();
 sg13g2_decap_8 FILLER_13_924 ();
 sg13g2_decap_8 FILLER_13_931 ();
 sg13g2_decap_8 FILLER_13_938 ();
 sg13g2_decap_8 FILLER_13_945 ();
 sg13g2_decap_8 FILLER_13_952 ();
 sg13g2_decap_8 FILLER_13_959 ();
 sg13g2_decap_8 FILLER_13_966 ();
 sg13g2_decap_8 FILLER_13_973 ();
 sg13g2_decap_8 FILLER_13_980 ();
 sg13g2_decap_8 FILLER_13_987 ();
 sg13g2_decap_8 FILLER_13_994 ();
 sg13g2_decap_8 FILLER_13_1001 ();
 sg13g2_decap_8 FILLER_13_1008 ();
 sg13g2_decap_8 FILLER_13_1015 ();
 sg13g2_decap_8 FILLER_13_1022 ();
 sg13g2_decap_8 FILLER_14_0 ();
 sg13g2_decap_8 FILLER_14_7 ();
 sg13g2_decap_8 FILLER_14_14 ();
 sg13g2_decap_8 FILLER_14_21 ();
 sg13g2_decap_8 FILLER_14_28 ();
 sg13g2_decap_8 FILLER_14_35 ();
 sg13g2_decap_8 FILLER_14_42 ();
 sg13g2_decap_8 FILLER_14_49 ();
 sg13g2_decap_8 FILLER_14_56 ();
 sg13g2_decap_8 FILLER_14_63 ();
 sg13g2_decap_8 FILLER_14_70 ();
 sg13g2_decap_8 FILLER_14_77 ();
 sg13g2_decap_8 FILLER_14_84 ();
 sg13g2_decap_8 FILLER_14_91 ();
 sg13g2_decap_8 FILLER_14_98 ();
 sg13g2_decap_8 FILLER_14_105 ();
 sg13g2_decap_8 FILLER_14_112 ();
 sg13g2_decap_8 FILLER_14_119 ();
 sg13g2_decap_8 FILLER_14_126 ();
 sg13g2_decap_8 FILLER_14_133 ();
 sg13g2_decap_8 FILLER_14_140 ();
 sg13g2_decap_8 FILLER_14_147 ();
 sg13g2_decap_8 FILLER_14_154 ();
 sg13g2_decap_8 FILLER_14_161 ();
 sg13g2_decap_8 FILLER_14_168 ();
 sg13g2_decap_8 FILLER_14_175 ();
 sg13g2_decap_8 FILLER_14_182 ();
 sg13g2_decap_8 FILLER_14_189 ();
 sg13g2_decap_8 FILLER_14_196 ();
 sg13g2_decap_8 FILLER_14_203 ();
 sg13g2_decap_8 FILLER_14_210 ();
 sg13g2_decap_8 FILLER_14_217 ();
 sg13g2_decap_8 FILLER_14_224 ();
 sg13g2_decap_8 FILLER_14_231 ();
 sg13g2_decap_8 FILLER_14_238 ();
 sg13g2_decap_8 FILLER_14_245 ();
 sg13g2_decap_8 FILLER_14_252 ();
 sg13g2_decap_8 FILLER_14_259 ();
 sg13g2_decap_8 FILLER_14_266 ();
 sg13g2_decap_8 FILLER_14_273 ();
 sg13g2_decap_8 FILLER_14_280 ();
 sg13g2_decap_8 FILLER_14_287 ();
 sg13g2_decap_8 FILLER_14_294 ();
 sg13g2_decap_8 FILLER_14_301 ();
 sg13g2_decap_8 FILLER_14_308 ();
 sg13g2_decap_8 FILLER_14_315 ();
 sg13g2_decap_8 FILLER_14_322 ();
 sg13g2_decap_8 FILLER_14_329 ();
 sg13g2_decap_8 FILLER_14_336 ();
 sg13g2_decap_8 FILLER_14_343 ();
 sg13g2_decap_8 FILLER_14_350 ();
 sg13g2_decap_8 FILLER_14_357 ();
 sg13g2_decap_8 FILLER_14_364 ();
 sg13g2_decap_8 FILLER_14_371 ();
 sg13g2_decap_8 FILLER_14_378 ();
 sg13g2_decap_8 FILLER_14_385 ();
 sg13g2_decap_8 FILLER_14_392 ();
 sg13g2_decap_8 FILLER_14_399 ();
 sg13g2_decap_8 FILLER_14_406 ();
 sg13g2_decap_8 FILLER_14_413 ();
 sg13g2_decap_8 FILLER_14_420 ();
 sg13g2_decap_8 FILLER_14_427 ();
 sg13g2_decap_8 FILLER_14_434 ();
 sg13g2_decap_8 FILLER_14_441 ();
 sg13g2_decap_8 FILLER_14_448 ();
 sg13g2_decap_8 FILLER_14_455 ();
 sg13g2_decap_8 FILLER_14_462 ();
 sg13g2_decap_8 FILLER_14_469 ();
 sg13g2_decap_8 FILLER_14_476 ();
 sg13g2_decap_8 FILLER_14_483 ();
 sg13g2_decap_8 FILLER_14_490 ();
 sg13g2_decap_8 FILLER_14_497 ();
 sg13g2_decap_8 FILLER_14_504 ();
 sg13g2_decap_8 FILLER_14_511 ();
 sg13g2_decap_8 FILLER_14_518 ();
 sg13g2_decap_8 FILLER_14_525 ();
 sg13g2_decap_8 FILLER_14_532 ();
 sg13g2_decap_8 FILLER_14_539 ();
 sg13g2_decap_8 FILLER_14_546 ();
 sg13g2_decap_8 FILLER_14_553 ();
 sg13g2_decap_8 FILLER_14_560 ();
 sg13g2_decap_8 FILLER_14_567 ();
 sg13g2_decap_8 FILLER_14_574 ();
 sg13g2_decap_8 FILLER_14_581 ();
 sg13g2_decap_8 FILLER_14_588 ();
 sg13g2_decap_8 FILLER_14_595 ();
 sg13g2_decap_8 FILLER_14_602 ();
 sg13g2_decap_8 FILLER_14_609 ();
 sg13g2_decap_8 FILLER_14_616 ();
 sg13g2_decap_8 FILLER_14_623 ();
 sg13g2_decap_8 FILLER_14_630 ();
 sg13g2_decap_8 FILLER_14_637 ();
 sg13g2_decap_8 FILLER_14_644 ();
 sg13g2_decap_8 FILLER_14_651 ();
 sg13g2_decap_8 FILLER_14_658 ();
 sg13g2_decap_8 FILLER_14_665 ();
 sg13g2_decap_8 FILLER_14_672 ();
 sg13g2_decap_8 FILLER_14_679 ();
 sg13g2_decap_8 FILLER_14_686 ();
 sg13g2_decap_8 FILLER_14_693 ();
 sg13g2_decap_8 FILLER_14_700 ();
 sg13g2_decap_8 FILLER_14_707 ();
 sg13g2_decap_8 FILLER_14_714 ();
 sg13g2_decap_8 FILLER_14_721 ();
 sg13g2_decap_8 FILLER_14_728 ();
 sg13g2_decap_8 FILLER_14_735 ();
 sg13g2_decap_8 FILLER_14_742 ();
 sg13g2_decap_8 FILLER_14_749 ();
 sg13g2_decap_8 FILLER_14_756 ();
 sg13g2_decap_8 FILLER_14_763 ();
 sg13g2_decap_8 FILLER_14_770 ();
 sg13g2_decap_8 FILLER_14_777 ();
 sg13g2_decap_8 FILLER_14_784 ();
 sg13g2_decap_8 FILLER_14_791 ();
 sg13g2_decap_8 FILLER_14_798 ();
 sg13g2_decap_8 FILLER_14_805 ();
 sg13g2_decap_8 FILLER_14_812 ();
 sg13g2_decap_8 FILLER_14_819 ();
 sg13g2_decap_8 FILLER_14_826 ();
 sg13g2_decap_8 FILLER_14_833 ();
 sg13g2_decap_8 FILLER_14_840 ();
 sg13g2_decap_8 FILLER_14_847 ();
 sg13g2_decap_8 FILLER_14_854 ();
 sg13g2_decap_8 FILLER_14_861 ();
 sg13g2_decap_8 FILLER_14_868 ();
 sg13g2_decap_8 FILLER_14_875 ();
 sg13g2_decap_8 FILLER_14_882 ();
 sg13g2_decap_8 FILLER_14_889 ();
 sg13g2_decap_8 FILLER_14_896 ();
 sg13g2_decap_8 FILLER_14_903 ();
 sg13g2_decap_8 FILLER_14_910 ();
 sg13g2_decap_8 FILLER_14_917 ();
 sg13g2_decap_8 FILLER_14_924 ();
 sg13g2_decap_8 FILLER_14_931 ();
 sg13g2_decap_8 FILLER_14_938 ();
 sg13g2_decap_8 FILLER_14_945 ();
 sg13g2_decap_8 FILLER_14_952 ();
 sg13g2_decap_8 FILLER_14_959 ();
 sg13g2_decap_8 FILLER_14_966 ();
 sg13g2_decap_8 FILLER_14_973 ();
 sg13g2_decap_8 FILLER_14_980 ();
 sg13g2_decap_8 FILLER_14_987 ();
 sg13g2_decap_8 FILLER_14_994 ();
 sg13g2_decap_8 FILLER_14_1001 ();
 sg13g2_decap_8 FILLER_14_1008 ();
 sg13g2_decap_8 FILLER_14_1015 ();
 sg13g2_decap_8 FILLER_14_1022 ();
 sg13g2_decap_8 FILLER_15_4 ();
 sg13g2_decap_8 FILLER_15_11 ();
 sg13g2_decap_8 FILLER_15_18 ();
 sg13g2_decap_8 FILLER_15_25 ();
 sg13g2_decap_8 FILLER_15_32 ();
 sg13g2_decap_8 FILLER_15_39 ();
 sg13g2_decap_8 FILLER_15_46 ();
 sg13g2_decap_8 FILLER_15_53 ();
 sg13g2_decap_8 FILLER_15_60 ();
 sg13g2_decap_8 FILLER_15_67 ();
 sg13g2_decap_8 FILLER_15_74 ();
 sg13g2_decap_8 FILLER_15_81 ();
 sg13g2_decap_8 FILLER_15_88 ();
 sg13g2_decap_8 FILLER_15_95 ();
 sg13g2_decap_8 FILLER_15_102 ();
 sg13g2_decap_8 FILLER_15_109 ();
 sg13g2_decap_8 FILLER_15_116 ();
 sg13g2_decap_8 FILLER_15_123 ();
 sg13g2_decap_8 FILLER_15_130 ();
 sg13g2_decap_8 FILLER_15_137 ();
 sg13g2_decap_8 FILLER_15_144 ();
 sg13g2_decap_8 FILLER_15_151 ();
 sg13g2_decap_8 FILLER_15_158 ();
 sg13g2_decap_8 FILLER_15_165 ();
 sg13g2_decap_8 FILLER_15_172 ();
 sg13g2_decap_8 FILLER_15_179 ();
 sg13g2_decap_8 FILLER_15_186 ();
 sg13g2_decap_8 FILLER_15_193 ();
 sg13g2_decap_8 FILLER_15_200 ();
 sg13g2_decap_8 FILLER_15_207 ();
 sg13g2_decap_8 FILLER_15_214 ();
 sg13g2_decap_8 FILLER_15_221 ();
 sg13g2_decap_8 FILLER_15_228 ();
 sg13g2_decap_8 FILLER_15_235 ();
 sg13g2_decap_8 FILLER_15_242 ();
 sg13g2_decap_8 FILLER_15_249 ();
 sg13g2_decap_8 FILLER_15_256 ();
 sg13g2_decap_8 FILLER_15_263 ();
 sg13g2_decap_8 FILLER_15_270 ();
 sg13g2_decap_8 FILLER_15_277 ();
 sg13g2_decap_8 FILLER_15_284 ();
 sg13g2_decap_8 FILLER_15_291 ();
 sg13g2_decap_8 FILLER_15_298 ();
 sg13g2_decap_8 FILLER_15_305 ();
 sg13g2_decap_8 FILLER_15_312 ();
 sg13g2_decap_8 FILLER_15_319 ();
 sg13g2_decap_8 FILLER_15_326 ();
 sg13g2_decap_8 FILLER_15_333 ();
 sg13g2_decap_8 FILLER_15_340 ();
 sg13g2_decap_8 FILLER_15_347 ();
 sg13g2_decap_8 FILLER_15_354 ();
 sg13g2_decap_8 FILLER_15_361 ();
 sg13g2_decap_8 FILLER_15_368 ();
 sg13g2_decap_8 FILLER_15_375 ();
 sg13g2_decap_8 FILLER_15_382 ();
 sg13g2_decap_8 FILLER_15_389 ();
 sg13g2_decap_8 FILLER_15_396 ();
 sg13g2_decap_8 FILLER_15_403 ();
 sg13g2_decap_8 FILLER_15_410 ();
 sg13g2_decap_8 FILLER_15_417 ();
 sg13g2_decap_8 FILLER_15_424 ();
 sg13g2_decap_8 FILLER_15_431 ();
 sg13g2_decap_8 FILLER_15_438 ();
 sg13g2_decap_8 FILLER_15_445 ();
 sg13g2_decap_8 FILLER_15_452 ();
 sg13g2_decap_8 FILLER_15_459 ();
 sg13g2_decap_8 FILLER_15_466 ();
 sg13g2_decap_8 FILLER_15_473 ();
 sg13g2_decap_8 FILLER_15_480 ();
 sg13g2_decap_8 FILLER_15_487 ();
 sg13g2_decap_8 FILLER_15_494 ();
 sg13g2_decap_8 FILLER_15_501 ();
 sg13g2_decap_8 FILLER_15_508 ();
 sg13g2_decap_8 FILLER_15_515 ();
 sg13g2_decap_8 FILLER_15_522 ();
 sg13g2_decap_8 FILLER_15_529 ();
 sg13g2_decap_8 FILLER_15_536 ();
 sg13g2_decap_8 FILLER_15_543 ();
 sg13g2_decap_8 FILLER_15_550 ();
 sg13g2_decap_8 FILLER_15_557 ();
 sg13g2_decap_8 FILLER_15_564 ();
 sg13g2_decap_8 FILLER_15_571 ();
 sg13g2_decap_8 FILLER_15_578 ();
 sg13g2_decap_8 FILLER_15_585 ();
 sg13g2_decap_8 FILLER_15_592 ();
 sg13g2_decap_8 FILLER_15_599 ();
 sg13g2_decap_8 FILLER_15_606 ();
 sg13g2_decap_8 FILLER_15_613 ();
 sg13g2_decap_8 FILLER_15_620 ();
 sg13g2_decap_8 FILLER_15_627 ();
 sg13g2_decap_8 FILLER_15_634 ();
 sg13g2_decap_8 FILLER_15_641 ();
 sg13g2_decap_8 FILLER_15_648 ();
 sg13g2_decap_8 FILLER_15_655 ();
 sg13g2_decap_8 FILLER_15_662 ();
 sg13g2_decap_8 FILLER_15_669 ();
 sg13g2_decap_8 FILLER_15_676 ();
 sg13g2_decap_8 FILLER_15_683 ();
 sg13g2_decap_8 FILLER_15_690 ();
 sg13g2_decap_8 FILLER_15_697 ();
 sg13g2_decap_8 FILLER_15_704 ();
 sg13g2_decap_8 FILLER_15_711 ();
 sg13g2_decap_8 FILLER_15_718 ();
 sg13g2_decap_8 FILLER_15_725 ();
 sg13g2_decap_8 FILLER_15_732 ();
 sg13g2_decap_8 FILLER_15_739 ();
 sg13g2_decap_8 FILLER_15_746 ();
 sg13g2_decap_8 FILLER_15_753 ();
 sg13g2_decap_8 FILLER_15_760 ();
 sg13g2_decap_8 FILLER_15_767 ();
 sg13g2_decap_8 FILLER_15_774 ();
 sg13g2_decap_8 FILLER_15_781 ();
 sg13g2_decap_8 FILLER_15_788 ();
 sg13g2_decap_8 FILLER_15_795 ();
 sg13g2_decap_8 FILLER_15_802 ();
 sg13g2_decap_8 FILLER_15_809 ();
 sg13g2_decap_8 FILLER_15_816 ();
 sg13g2_decap_8 FILLER_15_823 ();
 sg13g2_decap_8 FILLER_15_830 ();
 sg13g2_decap_8 FILLER_15_837 ();
 sg13g2_decap_8 FILLER_15_844 ();
 sg13g2_decap_8 FILLER_15_851 ();
 sg13g2_decap_8 FILLER_15_858 ();
 sg13g2_decap_8 FILLER_15_865 ();
 sg13g2_decap_8 FILLER_15_872 ();
 sg13g2_decap_8 FILLER_15_879 ();
 sg13g2_decap_8 FILLER_15_886 ();
 sg13g2_decap_8 FILLER_15_893 ();
 sg13g2_decap_8 FILLER_15_900 ();
 sg13g2_decap_8 FILLER_15_907 ();
 sg13g2_decap_8 FILLER_15_914 ();
 sg13g2_decap_8 FILLER_15_921 ();
 sg13g2_decap_8 FILLER_15_928 ();
 sg13g2_decap_8 FILLER_15_935 ();
 sg13g2_decap_8 FILLER_15_942 ();
 sg13g2_decap_8 FILLER_15_949 ();
 sg13g2_decap_8 FILLER_15_956 ();
 sg13g2_decap_8 FILLER_15_963 ();
 sg13g2_decap_8 FILLER_15_970 ();
 sg13g2_decap_8 FILLER_15_977 ();
 sg13g2_decap_8 FILLER_15_984 ();
 sg13g2_decap_8 FILLER_15_991 ();
 sg13g2_decap_8 FILLER_15_998 ();
 sg13g2_decap_8 FILLER_15_1005 ();
 sg13g2_decap_8 FILLER_15_1012 ();
 sg13g2_decap_8 FILLER_15_1019 ();
 sg13g2_fill_2 FILLER_15_1026 ();
 sg13g2_fill_1 FILLER_15_1028 ();
 sg13g2_decap_8 FILLER_16_0 ();
 sg13g2_decap_8 FILLER_16_7 ();
 sg13g2_decap_8 FILLER_16_14 ();
 sg13g2_decap_8 FILLER_16_21 ();
 sg13g2_decap_8 FILLER_16_28 ();
 sg13g2_decap_8 FILLER_16_35 ();
 sg13g2_decap_8 FILLER_16_42 ();
 sg13g2_decap_8 FILLER_16_49 ();
 sg13g2_decap_8 FILLER_16_56 ();
 sg13g2_decap_8 FILLER_16_63 ();
 sg13g2_decap_8 FILLER_16_70 ();
 sg13g2_decap_8 FILLER_16_77 ();
 sg13g2_decap_8 FILLER_16_84 ();
 sg13g2_decap_8 FILLER_16_91 ();
 sg13g2_decap_8 FILLER_16_98 ();
 sg13g2_decap_8 FILLER_16_105 ();
 sg13g2_decap_8 FILLER_16_112 ();
 sg13g2_decap_8 FILLER_16_119 ();
 sg13g2_decap_8 FILLER_16_126 ();
 sg13g2_decap_8 FILLER_16_133 ();
 sg13g2_decap_8 FILLER_16_140 ();
 sg13g2_decap_8 FILLER_16_147 ();
 sg13g2_decap_8 FILLER_16_154 ();
 sg13g2_decap_8 FILLER_16_161 ();
 sg13g2_decap_8 FILLER_16_168 ();
 sg13g2_decap_8 FILLER_16_175 ();
 sg13g2_decap_8 FILLER_16_182 ();
 sg13g2_decap_8 FILLER_16_189 ();
 sg13g2_decap_8 FILLER_16_196 ();
 sg13g2_decap_8 FILLER_16_203 ();
 sg13g2_decap_8 FILLER_16_210 ();
 sg13g2_decap_8 FILLER_16_217 ();
 sg13g2_decap_8 FILLER_16_224 ();
 sg13g2_decap_8 FILLER_16_231 ();
 sg13g2_decap_8 FILLER_16_238 ();
 sg13g2_decap_8 FILLER_16_245 ();
 sg13g2_decap_8 FILLER_16_252 ();
 sg13g2_decap_8 FILLER_16_259 ();
 sg13g2_decap_8 FILLER_16_266 ();
 sg13g2_decap_8 FILLER_16_273 ();
 sg13g2_decap_8 FILLER_16_280 ();
 sg13g2_decap_8 FILLER_16_287 ();
 sg13g2_decap_8 FILLER_16_294 ();
 sg13g2_decap_8 FILLER_16_301 ();
 sg13g2_decap_8 FILLER_16_308 ();
 sg13g2_decap_8 FILLER_16_315 ();
 sg13g2_decap_8 FILLER_16_322 ();
 sg13g2_decap_8 FILLER_16_329 ();
 sg13g2_decap_8 FILLER_16_336 ();
 sg13g2_decap_8 FILLER_16_343 ();
 sg13g2_decap_8 FILLER_16_350 ();
 sg13g2_decap_8 FILLER_16_357 ();
 sg13g2_decap_8 FILLER_16_364 ();
 sg13g2_decap_8 FILLER_16_371 ();
 sg13g2_decap_8 FILLER_16_378 ();
 sg13g2_decap_8 FILLER_16_385 ();
 sg13g2_decap_8 FILLER_16_392 ();
 sg13g2_decap_8 FILLER_16_399 ();
 sg13g2_decap_8 FILLER_16_406 ();
 sg13g2_decap_8 FILLER_16_413 ();
 sg13g2_decap_8 FILLER_16_420 ();
 sg13g2_decap_8 FILLER_16_427 ();
 sg13g2_decap_8 FILLER_16_434 ();
 sg13g2_decap_8 FILLER_16_441 ();
 sg13g2_decap_8 FILLER_16_448 ();
 sg13g2_decap_8 FILLER_16_455 ();
 sg13g2_decap_8 FILLER_16_462 ();
 sg13g2_decap_8 FILLER_16_469 ();
 sg13g2_decap_8 FILLER_16_476 ();
 sg13g2_decap_8 FILLER_16_483 ();
 sg13g2_decap_8 FILLER_16_490 ();
 sg13g2_decap_8 FILLER_16_497 ();
 sg13g2_decap_8 FILLER_16_504 ();
 sg13g2_decap_8 FILLER_16_511 ();
 sg13g2_decap_8 FILLER_16_518 ();
 sg13g2_decap_8 FILLER_16_525 ();
 sg13g2_decap_8 FILLER_16_532 ();
 sg13g2_decap_8 FILLER_16_539 ();
 sg13g2_decap_8 FILLER_16_546 ();
 sg13g2_decap_8 FILLER_16_553 ();
 sg13g2_decap_8 FILLER_16_560 ();
 sg13g2_decap_8 FILLER_16_567 ();
 sg13g2_decap_8 FILLER_16_574 ();
 sg13g2_decap_8 FILLER_16_581 ();
 sg13g2_decap_8 FILLER_16_588 ();
 sg13g2_decap_8 FILLER_16_595 ();
 sg13g2_decap_8 FILLER_16_602 ();
 sg13g2_decap_8 FILLER_16_609 ();
 sg13g2_decap_8 FILLER_16_616 ();
 sg13g2_decap_8 FILLER_16_623 ();
 sg13g2_decap_8 FILLER_16_630 ();
 sg13g2_decap_8 FILLER_16_637 ();
 sg13g2_decap_8 FILLER_16_644 ();
 sg13g2_decap_8 FILLER_16_651 ();
 sg13g2_decap_8 FILLER_16_658 ();
 sg13g2_decap_8 FILLER_16_665 ();
 sg13g2_decap_8 FILLER_16_672 ();
 sg13g2_decap_8 FILLER_16_679 ();
 sg13g2_decap_8 FILLER_16_686 ();
 sg13g2_decap_8 FILLER_16_693 ();
 sg13g2_decap_8 FILLER_16_700 ();
 sg13g2_decap_8 FILLER_16_707 ();
 sg13g2_decap_8 FILLER_16_714 ();
 sg13g2_decap_8 FILLER_16_721 ();
 sg13g2_decap_8 FILLER_16_728 ();
 sg13g2_decap_8 FILLER_16_735 ();
 sg13g2_decap_8 FILLER_16_742 ();
 sg13g2_decap_8 FILLER_16_749 ();
 sg13g2_decap_8 FILLER_16_756 ();
 sg13g2_decap_8 FILLER_16_763 ();
 sg13g2_decap_8 FILLER_16_770 ();
 sg13g2_decap_8 FILLER_16_777 ();
 sg13g2_decap_8 FILLER_16_784 ();
 sg13g2_decap_8 FILLER_16_791 ();
 sg13g2_decap_8 FILLER_16_798 ();
 sg13g2_decap_8 FILLER_16_805 ();
 sg13g2_decap_8 FILLER_16_812 ();
 sg13g2_decap_8 FILLER_16_819 ();
 sg13g2_decap_8 FILLER_16_826 ();
 sg13g2_decap_8 FILLER_16_833 ();
 sg13g2_decap_8 FILLER_16_840 ();
 sg13g2_decap_8 FILLER_16_847 ();
 sg13g2_decap_8 FILLER_16_854 ();
 sg13g2_decap_8 FILLER_16_861 ();
 sg13g2_decap_8 FILLER_16_868 ();
 sg13g2_decap_8 FILLER_16_875 ();
 sg13g2_decap_8 FILLER_16_882 ();
 sg13g2_decap_8 FILLER_16_889 ();
 sg13g2_decap_8 FILLER_16_896 ();
 sg13g2_decap_8 FILLER_16_903 ();
 sg13g2_decap_8 FILLER_16_910 ();
 sg13g2_decap_8 FILLER_16_917 ();
 sg13g2_decap_8 FILLER_16_924 ();
 sg13g2_decap_8 FILLER_16_931 ();
 sg13g2_decap_8 FILLER_16_938 ();
 sg13g2_decap_8 FILLER_16_945 ();
 sg13g2_decap_8 FILLER_16_952 ();
 sg13g2_decap_8 FILLER_16_959 ();
 sg13g2_decap_8 FILLER_16_966 ();
 sg13g2_decap_8 FILLER_16_973 ();
 sg13g2_decap_8 FILLER_16_980 ();
 sg13g2_decap_8 FILLER_16_987 ();
 sg13g2_decap_8 FILLER_16_994 ();
 sg13g2_decap_8 FILLER_16_1001 ();
 sg13g2_decap_8 FILLER_16_1008 ();
 sg13g2_decap_8 FILLER_16_1015 ();
 sg13g2_decap_8 FILLER_16_1022 ();
 sg13g2_decap_8 FILLER_17_4 ();
 sg13g2_decap_8 FILLER_17_11 ();
 sg13g2_decap_8 FILLER_17_18 ();
 sg13g2_decap_8 FILLER_17_25 ();
 sg13g2_decap_8 FILLER_17_32 ();
 sg13g2_decap_8 FILLER_17_39 ();
 sg13g2_decap_8 FILLER_17_46 ();
 sg13g2_decap_8 FILLER_17_53 ();
 sg13g2_decap_8 FILLER_17_60 ();
 sg13g2_decap_8 FILLER_17_67 ();
 sg13g2_decap_8 FILLER_17_74 ();
 sg13g2_decap_8 FILLER_17_81 ();
 sg13g2_decap_8 FILLER_17_88 ();
 sg13g2_decap_8 FILLER_17_95 ();
 sg13g2_decap_8 FILLER_17_102 ();
 sg13g2_decap_8 FILLER_17_109 ();
 sg13g2_decap_8 FILLER_17_116 ();
 sg13g2_decap_8 FILLER_17_123 ();
 sg13g2_decap_8 FILLER_17_130 ();
 sg13g2_decap_8 FILLER_17_137 ();
 sg13g2_decap_8 FILLER_17_144 ();
 sg13g2_decap_8 FILLER_17_151 ();
 sg13g2_decap_8 FILLER_17_158 ();
 sg13g2_decap_8 FILLER_17_165 ();
 sg13g2_decap_8 FILLER_17_172 ();
 sg13g2_decap_8 FILLER_17_179 ();
 sg13g2_decap_8 FILLER_17_186 ();
 sg13g2_decap_8 FILLER_17_193 ();
 sg13g2_decap_8 FILLER_17_200 ();
 sg13g2_decap_8 FILLER_17_207 ();
 sg13g2_decap_8 FILLER_17_214 ();
 sg13g2_decap_8 FILLER_17_221 ();
 sg13g2_decap_8 FILLER_17_228 ();
 sg13g2_decap_8 FILLER_17_235 ();
 sg13g2_decap_8 FILLER_17_242 ();
 sg13g2_decap_8 FILLER_17_249 ();
 sg13g2_decap_8 FILLER_17_256 ();
 sg13g2_decap_8 FILLER_17_263 ();
 sg13g2_decap_8 FILLER_17_270 ();
 sg13g2_decap_8 FILLER_17_277 ();
 sg13g2_decap_8 FILLER_17_284 ();
 sg13g2_decap_8 FILLER_17_291 ();
 sg13g2_decap_8 FILLER_17_298 ();
 sg13g2_decap_8 FILLER_17_305 ();
 sg13g2_decap_8 FILLER_17_312 ();
 sg13g2_decap_8 FILLER_17_319 ();
 sg13g2_decap_8 FILLER_17_326 ();
 sg13g2_decap_8 FILLER_17_333 ();
 sg13g2_decap_8 FILLER_17_340 ();
 sg13g2_decap_8 FILLER_17_347 ();
 sg13g2_decap_8 FILLER_17_354 ();
 sg13g2_decap_8 FILLER_17_361 ();
 sg13g2_decap_8 FILLER_17_368 ();
 sg13g2_decap_8 FILLER_17_375 ();
 sg13g2_decap_8 FILLER_17_382 ();
 sg13g2_decap_8 FILLER_17_389 ();
 sg13g2_decap_8 FILLER_17_396 ();
 sg13g2_decap_8 FILLER_17_403 ();
 sg13g2_decap_8 FILLER_17_410 ();
 sg13g2_decap_8 FILLER_17_417 ();
 sg13g2_decap_8 FILLER_17_424 ();
 sg13g2_decap_8 FILLER_17_431 ();
 sg13g2_decap_8 FILLER_17_438 ();
 sg13g2_decap_8 FILLER_17_445 ();
 sg13g2_decap_8 FILLER_17_452 ();
 sg13g2_decap_8 FILLER_17_459 ();
 sg13g2_decap_8 FILLER_17_466 ();
 sg13g2_decap_8 FILLER_17_473 ();
 sg13g2_decap_8 FILLER_17_480 ();
 sg13g2_decap_8 FILLER_17_487 ();
 sg13g2_decap_8 FILLER_17_494 ();
 sg13g2_decap_8 FILLER_17_501 ();
 sg13g2_decap_8 FILLER_17_508 ();
 sg13g2_decap_8 FILLER_17_515 ();
 sg13g2_decap_8 FILLER_17_522 ();
 sg13g2_decap_8 FILLER_17_529 ();
 sg13g2_decap_8 FILLER_17_536 ();
 sg13g2_decap_8 FILLER_17_543 ();
 sg13g2_decap_8 FILLER_17_550 ();
 sg13g2_decap_8 FILLER_17_557 ();
 sg13g2_decap_8 FILLER_17_564 ();
 sg13g2_decap_8 FILLER_17_571 ();
 sg13g2_decap_8 FILLER_17_578 ();
 sg13g2_decap_8 FILLER_17_585 ();
 sg13g2_decap_8 FILLER_17_592 ();
 sg13g2_decap_8 FILLER_17_599 ();
 sg13g2_decap_8 FILLER_17_606 ();
 sg13g2_decap_8 FILLER_17_613 ();
 sg13g2_decap_8 FILLER_17_620 ();
 sg13g2_decap_8 FILLER_17_627 ();
 sg13g2_decap_8 FILLER_17_634 ();
 sg13g2_decap_8 FILLER_17_641 ();
 sg13g2_decap_8 FILLER_17_648 ();
 sg13g2_decap_8 FILLER_17_655 ();
 sg13g2_decap_8 FILLER_17_662 ();
 sg13g2_decap_8 FILLER_17_669 ();
 sg13g2_decap_8 FILLER_17_676 ();
 sg13g2_decap_8 FILLER_17_683 ();
 sg13g2_decap_8 FILLER_17_690 ();
 sg13g2_decap_8 FILLER_17_697 ();
 sg13g2_decap_8 FILLER_17_704 ();
 sg13g2_decap_8 FILLER_17_711 ();
 sg13g2_decap_8 FILLER_17_718 ();
 sg13g2_decap_8 FILLER_17_725 ();
 sg13g2_decap_8 FILLER_17_732 ();
 sg13g2_decap_8 FILLER_17_739 ();
 sg13g2_decap_8 FILLER_17_746 ();
 sg13g2_decap_8 FILLER_17_753 ();
 sg13g2_decap_8 FILLER_17_760 ();
 sg13g2_decap_8 FILLER_17_767 ();
 sg13g2_decap_8 FILLER_17_774 ();
 sg13g2_decap_8 FILLER_17_781 ();
 sg13g2_decap_8 FILLER_17_788 ();
 sg13g2_decap_8 FILLER_17_795 ();
 sg13g2_decap_8 FILLER_17_802 ();
 sg13g2_decap_8 FILLER_17_809 ();
 sg13g2_decap_8 FILLER_17_816 ();
 sg13g2_decap_8 FILLER_17_823 ();
 sg13g2_decap_8 FILLER_17_830 ();
 sg13g2_decap_8 FILLER_17_837 ();
 sg13g2_decap_8 FILLER_17_844 ();
 sg13g2_decap_8 FILLER_17_851 ();
 sg13g2_decap_8 FILLER_17_858 ();
 sg13g2_decap_8 FILLER_17_865 ();
 sg13g2_decap_8 FILLER_17_872 ();
 sg13g2_decap_8 FILLER_17_879 ();
 sg13g2_decap_8 FILLER_17_886 ();
 sg13g2_decap_8 FILLER_17_893 ();
 sg13g2_decap_8 FILLER_17_900 ();
 sg13g2_decap_8 FILLER_17_907 ();
 sg13g2_decap_8 FILLER_17_914 ();
 sg13g2_decap_8 FILLER_17_921 ();
 sg13g2_decap_8 FILLER_17_928 ();
 sg13g2_decap_8 FILLER_17_935 ();
 sg13g2_decap_8 FILLER_17_942 ();
 sg13g2_decap_8 FILLER_17_949 ();
 sg13g2_decap_8 FILLER_17_956 ();
 sg13g2_decap_8 FILLER_17_963 ();
 sg13g2_decap_8 FILLER_17_970 ();
 sg13g2_decap_8 FILLER_17_977 ();
 sg13g2_decap_8 FILLER_17_984 ();
 sg13g2_decap_8 FILLER_17_991 ();
 sg13g2_decap_8 FILLER_17_998 ();
 sg13g2_decap_8 FILLER_17_1005 ();
 sg13g2_decap_8 FILLER_17_1012 ();
 sg13g2_decap_8 FILLER_17_1019 ();
 sg13g2_fill_2 FILLER_17_1026 ();
 sg13g2_fill_1 FILLER_17_1028 ();
 sg13g2_decap_8 FILLER_18_0 ();
 sg13g2_decap_8 FILLER_18_7 ();
 sg13g2_decap_8 FILLER_18_14 ();
 sg13g2_decap_8 FILLER_18_21 ();
 sg13g2_decap_8 FILLER_18_28 ();
 sg13g2_decap_8 FILLER_18_35 ();
 sg13g2_decap_8 FILLER_18_42 ();
 sg13g2_decap_8 FILLER_18_49 ();
 sg13g2_decap_8 FILLER_18_56 ();
 sg13g2_decap_8 FILLER_18_63 ();
 sg13g2_decap_8 FILLER_18_70 ();
 sg13g2_decap_8 FILLER_18_77 ();
 sg13g2_decap_8 FILLER_18_84 ();
 sg13g2_decap_8 FILLER_18_91 ();
 sg13g2_decap_8 FILLER_18_98 ();
 sg13g2_decap_8 FILLER_18_105 ();
 sg13g2_decap_8 FILLER_18_112 ();
 sg13g2_decap_8 FILLER_18_119 ();
 sg13g2_decap_8 FILLER_18_126 ();
 sg13g2_decap_8 FILLER_18_133 ();
 sg13g2_decap_8 FILLER_18_140 ();
 sg13g2_decap_8 FILLER_18_147 ();
 sg13g2_decap_8 FILLER_18_154 ();
 sg13g2_decap_8 FILLER_18_161 ();
 sg13g2_decap_8 FILLER_18_168 ();
 sg13g2_decap_8 FILLER_18_175 ();
 sg13g2_decap_8 FILLER_18_182 ();
 sg13g2_decap_8 FILLER_18_189 ();
 sg13g2_decap_8 FILLER_18_196 ();
 sg13g2_decap_8 FILLER_18_203 ();
 sg13g2_decap_8 FILLER_18_210 ();
 sg13g2_decap_8 FILLER_18_217 ();
 sg13g2_decap_8 FILLER_18_224 ();
 sg13g2_decap_8 FILLER_18_231 ();
 sg13g2_decap_8 FILLER_18_238 ();
 sg13g2_decap_8 FILLER_18_245 ();
 sg13g2_decap_8 FILLER_18_252 ();
 sg13g2_decap_8 FILLER_18_259 ();
 sg13g2_decap_8 FILLER_18_266 ();
 sg13g2_decap_8 FILLER_18_273 ();
 sg13g2_decap_8 FILLER_18_280 ();
 sg13g2_decap_8 FILLER_18_287 ();
 sg13g2_decap_8 FILLER_18_294 ();
 sg13g2_decap_8 FILLER_18_301 ();
 sg13g2_decap_8 FILLER_18_308 ();
 sg13g2_decap_8 FILLER_18_315 ();
 sg13g2_decap_8 FILLER_18_322 ();
 sg13g2_decap_8 FILLER_18_329 ();
 sg13g2_decap_8 FILLER_18_336 ();
 sg13g2_decap_8 FILLER_18_343 ();
 sg13g2_decap_8 FILLER_18_350 ();
 sg13g2_decap_8 FILLER_18_357 ();
 sg13g2_decap_8 FILLER_18_364 ();
 sg13g2_decap_8 FILLER_18_371 ();
 sg13g2_decap_8 FILLER_18_378 ();
 sg13g2_decap_8 FILLER_18_385 ();
 sg13g2_decap_8 FILLER_18_392 ();
 sg13g2_decap_8 FILLER_18_399 ();
 sg13g2_decap_8 FILLER_18_406 ();
 sg13g2_decap_8 FILLER_18_413 ();
 sg13g2_decap_8 FILLER_18_420 ();
 sg13g2_decap_8 FILLER_18_427 ();
 sg13g2_decap_8 FILLER_18_434 ();
 sg13g2_decap_8 FILLER_18_441 ();
 sg13g2_decap_8 FILLER_18_448 ();
 sg13g2_decap_8 FILLER_18_455 ();
 sg13g2_decap_8 FILLER_18_462 ();
 sg13g2_decap_8 FILLER_18_469 ();
 sg13g2_decap_8 FILLER_18_476 ();
 sg13g2_decap_8 FILLER_18_483 ();
 sg13g2_decap_8 FILLER_18_490 ();
 sg13g2_decap_8 FILLER_18_497 ();
 sg13g2_decap_8 FILLER_18_504 ();
 sg13g2_decap_8 FILLER_18_511 ();
 sg13g2_decap_8 FILLER_18_518 ();
 sg13g2_decap_8 FILLER_18_525 ();
 sg13g2_decap_8 FILLER_18_532 ();
 sg13g2_decap_8 FILLER_18_539 ();
 sg13g2_decap_8 FILLER_18_546 ();
 sg13g2_decap_8 FILLER_18_553 ();
 sg13g2_decap_8 FILLER_18_560 ();
 sg13g2_decap_8 FILLER_18_567 ();
 sg13g2_decap_8 FILLER_18_574 ();
 sg13g2_decap_8 FILLER_18_581 ();
 sg13g2_decap_8 FILLER_18_588 ();
 sg13g2_decap_8 FILLER_18_595 ();
 sg13g2_decap_8 FILLER_18_602 ();
 sg13g2_decap_8 FILLER_18_609 ();
 sg13g2_decap_8 FILLER_18_616 ();
 sg13g2_decap_8 FILLER_18_623 ();
 sg13g2_decap_8 FILLER_18_630 ();
 sg13g2_decap_8 FILLER_18_637 ();
 sg13g2_decap_8 FILLER_18_644 ();
 sg13g2_decap_8 FILLER_18_651 ();
 sg13g2_decap_8 FILLER_18_658 ();
 sg13g2_decap_8 FILLER_18_665 ();
 sg13g2_decap_8 FILLER_18_672 ();
 sg13g2_decap_8 FILLER_18_679 ();
 sg13g2_decap_8 FILLER_18_686 ();
 sg13g2_decap_8 FILLER_18_693 ();
 sg13g2_decap_8 FILLER_18_700 ();
 sg13g2_decap_8 FILLER_18_707 ();
 sg13g2_decap_8 FILLER_18_714 ();
 sg13g2_decap_8 FILLER_18_721 ();
 sg13g2_decap_8 FILLER_18_728 ();
 sg13g2_decap_8 FILLER_18_735 ();
 sg13g2_decap_8 FILLER_18_742 ();
 sg13g2_decap_8 FILLER_18_749 ();
 sg13g2_decap_8 FILLER_18_756 ();
 sg13g2_decap_8 FILLER_18_763 ();
 sg13g2_decap_8 FILLER_18_770 ();
 sg13g2_decap_8 FILLER_18_777 ();
 sg13g2_decap_8 FILLER_18_784 ();
 sg13g2_decap_8 FILLER_18_791 ();
 sg13g2_decap_8 FILLER_18_798 ();
 sg13g2_decap_8 FILLER_18_805 ();
 sg13g2_decap_8 FILLER_18_812 ();
 sg13g2_decap_8 FILLER_18_819 ();
 sg13g2_decap_8 FILLER_18_826 ();
 sg13g2_decap_8 FILLER_18_833 ();
 sg13g2_decap_8 FILLER_18_840 ();
 sg13g2_decap_8 FILLER_18_847 ();
 sg13g2_decap_8 FILLER_18_854 ();
 sg13g2_decap_8 FILLER_18_861 ();
 sg13g2_decap_8 FILLER_18_868 ();
 sg13g2_decap_8 FILLER_18_875 ();
 sg13g2_decap_8 FILLER_18_882 ();
 sg13g2_decap_8 FILLER_18_889 ();
 sg13g2_decap_8 FILLER_18_896 ();
 sg13g2_decap_8 FILLER_18_903 ();
 sg13g2_decap_8 FILLER_18_910 ();
 sg13g2_decap_8 FILLER_18_917 ();
 sg13g2_decap_8 FILLER_18_924 ();
 sg13g2_decap_8 FILLER_18_931 ();
 sg13g2_decap_8 FILLER_18_938 ();
 sg13g2_decap_8 FILLER_18_945 ();
 sg13g2_decap_8 FILLER_18_952 ();
 sg13g2_decap_8 FILLER_18_959 ();
 sg13g2_decap_8 FILLER_18_966 ();
 sg13g2_decap_8 FILLER_18_973 ();
 sg13g2_decap_8 FILLER_18_980 ();
 sg13g2_decap_8 FILLER_18_987 ();
 sg13g2_decap_8 FILLER_18_994 ();
 sg13g2_decap_8 FILLER_18_1001 ();
 sg13g2_decap_8 FILLER_18_1008 ();
 sg13g2_decap_8 FILLER_18_1015 ();
 sg13g2_decap_8 FILLER_18_1022 ();
 sg13g2_decap_8 FILLER_19_0 ();
 sg13g2_decap_8 FILLER_19_7 ();
 sg13g2_decap_8 FILLER_19_14 ();
 sg13g2_decap_8 FILLER_19_21 ();
 sg13g2_decap_8 FILLER_19_28 ();
 sg13g2_decap_8 FILLER_19_35 ();
 sg13g2_decap_8 FILLER_19_42 ();
 sg13g2_decap_8 FILLER_19_49 ();
 sg13g2_decap_8 FILLER_19_56 ();
 sg13g2_decap_8 FILLER_19_63 ();
 sg13g2_decap_8 FILLER_19_70 ();
 sg13g2_decap_8 FILLER_19_77 ();
 sg13g2_decap_8 FILLER_19_84 ();
 sg13g2_decap_8 FILLER_19_91 ();
 sg13g2_decap_8 FILLER_19_98 ();
 sg13g2_decap_8 FILLER_19_105 ();
 sg13g2_decap_8 FILLER_19_112 ();
 sg13g2_decap_8 FILLER_19_119 ();
 sg13g2_decap_8 FILLER_19_126 ();
 sg13g2_decap_8 FILLER_19_133 ();
 sg13g2_decap_8 FILLER_19_140 ();
 sg13g2_decap_8 FILLER_19_147 ();
 sg13g2_decap_8 FILLER_19_154 ();
 sg13g2_decap_8 FILLER_19_161 ();
 sg13g2_decap_8 FILLER_19_168 ();
 sg13g2_decap_8 FILLER_19_175 ();
 sg13g2_decap_8 FILLER_19_182 ();
 sg13g2_decap_8 FILLER_19_189 ();
 sg13g2_decap_8 FILLER_19_196 ();
 sg13g2_decap_8 FILLER_19_203 ();
 sg13g2_decap_8 FILLER_19_210 ();
 sg13g2_decap_8 FILLER_19_217 ();
 sg13g2_decap_8 FILLER_19_224 ();
 sg13g2_decap_8 FILLER_19_231 ();
 sg13g2_decap_8 FILLER_19_238 ();
 sg13g2_decap_8 FILLER_19_245 ();
 sg13g2_decap_8 FILLER_19_252 ();
 sg13g2_decap_8 FILLER_19_259 ();
 sg13g2_decap_8 FILLER_19_266 ();
 sg13g2_decap_8 FILLER_19_273 ();
 sg13g2_decap_8 FILLER_19_280 ();
 sg13g2_decap_8 FILLER_19_287 ();
 sg13g2_decap_8 FILLER_19_294 ();
 sg13g2_decap_8 FILLER_19_301 ();
 sg13g2_decap_8 FILLER_19_308 ();
 sg13g2_decap_8 FILLER_19_315 ();
 sg13g2_decap_8 FILLER_19_322 ();
 sg13g2_decap_8 FILLER_19_329 ();
 sg13g2_decap_8 FILLER_19_336 ();
 sg13g2_decap_8 FILLER_19_343 ();
 sg13g2_decap_8 FILLER_19_350 ();
 sg13g2_decap_8 FILLER_19_357 ();
 sg13g2_decap_8 FILLER_19_364 ();
 sg13g2_decap_8 FILLER_19_371 ();
 sg13g2_decap_8 FILLER_19_378 ();
 sg13g2_decap_8 FILLER_19_385 ();
 sg13g2_decap_8 FILLER_19_392 ();
 sg13g2_decap_8 FILLER_19_399 ();
 sg13g2_decap_8 FILLER_19_406 ();
 sg13g2_decap_8 FILLER_19_413 ();
 sg13g2_decap_8 FILLER_19_420 ();
 sg13g2_decap_8 FILLER_19_427 ();
 sg13g2_decap_8 FILLER_19_434 ();
 sg13g2_decap_8 FILLER_19_441 ();
 sg13g2_decap_8 FILLER_19_448 ();
 sg13g2_decap_8 FILLER_19_455 ();
 sg13g2_decap_8 FILLER_19_462 ();
 sg13g2_decap_8 FILLER_19_469 ();
 sg13g2_decap_8 FILLER_19_476 ();
 sg13g2_decap_8 FILLER_19_483 ();
 sg13g2_decap_8 FILLER_19_490 ();
 sg13g2_decap_8 FILLER_19_497 ();
 sg13g2_decap_8 FILLER_19_504 ();
 sg13g2_decap_8 FILLER_19_511 ();
 sg13g2_decap_8 FILLER_19_518 ();
 sg13g2_decap_8 FILLER_19_525 ();
 sg13g2_decap_8 FILLER_19_532 ();
 sg13g2_decap_8 FILLER_19_539 ();
 sg13g2_decap_8 FILLER_19_546 ();
 sg13g2_decap_8 FILLER_19_553 ();
 sg13g2_decap_8 FILLER_19_560 ();
 sg13g2_decap_8 FILLER_19_567 ();
 sg13g2_decap_8 FILLER_19_574 ();
 sg13g2_decap_8 FILLER_19_581 ();
 sg13g2_decap_8 FILLER_19_588 ();
 sg13g2_decap_8 FILLER_19_595 ();
 sg13g2_decap_8 FILLER_19_602 ();
 sg13g2_decap_8 FILLER_19_609 ();
 sg13g2_decap_8 FILLER_19_616 ();
 sg13g2_decap_8 FILLER_19_623 ();
 sg13g2_decap_8 FILLER_19_630 ();
 sg13g2_decap_8 FILLER_19_637 ();
 sg13g2_decap_8 FILLER_19_644 ();
 sg13g2_decap_8 FILLER_19_651 ();
 sg13g2_decap_8 FILLER_19_658 ();
 sg13g2_decap_8 FILLER_19_665 ();
 sg13g2_decap_8 FILLER_19_672 ();
 sg13g2_decap_8 FILLER_19_679 ();
 sg13g2_decap_8 FILLER_19_686 ();
 sg13g2_decap_8 FILLER_19_693 ();
 sg13g2_decap_8 FILLER_19_700 ();
 sg13g2_decap_8 FILLER_19_707 ();
 sg13g2_decap_8 FILLER_19_714 ();
 sg13g2_decap_8 FILLER_19_721 ();
 sg13g2_decap_8 FILLER_19_728 ();
 sg13g2_decap_8 FILLER_19_735 ();
 sg13g2_decap_8 FILLER_19_742 ();
 sg13g2_decap_8 FILLER_19_749 ();
 sg13g2_decap_8 FILLER_19_756 ();
 sg13g2_decap_8 FILLER_19_763 ();
 sg13g2_decap_8 FILLER_19_770 ();
 sg13g2_decap_8 FILLER_19_777 ();
 sg13g2_decap_8 FILLER_19_784 ();
 sg13g2_decap_8 FILLER_19_791 ();
 sg13g2_decap_8 FILLER_19_798 ();
 sg13g2_decap_8 FILLER_19_805 ();
 sg13g2_decap_8 FILLER_19_812 ();
 sg13g2_decap_8 FILLER_19_819 ();
 sg13g2_decap_8 FILLER_19_826 ();
 sg13g2_decap_8 FILLER_19_833 ();
 sg13g2_decap_8 FILLER_19_840 ();
 sg13g2_decap_8 FILLER_19_847 ();
 sg13g2_decap_8 FILLER_19_854 ();
 sg13g2_decap_8 FILLER_19_861 ();
 sg13g2_decap_8 FILLER_19_868 ();
 sg13g2_decap_8 FILLER_19_875 ();
 sg13g2_decap_8 FILLER_19_882 ();
 sg13g2_decap_8 FILLER_19_889 ();
 sg13g2_decap_8 FILLER_19_896 ();
 sg13g2_decap_8 FILLER_19_903 ();
 sg13g2_decap_8 FILLER_19_910 ();
 sg13g2_decap_8 FILLER_19_917 ();
 sg13g2_decap_8 FILLER_19_924 ();
 sg13g2_decap_8 FILLER_19_931 ();
 sg13g2_decap_8 FILLER_19_938 ();
 sg13g2_decap_8 FILLER_19_945 ();
 sg13g2_decap_8 FILLER_19_952 ();
 sg13g2_decap_8 FILLER_19_959 ();
 sg13g2_decap_8 FILLER_19_966 ();
 sg13g2_decap_8 FILLER_19_973 ();
 sg13g2_decap_8 FILLER_19_980 ();
 sg13g2_decap_8 FILLER_19_987 ();
 sg13g2_decap_8 FILLER_19_994 ();
 sg13g2_decap_8 FILLER_19_1001 ();
 sg13g2_decap_8 FILLER_19_1008 ();
 sg13g2_decap_8 FILLER_19_1015 ();
 sg13g2_decap_8 FILLER_19_1022 ();
 sg13g2_decap_8 FILLER_20_4 ();
 sg13g2_decap_8 FILLER_20_11 ();
 sg13g2_decap_8 FILLER_20_18 ();
 sg13g2_decap_8 FILLER_20_25 ();
 sg13g2_decap_8 FILLER_20_32 ();
 sg13g2_decap_8 FILLER_20_39 ();
 sg13g2_decap_8 FILLER_20_46 ();
 sg13g2_decap_8 FILLER_20_53 ();
 sg13g2_decap_8 FILLER_20_60 ();
 sg13g2_decap_8 FILLER_20_67 ();
 sg13g2_decap_8 FILLER_20_74 ();
 sg13g2_decap_8 FILLER_20_81 ();
 sg13g2_decap_8 FILLER_20_88 ();
 sg13g2_decap_8 FILLER_20_95 ();
 sg13g2_decap_8 FILLER_20_102 ();
 sg13g2_decap_8 FILLER_20_109 ();
 sg13g2_decap_8 FILLER_20_116 ();
 sg13g2_decap_8 FILLER_20_123 ();
 sg13g2_decap_8 FILLER_20_130 ();
 sg13g2_decap_8 FILLER_20_137 ();
 sg13g2_decap_8 FILLER_20_144 ();
 sg13g2_decap_8 FILLER_20_151 ();
 sg13g2_decap_8 FILLER_20_158 ();
 sg13g2_decap_8 FILLER_20_165 ();
 sg13g2_decap_8 FILLER_20_172 ();
 sg13g2_decap_8 FILLER_20_179 ();
 sg13g2_decap_8 FILLER_20_186 ();
 sg13g2_decap_8 FILLER_20_193 ();
 sg13g2_decap_8 FILLER_20_200 ();
 sg13g2_decap_8 FILLER_20_207 ();
 sg13g2_decap_8 FILLER_20_214 ();
 sg13g2_decap_8 FILLER_20_221 ();
 sg13g2_decap_8 FILLER_20_228 ();
 sg13g2_decap_8 FILLER_20_235 ();
 sg13g2_decap_8 FILLER_20_242 ();
 sg13g2_decap_8 FILLER_20_249 ();
 sg13g2_decap_8 FILLER_20_256 ();
 sg13g2_decap_8 FILLER_20_263 ();
 sg13g2_decap_8 FILLER_20_270 ();
 sg13g2_decap_8 FILLER_20_277 ();
 sg13g2_decap_8 FILLER_20_284 ();
 sg13g2_decap_8 FILLER_20_291 ();
 sg13g2_decap_8 FILLER_20_298 ();
 sg13g2_decap_8 FILLER_20_305 ();
 sg13g2_decap_8 FILLER_20_312 ();
 sg13g2_decap_8 FILLER_20_319 ();
 sg13g2_decap_8 FILLER_20_326 ();
 sg13g2_decap_8 FILLER_20_333 ();
 sg13g2_decap_8 FILLER_20_340 ();
 sg13g2_decap_8 FILLER_20_347 ();
 sg13g2_decap_8 FILLER_20_354 ();
 sg13g2_decap_8 FILLER_20_361 ();
 sg13g2_decap_8 FILLER_20_368 ();
 sg13g2_decap_8 FILLER_20_375 ();
 sg13g2_decap_8 FILLER_20_382 ();
 sg13g2_decap_8 FILLER_20_389 ();
 sg13g2_decap_8 FILLER_20_396 ();
 sg13g2_decap_8 FILLER_20_403 ();
 sg13g2_decap_8 FILLER_20_410 ();
 sg13g2_decap_8 FILLER_20_417 ();
 sg13g2_decap_8 FILLER_20_424 ();
 sg13g2_decap_8 FILLER_20_431 ();
 sg13g2_decap_8 FILLER_20_438 ();
 sg13g2_decap_8 FILLER_20_445 ();
 sg13g2_decap_8 FILLER_20_452 ();
 sg13g2_decap_8 FILLER_20_459 ();
 sg13g2_decap_8 FILLER_20_466 ();
 sg13g2_decap_8 FILLER_20_473 ();
 sg13g2_decap_8 FILLER_20_480 ();
 sg13g2_decap_8 FILLER_20_487 ();
 sg13g2_decap_8 FILLER_20_494 ();
 sg13g2_decap_8 FILLER_20_501 ();
 sg13g2_decap_8 FILLER_20_508 ();
 sg13g2_decap_8 FILLER_20_515 ();
 sg13g2_decap_8 FILLER_20_522 ();
 sg13g2_decap_8 FILLER_20_529 ();
 sg13g2_decap_8 FILLER_20_536 ();
 sg13g2_decap_8 FILLER_20_543 ();
 sg13g2_decap_8 FILLER_20_550 ();
 sg13g2_decap_8 FILLER_20_557 ();
 sg13g2_decap_8 FILLER_20_564 ();
 sg13g2_decap_8 FILLER_20_571 ();
 sg13g2_decap_8 FILLER_20_578 ();
 sg13g2_decap_8 FILLER_20_585 ();
 sg13g2_decap_8 FILLER_20_592 ();
 sg13g2_decap_8 FILLER_20_599 ();
 sg13g2_decap_8 FILLER_20_606 ();
 sg13g2_decap_8 FILLER_20_613 ();
 sg13g2_decap_8 FILLER_20_620 ();
 sg13g2_decap_8 FILLER_20_627 ();
 sg13g2_decap_8 FILLER_20_634 ();
 sg13g2_decap_8 FILLER_20_641 ();
 sg13g2_decap_8 FILLER_20_648 ();
 sg13g2_decap_8 FILLER_20_655 ();
 sg13g2_decap_8 FILLER_20_662 ();
 sg13g2_decap_8 FILLER_20_669 ();
 sg13g2_decap_8 FILLER_20_676 ();
 sg13g2_decap_8 FILLER_20_683 ();
 sg13g2_decap_8 FILLER_20_690 ();
 sg13g2_decap_8 FILLER_20_697 ();
 sg13g2_decap_8 FILLER_20_704 ();
 sg13g2_decap_8 FILLER_20_711 ();
 sg13g2_decap_8 FILLER_20_718 ();
 sg13g2_decap_8 FILLER_20_725 ();
 sg13g2_decap_8 FILLER_20_732 ();
 sg13g2_decap_8 FILLER_20_739 ();
 sg13g2_decap_8 FILLER_20_746 ();
 sg13g2_decap_8 FILLER_20_753 ();
 sg13g2_decap_8 FILLER_20_760 ();
 sg13g2_decap_8 FILLER_20_767 ();
 sg13g2_decap_8 FILLER_20_774 ();
 sg13g2_decap_8 FILLER_20_781 ();
 sg13g2_decap_8 FILLER_20_788 ();
 sg13g2_decap_8 FILLER_20_795 ();
 sg13g2_decap_8 FILLER_20_802 ();
 sg13g2_decap_8 FILLER_20_809 ();
 sg13g2_decap_8 FILLER_20_816 ();
 sg13g2_decap_8 FILLER_20_823 ();
 sg13g2_decap_8 FILLER_20_830 ();
 sg13g2_decap_8 FILLER_20_837 ();
 sg13g2_decap_8 FILLER_20_844 ();
 sg13g2_decap_8 FILLER_20_851 ();
 sg13g2_decap_8 FILLER_20_858 ();
 sg13g2_decap_8 FILLER_20_865 ();
 sg13g2_decap_8 FILLER_20_872 ();
 sg13g2_decap_8 FILLER_20_879 ();
 sg13g2_decap_8 FILLER_20_886 ();
 sg13g2_decap_8 FILLER_20_893 ();
 sg13g2_decap_8 FILLER_20_900 ();
 sg13g2_decap_8 FILLER_20_907 ();
 sg13g2_decap_8 FILLER_20_914 ();
 sg13g2_decap_8 FILLER_20_921 ();
 sg13g2_decap_8 FILLER_20_928 ();
 sg13g2_decap_8 FILLER_20_935 ();
 sg13g2_decap_8 FILLER_20_942 ();
 sg13g2_decap_8 FILLER_20_949 ();
 sg13g2_decap_8 FILLER_20_956 ();
 sg13g2_decap_8 FILLER_20_963 ();
 sg13g2_decap_8 FILLER_20_970 ();
 sg13g2_decap_8 FILLER_20_977 ();
 sg13g2_decap_8 FILLER_20_984 ();
 sg13g2_decap_8 FILLER_20_991 ();
 sg13g2_decap_8 FILLER_20_998 ();
 sg13g2_decap_8 FILLER_20_1005 ();
 sg13g2_decap_8 FILLER_20_1012 ();
 sg13g2_decap_8 FILLER_20_1019 ();
 sg13g2_fill_2 FILLER_20_1026 ();
 sg13g2_fill_1 FILLER_20_1028 ();
 sg13g2_decap_8 FILLER_21_0 ();
 sg13g2_decap_8 FILLER_21_7 ();
 sg13g2_decap_8 FILLER_21_14 ();
 sg13g2_decap_8 FILLER_21_21 ();
 sg13g2_decap_8 FILLER_21_28 ();
 sg13g2_decap_8 FILLER_21_35 ();
 sg13g2_decap_8 FILLER_21_42 ();
 sg13g2_decap_8 FILLER_21_49 ();
 sg13g2_decap_8 FILLER_21_56 ();
 sg13g2_decap_8 FILLER_21_63 ();
 sg13g2_decap_8 FILLER_21_70 ();
 sg13g2_decap_8 FILLER_21_77 ();
 sg13g2_decap_8 FILLER_21_84 ();
 sg13g2_decap_8 FILLER_21_91 ();
 sg13g2_decap_8 FILLER_21_98 ();
 sg13g2_decap_8 FILLER_21_105 ();
 sg13g2_decap_8 FILLER_21_112 ();
 sg13g2_decap_8 FILLER_21_119 ();
 sg13g2_decap_8 FILLER_21_126 ();
 sg13g2_decap_8 FILLER_21_133 ();
 sg13g2_decap_8 FILLER_21_140 ();
 sg13g2_decap_8 FILLER_21_147 ();
 sg13g2_decap_8 FILLER_21_154 ();
 sg13g2_decap_8 FILLER_21_161 ();
 sg13g2_decap_8 FILLER_21_168 ();
 sg13g2_decap_8 FILLER_21_175 ();
 sg13g2_decap_8 FILLER_21_182 ();
 sg13g2_decap_8 FILLER_21_189 ();
 sg13g2_decap_8 FILLER_21_196 ();
 sg13g2_decap_8 FILLER_21_203 ();
 sg13g2_decap_8 FILLER_21_210 ();
 sg13g2_decap_8 FILLER_21_217 ();
 sg13g2_decap_8 FILLER_21_224 ();
 sg13g2_decap_8 FILLER_21_231 ();
 sg13g2_decap_8 FILLER_21_238 ();
 sg13g2_decap_8 FILLER_21_245 ();
 sg13g2_decap_8 FILLER_21_252 ();
 sg13g2_decap_8 FILLER_21_259 ();
 sg13g2_decap_8 FILLER_21_266 ();
 sg13g2_decap_8 FILLER_21_273 ();
 sg13g2_decap_8 FILLER_21_280 ();
 sg13g2_decap_8 FILLER_21_287 ();
 sg13g2_decap_8 FILLER_21_294 ();
 sg13g2_decap_8 FILLER_21_301 ();
 sg13g2_decap_8 FILLER_21_308 ();
 sg13g2_decap_8 FILLER_21_315 ();
 sg13g2_decap_8 FILLER_21_322 ();
 sg13g2_decap_8 FILLER_21_329 ();
 sg13g2_decap_8 FILLER_21_336 ();
 sg13g2_decap_8 FILLER_21_343 ();
 sg13g2_decap_8 FILLER_21_350 ();
 sg13g2_decap_8 FILLER_21_357 ();
 sg13g2_decap_8 FILLER_21_364 ();
 sg13g2_decap_8 FILLER_21_371 ();
 sg13g2_decap_8 FILLER_21_378 ();
 sg13g2_decap_8 FILLER_21_385 ();
 sg13g2_decap_8 FILLER_21_392 ();
 sg13g2_decap_8 FILLER_21_399 ();
 sg13g2_decap_8 FILLER_21_406 ();
 sg13g2_decap_8 FILLER_21_413 ();
 sg13g2_decap_8 FILLER_21_420 ();
 sg13g2_decap_8 FILLER_21_427 ();
 sg13g2_decap_8 FILLER_21_434 ();
 sg13g2_decap_8 FILLER_21_441 ();
 sg13g2_decap_8 FILLER_21_448 ();
 sg13g2_decap_8 FILLER_21_455 ();
 sg13g2_decap_8 FILLER_21_462 ();
 sg13g2_decap_8 FILLER_21_469 ();
 sg13g2_decap_8 FILLER_21_476 ();
 sg13g2_decap_8 FILLER_21_483 ();
 sg13g2_decap_8 FILLER_21_490 ();
 sg13g2_decap_8 FILLER_21_497 ();
 sg13g2_decap_8 FILLER_21_504 ();
 sg13g2_decap_8 FILLER_21_511 ();
 sg13g2_decap_8 FILLER_21_518 ();
 sg13g2_decap_8 FILLER_21_525 ();
 sg13g2_decap_8 FILLER_21_532 ();
 sg13g2_decap_8 FILLER_21_539 ();
 sg13g2_decap_8 FILLER_21_546 ();
 sg13g2_decap_8 FILLER_21_553 ();
 sg13g2_decap_8 FILLER_21_560 ();
 sg13g2_decap_8 FILLER_21_567 ();
 sg13g2_decap_8 FILLER_21_574 ();
 sg13g2_decap_8 FILLER_21_581 ();
 sg13g2_decap_8 FILLER_21_588 ();
 sg13g2_decap_8 FILLER_21_595 ();
 sg13g2_decap_8 FILLER_21_602 ();
 sg13g2_decap_8 FILLER_21_609 ();
 sg13g2_decap_8 FILLER_21_616 ();
 sg13g2_decap_8 FILLER_21_623 ();
 sg13g2_decap_8 FILLER_21_630 ();
 sg13g2_decap_8 FILLER_21_637 ();
 sg13g2_decap_8 FILLER_21_644 ();
 sg13g2_decap_8 FILLER_21_651 ();
 sg13g2_decap_8 FILLER_21_658 ();
 sg13g2_decap_8 FILLER_21_665 ();
 sg13g2_decap_8 FILLER_21_672 ();
 sg13g2_decap_8 FILLER_21_679 ();
 sg13g2_decap_8 FILLER_21_686 ();
 sg13g2_decap_8 FILLER_21_693 ();
 sg13g2_decap_8 FILLER_21_700 ();
 sg13g2_decap_8 FILLER_21_707 ();
 sg13g2_decap_8 FILLER_21_714 ();
 sg13g2_decap_8 FILLER_21_721 ();
 sg13g2_decap_8 FILLER_21_728 ();
 sg13g2_decap_8 FILLER_21_735 ();
 sg13g2_decap_8 FILLER_21_742 ();
 sg13g2_decap_8 FILLER_21_749 ();
 sg13g2_decap_8 FILLER_21_756 ();
 sg13g2_decap_8 FILLER_21_763 ();
 sg13g2_decap_8 FILLER_21_770 ();
 sg13g2_decap_8 FILLER_21_777 ();
 sg13g2_decap_8 FILLER_21_784 ();
 sg13g2_decap_8 FILLER_21_791 ();
 sg13g2_decap_8 FILLER_21_798 ();
 sg13g2_decap_8 FILLER_21_805 ();
 sg13g2_decap_8 FILLER_21_812 ();
 sg13g2_decap_8 FILLER_21_819 ();
 sg13g2_decap_8 FILLER_21_826 ();
 sg13g2_decap_8 FILLER_21_833 ();
 sg13g2_decap_8 FILLER_21_840 ();
 sg13g2_decap_8 FILLER_21_847 ();
 sg13g2_decap_8 FILLER_21_854 ();
 sg13g2_decap_8 FILLER_21_861 ();
 sg13g2_decap_8 FILLER_21_868 ();
 sg13g2_decap_8 FILLER_21_875 ();
 sg13g2_decap_8 FILLER_21_882 ();
 sg13g2_decap_8 FILLER_21_889 ();
 sg13g2_decap_8 FILLER_21_896 ();
 sg13g2_decap_8 FILLER_21_903 ();
 sg13g2_decap_8 FILLER_21_910 ();
 sg13g2_decap_8 FILLER_21_917 ();
 sg13g2_decap_8 FILLER_21_924 ();
 sg13g2_decap_8 FILLER_21_931 ();
 sg13g2_decap_8 FILLER_21_938 ();
 sg13g2_decap_8 FILLER_21_945 ();
 sg13g2_decap_8 FILLER_21_952 ();
 sg13g2_decap_8 FILLER_21_959 ();
 sg13g2_decap_8 FILLER_21_966 ();
 sg13g2_decap_8 FILLER_21_973 ();
 sg13g2_decap_8 FILLER_21_980 ();
 sg13g2_decap_8 FILLER_21_987 ();
 sg13g2_decap_8 FILLER_21_994 ();
 sg13g2_decap_8 FILLER_21_1001 ();
 sg13g2_decap_8 FILLER_21_1008 ();
 sg13g2_decap_8 FILLER_21_1015 ();
 sg13g2_decap_8 FILLER_21_1022 ();
 sg13g2_decap_8 FILLER_22_4 ();
 sg13g2_decap_8 FILLER_22_11 ();
 sg13g2_decap_8 FILLER_22_18 ();
 sg13g2_decap_8 FILLER_22_25 ();
 sg13g2_decap_8 FILLER_22_32 ();
 sg13g2_decap_8 FILLER_22_39 ();
 sg13g2_decap_8 FILLER_22_46 ();
 sg13g2_decap_8 FILLER_22_53 ();
 sg13g2_decap_8 FILLER_22_60 ();
 sg13g2_decap_8 FILLER_22_67 ();
 sg13g2_decap_8 FILLER_22_74 ();
 sg13g2_decap_8 FILLER_22_81 ();
 sg13g2_decap_8 FILLER_22_88 ();
 sg13g2_decap_8 FILLER_22_95 ();
 sg13g2_decap_8 FILLER_22_102 ();
 sg13g2_decap_8 FILLER_22_109 ();
 sg13g2_decap_8 FILLER_22_116 ();
 sg13g2_decap_8 FILLER_22_123 ();
 sg13g2_decap_8 FILLER_22_130 ();
 sg13g2_decap_8 FILLER_22_137 ();
 sg13g2_decap_8 FILLER_22_144 ();
 sg13g2_decap_8 FILLER_22_151 ();
 sg13g2_decap_8 FILLER_22_158 ();
 sg13g2_decap_8 FILLER_22_165 ();
 sg13g2_decap_8 FILLER_22_172 ();
 sg13g2_decap_8 FILLER_22_179 ();
 sg13g2_decap_8 FILLER_22_186 ();
 sg13g2_decap_8 FILLER_22_193 ();
 sg13g2_decap_8 FILLER_22_200 ();
 sg13g2_decap_8 FILLER_22_207 ();
 sg13g2_decap_8 FILLER_22_214 ();
 sg13g2_decap_8 FILLER_22_221 ();
 sg13g2_decap_8 FILLER_22_228 ();
 sg13g2_decap_8 FILLER_22_235 ();
 sg13g2_decap_8 FILLER_22_242 ();
 sg13g2_decap_8 FILLER_22_249 ();
 sg13g2_decap_8 FILLER_22_256 ();
 sg13g2_decap_8 FILLER_22_263 ();
 sg13g2_decap_8 FILLER_22_270 ();
 sg13g2_decap_8 FILLER_22_277 ();
 sg13g2_decap_8 FILLER_22_284 ();
 sg13g2_decap_8 FILLER_22_291 ();
 sg13g2_decap_8 FILLER_22_298 ();
 sg13g2_decap_8 FILLER_22_305 ();
 sg13g2_decap_8 FILLER_22_312 ();
 sg13g2_decap_8 FILLER_22_319 ();
 sg13g2_decap_8 FILLER_22_326 ();
 sg13g2_decap_8 FILLER_22_333 ();
 sg13g2_decap_8 FILLER_22_340 ();
 sg13g2_decap_8 FILLER_22_347 ();
 sg13g2_decap_8 FILLER_22_354 ();
 sg13g2_decap_8 FILLER_22_361 ();
 sg13g2_decap_8 FILLER_22_368 ();
 sg13g2_decap_8 FILLER_22_375 ();
 sg13g2_decap_8 FILLER_22_382 ();
 sg13g2_decap_8 FILLER_22_389 ();
 sg13g2_decap_8 FILLER_22_396 ();
 sg13g2_decap_8 FILLER_22_403 ();
 sg13g2_decap_8 FILLER_22_410 ();
 sg13g2_decap_8 FILLER_22_417 ();
 sg13g2_decap_8 FILLER_22_424 ();
 sg13g2_decap_8 FILLER_22_431 ();
 sg13g2_decap_8 FILLER_22_438 ();
 sg13g2_decap_8 FILLER_22_445 ();
 sg13g2_decap_8 FILLER_22_452 ();
 sg13g2_decap_8 FILLER_22_459 ();
 sg13g2_decap_8 FILLER_22_466 ();
 sg13g2_decap_8 FILLER_22_473 ();
 sg13g2_decap_8 FILLER_22_480 ();
 sg13g2_decap_8 FILLER_22_487 ();
 sg13g2_decap_8 FILLER_22_494 ();
 sg13g2_decap_8 FILLER_22_501 ();
 sg13g2_decap_8 FILLER_22_508 ();
 sg13g2_decap_8 FILLER_22_515 ();
 sg13g2_decap_8 FILLER_22_522 ();
 sg13g2_decap_8 FILLER_22_529 ();
 sg13g2_decap_8 FILLER_22_536 ();
 sg13g2_decap_8 FILLER_22_543 ();
 sg13g2_decap_8 FILLER_22_550 ();
 sg13g2_decap_8 FILLER_22_557 ();
 sg13g2_decap_8 FILLER_22_564 ();
 sg13g2_decap_8 FILLER_22_571 ();
 sg13g2_decap_8 FILLER_22_578 ();
 sg13g2_decap_8 FILLER_22_585 ();
 sg13g2_decap_8 FILLER_22_592 ();
 sg13g2_decap_8 FILLER_22_599 ();
 sg13g2_decap_8 FILLER_22_606 ();
 sg13g2_decap_8 FILLER_22_613 ();
 sg13g2_decap_8 FILLER_22_620 ();
 sg13g2_decap_8 FILLER_22_627 ();
 sg13g2_decap_8 FILLER_22_634 ();
 sg13g2_decap_8 FILLER_22_641 ();
 sg13g2_decap_8 FILLER_22_648 ();
 sg13g2_decap_8 FILLER_22_655 ();
 sg13g2_decap_8 FILLER_22_662 ();
 sg13g2_decap_8 FILLER_22_669 ();
 sg13g2_decap_8 FILLER_22_676 ();
 sg13g2_decap_8 FILLER_22_683 ();
 sg13g2_decap_8 FILLER_22_690 ();
 sg13g2_decap_8 FILLER_22_697 ();
 sg13g2_decap_8 FILLER_22_704 ();
 sg13g2_decap_8 FILLER_22_711 ();
 sg13g2_decap_8 FILLER_22_718 ();
 sg13g2_decap_8 FILLER_22_725 ();
 sg13g2_decap_8 FILLER_22_732 ();
 sg13g2_decap_8 FILLER_22_739 ();
 sg13g2_decap_8 FILLER_22_746 ();
 sg13g2_decap_8 FILLER_22_753 ();
 sg13g2_decap_8 FILLER_22_760 ();
 sg13g2_decap_8 FILLER_22_767 ();
 sg13g2_decap_8 FILLER_22_774 ();
 sg13g2_decap_8 FILLER_22_781 ();
 sg13g2_decap_8 FILLER_22_788 ();
 sg13g2_decap_8 FILLER_22_795 ();
 sg13g2_decap_8 FILLER_22_802 ();
 sg13g2_decap_8 FILLER_22_809 ();
 sg13g2_decap_8 FILLER_22_816 ();
 sg13g2_decap_8 FILLER_22_823 ();
 sg13g2_decap_8 FILLER_22_830 ();
 sg13g2_decap_8 FILLER_22_837 ();
 sg13g2_decap_8 FILLER_22_844 ();
 sg13g2_decap_8 FILLER_22_851 ();
 sg13g2_decap_8 FILLER_22_858 ();
 sg13g2_decap_8 FILLER_22_865 ();
 sg13g2_decap_8 FILLER_22_872 ();
 sg13g2_decap_8 FILLER_22_879 ();
 sg13g2_decap_8 FILLER_22_886 ();
 sg13g2_decap_8 FILLER_22_893 ();
 sg13g2_decap_8 FILLER_22_900 ();
 sg13g2_decap_8 FILLER_22_907 ();
 sg13g2_decap_8 FILLER_22_914 ();
 sg13g2_decap_8 FILLER_22_921 ();
 sg13g2_decap_8 FILLER_22_928 ();
 sg13g2_decap_8 FILLER_22_935 ();
 sg13g2_decap_8 FILLER_22_942 ();
 sg13g2_decap_8 FILLER_22_949 ();
 sg13g2_decap_8 FILLER_22_956 ();
 sg13g2_decap_8 FILLER_22_963 ();
 sg13g2_decap_8 FILLER_22_970 ();
 sg13g2_decap_8 FILLER_22_977 ();
 sg13g2_decap_8 FILLER_22_984 ();
 sg13g2_decap_8 FILLER_22_991 ();
 sg13g2_decap_8 FILLER_22_998 ();
 sg13g2_decap_8 FILLER_22_1005 ();
 sg13g2_decap_8 FILLER_22_1012 ();
 sg13g2_decap_8 FILLER_22_1019 ();
 sg13g2_fill_2 FILLER_22_1026 ();
 sg13g2_fill_1 FILLER_22_1028 ();
 sg13g2_decap_8 FILLER_23_0 ();
 sg13g2_decap_8 FILLER_23_7 ();
 sg13g2_decap_8 FILLER_23_14 ();
 sg13g2_decap_8 FILLER_23_21 ();
 sg13g2_decap_8 FILLER_23_28 ();
 sg13g2_decap_8 FILLER_23_35 ();
 sg13g2_decap_8 FILLER_23_42 ();
 sg13g2_decap_8 FILLER_23_49 ();
 sg13g2_decap_8 FILLER_23_56 ();
 sg13g2_decap_8 FILLER_23_63 ();
 sg13g2_decap_8 FILLER_23_70 ();
 sg13g2_decap_8 FILLER_23_77 ();
 sg13g2_decap_8 FILLER_23_84 ();
 sg13g2_decap_8 FILLER_23_91 ();
 sg13g2_decap_8 FILLER_23_98 ();
 sg13g2_decap_8 FILLER_23_105 ();
 sg13g2_decap_8 FILLER_23_112 ();
 sg13g2_decap_8 FILLER_23_119 ();
 sg13g2_decap_8 FILLER_23_126 ();
 sg13g2_decap_8 FILLER_23_133 ();
 sg13g2_decap_8 FILLER_23_140 ();
 sg13g2_decap_8 FILLER_23_147 ();
 sg13g2_decap_8 FILLER_23_154 ();
 sg13g2_decap_8 FILLER_23_161 ();
 sg13g2_decap_8 FILLER_23_168 ();
 sg13g2_decap_8 FILLER_23_175 ();
 sg13g2_decap_8 FILLER_23_182 ();
 sg13g2_decap_8 FILLER_23_189 ();
 sg13g2_decap_8 FILLER_23_196 ();
 sg13g2_decap_8 FILLER_23_203 ();
 sg13g2_decap_8 FILLER_23_210 ();
 sg13g2_decap_8 FILLER_23_217 ();
 sg13g2_decap_8 FILLER_23_224 ();
 sg13g2_decap_8 FILLER_23_231 ();
 sg13g2_decap_8 FILLER_23_238 ();
 sg13g2_decap_8 FILLER_23_245 ();
 sg13g2_decap_8 FILLER_23_252 ();
 sg13g2_decap_8 FILLER_23_259 ();
 sg13g2_decap_8 FILLER_23_266 ();
 sg13g2_decap_8 FILLER_23_273 ();
 sg13g2_decap_8 FILLER_23_280 ();
 sg13g2_decap_8 FILLER_23_287 ();
 sg13g2_decap_8 FILLER_23_294 ();
 sg13g2_decap_8 FILLER_23_301 ();
 sg13g2_decap_8 FILLER_23_308 ();
 sg13g2_decap_8 FILLER_23_315 ();
 sg13g2_decap_8 FILLER_23_322 ();
 sg13g2_decap_8 FILLER_23_329 ();
 sg13g2_decap_8 FILLER_23_336 ();
 sg13g2_decap_8 FILLER_23_343 ();
 sg13g2_decap_8 FILLER_23_350 ();
 sg13g2_decap_8 FILLER_23_357 ();
 sg13g2_decap_8 FILLER_23_364 ();
 sg13g2_decap_8 FILLER_23_371 ();
 sg13g2_decap_8 FILLER_23_378 ();
 sg13g2_decap_8 FILLER_23_385 ();
 sg13g2_decap_8 FILLER_23_392 ();
 sg13g2_decap_8 FILLER_23_399 ();
 sg13g2_decap_8 FILLER_23_406 ();
 sg13g2_decap_8 FILLER_23_413 ();
 sg13g2_decap_8 FILLER_23_420 ();
 sg13g2_decap_8 FILLER_23_427 ();
 sg13g2_decap_8 FILLER_23_434 ();
 sg13g2_decap_8 FILLER_23_441 ();
 sg13g2_decap_8 FILLER_23_448 ();
 sg13g2_decap_8 FILLER_23_455 ();
 sg13g2_decap_8 FILLER_23_462 ();
 sg13g2_decap_8 FILLER_23_469 ();
 sg13g2_decap_8 FILLER_23_476 ();
 sg13g2_decap_8 FILLER_23_483 ();
 sg13g2_decap_8 FILLER_23_490 ();
 sg13g2_decap_8 FILLER_23_497 ();
 sg13g2_decap_8 FILLER_23_504 ();
 sg13g2_decap_8 FILLER_23_511 ();
 sg13g2_decap_8 FILLER_23_518 ();
 sg13g2_decap_8 FILLER_23_525 ();
 sg13g2_decap_8 FILLER_23_532 ();
 sg13g2_decap_8 FILLER_23_539 ();
 sg13g2_decap_8 FILLER_23_546 ();
 sg13g2_decap_8 FILLER_23_553 ();
 sg13g2_decap_8 FILLER_23_560 ();
 sg13g2_decap_8 FILLER_23_567 ();
 sg13g2_decap_8 FILLER_23_574 ();
 sg13g2_decap_8 FILLER_23_581 ();
 sg13g2_decap_8 FILLER_23_588 ();
 sg13g2_decap_8 FILLER_23_595 ();
 sg13g2_decap_8 FILLER_23_602 ();
 sg13g2_decap_8 FILLER_23_609 ();
 sg13g2_decap_8 FILLER_23_616 ();
 sg13g2_decap_8 FILLER_23_623 ();
 sg13g2_decap_8 FILLER_23_630 ();
 sg13g2_decap_8 FILLER_23_637 ();
 sg13g2_decap_8 FILLER_23_644 ();
 sg13g2_decap_8 FILLER_23_651 ();
 sg13g2_decap_8 FILLER_23_658 ();
 sg13g2_decap_8 FILLER_23_665 ();
 sg13g2_decap_8 FILLER_23_672 ();
 sg13g2_decap_8 FILLER_23_679 ();
 sg13g2_decap_8 FILLER_23_686 ();
 sg13g2_decap_8 FILLER_23_693 ();
 sg13g2_decap_8 FILLER_23_700 ();
 sg13g2_decap_8 FILLER_23_707 ();
 sg13g2_decap_8 FILLER_23_714 ();
 sg13g2_decap_8 FILLER_23_721 ();
 sg13g2_decap_8 FILLER_23_728 ();
 sg13g2_decap_8 FILLER_23_735 ();
 sg13g2_decap_8 FILLER_23_742 ();
 sg13g2_decap_8 FILLER_23_749 ();
 sg13g2_decap_8 FILLER_23_756 ();
 sg13g2_decap_8 FILLER_23_763 ();
 sg13g2_decap_8 FILLER_23_770 ();
 sg13g2_decap_8 FILLER_23_777 ();
 sg13g2_decap_8 FILLER_23_784 ();
 sg13g2_decap_8 FILLER_23_791 ();
 sg13g2_decap_8 FILLER_23_798 ();
 sg13g2_decap_8 FILLER_23_805 ();
 sg13g2_decap_8 FILLER_23_812 ();
 sg13g2_decap_8 FILLER_23_819 ();
 sg13g2_decap_8 FILLER_23_826 ();
 sg13g2_decap_8 FILLER_23_833 ();
 sg13g2_decap_8 FILLER_23_840 ();
 sg13g2_decap_8 FILLER_23_847 ();
 sg13g2_decap_8 FILLER_23_854 ();
 sg13g2_decap_8 FILLER_23_861 ();
 sg13g2_decap_8 FILLER_23_868 ();
 sg13g2_decap_8 FILLER_23_875 ();
 sg13g2_decap_8 FILLER_23_882 ();
 sg13g2_decap_8 FILLER_23_889 ();
 sg13g2_decap_8 FILLER_23_896 ();
 sg13g2_decap_8 FILLER_23_903 ();
 sg13g2_decap_8 FILLER_23_910 ();
 sg13g2_decap_8 FILLER_23_917 ();
 sg13g2_decap_8 FILLER_23_924 ();
 sg13g2_decap_8 FILLER_23_931 ();
 sg13g2_decap_8 FILLER_23_938 ();
 sg13g2_decap_8 FILLER_23_945 ();
 sg13g2_decap_8 FILLER_23_952 ();
 sg13g2_decap_8 FILLER_23_959 ();
 sg13g2_decap_8 FILLER_23_966 ();
 sg13g2_decap_8 FILLER_23_973 ();
 sg13g2_decap_8 FILLER_23_980 ();
 sg13g2_decap_8 FILLER_23_987 ();
 sg13g2_decap_8 FILLER_23_994 ();
 sg13g2_decap_8 FILLER_23_1001 ();
 sg13g2_decap_8 FILLER_23_1008 ();
 sg13g2_decap_8 FILLER_23_1015 ();
 sg13g2_decap_8 FILLER_23_1022 ();
 sg13g2_decap_8 FILLER_24_4 ();
 sg13g2_decap_8 FILLER_24_11 ();
 sg13g2_decap_8 FILLER_24_18 ();
 sg13g2_decap_8 FILLER_24_25 ();
 sg13g2_decap_8 FILLER_24_32 ();
 sg13g2_decap_8 FILLER_24_39 ();
 sg13g2_decap_8 FILLER_24_46 ();
 sg13g2_decap_8 FILLER_24_53 ();
 sg13g2_decap_8 FILLER_24_60 ();
 sg13g2_decap_8 FILLER_24_67 ();
 sg13g2_decap_8 FILLER_24_74 ();
 sg13g2_decap_8 FILLER_24_81 ();
 sg13g2_decap_8 FILLER_24_88 ();
 sg13g2_decap_8 FILLER_24_95 ();
 sg13g2_decap_8 FILLER_24_102 ();
 sg13g2_decap_8 FILLER_24_109 ();
 sg13g2_decap_8 FILLER_24_116 ();
 sg13g2_decap_8 FILLER_24_123 ();
 sg13g2_decap_8 FILLER_24_130 ();
 sg13g2_decap_8 FILLER_24_137 ();
 sg13g2_decap_8 FILLER_24_144 ();
 sg13g2_decap_8 FILLER_24_151 ();
 sg13g2_decap_8 FILLER_24_158 ();
 sg13g2_decap_8 FILLER_24_165 ();
 sg13g2_decap_8 FILLER_24_172 ();
 sg13g2_decap_8 FILLER_24_179 ();
 sg13g2_decap_8 FILLER_24_186 ();
 sg13g2_decap_8 FILLER_24_193 ();
 sg13g2_decap_8 FILLER_24_200 ();
 sg13g2_decap_8 FILLER_24_207 ();
 sg13g2_decap_8 FILLER_24_214 ();
 sg13g2_decap_8 FILLER_24_221 ();
 sg13g2_decap_8 FILLER_24_228 ();
 sg13g2_decap_8 FILLER_24_235 ();
 sg13g2_decap_8 FILLER_24_242 ();
 sg13g2_decap_8 FILLER_24_249 ();
 sg13g2_decap_8 FILLER_24_256 ();
 sg13g2_decap_8 FILLER_24_263 ();
 sg13g2_decap_8 FILLER_24_270 ();
 sg13g2_decap_8 FILLER_24_277 ();
 sg13g2_decap_8 FILLER_24_284 ();
 sg13g2_decap_8 FILLER_24_291 ();
 sg13g2_decap_8 FILLER_24_298 ();
 sg13g2_decap_8 FILLER_24_305 ();
 sg13g2_decap_8 FILLER_24_312 ();
 sg13g2_decap_8 FILLER_24_319 ();
 sg13g2_decap_8 FILLER_24_326 ();
 sg13g2_decap_8 FILLER_24_333 ();
 sg13g2_decap_8 FILLER_24_340 ();
 sg13g2_decap_8 FILLER_24_347 ();
 sg13g2_decap_8 FILLER_24_354 ();
 sg13g2_decap_8 FILLER_24_361 ();
 sg13g2_decap_8 FILLER_24_368 ();
 sg13g2_decap_8 FILLER_24_375 ();
 sg13g2_decap_8 FILLER_24_382 ();
 sg13g2_decap_8 FILLER_24_389 ();
 sg13g2_decap_8 FILLER_24_396 ();
 sg13g2_decap_8 FILLER_24_403 ();
 sg13g2_decap_8 FILLER_24_410 ();
 sg13g2_decap_8 FILLER_24_417 ();
 sg13g2_decap_8 FILLER_24_424 ();
 sg13g2_decap_8 FILLER_24_431 ();
 sg13g2_decap_8 FILLER_24_438 ();
 sg13g2_decap_8 FILLER_24_445 ();
 sg13g2_decap_8 FILLER_24_452 ();
 sg13g2_decap_8 FILLER_24_459 ();
 sg13g2_decap_8 FILLER_24_466 ();
 sg13g2_decap_8 FILLER_24_473 ();
 sg13g2_decap_8 FILLER_24_480 ();
 sg13g2_decap_8 FILLER_24_487 ();
 sg13g2_decap_8 FILLER_24_494 ();
 sg13g2_decap_8 FILLER_24_501 ();
 sg13g2_decap_8 FILLER_24_508 ();
 sg13g2_decap_8 FILLER_24_515 ();
 sg13g2_decap_8 FILLER_24_522 ();
 sg13g2_decap_8 FILLER_24_529 ();
 sg13g2_decap_8 FILLER_24_536 ();
 sg13g2_decap_8 FILLER_24_543 ();
 sg13g2_decap_8 FILLER_24_550 ();
 sg13g2_decap_8 FILLER_24_557 ();
 sg13g2_decap_8 FILLER_24_564 ();
 sg13g2_decap_8 FILLER_24_571 ();
 sg13g2_decap_8 FILLER_24_578 ();
 sg13g2_decap_8 FILLER_24_585 ();
 sg13g2_decap_8 FILLER_24_592 ();
 sg13g2_decap_8 FILLER_24_599 ();
 sg13g2_decap_8 FILLER_24_606 ();
 sg13g2_decap_8 FILLER_24_613 ();
 sg13g2_decap_8 FILLER_24_620 ();
 sg13g2_decap_8 FILLER_24_627 ();
 sg13g2_decap_8 FILLER_24_634 ();
 sg13g2_decap_8 FILLER_24_641 ();
 sg13g2_decap_8 FILLER_24_648 ();
 sg13g2_decap_8 FILLER_24_655 ();
 sg13g2_decap_8 FILLER_24_662 ();
 sg13g2_decap_8 FILLER_24_669 ();
 sg13g2_decap_8 FILLER_24_676 ();
 sg13g2_decap_8 FILLER_24_683 ();
 sg13g2_decap_8 FILLER_24_690 ();
 sg13g2_decap_8 FILLER_24_697 ();
 sg13g2_decap_8 FILLER_24_704 ();
 sg13g2_decap_8 FILLER_24_711 ();
 sg13g2_decap_8 FILLER_24_718 ();
 sg13g2_decap_8 FILLER_24_725 ();
 sg13g2_decap_8 FILLER_24_732 ();
 sg13g2_decap_8 FILLER_24_739 ();
 sg13g2_decap_8 FILLER_24_746 ();
 sg13g2_decap_8 FILLER_24_753 ();
 sg13g2_decap_8 FILLER_24_760 ();
 sg13g2_decap_8 FILLER_24_767 ();
 sg13g2_decap_8 FILLER_24_774 ();
 sg13g2_decap_8 FILLER_24_781 ();
 sg13g2_decap_8 FILLER_24_788 ();
 sg13g2_decap_8 FILLER_24_795 ();
 sg13g2_decap_8 FILLER_24_802 ();
 sg13g2_decap_8 FILLER_24_809 ();
 sg13g2_decap_8 FILLER_24_816 ();
 sg13g2_decap_8 FILLER_24_823 ();
 sg13g2_decap_8 FILLER_24_830 ();
 sg13g2_decap_8 FILLER_24_837 ();
 sg13g2_decap_8 FILLER_24_844 ();
 sg13g2_decap_8 FILLER_24_851 ();
 sg13g2_decap_8 FILLER_24_858 ();
 sg13g2_decap_8 FILLER_24_865 ();
 sg13g2_decap_8 FILLER_24_872 ();
 sg13g2_decap_8 FILLER_24_879 ();
 sg13g2_decap_8 FILLER_24_886 ();
 sg13g2_decap_8 FILLER_24_893 ();
 sg13g2_decap_8 FILLER_24_900 ();
 sg13g2_decap_8 FILLER_24_907 ();
 sg13g2_decap_8 FILLER_24_914 ();
 sg13g2_decap_8 FILLER_24_921 ();
 sg13g2_decap_8 FILLER_24_928 ();
 sg13g2_decap_8 FILLER_24_935 ();
 sg13g2_decap_8 FILLER_24_942 ();
 sg13g2_decap_8 FILLER_24_949 ();
 sg13g2_decap_8 FILLER_24_956 ();
 sg13g2_decap_8 FILLER_24_963 ();
 sg13g2_decap_8 FILLER_24_970 ();
 sg13g2_decap_8 FILLER_24_977 ();
 sg13g2_decap_8 FILLER_24_984 ();
 sg13g2_decap_8 FILLER_24_991 ();
 sg13g2_decap_8 FILLER_24_998 ();
 sg13g2_decap_8 FILLER_24_1005 ();
 sg13g2_decap_8 FILLER_24_1012 ();
 sg13g2_decap_8 FILLER_24_1019 ();
 sg13g2_fill_2 FILLER_24_1026 ();
 sg13g2_fill_1 FILLER_24_1028 ();
 sg13g2_decap_8 FILLER_25_0 ();
 sg13g2_decap_8 FILLER_25_7 ();
 sg13g2_decap_8 FILLER_25_14 ();
 sg13g2_decap_8 FILLER_25_21 ();
 sg13g2_decap_8 FILLER_25_28 ();
 sg13g2_decap_8 FILLER_25_35 ();
 sg13g2_decap_8 FILLER_25_42 ();
 sg13g2_decap_8 FILLER_25_49 ();
 sg13g2_decap_8 FILLER_25_56 ();
 sg13g2_decap_8 FILLER_25_63 ();
 sg13g2_decap_8 FILLER_25_70 ();
 sg13g2_decap_8 FILLER_25_77 ();
 sg13g2_decap_8 FILLER_25_84 ();
 sg13g2_decap_8 FILLER_25_91 ();
 sg13g2_decap_8 FILLER_25_98 ();
 sg13g2_decap_8 FILLER_25_105 ();
 sg13g2_decap_8 FILLER_25_112 ();
 sg13g2_decap_8 FILLER_25_119 ();
 sg13g2_decap_8 FILLER_25_126 ();
 sg13g2_decap_8 FILLER_25_133 ();
 sg13g2_decap_8 FILLER_25_140 ();
 sg13g2_decap_8 FILLER_25_147 ();
 sg13g2_decap_8 FILLER_25_154 ();
 sg13g2_decap_8 FILLER_25_161 ();
 sg13g2_decap_8 FILLER_25_168 ();
 sg13g2_decap_8 FILLER_25_175 ();
 sg13g2_decap_8 FILLER_25_182 ();
 sg13g2_decap_8 FILLER_25_189 ();
 sg13g2_decap_8 FILLER_25_196 ();
 sg13g2_decap_8 FILLER_25_203 ();
 sg13g2_decap_8 FILLER_25_210 ();
 sg13g2_decap_8 FILLER_25_217 ();
 sg13g2_decap_8 FILLER_25_224 ();
 sg13g2_decap_8 FILLER_25_231 ();
 sg13g2_decap_8 FILLER_25_238 ();
 sg13g2_decap_8 FILLER_25_245 ();
 sg13g2_decap_8 FILLER_25_252 ();
 sg13g2_decap_8 FILLER_25_259 ();
 sg13g2_decap_8 FILLER_25_266 ();
 sg13g2_decap_8 FILLER_25_273 ();
 sg13g2_decap_8 FILLER_25_280 ();
 sg13g2_decap_8 FILLER_25_287 ();
 sg13g2_decap_8 FILLER_25_294 ();
 sg13g2_decap_8 FILLER_25_301 ();
 sg13g2_decap_8 FILLER_25_308 ();
 sg13g2_decap_8 FILLER_25_315 ();
 sg13g2_decap_8 FILLER_25_322 ();
 sg13g2_decap_8 FILLER_25_329 ();
 sg13g2_decap_8 FILLER_25_336 ();
 sg13g2_decap_8 FILLER_25_343 ();
 sg13g2_decap_8 FILLER_25_350 ();
 sg13g2_decap_8 FILLER_25_357 ();
 sg13g2_decap_8 FILLER_25_364 ();
 sg13g2_decap_8 FILLER_25_371 ();
 sg13g2_decap_8 FILLER_25_378 ();
 sg13g2_decap_8 FILLER_25_385 ();
 sg13g2_decap_8 FILLER_25_392 ();
 sg13g2_decap_8 FILLER_25_399 ();
 sg13g2_decap_8 FILLER_25_406 ();
 sg13g2_decap_8 FILLER_25_413 ();
 sg13g2_decap_8 FILLER_25_420 ();
 sg13g2_decap_8 FILLER_25_427 ();
 sg13g2_decap_8 FILLER_25_434 ();
 sg13g2_decap_8 FILLER_25_441 ();
 sg13g2_decap_8 FILLER_25_448 ();
 sg13g2_decap_8 FILLER_25_455 ();
 sg13g2_decap_8 FILLER_25_462 ();
 sg13g2_decap_8 FILLER_25_469 ();
 sg13g2_decap_8 FILLER_25_476 ();
 sg13g2_decap_8 FILLER_25_483 ();
 sg13g2_decap_8 FILLER_25_490 ();
 sg13g2_decap_8 FILLER_25_497 ();
 sg13g2_decap_8 FILLER_25_504 ();
 sg13g2_decap_8 FILLER_25_511 ();
 sg13g2_decap_8 FILLER_25_518 ();
 sg13g2_decap_8 FILLER_25_525 ();
 sg13g2_decap_8 FILLER_25_532 ();
 sg13g2_decap_8 FILLER_25_539 ();
 sg13g2_decap_8 FILLER_25_546 ();
 sg13g2_decap_8 FILLER_25_553 ();
 sg13g2_decap_8 FILLER_25_560 ();
 sg13g2_decap_8 FILLER_25_567 ();
 sg13g2_decap_8 FILLER_25_574 ();
 sg13g2_decap_8 FILLER_25_581 ();
 sg13g2_decap_8 FILLER_25_588 ();
 sg13g2_decap_8 FILLER_25_595 ();
 sg13g2_decap_8 FILLER_25_602 ();
 sg13g2_decap_8 FILLER_25_609 ();
 sg13g2_decap_8 FILLER_25_616 ();
 sg13g2_decap_8 FILLER_25_623 ();
 sg13g2_decap_8 FILLER_25_630 ();
 sg13g2_decap_8 FILLER_25_637 ();
 sg13g2_decap_8 FILLER_25_644 ();
 sg13g2_decap_8 FILLER_25_651 ();
 sg13g2_decap_8 FILLER_25_658 ();
 sg13g2_decap_8 FILLER_25_665 ();
 sg13g2_decap_8 FILLER_25_672 ();
 sg13g2_decap_8 FILLER_25_679 ();
 sg13g2_decap_8 FILLER_25_686 ();
 sg13g2_decap_8 FILLER_25_693 ();
 sg13g2_decap_8 FILLER_25_700 ();
 sg13g2_decap_8 FILLER_25_707 ();
 sg13g2_decap_8 FILLER_25_714 ();
 sg13g2_decap_8 FILLER_25_721 ();
 sg13g2_decap_8 FILLER_25_728 ();
 sg13g2_decap_8 FILLER_25_735 ();
 sg13g2_decap_8 FILLER_25_742 ();
 sg13g2_decap_8 FILLER_25_749 ();
 sg13g2_decap_8 FILLER_25_756 ();
 sg13g2_decap_8 FILLER_25_763 ();
 sg13g2_decap_8 FILLER_25_770 ();
 sg13g2_decap_8 FILLER_25_777 ();
 sg13g2_decap_8 FILLER_25_784 ();
 sg13g2_decap_8 FILLER_25_791 ();
 sg13g2_decap_8 FILLER_25_798 ();
 sg13g2_decap_8 FILLER_25_805 ();
 sg13g2_decap_8 FILLER_25_812 ();
 sg13g2_decap_8 FILLER_25_819 ();
 sg13g2_decap_8 FILLER_25_826 ();
 sg13g2_decap_8 FILLER_25_833 ();
 sg13g2_decap_8 FILLER_25_840 ();
 sg13g2_decap_8 FILLER_25_847 ();
 sg13g2_decap_8 FILLER_25_854 ();
 sg13g2_decap_8 FILLER_25_861 ();
 sg13g2_decap_8 FILLER_25_868 ();
 sg13g2_decap_8 FILLER_25_875 ();
 sg13g2_decap_8 FILLER_25_882 ();
 sg13g2_decap_8 FILLER_25_889 ();
 sg13g2_decap_8 FILLER_25_896 ();
 sg13g2_decap_8 FILLER_25_903 ();
 sg13g2_decap_8 FILLER_25_910 ();
 sg13g2_decap_8 FILLER_25_917 ();
 sg13g2_decap_8 FILLER_25_924 ();
 sg13g2_decap_8 FILLER_25_931 ();
 sg13g2_decap_8 FILLER_25_938 ();
 sg13g2_decap_8 FILLER_25_945 ();
 sg13g2_decap_8 FILLER_25_952 ();
 sg13g2_decap_8 FILLER_25_959 ();
 sg13g2_decap_8 FILLER_25_966 ();
 sg13g2_decap_8 FILLER_25_973 ();
 sg13g2_decap_8 FILLER_25_980 ();
 sg13g2_decap_8 FILLER_25_987 ();
 sg13g2_decap_8 FILLER_25_994 ();
 sg13g2_decap_8 FILLER_25_1001 ();
 sg13g2_decap_8 FILLER_25_1008 ();
 sg13g2_decap_8 FILLER_25_1015 ();
 sg13g2_decap_8 FILLER_25_1022 ();
 sg13g2_decap_8 FILLER_26_0 ();
 sg13g2_decap_8 FILLER_26_7 ();
 sg13g2_decap_8 FILLER_26_14 ();
 sg13g2_decap_8 FILLER_26_21 ();
 sg13g2_decap_8 FILLER_26_28 ();
 sg13g2_decap_8 FILLER_26_35 ();
 sg13g2_decap_8 FILLER_26_42 ();
 sg13g2_decap_8 FILLER_26_49 ();
 sg13g2_decap_8 FILLER_26_56 ();
 sg13g2_decap_8 FILLER_26_63 ();
 sg13g2_decap_8 FILLER_26_70 ();
 sg13g2_decap_8 FILLER_26_77 ();
 sg13g2_decap_8 FILLER_26_84 ();
 sg13g2_decap_8 FILLER_26_91 ();
 sg13g2_decap_8 FILLER_26_98 ();
 sg13g2_decap_8 FILLER_26_105 ();
 sg13g2_decap_8 FILLER_26_112 ();
 sg13g2_decap_8 FILLER_26_119 ();
 sg13g2_decap_8 FILLER_26_126 ();
 sg13g2_decap_8 FILLER_26_133 ();
 sg13g2_decap_8 FILLER_26_140 ();
 sg13g2_decap_8 FILLER_26_147 ();
 sg13g2_decap_8 FILLER_26_154 ();
 sg13g2_decap_8 FILLER_26_161 ();
 sg13g2_decap_8 FILLER_26_168 ();
 sg13g2_decap_8 FILLER_26_175 ();
 sg13g2_decap_8 FILLER_26_182 ();
 sg13g2_decap_8 FILLER_26_189 ();
 sg13g2_decap_8 FILLER_26_196 ();
 sg13g2_decap_8 FILLER_26_203 ();
 sg13g2_decap_8 FILLER_26_210 ();
 sg13g2_decap_8 FILLER_26_217 ();
 sg13g2_decap_8 FILLER_26_224 ();
 sg13g2_decap_8 FILLER_26_231 ();
 sg13g2_decap_8 FILLER_26_238 ();
 sg13g2_decap_8 FILLER_26_245 ();
 sg13g2_decap_8 FILLER_26_252 ();
 sg13g2_decap_8 FILLER_26_259 ();
 sg13g2_decap_8 FILLER_26_266 ();
 sg13g2_decap_8 FILLER_26_273 ();
 sg13g2_decap_8 FILLER_26_280 ();
 sg13g2_decap_8 FILLER_26_287 ();
 sg13g2_decap_8 FILLER_26_294 ();
 sg13g2_decap_8 FILLER_26_301 ();
 sg13g2_decap_8 FILLER_26_308 ();
 sg13g2_decap_8 FILLER_26_315 ();
 sg13g2_decap_8 FILLER_26_322 ();
 sg13g2_decap_8 FILLER_26_329 ();
 sg13g2_decap_8 FILLER_26_336 ();
 sg13g2_decap_8 FILLER_26_343 ();
 sg13g2_decap_8 FILLER_26_350 ();
 sg13g2_decap_8 FILLER_26_357 ();
 sg13g2_decap_8 FILLER_26_364 ();
 sg13g2_decap_8 FILLER_26_371 ();
 sg13g2_decap_8 FILLER_26_378 ();
 sg13g2_decap_8 FILLER_26_385 ();
 sg13g2_decap_8 FILLER_26_392 ();
 sg13g2_decap_8 FILLER_26_399 ();
 sg13g2_decap_8 FILLER_26_406 ();
 sg13g2_decap_8 FILLER_26_413 ();
 sg13g2_decap_8 FILLER_26_420 ();
 sg13g2_decap_8 FILLER_26_427 ();
 sg13g2_decap_8 FILLER_26_434 ();
 sg13g2_decap_8 FILLER_26_441 ();
 sg13g2_decap_8 FILLER_26_448 ();
 sg13g2_decap_8 FILLER_26_455 ();
 sg13g2_decap_8 FILLER_26_462 ();
 sg13g2_decap_8 FILLER_26_469 ();
 sg13g2_decap_8 FILLER_26_476 ();
 sg13g2_decap_8 FILLER_26_483 ();
 sg13g2_decap_8 FILLER_26_490 ();
 sg13g2_decap_8 FILLER_26_497 ();
 sg13g2_decap_8 FILLER_26_504 ();
 sg13g2_decap_8 FILLER_26_511 ();
 sg13g2_decap_8 FILLER_26_518 ();
 sg13g2_decap_8 FILLER_26_525 ();
 sg13g2_decap_8 FILLER_26_532 ();
 sg13g2_decap_8 FILLER_26_539 ();
 sg13g2_decap_8 FILLER_26_546 ();
 sg13g2_decap_8 FILLER_26_553 ();
 sg13g2_decap_8 FILLER_26_560 ();
 sg13g2_decap_8 FILLER_26_567 ();
 sg13g2_decap_8 FILLER_26_574 ();
 sg13g2_decap_8 FILLER_26_581 ();
 sg13g2_decap_8 FILLER_26_588 ();
 sg13g2_decap_8 FILLER_26_595 ();
 sg13g2_decap_8 FILLER_26_602 ();
 sg13g2_decap_8 FILLER_26_609 ();
 sg13g2_decap_8 FILLER_26_616 ();
 sg13g2_decap_8 FILLER_26_623 ();
 sg13g2_decap_8 FILLER_26_630 ();
 sg13g2_decap_8 FILLER_26_637 ();
 sg13g2_decap_8 FILLER_26_644 ();
 sg13g2_decap_8 FILLER_26_651 ();
 sg13g2_decap_8 FILLER_26_658 ();
 sg13g2_decap_8 FILLER_26_665 ();
 sg13g2_decap_8 FILLER_26_672 ();
 sg13g2_decap_8 FILLER_26_679 ();
 sg13g2_decap_8 FILLER_26_686 ();
 sg13g2_decap_8 FILLER_26_693 ();
 sg13g2_decap_8 FILLER_26_700 ();
 sg13g2_decap_8 FILLER_26_707 ();
 sg13g2_decap_8 FILLER_26_714 ();
 sg13g2_decap_8 FILLER_26_721 ();
 sg13g2_decap_8 FILLER_26_728 ();
 sg13g2_decap_8 FILLER_26_735 ();
 sg13g2_decap_8 FILLER_26_742 ();
 sg13g2_decap_8 FILLER_26_749 ();
 sg13g2_decap_8 FILLER_26_756 ();
 sg13g2_decap_8 FILLER_26_763 ();
 sg13g2_decap_8 FILLER_26_770 ();
 sg13g2_decap_8 FILLER_26_777 ();
 sg13g2_decap_8 FILLER_26_784 ();
 sg13g2_decap_8 FILLER_26_791 ();
 sg13g2_decap_8 FILLER_26_798 ();
 sg13g2_decap_8 FILLER_26_805 ();
 sg13g2_decap_8 FILLER_26_812 ();
 sg13g2_decap_8 FILLER_26_819 ();
 sg13g2_decap_8 FILLER_26_826 ();
 sg13g2_decap_8 FILLER_26_833 ();
 sg13g2_decap_8 FILLER_26_840 ();
 sg13g2_decap_8 FILLER_26_847 ();
 sg13g2_decap_8 FILLER_26_854 ();
 sg13g2_decap_8 FILLER_26_861 ();
 sg13g2_decap_8 FILLER_26_868 ();
 sg13g2_decap_8 FILLER_26_875 ();
 sg13g2_decap_8 FILLER_26_882 ();
 sg13g2_decap_8 FILLER_26_889 ();
 sg13g2_decap_8 FILLER_26_896 ();
 sg13g2_decap_8 FILLER_26_903 ();
 sg13g2_decap_8 FILLER_26_910 ();
 sg13g2_decap_8 FILLER_26_917 ();
 sg13g2_decap_8 FILLER_26_924 ();
 sg13g2_decap_8 FILLER_26_931 ();
 sg13g2_decap_8 FILLER_26_938 ();
 sg13g2_decap_8 FILLER_26_945 ();
 sg13g2_decap_8 FILLER_26_952 ();
 sg13g2_decap_8 FILLER_26_959 ();
 sg13g2_decap_8 FILLER_26_966 ();
 sg13g2_decap_8 FILLER_26_973 ();
 sg13g2_decap_8 FILLER_26_980 ();
 sg13g2_decap_8 FILLER_26_987 ();
 sg13g2_decap_8 FILLER_26_994 ();
 sg13g2_decap_8 FILLER_26_1001 ();
 sg13g2_decap_8 FILLER_26_1008 ();
 sg13g2_decap_8 FILLER_26_1015 ();
 sg13g2_decap_8 FILLER_26_1022 ();
 sg13g2_decap_8 FILLER_27_4 ();
 sg13g2_decap_8 FILLER_27_11 ();
 sg13g2_decap_8 FILLER_27_18 ();
 sg13g2_decap_8 FILLER_27_25 ();
 sg13g2_decap_8 FILLER_27_32 ();
 sg13g2_decap_8 FILLER_27_39 ();
 sg13g2_decap_8 FILLER_27_46 ();
 sg13g2_decap_8 FILLER_27_53 ();
 sg13g2_decap_8 FILLER_27_60 ();
 sg13g2_decap_8 FILLER_27_67 ();
 sg13g2_decap_8 FILLER_27_74 ();
 sg13g2_decap_8 FILLER_27_81 ();
 sg13g2_decap_8 FILLER_27_88 ();
 sg13g2_decap_8 FILLER_27_95 ();
 sg13g2_decap_8 FILLER_27_102 ();
 sg13g2_decap_8 FILLER_27_109 ();
 sg13g2_decap_8 FILLER_27_116 ();
 sg13g2_decap_8 FILLER_27_123 ();
 sg13g2_decap_8 FILLER_27_130 ();
 sg13g2_decap_8 FILLER_27_137 ();
 sg13g2_decap_8 FILLER_27_144 ();
 sg13g2_decap_8 FILLER_27_151 ();
 sg13g2_decap_8 FILLER_27_158 ();
 sg13g2_decap_8 FILLER_27_165 ();
 sg13g2_decap_8 FILLER_27_172 ();
 sg13g2_decap_8 FILLER_27_179 ();
 sg13g2_decap_8 FILLER_27_186 ();
 sg13g2_decap_8 FILLER_27_193 ();
 sg13g2_decap_8 FILLER_27_200 ();
 sg13g2_decap_8 FILLER_27_207 ();
 sg13g2_decap_8 FILLER_27_214 ();
 sg13g2_decap_8 FILLER_27_221 ();
 sg13g2_decap_8 FILLER_27_228 ();
 sg13g2_decap_8 FILLER_27_235 ();
 sg13g2_decap_8 FILLER_27_242 ();
 sg13g2_decap_8 FILLER_27_249 ();
 sg13g2_decap_8 FILLER_27_256 ();
 sg13g2_decap_8 FILLER_27_263 ();
 sg13g2_decap_8 FILLER_27_270 ();
 sg13g2_decap_8 FILLER_27_277 ();
 sg13g2_decap_8 FILLER_27_284 ();
 sg13g2_decap_8 FILLER_27_291 ();
 sg13g2_decap_8 FILLER_27_298 ();
 sg13g2_decap_8 FILLER_27_305 ();
 sg13g2_decap_8 FILLER_27_312 ();
 sg13g2_decap_8 FILLER_27_319 ();
 sg13g2_decap_8 FILLER_27_326 ();
 sg13g2_decap_8 FILLER_27_333 ();
 sg13g2_decap_8 FILLER_27_340 ();
 sg13g2_decap_8 FILLER_27_347 ();
 sg13g2_decap_8 FILLER_27_354 ();
 sg13g2_decap_8 FILLER_27_361 ();
 sg13g2_decap_8 FILLER_27_368 ();
 sg13g2_decap_8 FILLER_27_375 ();
 sg13g2_decap_8 FILLER_27_382 ();
 sg13g2_decap_8 FILLER_27_389 ();
 sg13g2_decap_8 FILLER_27_396 ();
 sg13g2_decap_8 FILLER_27_403 ();
 sg13g2_decap_8 FILLER_27_410 ();
 sg13g2_decap_8 FILLER_27_417 ();
 sg13g2_decap_8 FILLER_27_424 ();
 sg13g2_decap_8 FILLER_27_431 ();
 sg13g2_decap_8 FILLER_27_438 ();
 sg13g2_decap_8 FILLER_27_445 ();
 sg13g2_decap_8 FILLER_27_452 ();
 sg13g2_decap_8 FILLER_27_459 ();
 sg13g2_decap_8 FILLER_27_466 ();
 sg13g2_decap_8 FILLER_27_473 ();
 sg13g2_decap_8 FILLER_27_480 ();
 sg13g2_decap_8 FILLER_27_487 ();
 sg13g2_decap_8 FILLER_27_494 ();
 sg13g2_decap_8 FILLER_27_501 ();
 sg13g2_decap_8 FILLER_27_508 ();
 sg13g2_decap_8 FILLER_27_515 ();
 sg13g2_decap_8 FILLER_27_522 ();
 sg13g2_decap_8 FILLER_27_529 ();
 sg13g2_decap_8 FILLER_27_536 ();
 sg13g2_decap_8 FILLER_27_543 ();
 sg13g2_decap_8 FILLER_27_550 ();
 sg13g2_decap_8 FILLER_27_557 ();
 sg13g2_decap_8 FILLER_27_564 ();
 sg13g2_decap_8 FILLER_27_571 ();
 sg13g2_decap_8 FILLER_27_578 ();
 sg13g2_decap_8 FILLER_27_585 ();
 sg13g2_decap_8 FILLER_27_592 ();
 sg13g2_decap_8 FILLER_27_599 ();
 sg13g2_decap_8 FILLER_27_606 ();
 sg13g2_decap_8 FILLER_27_613 ();
 sg13g2_decap_8 FILLER_27_620 ();
 sg13g2_decap_8 FILLER_27_627 ();
 sg13g2_decap_8 FILLER_27_634 ();
 sg13g2_decap_8 FILLER_27_641 ();
 sg13g2_decap_8 FILLER_27_648 ();
 sg13g2_decap_8 FILLER_27_655 ();
 sg13g2_decap_8 FILLER_27_662 ();
 sg13g2_decap_8 FILLER_27_669 ();
 sg13g2_decap_8 FILLER_27_676 ();
 sg13g2_decap_8 FILLER_27_683 ();
 sg13g2_decap_8 FILLER_27_690 ();
 sg13g2_decap_8 FILLER_27_697 ();
 sg13g2_decap_8 FILLER_27_704 ();
 sg13g2_decap_8 FILLER_27_711 ();
 sg13g2_decap_8 FILLER_27_718 ();
 sg13g2_decap_8 FILLER_27_725 ();
 sg13g2_decap_8 FILLER_27_732 ();
 sg13g2_decap_8 FILLER_27_739 ();
 sg13g2_decap_8 FILLER_27_746 ();
 sg13g2_decap_8 FILLER_27_753 ();
 sg13g2_decap_8 FILLER_27_760 ();
 sg13g2_decap_8 FILLER_27_767 ();
 sg13g2_decap_8 FILLER_27_774 ();
 sg13g2_decap_8 FILLER_27_781 ();
 sg13g2_decap_8 FILLER_27_788 ();
 sg13g2_decap_8 FILLER_27_795 ();
 sg13g2_decap_8 FILLER_27_802 ();
 sg13g2_decap_8 FILLER_27_809 ();
 sg13g2_decap_8 FILLER_27_816 ();
 sg13g2_decap_8 FILLER_27_823 ();
 sg13g2_decap_8 FILLER_27_830 ();
 sg13g2_decap_8 FILLER_27_837 ();
 sg13g2_decap_8 FILLER_27_844 ();
 sg13g2_decap_8 FILLER_27_851 ();
 sg13g2_decap_8 FILLER_27_858 ();
 sg13g2_decap_8 FILLER_27_865 ();
 sg13g2_decap_8 FILLER_27_872 ();
 sg13g2_decap_8 FILLER_27_879 ();
 sg13g2_decap_8 FILLER_27_886 ();
 sg13g2_decap_8 FILLER_27_893 ();
 sg13g2_decap_8 FILLER_27_900 ();
 sg13g2_decap_8 FILLER_27_907 ();
 sg13g2_decap_8 FILLER_27_914 ();
 sg13g2_decap_8 FILLER_27_921 ();
 sg13g2_decap_8 FILLER_27_928 ();
 sg13g2_decap_8 FILLER_27_935 ();
 sg13g2_decap_8 FILLER_27_942 ();
 sg13g2_decap_8 FILLER_27_949 ();
 sg13g2_decap_8 FILLER_27_956 ();
 sg13g2_decap_8 FILLER_27_963 ();
 sg13g2_decap_8 FILLER_27_970 ();
 sg13g2_decap_8 FILLER_27_977 ();
 sg13g2_decap_8 FILLER_27_984 ();
 sg13g2_decap_8 FILLER_27_991 ();
 sg13g2_decap_8 FILLER_27_998 ();
 sg13g2_decap_8 FILLER_27_1005 ();
 sg13g2_decap_8 FILLER_27_1012 ();
 sg13g2_decap_8 FILLER_27_1019 ();
 sg13g2_fill_2 FILLER_27_1026 ();
 sg13g2_fill_1 FILLER_27_1028 ();
 sg13g2_decap_8 FILLER_28_0 ();
 sg13g2_decap_8 FILLER_28_7 ();
 sg13g2_decap_8 FILLER_28_14 ();
 sg13g2_decap_8 FILLER_28_21 ();
 sg13g2_decap_8 FILLER_28_28 ();
 sg13g2_decap_8 FILLER_28_35 ();
 sg13g2_decap_8 FILLER_28_42 ();
 sg13g2_decap_8 FILLER_28_49 ();
 sg13g2_decap_8 FILLER_28_56 ();
 sg13g2_decap_8 FILLER_28_63 ();
 sg13g2_decap_8 FILLER_28_70 ();
 sg13g2_decap_8 FILLER_28_77 ();
 sg13g2_decap_8 FILLER_28_84 ();
 sg13g2_decap_8 FILLER_28_91 ();
 sg13g2_decap_8 FILLER_28_98 ();
 sg13g2_decap_8 FILLER_28_105 ();
 sg13g2_decap_8 FILLER_28_112 ();
 sg13g2_decap_8 FILLER_28_119 ();
 sg13g2_decap_8 FILLER_28_126 ();
 sg13g2_decap_8 FILLER_28_133 ();
 sg13g2_decap_8 FILLER_28_140 ();
 sg13g2_decap_8 FILLER_28_147 ();
 sg13g2_decap_8 FILLER_28_154 ();
 sg13g2_decap_8 FILLER_28_161 ();
 sg13g2_decap_8 FILLER_28_168 ();
 sg13g2_decap_8 FILLER_28_175 ();
 sg13g2_decap_8 FILLER_28_182 ();
 sg13g2_decap_8 FILLER_28_189 ();
 sg13g2_decap_8 FILLER_28_196 ();
 sg13g2_decap_8 FILLER_28_203 ();
 sg13g2_decap_8 FILLER_28_210 ();
 sg13g2_decap_8 FILLER_28_217 ();
 sg13g2_decap_8 FILLER_28_224 ();
 sg13g2_decap_8 FILLER_28_231 ();
 sg13g2_decap_8 FILLER_28_238 ();
 sg13g2_decap_8 FILLER_28_245 ();
 sg13g2_decap_8 FILLER_28_252 ();
 sg13g2_decap_8 FILLER_28_259 ();
 sg13g2_decap_8 FILLER_28_266 ();
 sg13g2_decap_8 FILLER_28_273 ();
 sg13g2_decap_8 FILLER_28_280 ();
 sg13g2_decap_8 FILLER_28_287 ();
 sg13g2_decap_8 FILLER_28_294 ();
 sg13g2_decap_8 FILLER_28_301 ();
 sg13g2_decap_8 FILLER_28_308 ();
 sg13g2_decap_8 FILLER_28_315 ();
 sg13g2_decap_8 FILLER_28_322 ();
 sg13g2_decap_8 FILLER_28_329 ();
 sg13g2_decap_8 FILLER_28_336 ();
 sg13g2_decap_8 FILLER_28_343 ();
 sg13g2_decap_8 FILLER_28_350 ();
 sg13g2_decap_8 FILLER_28_357 ();
 sg13g2_decap_8 FILLER_28_364 ();
 sg13g2_decap_8 FILLER_28_371 ();
 sg13g2_decap_8 FILLER_28_378 ();
 sg13g2_decap_8 FILLER_28_385 ();
 sg13g2_decap_8 FILLER_28_392 ();
 sg13g2_decap_8 FILLER_28_399 ();
 sg13g2_decap_8 FILLER_28_406 ();
 sg13g2_decap_8 FILLER_28_413 ();
 sg13g2_decap_8 FILLER_28_420 ();
 sg13g2_decap_8 FILLER_28_427 ();
 sg13g2_decap_8 FILLER_28_434 ();
 sg13g2_decap_8 FILLER_28_441 ();
 sg13g2_decap_8 FILLER_28_448 ();
 sg13g2_decap_8 FILLER_28_455 ();
 sg13g2_decap_8 FILLER_28_462 ();
 sg13g2_decap_8 FILLER_28_469 ();
 sg13g2_decap_8 FILLER_28_476 ();
 sg13g2_decap_8 FILLER_28_483 ();
 sg13g2_decap_8 FILLER_28_490 ();
 sg13g2_decap_8 FILLER_28_497 ();
 sg13g2_decap_8 FILLER_28_504 ();
 sg13g2_decap_8 FILLER_28_511 ();
 sg13g2_decap_8 FILLER_28_518 ();
 sg13g2_decap_8 FILLER_28_525 ();
 sg13g2_decap_8 FILLER_28_532 ();
 sg13g2_decap_8 FILLER_28_539 ();
 sg13g2_decap_8 FILLER_28_546 ();
 sg13g2_decap_8 FILLER_28_553 ();
 sg13g2_decap_8 FILLER_28_560 ();
 sg13g2_decap_8 FILLER_28_567 ();
 sg13g2_decap_8 FILLER_28_574 ();
 sg13g2_decap_8 FILLER_28_581 ();
 sg13g2_decap_8 FILLER_28_588 ();
 sg13g2_decap_8 FILLER_28_595 ();
 sg13g2_decap_8 FILLER_28_602 ();
 sg13g2_decap_8 FILLER_28_609 ();
 sg13g2_decap_8 FILLER_28_616 ();
 sg13g2_decap_8 FILLER_28_623 ();
 sg13g2_decap_8 FILLER_28_630 ();
 sg13g2_decap_8 FILLER_28_637 ();
 sg13g2_decap_8 FILLER_28_644 ();
 sg13g2_decap_8 FILLER_28_651 ();
 sg13g2_decap_8 FILLER_28_658 ();
 sg13g2_decap_8 FILLER_28_665 ();
 sg13g2_decap_8 FILLER_28_672 ();
 sg13g2_decap_8 FILLER_28_679 ();
 sg13g2_decap_8 FILLER_28_686 ();
 sg13g2_decap_8 FILLER_28_693 ();
 sg13g2_decap_8 FILLER_28_700 ();
 sg13g2_decap_8 FILLER_28_707 ();
 sg13g2_decap_8 FILLER_28_714 ();
 sg13g2_decap_8 FILLER_28_721 ();
 sg13g2_decap_8 FILLER_28_728 ();
 sg13g2_decap_8 FILLER_28_735 ();
 sg13g2_decap_8 FILLER_28_742 ();
 sg13g2_decap_8 FILLER_28_749 ();
 sg13g2_decap_8 FILLER_28_756 ();
 sg13g2_decap_8 FILLER_28_763 ();
 sg13g2_decap_8 FILLER_28_770 ();
 sg13g2_decap_8 FILLER_28_777 ();
 sg13g2_decap_8 FILLER_28_784 ();
 sg13g2_decap_8 FILLER_28_791 ();
 sg13g2_decap_8 FILLER_28_798 ();
 sg13g2_decap_8 FILLER_28_805 ();
 sg13g2_decap_8 FILLER_28_812 ();
 sg13g2_decap_8 FILLER_28_819 ();
 sg13g2_decap_8 FILLER_28_826 ();
 sg13g2_decap_8 FILLER_28_833 ();
 sg13g2_decap_8 FILLER_28_840 ();
 sg13g2_decap_8 FILLER_28_847 ();
 sg13g2_decap_8 FILLER_28_854 ();
 sg13g2_decap_8 FILLER_28_861 ();
 sg13g2_decap_8 FILLER_28_868 ();
 sg13g2_decap_8 FILLER_28_875 ();
 sg13g2_decap_8 FILLER_28_882 ();
 sg13g2_decap_8 FILLER_28_889 ();
 sg13g2_decap_8 FILLER_28_896 ();
 sg13g2_decap_8 FILLER_28_903 ();
 sg13g2_decap_8 FILLER_28_910 ();
 sg13g2_decap_8 FILLER_28_917 ();
 sg13g2_decap_8 FILLER_28_924 ();
 sg13g2_decap_8 FILLER_28_931 ();
 sg13g2_decap_8 FILLER_28_938 ();
 sg13g2_decap_8 FILLER_28_945 ();
 sg13g2_decap_8 FILLER_28_952 ();
 sg13g2_decap_8 FILLER_28_959 ();
 sg13g2_decap_8 FILLER_28_966 ();
 sg13g2_decap_8 FILLER_28_973 ();
 sg13g2_decap_8 FILLER_28_980 ();
 sg13g2_decap_8 FILLER_28_987 ();
 sg13g2_decap_8 FILLER_28_994 ();
 sg13g2_decap_8 FILLER_28_1001 ();
 sg13g2_decap_8 FILLER_28_1008 ();
 sg13g2_decap_8 FILLER_28_1015 ();
 sg13g2_decap_8 FILLER_28_1022 ();
 sg13g2_decap_8 FILLER_29_4 ();
 sg13g2_decap_8 FILLER_29_11 ();
 sg13g2_decap_8 FILLER_29_18 ();
 sg13g2_decap_8 FILLER_29_25 ();
 sg13g2_decap_8 FILLER_29_32 ();
 sg13g2_decap_8 FILLER_29_39 ();
 sg13g2_decap_8 FILLER_29_46 ();
 sg13g2_decap_8 FILLER_29_53 ();
 sg13g2_decap_8 FILLER_29_60 ();
 sg13g2_decap_8 FILLER_29_67 ();
 sg13g2_decap_8 FILLER_29_74 ();
 sg13g2_decap_8 FILLER_29_81 ();
 sg13g2_decap_8 FILLER_29_88 ();
 sg13g2_decap_8 FILLER_29_95 ();
 sg13g2_decap_8 FILLER_29_102 ();
 sg13g2_decap_8 FILLER_29_109 ();
 sg13g2_decap_8 FILLER_29_116 ();
 sg13g2_decap_8 FILLER_29_123 ();
 sg13g2_decap_8 FILLER_29_130 ();
 sg13g2_decap_8 FILLER_29_137 ();
 sg13g2_decap_8 FILLER_29_144 ();
 sg13g2_decap_8 FILLER_29_151 ();
 sg13g2_decap_8 FILLER_29_158 ();
 sg13g2_decap_8 FILLER_29_165 ();
 sg13g2_decap_8 FILLER_29_172 ();
 sg13g2_decap_8 FILLER_29_179 ();
 sg13g2_decap_8 FILLER_29_186 ();
 sg13g2_decap_8 FILLER_29_193 ();
 sg13g2_decap_8 FILLER_29_200 ();
 sg13g2_decap_8 FILLER_29_207 ();
 sg13g2_decap_8 FILLER_29_214 ();
 sg13g2_decap_8 FILLER_29_221 ();
 sg13g2_decap_8 FILLER_29_228 ();
 sg13g2_decap_8 FILLER_29_235 ();
 sg13g2_decap_8 FILLER_29_242 ();
 sg13g2_decap_8 FILLER_29_249 ();
 sg13g2_decap_8 FILLER_29_256 ();
 sg13g2_decap_8 FILLER_29_263 ();
 sg13g2_decap_8 FILLER_29_270 ();
 sg13g2_decap_8 FILLER_29_277 ();
 sg13g2_decap_8 FILLER_29_284 ();
 sg13g2_decap_8 FILLER_29_291 ();
 sg13g2_decap_8 FILLER_29_298 ();
 sg13g2_decap_8 FILLER_29_305 ();
 sg13g2_decap_8 FILLER_29_312 ();
 sg13g2_decap_8 FILLER_29_319 ();
 sg13g2_decap_8 FILLER_29_326 ();
 sg13g2_decap_8 FILLER_29_333 ();
 sg13g2_decap_8 FILLER_29_340 ();
 sg13g2_decap_8 FILLER_29_347 ();
 sg13g2_decap_8 FILLER_29_354 ();
 sg13g2_decap_8 FILLER_29_361 ();
 sg13g2_decap_8 FILLER_29_368 ();
 sg13g2_decap_8 FILLER_29_375 ();
 sg13g2_decap_8 FILLER_29_382 ();
 sg13g2_decap_8 FILLER_29_389 ();
 sg13g2_decap_8 FILLER_29_396 ();
 sg13g2_decap_8 FILLER_29_403 ();
 sg13g2_decap_8 FILLER_29_410 ();
 sg13g2_decap_8 FILLER_29_417 ();
 sg13g2_decap_8 FILLER_29_424 ();
 sg13g2_decap_8 FILLER_29_431 ();
 sg13g2_decap_8 FILLER_29_438 ();
 sg13g2_decap_8 FILLER_29_445 ();
 sg13g2_decap_8 FILLER_29_452 ();
 sg13g2_decap_8 FILLER_29_459 ();
 sg13g2_decap_8 FILLER_29_466 ();
 sg13g2_decap_8 FILLER_29_473 ();
 sg13g2_decap_8 FILLER_29_480 ();
 sg13g2_decap_8 FILLER_29_487 ();
 sg13g2_decap_8 FILLER_29_494 ();
 sg13g2_decap_8 FILLER_29_501 ();
 sg13g2_decap_8 FILLER_29_508 ();
 sg13g2_decap_8 FILLER_29_515 ();
 sg13g2_decap_8 FILLER_29_522 ();
 sg13g2_decap_8 FILLER_29_529 ();
 sg13g2_decap_8 FILLER_29_536 ();
 sg13g2_decap_8 FILLER_29_543 ();
 sg13g2_decap_8 FILLER_29_550 ();
 sg13g2_decap_8 FILLER_29_557 ();
 sg13g2_decap_8 FILLER_29_564 ();
 sg13g2_decap_8 FILLER_29_571 ();
 sg13g2_decap_8 FILLER_29_578 ();
 sg13g2_decap_8 FILLER_29_585 ();
 sg13g2_decap_8 FILLER_29_592 ();
 sg13g2_decap_8 FILLER_29_599 ();
 sg13g2_decap_8 FILLER_29_606 ();
 sg13g2_decap_8 FILLER_29_613 ();
 sg13g2_decap_8 FILLER_29_620 ();
 sg13g2_decap_8 FILLER_29_627 ();
 sg13g2_decap_8 FILLER_29_634 ();
 sg13g2_decap_8 FILLER_29_641 ();
 sg13g2_decap_8 FILLER_29_648 ();
 sg13g2_decap_8 FILLER_29_655 ();
 sg13g2_decap_8 FILLER_29_662 ();
 sg13g2_decap_8 FILLER_29_669 ();
 sg13g2_decap_8 FILLER_29_676 ();
 sg13g2_decap_8 FILLER_29_683 ();
 sg13g2_decap_8 FILLER_29_690 ();
 sg13g2_decap_8 FILLER_29_697 ();
 sg13g2_decap_8 FILLER_29_704 ();
 sg13g2_decap_8 FILLER_29_711 ();
 sg13g2_decap_8 FILLER_29_718 ();
 sg13g2_decap_8 FILLER_29_725 ();
 sg13g2_decap_8 FILLER_29_732 ();
 sg13g2_decap_8 FILLER_29_739 ();
 sg13g2_decap_8 FILLER_29_746 ();
 sg13g2_decap_8 FILLER_29_753 ();
 sg13g2_decap_8 FILLER_29_760 ();
 sg13g2_decap_8 FILLER_29_767 ();
 sg13g2_decap_8 FILLER_29_774 ();
 sg13g2_decap_8 FILLER_29_781 ();
 sg13g2_decap_8 FILLER_29_788 ();
 sg13g2_decap_8 FILLER_29_795 ();
 sg13g2_decap_8 FILLER_29_802 ();
 sg13g2_decap_8 FILLER_29_809 ();
 sg13g2_decap_8 FILLER_29_816 ();
 sg13g2_decap_8 FILLER_29_823 ();
 sg13g2_decap_8 FILLER_29_830 ();
 sg13g2_decap_8 FILLER_29_837 ();
 sg13g2_decap_8 FILLER_29_844 ();
 sg13g2_decap_8 FILLER_29_851 ();
 sg13g2_decap_8 FILLER_29_858 ();
 sg13g2_decap_8 FILLER_29_865 ();
 sg13g2_decap_8 FILLER_29_872 ();
 sg13g2_decap_8 FILLER_29_879 ();
 sg13g2_decap_8 FILLER_29_886 ();
 sg13g2_decap_8 FILLER_29_893 ();
 sg13g2_decap_8 FILLER_29_900 ();
 sg13g2_decap_8 FILLER_29_907 ();
 sg13g2_decap_8 FILLER_29_914 ();
 sg13g2_decap_8 FILLER_29_921 ();
 sg13g2_decap_8 FILLER_29_928 ();
 sg13g2_decap_8 FILLER_29_935 ();
 sg13g2_decap_8 FILLER_29_942 ();
 sg13g2_decap_8 FILLER_29_949 ();
 sg13g2_decap_8 FILLER_29_956 ();
 sg13g2_decap_8 FILLER_29_963 ();
 sg13g2_decap_8 FILLER_29_970 ();
 sg13g2_decap_8 FILLER_29_977 ();
 sg13g2_decap_8 FILLER_29_984 ();
 sg13g2_decap_8 FILLER_29_991 ();
 sg13g2_decap_8 FILLER_29_998 ();
 sg13g2_decap_8 FILLER_29_1005 ();
 sg13g2_decap_8 FILLER_29_1012 ();
 sg13g2_decap_8 FILLER_29_1019 ();
 sg13g2_fill_2 FILLER_29_1026 ();
 sg13g2_fill_1 FILLER_29_1028 ();
 sg13g2_decap_8 FILLER_30_0 ();
 sg13g2_decap_8 FILLER_30_7 ();
 sg13g2_decap_8 FILLER_30_14 ();
 sg13g2_decap_8 FILLER_30_21 ();
 sg13g2_decap_8 FILLER_30_28 ();
 sg13g2_decap_8 FILLER_30_35 ();
 sg13g2_decap_8 FILLER_30_42 ();
 sg13g2_decap_8 FILLER_30_49 ();
 sg13g2_decap_8 FILLER_30_56 ();
 sg13g2_decap_8 FILLER_30_63 ();
 sg13g2_decap_8 FILLER_30_70 ();
 sg13g2_decap_8 FILLER_30_77 ();
 sg13g2_decap_8 FILLER_30_84 ();
 sg13g2_decap_8 FILLER_30_91 ();
 sg13g2_decap_8 FILLER_30_98 ();
 sg13g2_decap_8 FILLER_30_105 ();
 sg13g2_decap_8 FILLER_30_112 ();
 sg13g2_decap_8 FILLER_30_119 ();
 sg13g2_decap_8 FILLER_30_126 ();
 sg13g2_decap_8 FILLER_30_133 ();
 sg13g2_decap_8 FILLER_30_140 ();
 sg13g2_decap_8 FILLER_30_147 ();
 sg13g2_decap_8 FILLER_30_154 ();
 sg13g2_decap_8 FILLER_30_161 ();
 sg13g2_decap_8 FILLER_30_168 ();
 sg13g2_decap_8 FILLER_30_175 ();
 sg13g2_decap_8 FILLER_30_182 ();
 sg13g2_decap_8 FILLER_30_189 ();
 sg13g2_decap_8 FILLER_30_196 ();
 sg13g2_decap_8 FILLER_30_203 ();
 sg13g2_decap_8 FILLER_30_210 ();
 sg13g2_decap_8 FILLER_30_217 ();
 sg13g2_decap_8 FILLER_30_224 ();
 sg13g2_decap_8 FILLER_30_231 ();
 sg13g2_decap_8 FILLER_30_238 ();
 sg13g2_decap_8 FILLER_30_245 ();
 sg13g2_decap_8 FILLER_30_252 ();
 sg13g2_decap_8 FILLER_30_259 ();
 sg13g2_decap_8 FILLER_30_266 ();
 sg13g2_decap_8 FILLER_30_273 ();
 sg13g2_decap_8 FILLER_30_280 ();
 sg13g2_decap_8 FILLER_30_287 ();
 sg13g2_decap_8 FILLER_30_294 ();
 sg13g2_decap_8 FILLER_30_301 ();
 sg13g2_decap_8 FILLER_30_308 ();
 sg13g2_decap_8 FILLER_30_315 ();
 sg13g2_decap_8 FILLER_30_322 ();
 sg13g2_decap_8 FILLER_30_329 ();
 sg13g2_decap_8 FILLER_30_336 ();
 sg13g2_decap_8 FILLER_30_343 ();
 sg13g2_decap_8 FILLER_30_350 ();
 sg13g2_decap_8 FILLER_30_357 ();
 sg13g2_decap_8 FILLER_30_364 ();
 sg13g2_decap_8 FILLER_30_371 ();
 sg13g2_decap_8 FILLER_30_378 ();
 sg13g2_decap_8 FILLER_30_385 ();
 sg13g2_decap_8 FILLER_30_392 ();
 sg13g2_decap_8 FILLER_30_399 ();
 sg13g2_decap_8 FILLER_30_406 ();
 sg13g2_decap_8 FILLER_30_413 ();
 sg13g2_decap_8 FILLER_30_420 ();
 sg13g2_decap_8 FILLER_30_427 ();
 sg13g2_decap_8 FILLER_30_434 ();
 sg13g2_decap_8 FILLER_30_441 ();
 sg13g2_decap_8 FILLER_30_448 ();
 sg13g2_decap_8 FILLER_30_455 ();
 sg13g2_decap_8 FILLER_30_462 ();
 sg13g2_decap_8 FILLER_30_469 ();
 sg13g2_decap_8 FILLER_30_476 ();
 sg13g2_decap_8 FILLER_30_483 ();
 sg13g2_decap_8 FILLER_30_490 ();
 sg13g2_decap_8 FILLER_30_497 ();
 sg13g2_decap_8 FILLER_30_504 ();
 sg13g2_decap_8 FILLER_30_511 ();
 sg13g2_decap_8 FILLER_30_518 ();
 sg13g2_decap_8 FILLER_30_525 ();
 sg13g2_decap_8 FILLER_30_532 ();
 sg13g2_decap_8 FILLER_30_539 ();
 sg13g2_decap_8 FILLER_30_546 ();
 sg13g2_decap_8 FILLER_30_553 ();
 sg13g2_decap_8 FILLER_30_560 ();
 sg13g2_decap_8 FILLER_30_567 ();
 sg13g2_decap_8 FILLER_30_574 ();
 sg13g2_decap_8 FILLER_30_581 ();
 sg13g2_decap_8 FILLER_30_588 ();
 sg13g2_decap_8 FILLER_30_595 ();
 sg13g2_decap_8 FILLER_30_602 ();
 sg13g2_decap_8 FILLER_30_609 ();
 sg13g2_decap_8 FILLER_30_616 ();
 sg13g2_decap_8 FILLER_30_623 ();
 sg13g2_decap_8 FILLER_30_630 ();
 sg13g2_decap_8 FILLER_30_637 ();
 sg13g2_decap_8 FILLER_30_644 ();
 sg13g2_decap_8 FILLER_30_651 ();
 sg13g2_decap_8 FILLER_30_658 ();
 sg13g2_decap_8 FILLER_30_665 ();
 sg13g2_decap_8 FILLER_30_672 ();
 sg13g2_decap_8 FILLER_30_679 ();
 sg13g2_decap_8 FILLER_30_686 ();
 sg13g2_decap_8 FILLER_30_693 ();
 sg13g2_decap_8 FILLER_30_700 ();
 sg13g2_decap_8 FILLER_30_707 ();
 sg13g2_decap_8 FILLER_30_714 ();
 sg13g2_decap_8 FILLER_30_721 ();
 sg13g2_decap_8 FILLER_30_728 ();
 sg13g2_decap_8 FILLER_30_735 ();
 sg13g2_decap_8 FILLER_30_742 ();
 sg13g2_decap_8 FILLER_30_749 ();
 sg13g2_decap_8 FILLER_30_756 ();
 sg13g2_decap_8 FILLER_30_763 ();
 sg13g2_decap_8 FILLER_30_770 ();
 sg13g2_decap_8 FILLER_30_777 ();
 sg13g2_decap_8 FILLER_30_784 ();
 sg13g2_decap_8 FILLER_30_791 ();
 sg13g2_decap_8 FILLER_30_798 ();
 sg13g2_decap_8 FILLER_30_805 ();
 sg13g2_decap_8 FILLER_30_812 ();
 sg13g2_decap_8 FILLER_30_819 ();
 sg13g2_decap_8 FILLER_30_826 ();
 sg13g2_decap_8 FILLER_30_833 ();
 sg13g2_decap_8 FILLER_30_840 ();
 sg13g2_decap_8 FILLER_30_847 ();
 sg13g2_decap_8 FILLER_30_854 ();
 sg13g2_decap_8 FILLER_30_861 ();
 sg13g2_decap_8 FILLER_30_868 ();
 sg13g2_decap_8 FILLER_30_875 ();
 sg13g2_decap_8 FILLER_30_882 ();
 sg13g2_decap_8 FILLER_30_889 ();
 sg13g2_decap_8 FILLER_30_896 ();
 sg13g2_decap_8 FILLER_30_903 ();
 sg13g2_decap_8 FILLER_30_910 ();
 sg13g2_decap_8 FILLER_30_917 ();
 sg13g2_decap_8 FILLER_30_924 ();
 sg13g2_decap_8 FILLER_30_931 ();
 sg13g2_decap_8 FILLER_30_938 ();
 sg13g2_decap_8 FILLER_30_945 ();
 sg13g2_decap_8 FILLER_30_952 ();
 sg13g2_decap_8 FILLER_30_959 ();
 sg13g2_decap_8 FILLER_30_966 ();
 sg13g2_decap_8 FILLER_30_973 ();
 sg13g2_decap_8 FILLER_30_980 ();
 sg13g2_decap_8 FILLER_30_987 ();
 sg13g2_decap_8 FILLER_30_994 ();
 sg13g2_decap_8 FILLER_30_1001 ();
 sg13g2_decap_8 FILLER_30_1008 ();
 sg13g2_decap_8 FILLER_30_1015 ();
 sg13g2_decap_8 FILLER_30_1022 ();
 sg13g2_decap_8 FILLER_31_0 ();
 sg13g2_decap_8 FILLER_31_7 ();
 sg13g2_decap_8 FILLER_31_14 ();
 sg13g2_decap_8 FILLER_31_21 ();
 sg13g2_decap_8 FILLER_31_28 ();
 sg13g2_decap_8 FILLER_31_35 ();
 sg13g2_decap_8 FILLER_31_42 ();
 sg13g2_decap_8 FILLER_31_49 ();
 sg13g2_decap_8 FILLER_31_56 ();
 sg13g2_decap_8 FILLER_31_63 ();
 sg13g2_decap_8 FILLER_31_70 ();
 sg13g2_decap_8 FILLER_31_77 ();
 sg13g2_decap_8 FILLER_31_84 ();
 sg13g2_decap_8 FILLER_31_91 ();
 sg13g2_decap_8 FILLER_31_98 ();
 sg13g2_decap_8 FILLER_31_105 ();
 sg13g2_decap_8 FILLER_31_112 ();
 sg13g2_decap_8 FILLER_31_119 ();
 sg13g2_decap_8 FILLER_31_126 ();
 sg13g2_decap_8 FILLER_31_133 ();
 sg13g2_decap_8 FILLER_31_140 ();
 sg13g2_decap_8 FILLER_31_147 ();
 sg13g2_decap_8 FILLER_31_154 ();
 sg13g2_decap_8 FILLER_31_161 ();
 sg13g2_decap_8 FILLER_31_168 ();
 sg13g2_decap_8 FILLER_31_175 ();
 sg13g2_decap_8 FILLER_31_182 ();
 sg13g2_decap_8 FILLER_31_189 ();
 sg13g2_decap_8 FILLER_31_196 ();
 sg13g2_decap_8 FILLER_31_203 ();
 sg13g2_decap_8 FILLER_31_210 ();
 sg13g2_decap_8 FILLER_31_217 ();
 sg13g2_decap_8 FILLER_31_224 ();
 sg13g2_decap_8 FILLER_31_231 ();
 sg13g2_decap_8 FILLER_31_238 ();
 sg13g2_decap_8 FILLER_31_245 ();
 sg13g2_decap_8 FILLER_31_252 ();
 sg13g2_decap_8 FILLER_31_259 ();
 sg13g2_decap_8 FILLER_31_266 ();
 sg13g2_decap_8 FILLER_31_273 ();
 sg13g2_decap_8 FILLER_31_280 ();
 sg13g2_decap_8 FILLER_31_287 ();
 sg13g2_decap_8 FILLER_31_294 ();
 sg13g2_decap_8 FILLER_31_301 ();
 sg13g2_decap_8 FILLER_31_308 ();
 sg13g2_decap_8 FILLER_31_315 ();
 sg13g2_decap_8 FILLER_31_322 ();
 sg13g2_decap_8 FILLER_31_329 ();
 sg13g2_decap_8 FILLER_31_336 ();
 sg13g2_decap_8 FILLER_31_343 ();
 sg13g2_decap_8 FILLER_31_350 ();
 sg13g2_decap_8 FILLER_31_357 ();
 sg13g2_decap_8 FILLER_31_364 ();
 sg13g2_decap_8 FILLER_31_371 ();
 sg13g2_decap_8 FILLER_31_378 ();
 sg13g2_decap_8 FILLER_31_385 ();
 sg13g2_decap_8 FILLER_31_392 ();
 sg13g2_decap_8 FILLER_31_399 ();
 sg13g2_decap_8 FILLER_31_406 ();
 sg13g2_decap_8 FILLER_31_413 ();
 sg13g2_decap_8 FILLER_31_420 ();
 sg13g2_decap_8 FILLER_31_427 ();
 sg13g2_decap_8 FILLER_31_434 ();
 sg13g2_decap_8 FILLER_31_441 ();
 sg13g2_decap_8 FILLER_31_448 ();
 sg13g2_decap_8 FILLER_31_455 ();
 sg13g2_decap_8 FILLER_31_462 ();
 sg13g2_decap_8 FILLER_31_469 ();
 sg13g2_decap_8 FILLER_31_476 ();
 sg13g2_decap_8 FILLER_31_483 ();
 sg13g2_decap_8 FILLER_31_490 ();
 sg13g2_decap_8 FILLER_31_497 ();
 sg13g2_decap_8 FILLER_31_504 ();
 sg13g2_decap_8 FILLER_31_511 ();
 sg13g2_decap_8 FILLER_31_518 ();
 sg13g2_decap_8 FILLER_31_525 ();
 sg13g2_decap_8 FILLER_31_532 ();
 sg13g2_decap_8 FILLER_31_539 ();
 sg13g2_decap_8 FILLER_31_546 ();
 sg13g2_decap_8 FILLER_31_553 ();
 sg13g2_decap_8 FILLER_31_560 ();
 sg13g2_decap_8 FILLER_31_567 ();
 sg13g2_decap_8 FILLER_31_574 ();
 sg13g2_decap_8 FILLER_31_581 ();
 sg13g2_decap_8 FILLER_31_588 ();
 sg13g2_decap_8 FILLER_31_595 ();
 sg13g2_decap_8 FILLER_31_602 ();
 sg13g2_decap_8 FILLER_31_609 ();
 sg13g2_decap_8 FILLER_31_616 ();
 sg13g2_decap_8 FILLER_31_623 ();
 sg13g2_decap_8 FILLER_31_630 ();
 sg13g2_decap_8 FILLER_31_637 ();
 sg13g2_decap_8 FILLER_31_644 ();
 sg13g2_decap_8 FILLER_31_651 ();
 sg13g2_decap_8 FILLER_31_658 ();
 sg13g2_decap_8 FILLER_31_665 ();
 sg13g2_decap_8 FILLER_31_672 ();
 sg13g2_decap_8 FILLER_31_679 ();
 sg13g2_decap_8 FILLER_31_686 ();
 sg13g2_decap_8 FILLER_31_693 ();
 sg13g2_decap_8 FILLER_31_700 ();
 sg13g2_decap_8 FILLER_31_707 ();
 sg13g2_decap_8 FILLER_31_714 ();
 sg13g2_decap_8 FILLER_31_721 ();
 sg13g2_decap_8 FILLER_31_728 ();
 sg13g2_decap_8 FILLER_31_735 ();
 sg13g2_decap_8 FILLER_31_742 ();
 sg13g2_decap_8 FILLER_31_749 ();
 sg13g2_decap_8 FILLER_31_756 ();
 sg13g2_decap_8 FILLER_31_763 ();
 sg13g2_decap_8 FILLER_31_770 ();
 sg13g2_decap_8 FILLER_31_777 ();
 sg13g2_decap_8 FILLER_31_784 ();
 sg13g2_decap_8 FILLER_31_791 ();
 sg13g2_decap_8 FILLER_31_798 ();
 sg13g2_decap_8 FILLER_31_805 ();
 sg13g2_decap_8 FILLER_31_812 ();
 sg13g2_decap_8 FILLER_31_819 ();
 sg13g2_decap_8 FILLER_31_826 ();
 sg13g2_decap_8 FILLER_31_833 ();
 sg13g2_decap_8 FILLER_31_840 ();
 sg13g2_decap_8 FILLER_31_847 ();
 sg13g2_decap_8 FILLER_31_854 ();
 sg13g2_decap_8 FILLER_31_861 ();
 sg13g2_decap_8 FILLER_31_868 ();
 sg13g2_decap_8 FILLER_31_875 ();
 sg13g2_decap_8 FILLER_31_882 ();
 sg13g2_decap_8 FILLER_31_889 ();
 sg13g2_decap_8 FILLER_31_896 ();
 sg13g2_decap_8 FILLER_31_903 ();
 sg13g2_decap_8 FILLER_31_910 ();
 sg13g2_decap_8 FILLER_31_917 ();
 sg13g2_decap_8 FILLER_31_924 ();
 sg13g2_decap_8 FILLER_31_931 ();
 sg13g2_decap_8 FILLER_31_938 ();
 sg13g2_decap_8 FILLER_31_945 ();
 sg13g2_decap_8 FILLER_31_952 ();
 sg13g2_decap_8 FILLER_31_959 ();
 sg13g2_decap_8 FILLER_31_966 ();
 sg13g2_decap_8 FILLER_31_973 ();
 sg13g2_decap_8 FILLER_31_980 ();
 sg13g2_decap_8 FILLER_31_987 ();
 sg13g2_decap_8 FILLER_31_994 ();
 sg13g2_decap_8 FILLER_31_1001 ();
 sg13g2_decap_8 FILLER_31_1008 ();
 sg13g2_decap_8 FILLER_31_1015 ();
 sg13g2_decap_8 FILLER_31_1022 ();
 sg13g2_decap_8 FILLER_32_4 ();
 sg13g2_decap_8 FILLER_32_11 ();
 sg13g2_decap_8 FILLER_32_18 ();
 sg13g2_decap_8 FILLER_32_25 ();
 sg13g2_decap_8 FILLER_32_32 ();
 sg13g2_decap_8 FILLER_32_39 ();
 sg13g2_decap_8 FILLER_32_46 ();
 sg13g2_decap_8 FILLER_32_53 ();
 sg13g2_decap_8 FILLER_32_60 ();
 sg13g2_decap_8 FILLER_32_67 ();
 sg13g2_decap_8 FILLER_32_74 ();
 sg13g2_decap_8 FILLER_32_81 ();
 sg13g2_decap_8 FILLER_32_88 ();
 sg13g2_decap_8 FILLER_32_95 ();
 sg13g2_decap_8 FILLER_32_102 ();
 sg13g2_decap_8 FILLER_32_109 ();
 sg13g2_decap_8 FILLER_32_116 ();
 sg13g2_decap_8 FILLER_32_123 ();
 sg13g2_decap_8 FILLER_32_130 ();
 sg13g2_decap_8 FILLER_32_137 ();
 sg13g2_decap_8 FILLER_32_144 ();
 sg13g2_decap_8 FILLER_32_151 ();
 sg13g2_decap_8 FILLER_32_158 ();
 sg13g2_decap_8 FILLER_32_165 ();
 sg13g2_decap_8 FILLER_32_172 ();
 sg13g2_decap_8 FILLER_32_179 ();
 sg13g2_decap_8 FILLER_32_186 ();
 sg13g2_decap_8 FILLER_32_193 ();
 sg13g2_decap_8 FILLER_32_200 ();
 sg13g2_decap_8 FILLER_32_207 ();
 sg13g2_decap_8 FILLER_32_214 ();
 sg13g2_decap_8 FILLER_32_221 ();
 sg13g2_decap_8 FILLER_32_228 ();
 sg13g2_decap_8 FILLER_32_235 ();
 sg13g2_decap_8 FILLER_32_242 ();
 sg13g2_decap_8 FILLER_32_249 ();
 sg13g2_decap_8 FILLER_32_256 ();
 sg13g2_decap_8 FILLER_32_263 ();
 sg13g2_decap_8 FILLER_32_270 ();
 sg13g2_decap_8 FILLER_32_277 ();
 sg13g2_decap_8 FILLER_32_284 ();
 sg13g2_decap_8 FILLER_32_291 ();
 sg13g2_decap_8 FILLER_32_298 ();
 sg13g2_decap_8 FILLER_32_305 ();
 sg13g2_decap_8 FILLER_32_312 ();
 sg13g2_decap_8 FILLER_32_319 ();
 sg13g2_decap_8 FILLER_32_326 ();
 sg13g2_decap_8 FILLER_32_333 ();
 sg13g2_decap_8 FILLER_32_340 ();
 sg13g2_decap_8 FILLER_32_347 ();
 sg13g2_decap_8 FILLER_32_354 ();
 sg13g2_decap_8 FILLER_32_361 ();
 sg13g2_decap_8 FILLER_32_368 ();
 sg13g2_decap_8 FILLER_32_375 ();
 sg13g2_decap_8 FILLER_32_382 ();
 sg13g2_decap_8 FILLER_32_389 ();
 sg13g2_decap_8 FILLER_32_396 ();
 sg13g2_decap_8 FILLER_32_403 ();
 sg13g2_decap_8 FILLER_32_410 ();
 sg13g2_decap_8 FILLER_32_417 ();
 sg13g2_decap_8 FILLER_32_424 ();
 sg13g2_decap_8 FILLER_32_431 ();
 sg13g2_decap_8 FILLER_32_438 ();
 sg13g2_decap_8 FILLER_32_445 ();
 sg13g2_decap_8 FILLER_32_452 ();
 sg13g2_decap_8 FILLER_32_459 ();
 sg13g2_decap_8 FILLER_32_466 ();
 sg13g2_decap_8 FILLER_32_473 ();
 sg13g2_decap_8 FILLER_32_480 ();
 sg13g2_decap_8 FILLER_32_487 ();
 sg13g2_decap_8 FILLER_32_494 ();
 sg13g2_decap_8 FILLER_32_501 ();
 sg13g2_decap_8 FILLER_32_508 ();
 sg13g2_decap_8 FILLER_32_515 ();
 sg13g2_decap_8 FILLER_32_522 ();
 sg13g2_decap_8 FILLER_32_529 ();
 sg13g2_decap_8 FILLER_32_536 ();
 sg13g2_decap_8 FILLER_32_543 ();
 sg13g2_decap_8 FILLER_32_550 ();
 sg13g2_decap_8 FILLER_32_557 ();
 sg13g2_decap_8 FILLER_32_564 ();
 sg13g2_decap_8 FILLER_32_571 ();
 sg13g2_decap_8 FILLER_32_578 ();
 sg13g2_decap_8 FILLER_32_585 ();
 sg13g2_decap_8 FILLER_32_592 ();
 sg13g2_decap_8 FILLER_32_599 ();
 sg13g2_decap_8 FILLER_32_606 ();
 sg13g2_decap_8 FILLER_32_613 ();
 sg13g2_decap_8 FILLER_32_620 ();
 sg13g2_decap_8 FILLER_32_627 ();
 sg13g2_decap_8 FILLER_32_634 ();
 sg13g2_decap_8 FILLER_32_641 ();
 sg13g2_decap_8 FILLER_32_648 ();
 sg13g2_decap_8 FILLER_32_655 ();
 sg13g2_decap_8 FILLER_32_662 ();
 sg13g2_decap_8 FILLER_32_669 ();
 sg13g2_decap_8 FILLER_32_676 ();
 sg13g2_decap_8 FILLER_32_683 ();
 sg13g2_decap_8 FILLER_32_690 ();
 sg13g2_decap_8 FILLER_32_697 ();
 sg13g2_decap_8 FILLER_32_704 ();
 sg13g2_decap_8 FILLER_32_711 ();
 sg13g2_decap_8 FILLER_32_718 ();
 sg13g2_decap_8 FILLER_32_725 ();
 sg13g2_decap_8 FILLER_32_732 ();
 sg13g2_decap_8 FILLER_32_739 ();
 sg13g2_decap_8 FILLER_32_746 ();
 sg13g2_decap_8 FILLER_32_753 ();
 sg13g2_decap_8 FILLER_32_760 ();
 sg13g2_decap_8 FILLER_32_767 ();
 sg13g2_decap_8 FILLER_32_774 ();
 sg13g2_decap_8 FILLER_32_781 ();
 sg13g2_decap_8 FILLER_32_788 ();
 sg13g2_decap_8 FILLER_32_795 ();
 sg13g2_decap_8 FILLER_32_802 ();
 sg13g2_decap_8 FILLER_32_809 ();
 sg13g2_decap_8 FILLER_32_816 ();
 sg13g2_decap_8 FILLER_32_823 ();
 sg13g2_decap_8 FILLER_32_830 ();
 sg13g2_decap_8 FILLER_32_837 ();
 sg13g2_decap_8 FILLER_32_844 ();
 sg13g2_decap_8 FILLER_32_851 ();
 sg13g2_decap_8 FILLER_32_858 ();
 sg13g2_decap_8 FILLER_32_865 ();
 sg13g2_decap_8 FILLER_32_872 ();
 sg13g2_decap_8 FILLER_32_879 ();
 sg13g2_decap_8 FILLER_32_886 ();
 sg13g2_decap_8 FILLER_32_893 ();
 sg13g2_decap_8 FILLER_32_900 ();
 sg13g2_decap_8 FILLER_32_907 ();
 sg13g2_decap_8 FILLER_32_914 ();
 sg13g2_decap_8 FILLER_32_921 ();
 sg13g2_decap_8 FILLER_32_928 ();
 sg13g2_decap_8 FILLER_32_935 ();
 sg13g2_decap_8 FILLER_32_942 ();
 sg13g2_decap_8 FILLER_32_949 ();
 sg13g2_decap_8 FILLER_32_956 ();
 sg13g2_decap_8 FILLER_32_963 ();
 sg13g2_decap_8 FILLER_32_970 ();
 sg13g2_decap_8 FILLER_32_977 ();
 sg13g2_decap_8 FILLER_32_984 ();
 sg13g2_decap_8 FILLER_32_991 ();
 sg13g2_decap_8 FILLER_32_998 ();
 sg13g2_decap_8 FILLER_32_1005 ();
 sg13g2_decap_8 FILLER_32_1012 ();
 sg13g2_decap_8 FILLER_32_1019 ();
 sg13g2_fill_2 FILLER_32_1026 ();
 sg13g2_fill_1 FILLER_32_1028 ();
 sg13g2_decap_8 FILLER_33_0 ();
 sg13g2_decap_8 FILLER_33_7 ();
 sg13g2_decap_8 FILLER_33_14 ();
 sg13g2_decap_8 FILLER_33_21 ();
 sg13g2_decap_8 FILLER_33_28 ();
 sg13g2_decap_8 FILLER_33_35 ();
 sg13g2_decap_8 FILLER_33_42 ();
 sg13g2_decap_8 FILLER_33_49 ();
 sg13g2_decap_8 FILLER_33_56 ();
 sg13g2_decap_8 FILLER_33_63 ();
 sg13g2_decap_8 FILLER_33_70 ();
 sg13g2_decap_8 FILLER_33_77 ();
 sg13g2_decap_8 FILLER_33_84 ();
 sg13g2_decap_8 FILLER_33_91 ();
 sg13g2_decap_8 FILLER_33_98 ();
 sg13g2_decap_8 FILLER_33_105 ();
 sg13g2_decap_8 FILLER_33_112 ();
 sg13g2_decap_8 FILLER_33_119 ();
 sg13g2_decap_8 FILLER_33_126 ();
 sg13g2_decap_8 FILLER_33_133 ();
 sg13g2_decap_8 FILLER_33_140 ();
 sg13g2_decap_8 FILLER_33_147 ();
 sg13g2_decap_8 FILLER_33_154 ();
 sg13g2_decap_8 FILLER_33_161 ();
 sg13g2_decap_8 FILLER_33_168 ();
 sg13g2_decap_8 FILLER_33_175 ();
 sg13g2_decap_8 FILLER_33_182 ();
 sg13g2_decap_8 FILLER_33_189 ();
 sg13g2_decap_8 FILLER_33_196 ();
 sg13g2_decap_8 FILLER_33_203 ();
 sg13g2_decap_8 FILLER_33_210 ();
 sg13g2_decap_8 FILLER_33_217 ();
 sg13g2_decap_8 FILLER_33_224 ();
 sg13g2_decap_8 FILLER_33_231 ();
 sg13g2_decap_8 FILLER_33_238 ();
 sg13g2_decap_8 FILLER_33_245 ();
 sg13g2_decap_8 FILLER_33_252 ();
 sg13g2_decap_8 FILLER_33_259 ();
 sg13g2_decap_8 FILLER_33_266 ();
 sg13g2_decap_8 FILLER_33_273 ();
 sg13g2_decap_8 FILLER_33_280 ();
 sg13g2_decap_8 FILLER_33_287 ();
 sg13g2_decap_8 FILLER_33_294 ();
 sg13g2_decap_8 FILLER_33_301 ();
 sg13g2_decap_8 FILLER_33_308 ();
 sg13g2_decap_8 FILLER_33_315 ();
 sg13g2_decap_8 FILLER_33_322 ();
 sg13g2_decap_8 FILLER_33_329 ();
 sg13g2_decap_8 FILLER_33_336 ();
 sg13g2_decap_8 FILLER_33_343 ();
 sg13g2_decap_8 FILLER_33_350 ();
 sg13g2_decap_8 FILLER_33_357 ();
 sg13g2_decap_8 FILLER_33_364 ();
 sg13g2_decap_8 FILLER_33_371 ();
 sg13g2_decap_8 FILLER_33_378 ();
 sg13g2_decap_8 FILLER_33_385 ();
 sg13g2_decap_8 FILLER_33_392 ();
 sg13g2_decap_8 FILLER_33_399 ();
 sg13g2_decap_8 FILLER_33_406 ();
 sg13g2_decap_8 FILLER_33_413 ();
 sg13g2_decap_8 FILLER_33_420 ();
 sg13g2_decap_8 FILLER_33_427 ();
 sg13g2_decap_8 FILLER_33_434 ();
 sg13g2_decap_8 FILLER_33_441 ();
 sg13g2_decap_8 FILLER_33_448 ();
 sg13g2_decap_8 FILLER_33_455 ();
 sg13g2_decap_8 FILLER_33_462 ();
 sg13g2_decap_8 FILLER_33_469 ();
 sg13g2_decap_8 FILLER_33_476 ();
 sg13g2_decap_8 FILLER_33_483 ();
 sg13g2_decap_8 FILLER_33_490 ();
 sg13g2_decap_8 FILLER_33_497 ();
 sg13g2_decap_8 FILLER_33_504 ();
 sg13g2_decap_8 FILLER_33_511 ();
 sg13g2_decap_8 FILLER_33_518 ();
 sg13g2_decap_8 FILLER_33_525 ();
 sg13g2_decap_8 FILLER_33_532 ();
 sg13g2_decap_8 FILLER_33_539 ();
 sg13g2_decap_8 FILLER_33_546 ();
 sg13g2_decap_8 FILLER_33_553 ();
 sg13g2_decap_8 FILLER_33_560 ();
 sg13g2_decap_8 FILLER_33_567 ();
 sg13g2_decap_8 FILLER_33_574 ();
 sg13g2_decap_8 FILLER_33_581 ();
 sg13g2_decap_8 FILLER_33_588 ();
 sg13g2_decap_8 FILLER_33_595 ();
 sg13g2_decap_8 FILLER_33_602 ();
 sg13g2_decap_8 FILLER_33_609 ();
 sg13g2_decap_8 FILLER_33_616 ();
 sg13g2_decap_8 FILLER_33_623 ();
 sg13g2_decap_8 FILLER_33_630 ();
 sg13g2_decap_8 FILLER_33_637 ();
 sg13g2_decap_8 FILLER_33_644 ();
 sg13g2_decap_8 FILLER_33_651 ();
 sg13g2_decap_8 FILLER_33_658 ();
 sg13g2_decap_8 FILLER_33_665 ();
 sg13g2_decap_8 FILLER_33_672 ();
 sg13g2_decap_8 FILLER_33_679 ();
 sg13g2_decap_8 FILLER_33_686 ();
 sg13g2_decap_8 FILLER_33_693 ();
 sg13g2_decap_8 FILLER_33_700 ();
 sg13g2_decap_8 FILLER_33_707 ();
 sg13g2_decap_8 FILLER_33_714 ();
 sg13g2_decap_8 FILLER_33_721 ();
 sg13g2_decap_8 FILLER_33_728 ();
 sg13g2_decap_8 FILLER_33_735 ();
 sg13g2_decap_8 FILLER_33_742 ();
 sg13g2_decap_8 FILLER_33_749 ();
 sg13g2_decap_8 FILLER_33_756 ();
 sg13g2_decap_8 FILLER_33_763 ();
 sg13g2_decap_8 FILLER_33_770 ();
 sg13g2_decap_8 FILLER_33_777 ();
 sg13g2_decap_8 FILLER_33_784 ();
 sg13g2_decap_8 FILLER_33_791 ();
 sg13g2_decap_8 FILLER_33_798 ();
 sg13g2_decap_8 FILLER_33_805 ();
 sg13g2_decap_8 FILLER_33_812 ();
 sg13g2_decap_8 FILLER_33_819 ();
 sg13g2_decap_8 FILLER_33_826 ();
 sg13g2_decap_8 FILLER_33_833 ();
 sg13g2_decap_8 FILLER_33_840 ();
 sg13g2_decap_8 FILLER_33_847 ();
 sg13g2_decap_8 FILLER_33_854 ();
 sg13g2_decap_8 FILLER_33_861 ();
 sg13g2_decap_8 FILLER_33_868 ();
 sg13g2_decap_8 FILLER_33_875 ();
 sg13g2_decap_8 FILLER_33_882 ();
 sg13g2_decap_8 FILLER_33_889 ();
 sg13g2_decap_8 FILLER_33_896 ();
 sg13g2_decap_8 FILLER_33_903 ();
 sg13g2_decap_8 FILLER_33_910 ();
 sg13g2_decap_8 FILLER_33_917 ();
 sg13g2_decap_8 FILLER_33_924 ();
 sg13g2_decap_8 FILLER_33_931 ();
 sg13g2_decap_8 FILLER_33_938 ();
 sg13g2_decap_8 FILLER_33_945 ();
 sg13g2_decap_8 FILLER_33_952 ();
 sg13g2_decap_8 FILLER_33_959 ();
 sg13g2_decap_8 FILLER_33_966 ();
 sg13g2_decap_8 FILLER_33_973 ();
 sg13g2_decap_8 FILLER_33_980 ();
 sg13g2_decap_8 FILLER_33_987 ();
 sg13g2_decap_8 FILLER_33_994 ();
 sg13g2_decap_8 FILLER_33_1001 ();
 sg13g2_decap_8 FILLER_33_1008 ();
 sg13g2_decap_8 FILLER_33_1015 ();
 sg13g2_decap_8 FILLER_33_1022 ();
 sg13g2_decap_8 FILLER_34_4 ();
 sg13g2_decap_8 FILLER_34_11 ();
 sg13g2_decap_8 FILLER_34_18 ();
 sg13g2_decap_8 FILLER_34_25 ();
 sg13g2_decap_8 FILLER_34_32 ();
 sg13g2_decap_8 FILLER_34_39 ();
 sg13g2_decap_8 FILLER_34_46 ();
 sg13g2_decap_8 FILLER_34_53 ();
 sg13g2_decap_8 FILLER_34_60 ();
 sg13g2_decap_8 FILLER_34_67 ();
 sg13g2_decap_8 FILLER_34_74 ();
 sg13g2_decap_8 FILLER_34_81 ();
 sg13g2_decap_8 FILLER_34_88 ();
 sg13g2_decap_8 FILLER_34_95 ();
 sg13g2_decap_8 FILLER_34_102 ();
 sg13g2_decap_8 FILLER_34_109 ();
 sg13g2_decap_8 FILLER_34_116 ();
 sg13g2_decap_8 FILLER_34_123 ();
 sg13g2_decap_8 FILLER_34_130 ();
 sg13g2_decap_8 FILLER_34_137 ();
 sg13g2_decap_8 FILLER_34_144 ();
 sg13g2_decap_8 FILLER_34_151 ();
 sg13g2_decap_8 FILLER_34_158 ();
 sg13g2_decap_8 FILLER_34_165 ();
 sg13g2_decap_8 FILLER_34_172 ();
 sg13g2_decap_8 FILLER_34_179 ();
 sg13g2_decap_8 FILLER_34_186 ();
 sg13g2_decap_8 FILLER_34_193 ();
 sg13g2_decap_8 FILLER_34_200 ();
 sg13g2_decap_8 FILLER_34_207 ();
 sg13g2_decap_8 FILLER_34_214 ();
 sg13g2_decap_8 FILLER_34_221 ();
 sg13g2_decap_8 FILLER_34_228 ();
 sg13g2_decap_8 FILLER_34_235 ();
 sg13g2_decap_8 FILLER_34_242 ();
 sg13g2_decap_8 FILLER_34_249 ();
 sg13g2_decap_8 FILLER_34_256 ();
 sg13g2_decap_8 FILLER_34_263 ();
 sg13g2_decap_8 FILLER_34_270 ();
 sg13g2_decap_8 FILLER_34_277 ();
 sg13g2_decap_8 FILLER_34_284 ();
 sg13g2_decap_8 FILLER_34_291 ();
 sg13g2_decap_8 FILLER_34_298 ();
 sg13g2_decap_8 FILLER_34_305 ();
 sg13g2_decap_8 FILLER_34_312 ();
 sg13g2_decap_8 FILLER_34_319 ();
 sg13g2_decap_8 FILLER_34_326 ();
 sg13g2_decap_8 FILLER_34_333 ();
 sg13g2_decap_8 FILLER_34_340 ();
 sg13g2_decap_8 FILLER_34_347 ();
 sg13g2_decap_8 FILLER_34_354 ();
 sg13g2_decap_8 FILLER_34_361 ();
 sg13g2_decap_8 FILLER_34_368 ();
 sg13g2_decap_8 FILLER_34_375 ();
 sg13g2_decap_8 FILLER_34_382 ();
 sg13g2_decap_8 FILLER_34_389 ();
 sg13g2_decap_8 FILLER_34_396 ();
 sg13g2_decap_8 FILLER_34_403 ();
 sg13g2_decap_8 FILLER_34_410 ();
 sg13g2_decap_8 FILLER_34_417 ();
 sg13g2_decap_8 FILLER_34_424 ();
 sg13g2_decap_8 FILLER_34_431 ();
 sg13g2_decap_8 FILLER_34_438 ();
 sg13g2_decap_8 FILLER_34_445 ();
 sg13g2_decap_8 FILLER_34_452 ();
 sg13g2_decap_8 FILLER_34_459 ();
 sg13g2_decap_8 FILLER_34_466 ();
 sg13g2_decap_8 FILLER_34_473 ();
 sg13g2_decap_8 FILLER_34_480 ();
 sg13g2_decap_8 FILLER_34_487 ();
 sg13g2_decap_8 FILLER_34_494 ();
 sg13g2_decap_8 FILLER_34_501 ();
 sg13g2_decap_8 FILLER_34_508 ();
 sg13g2_decap_8 FILLER_34_515 ();
 sg13g2_decap_8 FILLER_34_522 ();
 sg13g2_decap_8 FILLER_34_529 ();
 sg13g2_decap_8 FILLER_34_536 ();
 sg13g2_decap_8 FILLER_34_543 ();
 sg13g2_decap_8 FILLER_34_550 ();
 sg13g2_decap_8 FILLER_34_557 ();
 sg13g2_decap_8 FILLER_34_564 ();
 sg13g2_decap_8 FILLER_34_571 ();
 sg13g2_decap_8 FILLER_34_578 ();
 sg13g2_decap_8 FILLER_34_585 ();
 sg13g2_decap_8 FILLER_34_592 ();
 sg13g2_decap_8 FILLER_34_599 ();
 sg13g2_decap_8 FILLER_34_606 ();
 sg13g2_decap_8 FILLER_34_613 ();
 sg13g2_decap_8 FILLER_34_620 ();
 sg13g2_decap_8 FILLER_34_627 ();
 sg13g2_decap_8 FILLER_34_634 ();
 sg13g2_decap_8 FILLER_34_641 ();
 sg13g2_decap_8 FILLER_34_648 ();
 sg13g2_decap_8 FILLER_34_655 ();
 sg13g2_decap_8 FILLER_34_662 ();
 sg13g2_decap_8 FILLER_34_669 ();
 sg13g2_decap_8 FILLER_34_676 ();
 sg13g2_decap_8 FILLER_34_683 ();
 sg13g2_decap_8 FILLER_34_690 ();
 sg13g2_decap_8 FILLER_34_697 ();
 sg13g2_decap_8 FILLER_34_704 ();
 sg13g2_decap_8 FILLER_34_711 ();
 sg13g2_decap_8 FILLER_34_718 ();
 sg13g2_decap_8 FILLER_34_725 ();
 sg13g2_decap_8 FILLER_34_732 ();
 sg13g2_decap_8 FILLER_34_739 ();
 sg13g2_decap_8 FILLER_34_746 ();
 sg13g2_decap_8 FILLER_34_753 ();
 sg13g2_decap_8 FILLER_34_760 ();
 sg13g2_decap_8 FILLER_34_767 ();
 sg13g2_decap_8 FILLER_34_774 ();
 sg13g2_decap_8 FILLER_34_781 ();
 sg13g2_decap_8 FILLER_34_788 ();
 sg13g2_decap_8 FILLER_34_795 ();
 sg13g2_decap_8 FILLER_34_802 ();
 sg13g2_decap_8 FILLER_34_809 ();
 sg13g2_decap_8 FILLER_34_816 ();
 sg13g2_decap_8 FILLER_34_823 ();
 sg13g2_decap_8 FILLER_34_830 ();
 sg13g2_decap_8 FILLER_34_837 ();
 sg13g2_decap_8 FILLER_34_844 ();
 sg13g2_decap_8 FILLER_34_851 ();
 sg13g2_decap_8 FILLER_34_858 ();
 sg13g2_decap_8 FILLER_34_865 ();
 sg13g2_decap_8 FILLER_34_872 ();
 sg13g2_decap_8 FILLER_34_879 ();
 sg13g2_decap_8 FILLER_34_886 ();
 sg13g2_decap_8 FILLER_34_893 ();
 sg13g2_decap_8 FILLER_34_900 ();
 sg13g2_decap_8 FILLER_34_907 ();
 sg13g2_decap_8 FILLER_34_914 ();
 sg13g2_decap_8 FILLER_34_921 ();
 sg13g2_decap_8 FILLER_34_928 ();
 sg13g2_decap_8 FILLER_34_935 ();
 sg13g2_decap_8 FILLER_34_942 ();
 sg13g2_decap_8 FILLER_34_949 ();
 sg13g2_decap_8 FILLER_34_956 ();
 sg13g2_decap_8 FILLER_34_963 ();
 sg13g2_decap_8 FILLER_34_970 ();
 sg13g2_decap_8 FILLER_34_977 ();
 sg13g2_decap_8 FILLER_34_984 ();
 sg13g2_decap_8 FILLER_34_991 ();
 sg13g2_decap_8 FILLER_34_998 ();
 sg13g2_decap_8 FILLER_34_1005 ();
 sg13g2_decap_8 FILLER_34_1012 ();
 sg13g2_decap_8 FILLER_34_1019 ();
 sg13g2_fill_2 FILLER_34_1026 ();
 sg13g2_fill_1 FILLER_34_1028 ();
 sg13g2_decap_8 FILLER_35_0 ();
 sg13g2_decap_8 FILLER_35_7 ();
 sg13g2_decap_8 FILLER_35_14 ();
 sg13g2_decap_8 FILLER_35_21 ();
 sg13g2_decap_8 FILLER_35_28 ();
 sg13g2_decap_8 FILLER_35_35 ();
 sg13g2_decap_8 FILLER_35_42 ();
 sg13g2_decap_8 FILLER_35_49 ();
 sg13g2_decap_8 FILLER_35_56 ();
 sg13g2_decap_8 FILLER_35_63 ();
 sg13g2_decap_8 FILLER_35_70 ();
 sg13g2_decap_8 FILLER_35_77 ();
 sg13g2_decap_8 FILLER_35_84 ();
 sg13g2_decap_8 FILLER_35_91 ();
 sg13g2_decap_8 FILLER_35_98 ();
 sg13g2_decap_8 FILLER_35_105 ();
 sg13g2_decap_8 FILLER_35_112 ();
 sg13g2_decap_8 FILLER_35_119 ();
 sg13g2_decap_8 FILLER_35_126 ();
 sg13g2_decap_8 FILLER_35_133 ();
 sg13g2_decap_8 FILLER_35_140 ();
 sg13g2_decap_8 FILLER_35_147 ();
 sg13g2_decap_8 FILLER_35_154 ();
 sg13g2_decap_8 FILLER_35_161 ();
 sg13g2_decap_8 FILLER_35_168 ();
 sg13g2_decap_8 FILLER_35_175 ();
 sg13g2_decap_8 FILLER_35_182 ();
 sg13g2_decap_8 FILLER_35_189 ();
 sg13g2_decap_8 FILLER_35_196 ();
 sg13g2_decap_8 FILLER_35_203 ();
 sg13g2_decap_8 FILLER_35_210 ();
 sg13g2_decap_8 FILLER_35_217 ();
 sg13g2_decap_8 FILLER_35_224 ();
 sg13g2_decap_8 FILLER_35_231 ();
 sg13g2_decap_8 FILLER_35_238 ();
 sg13g2_decap_8 FILLER_35_245 ();
 sg13g2_decap_8 FILLER_35_252 ();
 sg13g2_decap_8 FILLER_35_259 ();
 sg13g2_decap_8 FILLER_35_266 ();
 sg13g2_decap_8 FILLER_35_273 ();
 sg13g2_decap_8 FILLER_35_280 ();
 sg13g2_decap_8 FILLER_35_287 ();
 sg13g2_decap_8 FILLER_35_294 ();
 sg13g2_decap_8 FILLER_35_301 ();
 sg13g2_decap_8 FILLER_35_308 ();
 sg13g2_decap_8 FILLER_35_315 ();
 sg13g2_decap_8 FILLER_35_322 ();
 sg13g2_decap_8 FILLER_35_329 ();
 sg13g2_decap_8 FILLER_35_336 ();
 sg13g2_decap_8 FILLER_35_343 ();
 sg13g2_decap_8 FILLER_35_350 ();
 sg13g2_decap_8 FILLER_35_357 ();
 sg13g2_decap_8 FILLER_35_364 ();
 sg13g2_decap_8 FILLER_35_371 ();
 sg13g2_decap_8 FILLER_35_378 ();
 sg13g2_decap_8 FILLER_35_385 ();
 sg13g2_decap_8 FILLER_35_392 ();
 sg13g2_decap_8 FILLER_35_399 ();
 sg13g2_decap_8 FILLER_35_406 ();
 sg13g2_decap_8 FILLER_35_413 ();
 sg13g2_decap_8 FILLER_35_420 ();
 sg13g2_decap_8 FILLER_35_427 ();
 sg13g2_decap_8 FILLER_35_434 ();
 sg13g2_decap_8 FILLER_35_441 ();
 sg13g2_decap_8 FILLER_35_448 ();
 sg13g2_decap_8 FILLER_35_455 ();
 sg13g2_decap_8 FILLER_35_462 ();
 sg13g2_decap_8 FILLER_35_469 ();
 sg13g2_decap_8 FILLER_35_476 ();
 sg13g2_decap_8 FILLER_35_483 ();
 sg13g2_decap_8 FILLER_35_490 ();
 sg13g2_decap_8 FILLER_35_497 ();
 sg13g2_decap_8 FILLER_35_504 ();
 sg13g2_decap_8 FILLER_35_511 ();
 sg13g2_decap_8 FILLER_35_518 ();
 sg13g2_decap_8 FILLER_35_525 ();
 sg13g2_decap_8 FILLER_35_532 ();
 sg13g2_decap_8 FILLER_35_539 ();
 sg13g2_decap_8 FILLER_35_546 ();
 sg13g2_decap_8 FILLER_35_553 ();
 sg13g2_decap_8 FILLER_35_560 ();
 sg13g2_decap_8 FILLER_35_567 ();
 sg13g2_decap_8 FILLER_35_574 ();
 sg13g2_decap_8 FILLER_35_581 ();
 sg13g2_decap_8 FILLER_35_588 ();
 sg13g2_decap_8 FILLER_35_595 ();
 sg13g2_decap_8 FILLER_35_602 ();
 sg13g2_decap_8 FILLER_35_609 ();
 sg13g2_decap_8 FILLER_35_616 ();
 sg13g2_decap_8 FILLER_35_623 ();
 sg13g2_decap_8 FILLER_35_630 ();
 sg13g2_decap_8 FILLER_35_637 ();
 sg13g2_decap_8 FILLER_35_644 ();
 sg13g2_decap_8 FILLER_35_651 ();
 sg13g2_decap_8 FILLER_35_658 ();
 sg13g2_decap_8 FILLER_35_665 ();
 sg13g2_decap_8 FILLER_35_672 ();
 sg13g2_decap_8 FILLER_35_679 ();
 sg13g2_decap_8 FILLER_35_686 ();
 sg13g2_decap_8 FILLER_35_693 ();
 sg13g2_decap_8 FILLER_35_700 ();
 sg13g2_decap_8 FILLER_35_707 ();
 sg13g2_decap_8 FILLER_35_714 ();
 sg13g2_decap_8 FILLER_35_721 ();
 sg13g2_decap_8 FILLER_35_728 ();
 sg13g2_decap_8 FILLER_35_735 ();
 sg13g2_decap_8 FILLER_35_742 ();
 sg13g2_decap_8 FILLER_35_749 ();
 sg13g2_decap_8 FILLER_35_756 ();
 sg13g2_decap_8 FILLER_35_763 ();
 sg13g2_decap_8 FILLER_35_770 ();
 sg13g2_decap_8 FILLER_35_777 ();
 sg13g2_decap_8 FILLER_35_784 ();
 sg13g2_decap_8 FILLER_35_791 ();
 sg13g2_decap_8 FILLER_35_798 ();
 sg13g2_decap_8 FILLER_35_805 ();
 sg13g2_decap_8 FILLER_35_812 ();
 sg13g2_decap_8 FILLER_35_819 ();
 sg13g2_decap_8 FILLER_35_826 ();
 sg13g2_decap_8 FILLER_35_833 ();
 sg13g2_decap_8 FILLER_35_840 ();
 sg13g2_decap_8 FILLER_35_847 ();
 sg13g2_decap_8 FILLER_35_854 ();
 sg13g2_decap_8 FILLER_35_861 ();
 sg13g2_decap_8 FILLER_35_868 ();
 sg13g2_decap_8 FILLER_35_875 ();
 sg13g2_decap_8 FILLER_35_882 ();
 sg13g2_decap_8 FILLER_35_889 ();
 sg13g2_decap_8 FILLER_35_896 ();
 sg13g2_decap_8 FILLER_35_903 ();
 sg13g2_decap_8 FILLER_35_910 ();
 sg13g2_decap_8 FILLER_35_917 ();
 sg13g2_decap_8 FILLER_35_924 ();
 sg13g2_decap_8 FILLER_35_931 ();
 sg13g2_decap_8 FILLER_35_938 ();
 sg13g2_decap_8 FILLER_35_945 ();
 sg13g2_decap_8 FILLER_35_952 ();
 sg13g2_decap_8 FILLER_35_959 ();
 sg13g2_decap_8 FILLER_35_966 ();
 sg13g2_decap_8 FILLER_35_973 ();
 sg13g2_decap_8 FILLER_35_980 ();
 sg13g2_decap_8 FILLER_35_987 ();
 sg13g2_decap_8 FILLER_35_994 ();
 sg13g2_decap_8 FILLER_35_1001 ();
 sg13g2_decap_8 FILLER_35_1008 ();
 sg13g2_decap_8 FILLER_35_1015 ();
 sg13g2_decap_8 FILLER_35_1022 ();
 sg13g2_decap_8 FILLER_36_0 ();
 sg13g2_decap_8 FILLER_36_7 ();
 sg13g2_decap_8 FILLER_36_14 ();
 sg13g2_decap_8 FILLER_36_21 ();
 sg13g2_decap_8 FILLER_36_28 ();
 sg13g2_decap_8 FILLER_36_35 ();
 sg13g2_decap_8 FILLER_36_42 ();
 sg13g2_decap_8 FILLER_36_49 ();
 sg13g2_decap_8 FILLER_36_56 ();
 sg13g2_decap_8 FILLER_36_63 ();
 sg13g2_decap_8 FILLER_36_70 ();
 sg13g2_decap_8 FILLER_36_77 ();
 sg13g2_decap_8 FILLER_36_84 ();
 sg13g2_decap_8 FILLER_36_91 ();
 sg13g2_decap_8 FILLER_36_98 ();
 sg13g2_decap_8 FILLER_36_105 ();
 sg13g2_decap_8 FILLER_36_112 ();
 sg13g2_decap_8 FILLER_36_119 ();
 sg13g2_decap_8 FILLER_36_126 ();
 sg13g2_decap_8 FILLER_36_133 ();
 sg13g2_decap_8 FILLER_36_140 ();
 sg13g2_decap_8 FILLER_36_147 ();
 sg13g2_decap_8 FILLER_36_154 ();
 sg13g2_decap_8 FILLER_36_161 ();
 sg13g2_decap_8 FILLER_36_168 ();
 sg13g2_decap_8 FILLER_36_175 ();
 sg13g2_decap_8 FILLER_36_182 ();
 sg13g2_decap_8 FILLER_36_189 ();
 sg13g2_decap_8 FILLER_36_196 ();
 sg13g2_decap_8 FILLER_36_203 ();
 sg13g2_decap_8 FILLER_36_210 ();
 sg13g2_decap_8 FILLER_36_217 ();
 sg13g2_decap_8 FILLER_36_224 ();
 sg13g2_decap_8 FILLER_36_231 ();
 sg13g2_decap_8 FILLER_36_238 ();
 sg13g2_decap_8 FILLER_36_245 ();
 sg13g2_decap_8 FILLER_36_252 ();
 sg13g2_decap_8 FILLER_36_259 ();
 sg13g2_decap_8 FILLER_36_266 ();
 sg13g2_decap_8 FILLER_36_273 ();
 sg13g2_decap_8 FILLER_36_280 ();
 sg13g2_decap_8 FILLER_36_287 ();
 sg13g2_decap_8 FILLER_36_294 ();
 sg13g2_decap_8 FILLER_36_301 ();
 sg13g2_decap_8 FILLER_36_308 ();
 sg13g2_decap_8 FILLER_36_315 ();
 sg13g2_decap_8 FILLER_36_322 ();
 sg13g2_decap_8 FILLER_36_329 ();
 sg13g2_decap_8 FILLER_36_336 ();
 sg13g2_decap_8 FILLER_36_343 ();
 sg13g2_decap_8 FILLER_36_350 ();
 sg13g2_decap_8 FILLER_36_357 ();
 sg13g2_decap_8 FILLER_36_364 ();
 sg13g2_decap_8 FILLER_36_371 ();
 sg13g2_decap_8 FILLER_36_378 ();
 sg13g2_decap_8 FILLER_36_385 ();
 sg13g2_decap_8 FILLER_36_392 ();
 sg13g2_decap_8 FILLER_36_399 ();
 sg13g2_decap_8 FILLER_36_406 ();
 sg13g2_decap_8 FILLER_36_413 ();
 sg13g2_decap_8 FILLER_36_420 ();
 sg13g2_decap_8 FILLER_36_427 ();
 sg13g2_decap_8 FILLER_36_434 ();
 sg13g2_decap_8 FILLER_36_441 ();
 sg13g2_decap_8 FILLER_36_448 ();
 sg13g2_decap_8 FILLER_36_455 ();
 sg13g2_decap_8 FILLER_36_462 ();
 sg13g2_decap_8 FILLER_36_469 ();
 sg13g2_decap_8 FILLER_36_476 ();
 sg13g2_decap_8 FILLER_36_483 ();
 sg13g2_decap_8 FILLER_36_490 ();
 sg13g2_decap_8 FILLER_36_497 ();
 sg13g2_decap_8 FILLER_36_504 ();
 sg13g2_decap_8 FILLER_36_511 ();
 sg13g2_decap_8 FILLER_36_518 ();
 sg13g2_decap_8 FILLER_36_525 ();
 sg13g2_decap_8 FILLER_36_532 ();
 sg13g2_decap_8 FILLER_36_539 ();
 sg13g2_decap_8 FILLER_36_546 ();
 sg13g2_decap_8 FILLER_36_553 ();
 sg13g2_decap_8 FILLER_36_560 ();
 sg13g2_decap_8 FILLER_36_567 ();
 sg13g2_decap_8 FILLER_36_574 ();
 sg13g2_decap_8 FILLER_36_581 ();
 sg13g2_decap_8 FILLER_36_588 ();
 sg13g2_decap_8 FILLER_36_595 ();
 sg13g2_decap_8 FILLER_36_602 ();
 sg13g2_decap_8 FILLER_36_609 ();
 sg13g2_decap_8 FILLER_36_616 ();
 sg13g2_decap_8 FILLER_36_623 ();
 sg13g2_decap_8 FILLER_36_630 ();
 sg13g2_decap_8 FILLER_36_637 ();
 sg13g2_decap_8 FILLER_36_644 ();
 sg13g2_decap_8 FILLER_36_651 ();
 sg13g2_decap_8 FILLER_36_658 ();
 sg13g2_decap_8 FILLER_36_665 ();
 sg13g2_decap_8 FILLER_36_672 ();
 sg13g2_decap_8 FILLER_36_679 ();
 sg13g2_decap_8 FILLER_36_686 ();
 sg13g2_decap_8 FILLER_36_693 ();
 sg13g2_decap_8 FILLER_36_700 ();
 sg13g2_decap_8 FILLER_36_707 ();
 sg13g2_decap_8 FILLER_36_714 ();
 sg13g2_decap_8 FILLER_36_721 ();
 sg13g2_decap_8 FILLER_36_728 ();
 sg13g2_decap_8 FILLER_36_735 ();
 sg13g2_decap_8 FILLER_36_742 ();
 sg13g2_decap_8 FILLER_36_749 ();
 sg13g2_decap_8 FILLER_36_756 ();
 sg13g2_decap_8 FILLER_36_763 ();
 sg13g2_decap_8 FILLER_36_770 ();
 sg13g2_decap_8 FILLER_36_777 ();
 sg13g2_decap_8 FILLER_36_784 ();
 sg13g2_decap_8 FILLER_36_791 ();
 sg13g2_decap_8 FILLER_36_798 ();
 sg13g2_decap_8 FILLER_36_805 ();
 sg13g2_decap_8 FILLER_36_812 ();
 sg13g2_decap_8 FILLER_36_819 ();
 sg13g2_decap_8 FILLER_36_826 ();
 sg13g2_decap_8 FILLER_36_833 ();
 sg13g2_decap_8 FILLER_36_840 ();
 sg13g2_decap_8 FILLER_36_847 ();
 sg13g2_decap_8 FILLER_36_854 ();
 sg13g2_decap_8 FILLER_36_861 ();
 sg13g2_decap_8 FILLER_36_868 ();
 sg13g2_decap_8 FILLER_36_875 ();
 sg13g2_decap_8 FILLER_36_882 ();
 sg13g2_decap_8 FILLER_36_889 ();
 sg13g2_decap_8 FILLER_36_896 ();
 sg13g2_decap_8 FILLER_36_903 ();
 sg13g2_decap_8 FILLER_36_910 ();
 sg13g2_decap_8 FILLER_36_917 ();
 sg13g2_decap_8 FILLER_36_924 ();
 sg13g2_decap_8 FILLER_36_931 ();
 sg13g2_decap_8 FILLER_36_938 ();
 sg13g2_decap_8 FILLER_36_945 ();
 sg13g2_decap_8 FILLER_36_952 ();
 sg13g2_decap_8 FILLER_36_959 ();
 sg13g2_decap_8 FILLER_36_966 ();
 sg13g2_decap_8 FILLER_36_973 ();
 sg13g2_decap_8 FILLER_36_980 ();
 sg13g2_decap_8 FILLER_36_987 ();
 sg13g2_decap_8 FILLER_36_994 ();
 sg13g2_decap_8 FILLER_36_1001 ();
 sg13g2_decap_8 FILLER_36_1008 ();
 sg13g2_decap_8 FILLER_36_1015 ();
 sg13g2_decap_8 FILLER_36_1022 ();
 sg13g2_decap_8 FILLER_37_4 ();
 sg13g2_decap_8 FILLER_37_11 ();
 sg13g2_decap_8 FILLER_37_18 ();
 sg13g2_decap_8 FILLER_37_25 ();
 sg13g2_decap_8 FILLER_37_32 ();
 sg13g2_decap_8 FILLER_37_39 ();
 sg13g2_decap_8 FILLER_37_46 ();
 sg13g2_decap_8 FILLER_37_53 ();
 sg13g2_decap_8 FILLER_37_60 ();
 sg13g2_decap_8 FILLER_37_67 ();
 sg13g2_decap_8 FILLER_37_74 ();
 sg13g2_decap_8 FILLER_37_81 ();
 sg13g2_decap_8 FILLER_37_88 ();
 sg13g2_decap_8 FILLER_37_95 ();
 sg13g2_decap_8 FILLER_37_102 ();
 sg13g2_decap_8 FILLER_37_109 ();
 sg13g2_decap_8 FILLER_37_116 ();
 sg13g2_decap_8 FILLER_37_123 ();
 sg13g2_decap_8 FILLER_37_130 ();
 sg13g2_decap_8 FILLER_37_137 ();
 sg13g2_decap_8 FILLER_37_144 ();
 sg13g2_decap_8 FILLER_37_151 ();
 sg13g2_decap_8 FILLER_37_158 ();
 sg13g2_decap_8 FILLER_37_165 ();
 sg13g2_decap_8 FILLER_37_172 ();
 sg13g2_decap_8 FILLER_37_179 ();
 sg13g2_decap_8 FILLER_37_186 ();
 sg13g2_decap_8 FILLER_37_193 ();
 sg13g2_decap_8 FILLER_37_200 ();
 sg13g2_decap_8 FILLER_37_207 ();
 sg13g2_decap_8 FILLER_37_214 ();
 sg13g2_decap_8 FILLER_37_221 ();
 sg13g2_decap_8 FILLER_37_228 ();
 sg13g2_decap_8 FILLER_37_235 ();
 sg13g2_decap_8 FILLER_37_242 ();
 sg13g2_decap_8 FILLER_37_249 ();
 sg13g2_decap_8 FILLER_37_256 ();
 sg13g2_decap_8 FILLER_37_263 ();
 sg13g2_decap_8 FILLER_37_270 ();
 sg13g2_decap_8 FILLER_37_277 ();
 sg13g2_decap_8 FILLER_37_284 ();
 sg13g2_decap_8 FILLER_37_291 ();
 sg13g2_decap_8 FILLER_37_298 ();
 sg13g2_decap_8 FILLER_37_305 ();
 sg13g2_decap_8 FILLER_37_312 ();
 sg13g2_decap_8 FILLER_37_319 ();
 sg13g2_decap_8 FILLER_37_326 ();
 sg13g2_decap_8 FILLER_37_333 ();
 sg13g2_decap_8 FILLER_37_340 ();
 sg13g2_decap_8 FILLER_37_347 ();
 sg13g2_decap_8 FILLER_37_354 ();
 sg13g2_decap_8 FILLER_37_361 ();
 sg13g2_decap_8 FILLER_37_368 ();
 sg13g2_decap_8 FILLER_37_375 ();
 sg13g2_decap_8 FILLER_37_382 ();
 sg13g2_decap_8 FILLER_37_389 ();
 sg13g2_decap_8 FILLER_37_396 ();
 sg13g2_decap_8 FILLER_37_403 ();
 sg13g2_decap_8 FILLER_37_410 ();
 sg13g2_decap_8 FILLER_37_417 ();
 sg13g2_decap_8 FILLER_37_424 ();
 sg13g2_decap_8 FILLER_37_431 ();
 sg13g2_decap_8 FILLER_37_438 ();
 sg13g2_decap_8 FILLER_37_445 ();
 sg13g2_decap_8 FILLER_37_452 ();
 sg13g2_decap_8 FILLER_37_459 ();
 sg13g2_decap_8 FILLER_37_466 ();
 sg13g2_decap_8 FILLER_37_473 ();
 sg13g2_decap_8 FILLER_37_480 ();
 sg13g2_decap_8 FILLER_37_487 ();
 sg13g2_decap_8 FILLER_37_494 ();
 sg13g2_decap_8 FILLER_37_501 ();
 sg13g2_decap_8 FILLER_37_508 ();
 sg13g2_decap_8 FILLER_37_515 ();
 sg13g2_decap_8 FILLER_37_522 ();
 sg13g2_decap_8 FILLER_37_529 ();
 sg13g2_decap_8 FILLER_37_536 ();
 sg13g2_decap_8 FILLER_37_543 ();
 sg13g2_decap_8 FILLER_37_550 ();
 sg13g2_decap_8 FILLER_37_557 ();
 sg13g2_decap_8 FILLER_37_564 ();
 sg13g2_decap_8 FILLER_37_571 ();
 sg13g2_decap_8 FILLER_37_578 ();
 sg13g2_decap_8 FILLER_37_585 ();
 sg13g2_decap_8 FILLER_37_592 ();
 sg13g2_decap_8 FILLER_37_599 ();
 sg13g2_decap_8 FILLER_37_606 ();
 sg13g2_decap_8 FILLER_37_613 ();
 sg13g2_decap_8 FILLER_37_620 ();
 sg13g2_decap_8 FILLER_37_627 ();
 sg13g2_decap_8 FILLER_37_634 ();
 sg13g2_decap_8 FILLER_37_641 ();
 sg13g2_decap_8 FILLER_37_648 ();
 sg13g2_decap_8 FILLER_37_655 ();
 sg13g2_decap_8 FILLER_37_662 ();
 sg13g2_decap_8 FILLER_37_669 ();
 sg13g2_decap_8 FILLER_37_676 ();
 sg13g2_decap_8 FILLER_37_683 ();
 sg13g2_decap_8 FILLER_37_690 ();
 sg13g2_decap_8 FILLER_37_697 ();
 sg13g2_decap_8 FILLER_37_704 ();
 sg13g2_decap_8 FILLER_37_711 ();
 sg13g2_decap_8 FILLER_37_718 ();
 sg13g2_decap_8 FILLER_37_725 ();
 sg13g2_decap_8 FILLER_37_732 ();
 sg13g2_decap_8 FILLER_37_739 ();
 sg13g2_decap_8 FILLER_37_746 ();
 sg13g2_decap_8 FILLER_37_753 ();
 sg13g2_decap_8 FILLER_37_760 ();
 sg13g2_decap_8 FILLER_37_767 ();
 sg13g2_decap_8 FILLER_37_774 ();
 sg13g2_decap_8 FILLER_37_781 ();
 sg13g2_decap_8 FILLER_37_788 ();
 sg13g2_decap_8 FILLER_37_795 ();
 sg13g2_decap_8 FILLER_37_802 ();
 sg13g2_decap_8 FILLER_37_809 ();
 sg13g2_decap_8 FILLER_37_816 ();
 sg13g2_decap_8 FILLER_37_823 ();
 sg13g2_decap_8 FILLER_37_830 ();
 sg13g2_decap_8 FILLER_37_837 ();
 sg13g2_decap_8 FILLER_37_844 ();
 sg13g2_decap_8 FILLER_37_851 ();
 sg13g2_decap_8 FILLER_37_858 ();
 sg13g2_decap_8 FILLER_37_865 ();
 sg13g2_decap_8 FILLER_37_872 ();
 sg13g2_decap_8 FILLER_37_879 ();
 sg13g2_decap_8 FILLER_37_886 ();
 sg13g2_decap_8 FILLER_37_893 ();
 sg13g2_decap_8 FILLER_37_900 ();
 sg13g2_decap_8 FILLER_37_907 ();
 sg13g2_decap_8 FILLER_37_914 ();
 sg13g2_decap_8 FILLER_37_921 ();
 sg13g2_decap_8 FILLER_37_928 ();
 sg13g2_decap_8 FILLER_37_935 ();
 sg13g2_decap_8 FILLER_37_942 ();
 sg13g2_decap_8 FILLER_37_949 ();
 sg13g2_decap_8 FILLER_37_956 ();
 sg13g2_decap_8 FILLER_37_963 ();
 sg13g2_decap_8 FILLER_37_970 ();
 sg13g2_decap_8 FILLER_37_977 ();
 sg13g2_decap_8 FILLER_37_984 ();
 sg13g2_decap_8 FILLER_37_991 ();
 sg13g2_decap_8 FILLER_37_998 ();
 sg13g2_decap_8 FILLER_37_1005 ();
 sg13g2_decap_8 FILLER_37_1012 ();
 sg13g2_decap_8 FILLER_37_1019 ();
 sg13g2_fill_2 FILLER_37_1026 ();
 sg13g2_fill_1 FILLER_37_1028 ();
 sg13g2_decap_8 FILLER_38_0 ();
 sg13g2_decap_8 FILLER_38_7 ();
 sg13g2_decap_8 FILLER_38_14 ();
 sg13g2_decap_8 FILLER_38_21 ();
 sg13g2_decap_8 FILLER_38_28 ();
 sg13g2_decap_8 FILLER_38_35 ();
 sg13g2_decap_8 FILLER_38_42 ();
 sg13g2_decap_8 FILLER_38_49 ();
 sg13g2_decap_8 FILLER_38_56 ();
 sg13g2_decap_8 FILLER_38_63 ();
 sg13g2_decap_8 FILLER_38_70 ();
 sg13g2_decap_8 FILLER_38_77 ();
 sg13g2_decap_8 FILLER_38_84 ();
 sg13g2_decap_8 FILLER_38_91 ();
 sg13g2_decap_8 FILLER_38_98 ();
 sg13g2_decap_8 FILLER_38_105 ();
 sg13g2_decap_8 FILLER_38_112 ();
 sg13g2_decap_8 FILLER_38_119 ();
 sg13g2_decap_8 FILLER_38_126 ();
 sg13g2_decap_8 FILLER_38_133 ();
 sg13g2_decap_8 FILLER_38_140 ();
 sg13g2_decap_8 FILLER_38_147 ();
 sg13g2_decap_8 FILLER_38_154 ();
 sg13g2_decap_8 FILLER_38_161 ();
 sg13g2_decap_8 FILLER_38_168 ();
 sg13g2_decap_8 FILLER_38_175 ();
 sg13g2_decap_8 FILLER_38_182 ();
 sg13g2_decap_8 FILLER_38_189 ();
 sg13g2_decap_8 FILLER_38_196 ();
 sg13g2_decap_8 FILLER_38_203 ();
 sg13g2_decap_8 FILLER_38_210 ();
 sg13g2_decap_8 FILLER_38_217 ();
 sg13g2_decap_8 FILLER_38_224 ();
 sg13g2_decap_8 FILLER_38_231 ();
 sg13g2_decap_8 FILLER_38_238 ();
 sg13g2_decap_8 FILLER_38_245 ();
 sg13g2_decap_8 FILLER_38_252 ();
 sg13g2_decap_8 FILLER_38_259 ();
 sg13g2_decap_8 FILLER_38_266 ();
 sg13g2_decap_8 FILLER_38_273 ();
 sg13g2_decap_8 FILLER_38_280 ();
 sg13g2_decap_8 FILLER_38_287 ();
 sg13g2_decap_8 FILLER_38_294 ();
 sg13g2_decap_8 FILLER_38_301 ();
 sg13g2_decap_8 FILLER_38_308 ();
 sg13g2_decap_8 FILLER_38_315 ();
 sg13g2_decap_8 FILLER_38_322 ();
 sg13g2_decap_8 FILLER_38_329 ();
 sg13g2_decap_8 FILLER_38_336 ();
 sg13g2_decap_8 FILLER_38_343 ();
 sg13g2_decap_8 FILLER_38_350 ();
 sg13g2_decap_8 FILLER_38_357 ();
 sg13g2_decap_8 FILLER_38_364 ();
 sg13g2_decap_8 FILLER_38_371 ();
 sg13g2_decap_8 FILLER_38_378 ();
 sg13g2_decap_8 FILLER_38_385 ();
 sg13g2_decap_8 FILLER_38_392 ();
 sg13g2_decap_8 FILLER_38_399 ();
 sg13g2_decap_8 FILLER_38_406 ();
 sg13g2_decap_8 FILLER_38_413 ();
 sg13g2_decap_8 FILLER_38_420 ();
 sg13g2_decap_8 FILLER_38_427 ();
 sg13g2_decap_8 FILLER_38_434 ();
 sg13g2_decap_8 FILLER_38_441 ();
 sg13g2_decap_8 FILLER_38_448 ();
 sg13g2_decap_8 FILLER_38_455 ();
 sg13g2_decap_8 FILLER_38_462 ();
 sg13g2_decap_8 FILLER_38_469 ();
 sg13g2_decap_8 FILLER_38_476 ();
 sg13g2_decap_8 FILLER_38_483 ();
 sg13g2_decap_8 FILLER_38_490 ();
 sg13g2_decap_8 FILLER_38_497 ();
 sg13g2_decap_8 FILLER_38_504 ();
 sg13g2_decap_8 FILLER_38_511 ();
 sg13g2_decap_8 FILLER_38_518 ();
 sg13g2_decap_8 FILLER_38_525 ();
 sg13g2_decap_8 FILLER_38_532 ();
 sg13g2_decap_8 FILLER_38_539 ();
 sg13g2_decap_8 FILLER_38_546 ();
 sg13g2_decap_8 FILLER_38_553 ();
 sg13g2_decap_8 FILLER_38_560 ();
 sg13g2_decap_8 FILLER_38_567 ();
 sg13g2_decap_8 FILLER_38_574 ();
 sg13g2_decap_8 FILLER_38_581 ();
 sg13g2_decap_8 FILLER_38_588 ();
 sg13g2_decap_8 FILLER_38_595 ();
 sg13g2_decap_8 FILLER_38_602 ();
 sg13g2_decap_8 FILLER_38_609 ();
 sg13g2_decap_8 FILLER_38_616 ();
 sg13g2_decap_8 FILLER_38_623 ();
 sg13g2_decap_8 FILLER_38_630 ();
 sg13g2_decap_8 FILLER_38_637 ();
 sg13g2_decap_8 FILLER_38_644 ();
 sg13g2_decap_8 FILLER_38_651 ();
 sg13g2_decap_8 FILLER_38_658 ();
 sg13g2_decap_8 FILLER_38_665 ();
 sg13g2_decap_8 FILLER_38_672 ();
 sg13g2_decap_8 FILLER_38_679 ();
 sg13g2_decap_8 FILLER_38_686 ();
 sg13g2_decap_8 FILLER_38_693 ();
 sg13g2_decap_8 FILLER_38_700 ();
 sg13g2_decap_8 FILLER_38_707 ();
 sg13g2_decap_8 FILLER_38_714 ();
 sg13g2_decap_8 FILLER_38_721 ();
 sg13g2_decap_8 FILLER_38_728 ();
 sg13g2_decap_8 FILLER_38_735 ();
 sg13g2_decap_8 FILLER_38_742 ();
 sg13g2_decap_8 FILLER_38_749 ();
 sg13g2_decap_8 FILLER_38_756 ();
 sg13g2_decap_8 FILLER_38_763 ();
 sg13g2_decap_8 FILLER_38_770 ();
 sg13g2_decap_8 FILLER_38_777 ();
 sg13g2_decap_8 FILLER_38_784 ();
 sg13g2_decap_8 FILLER_38_791 ();
 sg13g2_decap_8 FILLER_38_798 ();
 sg13g2_decap_8 FILLER_38_805 ();
 sg13g2_decap_8 FILLER_38_812 ();
 sg13g2_decap_8 FILLER_38_819 ();
 sg13g2_decap_8 FILLER_38_826 ();
 sg13g2_decap_8 FILLER_38_833 ();
 sg13g2_decap_8 FILLER_38_840 ();
 sg13g2_decap_8 FILLER_38_847 ();
 sg13g2_decap_8 FILLER_38_854 ();
 sg13g2_decap_8 FILLER_38_861 ();
 sg13g2_decap_8 FILLER_38_868 ();
 sg13g2_decap_8 FILLER_38_875 ();
 sg13g2_decap_8 FILLER_38_882 ();
 sg13g2_decap_8 FILLER_38_889 ();
 sg13g2_decap_8 FILLER_38_896 ();
 sg13g2_decap_8 FILLER_38_903 ();
 sg13g2_decap_8 FILLER_38_910 ();
 sg13g2_decap_8 FILLER_38_917 ();
 sg13g2_decap_8 FILLER_38_924 ();
 sg13g2_decap_8 FILLER_38_931 ();
 sg13g2_decap_8 FILLER_38_938 ();
 sg13g2_decap_8 FILLER_38_945 ();
 sg13g2_decap_8 FILLER_38_952 ();
 sg13g2_decap_8 FILLER_38_959 ();
 sg13g2_decap_8 FILLER_38_966 ();
 sg13g2_decap_8 FILLER_38_973 ();
 sg13g2_decap_8 FILLER_38_980 ();
 sg13g2_decap_8 FILLER_38_987 ();
 sg13g2_decap_8 FILLER_38_994 ();
 sg13g2_decap_8 FILLER_38_1001 ();
 sg13g2_decap_8 FILLER_38_1008 ();
 sg13g2_decap_8 FILLER_38_1015 ();
 sg13g2_decap_8 FILLER_38_1022 ();
 sg13g2_decap_8 FILLER_39_4 ();
 sg13g2_decap_8 FILLER_39_11 ();
 sg13g2_decap_8 FILLER_39_18 ();
 sg13g2_decap_8 FILLER_39_25 ();
 sg13g2_decap_8 FILLER_39_32 ();
 sg13g2_decap_8 FILLER_39_39 ();
 sg13g2_decap_8 FILLER_39_46 ();
 sg13g2_decap_8 FILLER_39_53 ();
 sg13g2_decap_8 FILLER_39_60 ();
 sg13g2_decap_8 FILLER_39_67 ();
 sg13g2_decap_8 FILLER_39_74 ();
 sg13g2_decap_8 FILLER_39_81 ();
 sg13g2_decap_8 FILLER_39_88 ();
 sg13g2_decap_8 FILLER_39_95 ();
 sg13g2_decap_8 FILLER_39_102 ();
 sg13g2_decap_8 FILLER_39_109 ();
 sg13g2_decap_8 FILLER_39_116 ();
 sg13g2_decap_8 FILLER_39_123 ();
 sg13g2_decap_8 FILLER_39_130 ();
 sg13g2_decap_8 FILLER_39_137 ();
 sg13g2_decap_8 FILLER_39_144 ();
 sg13g2_decap_8 FILLER_39_151 ();
 sg13g2_decap_8 FILLER_39_158 ();
 sg13g2_decap_8 FILLER_39_165 ();
 sg13g2_decap_8 FILLER_39_172 ();
 sg13g2_decap_8 FILLER_39_179 ();
 sg13g2_decap_8 FILLER_39_186 ();
 sg13g2_decap_8 FILLER_39_193 ();
 sg13g2_decap_8 FILLER_39_200 ();
 sg13g2_decap_8 FILLER_39_207 ();
 sg13g2_decap_8 FILLER_39_214 ();
 sg13g2_decap_8 FILLER_39_221 ();
 sg13g2_decap_8 FILLER_39_228 ();
 sg13g2_decap_8 FILLER_39_235 ();
 sg13g2_decap_8 FILLER_39_242 ();
 sg13g2_decap_8 FILLER_39_249 ();
 sg13g2_decap_8 FILLER_39_256 ();
 sg13g2_decap_8 FILLER_39_263 ();
 sg13g2_decap_8 FILLER_39_270 ();
 sg13g2_decap_8 FILLER_39_277 ();
 sg13g2_decap_8 FILLER_39_284 ();
 sg13g2_decap_8 FILLER_39_291 ();
 sg13g2_decap_8 FILLER_39_298 ();
 sg13g2_decap_8 FILLER_39_305 ();
 sg13g2_decap_8 FILLER_39_312 ();
 sg13g2_decap_8 FILLER_39_319 ();
 sg13g2_decap_8 FILLER_39_326 ();
 sg13g2_decap_8 FILLER_39_333 ();
 sg13g2_decap_8 FILLER_39_340 ();
 sg13g2_decap_8 FILLER_39_347 ();
 sg13g2_decap_8 FILLER_39_354 ();
 sg13g2_decap_8 FILLER_39_361 ();
 sg13g2_decap_8 FILLER_39_368 ();
 sg13g2_decap_8 FILLER_39_375 ();
 sg13g2_decap_8 FILLER_39_382 ();
 sg13g2_decap_8 FILLER_39_389 ();
 sg13g2_decap_8 FILLER_39_396 ();
 sg13g2_decap_8 FILLER_39_403 ();
 sg13g2_decap_8 FILLER_39_410 ();
 sg13g2_decap_8 FILLER_39_417 ();
 sg13g2_decap_8 FILLER_39_424 ();
 sg13g2_decap_8 FILLER_39_431 ();
 sg13g2_decap_8 FILLER_39_438 ();
 sg13g2_decap_8 FILLER_39_445 ();
 sg13g2_decap_8 FILLER_39_452 ();
 sg13g2_decap_8 FILLER_39_459 ();
 sg13g2_decap_8 FILLER_39_466 ();
 sg13g2_decap_8 FILLER_39_473 ();
 sg13g2_decap_8 FILLER_39_480 ();
 sg13g2_decap_8 FILLER_39_487 ();
 sg13g2_decap_8 FILLER_39_494 ();
 sg13g2_decap_8 FILLER_39_501 ();
 sg13g2_decap_8 FILLER_39_508 ();
 sg13g2_decap_8 FILLER_39_515 ();
 sg13g2_decap_8 FILLER_39_522 ();
 sg13g2_decap_8 FILLER_39_529 ();
 sg13g2_decap_8 FILLER_39_536 ();
 sg13g2_decap_8 FILLER_39_543 ();
 sg13g2_decap_8 FILLER_39_550 ();
 sg13g2_decap_8 FILLER_39_557 ();
 sg13g2_decap_8 FILLER_39_564 ();
 sg13g2_decap_8 FILLER_39_571 ();
 sg13g2_decap_8 FILLER_39_578 ();
 sg13g2_decap_8 FILLER_39_585 ();
 sg13g2_decap_8 FILLER_39_592 ();
 sg13g2_decap_8 FILLER_39_599 ();
 sg13g2_decap_8 FILLER_39_606 ();
 sg13g2_decap_8 FILLER_39_613 ();
 sg13g2_decap_8 FILLER_39_620 ();
 sg13g2_decap_8 FILLER_39_627 ();
 sg13g2_decap_8 FILLER_39_634 ();
 sg13g2_decap_8 FILLER_39_641 ();
 sg13g2_decap_8 FILLER_39_648 ();
 sg13g2_decap_8 FILLER_39_655 ();
 sg13g2_decap_8 FILLER_39_662 ();
 sg13g2_decap_8 FILLER_39_669 ();
 sg13g2_decap_8 FILLER_39_676 ();
 sg13g2_decap_8 FILLER_39_683 ();
 sg13g2_decap_8 FILLER_39_690 ();
 sg13g2_decap_8 FILLER_39_697 ();
 sg13g2_decap_8 FILLER_39_704 ();
 sg13g2_decap_8 FILLER_39_711 ();
 sg13g2_decap_8 FILLER_39_718 ();
 sg13g2_decap_8 FILLER_39_725 ();
 sg13g2_decap_8 FILLER_39_732 ();
 sg13g2_decap_8 FILLER_39_739 ();
 sg13g2_decap_8 FILLER_39_746 ();
 sg13g2_decap_8 FILLER_39_753 ();
 sg13g2_decap_8 FILLER_39_760 ();
 sg13g2_decap_8 FILLER_39_767 ();
 sg13g2_decap_8 FILLER_39_774 ();
 sg13g2_decap_8 FILLER_39_781 ();
 sg13g2_decap_8 FILLER_39_788 ();
 sg13g2_decap_8 FILLER_39_795 ();
 sg13g2_decap_8 FILLER_39_802 ();
 sg13g2_decap_8 FILLER_39_809 ();
 sg13g2_decap_8 FILLER_39_816 ();
 sg13g2_decap_8 FILLER_39_823 ();
 sg13g2_decap_8 FILLER_39_830 ();
 sg13g2_decap_8 FILLER_39_837 ();
 sg13g2_decap_8 FILLER_39_844 ();
 sg13g2_decap_8 FILLER_39_851 ();
 sg13g2_decap_8 FILLER_39_858 ();
 sg13g2_decap_8 FILLER_39_865 ();
 sg13g2_decap_8 FILLER_39_872 ();
 sg13g2_decap_8 FILLER_39_879 ();
 sg13g2_decap_8 FILLER_39_886 ();
 sg13g2_decap_8 FILLER_39_893 ();
 sg13g2_decap_8 FILLER_39_900 ();
 sg13g2_decap_8 FILLER_39_907 ();
 sg13g2_decap_8 FILLER_39_914 ();
 sg13g2_decap_8 FILLER_39_921 ();
 sg13g2_decap_8 FILLER_39_928 ();
 sg13g2_decap_8 FILLER_39_935 ();
 sg13g2_decap_8 FILLER_39_942 ();
 sg13g2_decap_8 FILLER_39_949 ();
 sg13g2_decap_8 FILLER_39_956 ();
 sg13g2_decap_8 FILLER_39_963 ();
 sg13g2_decap_8 FILLER_39_970 ();
 sg13g2_decap_8 FILLER_39_977 ();
 sg13g2_decap_8 FILLER_39_984 ();
 sg13g2_decap_8 FILLER_39_991 ();
 sg13g2_decap_8 FILLER_39_998 ();
 sg13g2_decap_8 FILLER_39_1005 ();
 sg13g2_decap_8 FILLER_39_1012 ();
 sg13g2_decap_8 FILLER_39_1019 ();
 sg13g2_fill_2 FILLER_39_1026 ();
 sg13g2_fill_1 FILLER_39_1028 ();
 sg13g2_decap_8 FILLER_40_0 ();
 sg13g2_decap_8 FILLER_40_7 ();
 sg13g2_decap_8 FILLER_40_14 ();
 sg13g2_decap_8 FILLER_40_21 ();
 sg13g2_decap_8 FILLER_40_28 ();
 sg13g2_decap_8 FILLER_40_35 ();
 sg13g2_decap_8 FILLER_40_42 ();
 sg13g2_decap_8 FILLER_40_49 ();
 sg13g2_decap_8 FILLER_40_56 ();
 sg13g2_decap_8 FILLER_40_63 ();
 sg13g2_decap_8 FILLER_40_70 ();
 sg13g2_decap_8 FILLER_40_77 ();
 sg13g2_decap_8 FILLER_40_84 ();
 sg13g2_decap_8 FILLER_40_91 ();
 sg13g2_decap_8 FILLER_40_98 ();
 sg13g2_decap_8 FILLER_40_105 ();
 sg13g2_decap_8 FILLER_40_112 ();
 sg13g2_decap_8 FILLER_40_119 ();
 sg13g2_decap_8 FILLER_40_126 ();
 sg13g2_decap_8 FILLER_40_133 ();
 sg13g2_decap_8 FILLER_40_140 ();
 sg13g2_decap_8 FILLER_40_147 ();
 sg13g2_decap_8 FILLER_40_154 ();
 sg13g2_decap_8 FILLER_40_161 ();
 sg13g2_decap_8 FILLER_40_168 ();
 sg13g2_decap_8 FILLER_40_175 ();
 sg13g2_decap_8 FILLER_40_182 ();
 sg13g2_decap_8 FILLER_40_189 ();
 sg13g2_decap_8 FILLER_40_196 ();
 sg13g2_decap_8 FILLER_40_203 ();
 sg13g2_decap_8 FILLER_40_210 ();
 sg13g2_decap_8 FILLER_40_217 ();
 sg13g2_decap_8 FILLER_40_224 ();
 sg13g2_decap_8 FILLER_40_231 ();
 sg13g2_decap_8 FILLER_40_238 ();
 sg13g2_decap_8 FILLER_40_245 ();
 sg13g2_decap_8 FILLER_40_252 ();
 sg13g2_decap_8 FILLER_40_259 ();
 sg13g2_decap_8 FILLER_40_266 ();
 sg13g2_decap_8 FILLER_40_273 ();
 sg13g2_decap_8 FILLER_40_280 ();
 sg13g2_decap_8 FILLER_40_287 ();
 sg13g2_decap_8 FILLER_40_294 ();
 sg13g2_decap_8 FILLER_40_301 ();
 sg13g2_decap_8 FILLER_40_308 ();
 sg13g2_decap_8 FILLER_40_315 ();
 sg13g2_decap_8 FILLER_40_322 ();
 sg13g2_decap_8 FILLER_40_329 ();
 sg13g2_decap_8 FILLER_40_336 ();
 sg13g2_decap_8 FILLER_40_343 ();
 sg13g2_decap_8 FILLER_40_350 ();
 sg13g2_decap_8 FILLER_40_357 ();
 sg13g2_decap_8 FILLER_40_364 ();
 sg13g2_decap_8 FILLER_40_371 ();
 sg13g2_decap_8 FILLER_40_378 ();
 sg13g2_decap_8 FILLER_40_385 ();
 sg13g2_decap_8 FILLER_40_392 ();
 sg13g2_decap_8 FILLER_40_399 ();
 sg13g2_decap_8 FILLER_40_406 ();
 sg13g2_decap_8 FILLER_40_413 ();
 sg13g2_decap_8 FILLER_40_420 ();
 sg13g2_decap_8 FILLER_40_427 ();
 sg13g2_decap_8 FILLER_40_434 ();
 sg13g2_decap_8 FILLER_40_441 ();
 sg13g2_decap_8 FILLER_40_448 ();
 sg13g2_decap_8 FILLER_40_455 ();
 sg13g2_decap_8 FILLER_40_462 ();
 sg13g2_decap_8 FILLER_40_469 ();
 sg13g2_decap_8 FILLER_40_476 ();
 sg13g2_decap_8 FILLER_40_483 ();
 sg13g2_decap_8 FILLER_40_490 ();
 sg13g2_decap_8 FILLER_40_497 ();
 sg13g2_decap_8 FILLER_40_504 ();
 sg13g2_decap_8 FILLER_40_511 ();
 sg13g2_decap_8 FILLER_40_518 ();
 sg13g2_decap_8 FILLER_40_525 ();
 sg13g2_decap_8 FILLER_40_532 ();
 sg13g2_decap_8 FILLER_40_539 ();
 sg13g2_decap_8 FILLER_40_546 ();
 sg13g2_decap_8 FILLER_40_553 ();
 sg13g2_decap_8 FILLER_40_560 ();
 sg13g2_decap_8 FILLER_40_567 ();
 sg13g2_decap_8 FILLER_40_574 ();
 sg13g2_decap_8 FILLER_40_581 ();
 sg13g2_decap_8 FILLER_40_588 ();
 sg13g2_decap_8 FILLER_40_595 ();
 sg13g2_decap_8 FILLER_40_602 ();
 sg13g2_decap_8 FILLER_40_609 ();
 sg13g2_decap_8 FILLER_40_616 ();
 sg13g2_decap_8 FILLER_40_623 ();
 sg13g2_decap_8 FILLER_40_630 ();
 sg13g2_decap_8 FILLER_40_637 ();
 sg13g2_decap_8 FILLER_40_644 ();
 sg13g2_decap_8 FILLER_40_651 ();
 sg13g2_decap_8 FILLER_40_658 ();
 sg13g2_decap_8 FILLER_40_665 ();
 sg13g2_decap_8 FILLER_40_672 ();
 sg13g2_decap_8 FILLER_40_679 ();
 sg13g2_decap_8 FILLER_40_686 ();
 sg13g2_decap_8 FILLER_40_693 ();
 sg13g2_decap_8 FILLER_40_700 ();
 sg13g2_decap_8 FILLER_40_707 ();
 sg13g2_decap_8 FILLER_40_714 ();
 sg13g2_decap_8 FILLER_40_721 ();
 sg13g2_decap_8 FILLER_40_728 ();
 sg13g2_decap_8 FILLER_40_735 ();
 sg13g2_decap_8 FILLER_40_742 ();
 sg13g2_decap_8 FILLER_40_749 ();
 sg13g2_decap_8 FILLER_40_756 ();
 sg13g2_decap_8 FILLER_40_763 ();
 sg13g2_decap_8 FILLER_40_770 ();
 sg13g2_decap_8 FILLER_40_777 ();
 sg13g2_decap_8 FILLER_40_784 ();
 sg13g2_decap_8 FILLER_40_791 ();
 sg13g2_decap_8 FILLER_40_798 ();
 sg13g2_decap_8 FILLER_40_805 ();
 sg13g2_decap_8 FILLER_40_812 ();
 sg13g2_decap_8 FILLER_40_819 ();
 sg13g2_decap_8 FILLER_40_826 ();
 sg13g2_decap_8 FILLER_40_833 ();
 sg13g2_decap_8 FILLER_40_840 ();
 sg13g2_decap_8 FILLER_40_847 ();
 sg13g2_decap_8 FILLER_40_854 ();
 sg13g2_decap_8 FILLER_40_861 ();
 sg13g2_decap_8 FILLER_40_868 ();
 sg13g2_decap_8 FILLER_40_875 ();
 sg13g2_decap_8 FILLER_40_882 ();
 sg13g2_decap_8 FILLER_40_889 ();
 sg13g2_decap_8 FILLER_40_896 ();
 sg13g2_decap_8 FILLER_40_903 ();
 sg13g2_decap_8 FILLER_40_910 ();
 sg13g2_decap_8 FILLER_40_917 ();
 sg13g2_decap_8 FILLER_40_924 ();
 sg13g2_decap_8 FILLER_40_931 ();
 sg13g2_decap_8 FILLER_40_938 ();
 sg13g2_decap_8 FILLER_40_945 ();
 sg13g2_decap_8 FILLER_40_952 ();
 sg13g2_decap_8 FILLER_40_959 ();
 sg13g2_decap_8 FILLER_40_966 ();
 sg13g2_decap_8 FILLER_40_973 ();
 sg13g2_decap_8 FILLER_40_980 ();
 sg13g2_decap_8 FILLER_40_987 ();
 sg13g2_decap_8 FILLER_40_994 ();
 sg13g2_decap_8 FILLER_40_1001 ();
 sg13g2_decap_8 FILLER_40_1008 ();
 sg13g2_decap_8 FILLER_40_1015 ();
 sg13g2_decap_8 FILLER_40_1022 ();
 sg13g2_decap_8 FILLER_41_0 ();
 sg13g2_decap_8 FILLER_41_7 ();
 sg13g2_decap_8 FILLER_41_14 ();
 sg13g2_decap_8 FILLER_41_21 ();
 sg13g2_decap_8 FILLER_41_28 ();
 sg13g2_decap_8 FILLER_41_35 ();
 sg13g2_decap_8 FILLER_41_42 ();
 sg13g2_decap_8 FILLER_41_49 ();
 sg13g2_decap_8 FILLER_41_56 ();
 sg13g2_decap_8 FILLER_41_63 ();
 sg13g2_decap_8 FILLER_41_70 ();
 sg13g2_decap_8 FILLER_41_77 ();
 sg13g2_decap_8 FILLER_41_84 ();
 sg13g2_decap_8 FILLER_41_91 ();
 sg13g2_decap_8 FILLER_41_98 ();
 sg13g2_decap_8 FILLER_41_105 ();
 sg13g2_decap_8 FILLER_41_112 ();
 sg13g2_decap_8 FILLER_41_119 ();
 sg13g2_decap_8 FILLER_41_126 ();
 sg13g2_decap_8 FILLER_41_133 ();
 sg13g2_decap_8 FILLER_41_140 ();
 sg13g2_decap_8 FILLER_41_147 ();
 sg13g2_decap_8 FILLER_41_154 ();
 sg13g2_decap_8 FILLER_41_161 ();
 sg13g2_decap_8 FILLER_41_168 ();
 sg13g2_decap_8 FILLER_41_175 ();
 sg13g2_decap_8 FILLER_41_182 ();
 sg13g2_decap_8 FILLER_41_189 ();
 sg13g2_decap_8 FILLER_41_196 ();
 sg13g2_decap_8 FILLER_41_203 ();
 sg13g2_decap_8 FILLER_41_210 ();
 sg13g2_decap_8 FILLER_41_217 ();
 sg13g2_decap_8 FILLER_41_224 ();
 sg13g2_decap_8 FILLER_41_231 ();
 sg13g2_decap_8 FILLER_41_238 ();
 sg13g2_decap_8 FILLER_41_245 ();
 sg13g2_decap_8 FILLER_41_252 ();
 sg13g2_decap_8 FILLER_41_259 ();
 sg13g2_decap_8 FILLER_41_266 ();
 sg13g2_decap_8 FILLER_41_273 ();
 sg13g2_decap_8 FILLER_41_280 ();
 sg13g2_decap_8 FILLER_41_287 ();
 sg13g2_decap_8 FILLER_41_294 ();
 sg13g2_decap_8 FILLER_41_301 ();
 sg13g2_decap_8 FILLER_41_308 ();
 sg13g2_decap_8 FILLER_41_315 ();
 sg13g2_decap_8 FILLER_41_322 ();
 sg13g2_decap_8 FILLER_41_329 ();
 sg13g2_decap_8 FILLER_41_336 ();
 sg13g2_decap_8 FILLER_41_343 ();
 sg13g2_decap_8 FILLER_41_350 ();
 sg13g2_decap_8 FILLER_41_357 ();
 sg13g2_decap_8 FILLER_41_364 ();
 sg13g2_decap_8 FILLER_41_371 ();
 sg13g2_decap_8 FILLER_41_378 ();
 sg13g2_decap_8 FILLER_41_385 ();
 sg13g2_decap_8 FILLER_41_392 ();
 sg13g2_decap_8 FILLER_41_399 ();
 sg13g2_decap_8 FILLER_41_406 ();
 sg13g2_decap_8 FILLER_41_413 ();
 sg13g2_decap_8 FILLER_41_420 ();
 sg13g2_decap_8 FILLER_41_427 ();
 sg13g2_decap_8 FILLER_41_434 ();
 sg13g2_decap_8 FILLER_41_441 ();
 sg13g2_decap_8 FILLER_41_448 ();
 sg13g2_decap_8 FILLER_41_455 ();
 sg13g2_decap_8 FILLER_41_462 ();
 sg13g2_decap_8 FILLER_41_469 ();
 sg13g2_decap_8 FILLER_41_476 ();
 sg13g2_decap_8 FILLER_41_483 ();
 sg13g2_decap_8 FILLER_41_490 ();
 sg13g2_decap_8 FILLER_41_497 ();
 sg13g2_decap_8 FILLER_41_504 ();
 sg13g2_decap_8 FILLER_41_511 ();
 sg13g2_decap_8 FILLER_41_518 ();
 sg13g2_decap_8 FILLER_41_525 ();
 sg13g2_decap_8 FILLER_41_532 ();
 sg13g2_decap_8 FILLER_41_539 ();
 sg13g2_decap_8 FILLER_41_546 ();
 sg13g2_decap_8 FILLER_41_553 ();
 sg13g2_decap_8 FILLER_41_560 ();
 sg13g2_decap_8 FILLER_41_567 ();
 sg13g2_decap_8 FILLER_41_574 ();
 sg13g2_decap_8 FILLER_41_581 ();
 sg13g2_decap_8 FILLER_41_588 ();
 sg13g2_decap_8 FILLER_41_595 ();
 sg13g2_decap_8 FILLER_41_602 ();
 sg13g2_decap_8 FILLER_41_609 ();
 sg13g2_decap_8 FILLER_41_616 ();
 sg13g2_decap_8 FILLER_41_623 ();
 sg13g2_decap_8 FILLER_41_630 ();
 sg13g2_decap_8 FILLER_41_637 ();
 sg13g2_decap_8 FILLER_41_644 ();
 sg13g2_decap_8 FILLER_41_651 ();
 sg13g2_decap_8 FILLER_41_658 ();
 sg13g2_decap_8 FILLER_41_665 ();
 sg13g2_decap_8 FILLER_41_672 ();
 sg13g2_decap_8 FILLER_41_679 ();
 sg13g2_decap_8 FILLER_41_686 ();
 sg13g2_decap_8 FILLER_41_693 ();
 sg13g2_decap_8 FILLER_41_700 ();
 sg13g2_decap_8 FILLER_41_707 ();
 sg13g2_decap_8 FILLER_41_714 ();
 sg13g2_decap_8 FILLER_41_721 ();
 sg13g2_decap_8 FILLER_41_728 ();
 sg13g2_decap_8 FILLER_41_735 ();
 sg13g2_decap_8 FILLER_41_742 ();
 sg13g2_decap_8 FILLER_41_749 ();
 sg13g2_decap_8 FILLER_41_756 ();
 sg13g2_decap_8 FILLER_41_763 ();
 sg13g2_decap_8 FILLER_41_770 ();
 sg13g2_decap_8 FILLER_41_777 ();
 sg13g2_decap_8 FILLER_41_784 ();
 sg13g2_decap_8 FILLER_41_791 ();
 sg13g2_decap_8 FILLER_41_798 ();
 sg13g2_decap_8 FILLER_41_805 ();
 sg13g2_decap_8 FILLER_41_812 ();
 sg13g2_decap_8 FILLER_41_819 ();
 sg13g2_decap_8 FILLER_41_826 ();
 sg13g2_decap_8 FILLER_41_833 ();
 sg13g2_decap_8 FILLER_41_840 ();
 sg13g2_decap_8 FILLER_41_847 ();
 sg13g2_decap_8 FILLER_41_854 ();
 sg13g2_decap_8 FILLER_41_861 ();
 sg13g2_decap_8 FILLER_41_868 ();
 sg13g2_decap_8 FILLER_41_875 ();
 sg13g2_decap_8 FILLER_41_882 ();
 sg13g2_decap_8 FILLER_41_889 ();
 sg13g2_decap_8 FILLER_41_896 ();
 sg13g2_decap_8 FILLER_41_903 ();
 sg13g2_decap_8 FILLER_41_910 ();
 sg13g2_decap_8 FILLER_41_917 ();
 sg13g2_decap_8 FILLER_41_924 ();
 sg13g2_decap_8 FILLER_41_931 ();
 sg13g2_decap_8 FILLER_41_938 ();
 sg13g2_decap_8 FILLER_41_945 ();
 sg13g2_decap_8 FILLER_41_952 ();
 sg13g2_decap_8 FILLER_41_959 ();
 sg13g2_decap_8 FILLER_41_966 ();
 sg13g2_decap_8 FILLER_41_973 ();
 sg13g2_decap_8 FILLER_41_980 ();
 sg13g2_decap_8 FILLER_41_987 ();
 sg13g2_decap_8 FILLER_41_994 ();
 sg13g2_decap_8 FILLER_41_1001 ();
 sg13g2_decap_8 FILLER_41_1008 ();
 sg13g2_decap_8 FILLER_41_1015 ();
 sg13g2_decap_8 FILLER_41_1022 ();
 sg13g2_decap_8 FILLER_42_4 ();
 sg13g2_decap_8 FILLER_42_11 ();
 sg13g2_decap_8 FILLER_42_18 ();
 sg13g2_decap_8 FILLER_42_25 ();
 sg13g2_decap_8 FILLER_42_32 ();
 sg13g2_decap_8 FILLER_42_39 ();
 sg13g2_decap_8 FILLER_42_46 ();
 sg13g2_decap_8 FILLER_42_53 ();
 sg13g2_decap_8 FILLER_42_60 ();
 sg13g2_decap_8 FILLER_42_67 ();
 sg13g2_decap_8 FILLER_42_74 ();
 sg13g2_decap_8 FILLER_42_81 ();
 sg13g2_decap_8 FILLER_42_88 ();
 sg13g2_decap_8 FILLER_42_95 ();
 sg13g2_decap_8 FILLER_42_102 ();
 sg13g2_decap_8 FILLER_42_109 ();
 sg13g2_decap_8 FILLER_42_116 ();
 sg13g2_decap_8 FILLER_42_123 ();
 sg13g2_decap_8 FILLER_42_130 ();
 sg13g2_decap_8 FILLER_42_137 ();
 sg13g2_decap_8 FILLER_42_144 ();
 sg13g2_decap_8 FILLER_42_151 ();
 sg13g2_decap_8 FILLER_42_158 ();
 sg13g2_decap_8 FILLER_42_165 ();
 sg13g2_decap_8 FILLER_42_172 ();
 sg13g2_decap_8 FILLER_42_179 ();
 sg13g2_decap_8 FILLER_42_186 ();
 sg13g2_decap_8 FILLER_42_193 ();
 sg13g2_decap_8 FILLER_42_200 ();
 sg13g2_decap_8 FILLER_42_207 ();
 sg13g2_decap_8 FILLER_42_214 ();
 sg13g2_decap_8 FILLER_42_221 ();
 sg13g2_decap_8 FILLER_42_228 ();
 sg13g2_decap_8 FILLER_42_235 ();
 sg13g2_decap_8 FILLER_42_242 ();
 sg13g2_decap_8 FILLER_42_249 ();
 sg13g2_decap_8 FILLER_42_256 ();
 sg13g2_decap_8 FILLER_42_263 ();
 sg13g2_decap_8 FILLER_42_270 ();
 sg13g2_decap_8 FILLER_42_277 ();
 sg13g2_decap_8 FILLER_42_284 ();
 sg13g2_decap_8 FILLER_42_291 ();
 sg13g2_decap_8 FILLER_42_298 ();
 sg13g2_decap_8 FILLER_42_305 ();
 sg13g2_decap_8 FILLER_42_312 ();
 sg13g2_decap_8 FILLER_42_319 ();
 sg13g2_decap_8 FILLER_42_326 ();
 sg13g2_decap_8 FILLER_42_333 ();
 sg13g2_decap_8 FILLER_42_340 ();
 sg13g2_decap_8 FILLER_42_347 ();
 sg13g2_decap_8 FILLER_42_354 ();
 sg13g2_decap_8 FILLER_42_361 ();
 sg13g2_decap_8 FILLER_42_368 ();
 sg13g2_decap_8 FILLER_42_375 ();
 sg13g2_decap_8 FILLER_42_382 ();
 sg13g2_decap_8 FILLER_42_389 ();
 sg13g2_decap_8 FILLER_42_396 ();
 sg13g2_decap_8 FILLER_42_403 ();
 sg13g2_decap_8 FILLER_42_410 ();
 sg13g2_decap_8 FILLER_42_417 ();
 sg13g2_decap_8 FILLER_42_424 ();
 sg13g2_decap_8 FILLER_42_431 ();
 sg13g2_decap_8 FILLER_42_438 ();
 sg13g2_decap_8 FILLER_42_445 ();
 sg13g2_decap_8 FILLER_42_452 ();
 sg13g2_decap_8 FILLER_42_459 ();
 sg13g2_decap_8 FILLER_42_466 ();
 sg13g2_decap_8 FILLER_42_473 ();
 sg13g2_decap_8 FILLER_42_480 ();
 sg13g2_decap_8 FILLER_42_487 ();
 sg13g2_decap_8 FILLER_42_494 ();
 sg13g2_decap_8 FILLER_42_501 ();
 sg13g2_decap_8 FILLER_42_508 ();
 sg13g2_decap_8 FILLER_42_515 ();
 sg13g2_decap_8 FILLER_42_522 ();
 sg13g2_decap_8 FILLER_42_529 ();
 sg13g2_decap_8 FILLER_42_536 ();
 sg13g2_decap_8 FILLER_42_543 ();
 sg13g2_decap_8 FILLER_42_550 ();
 sg13g2_decap_8 FILLER_42_557 ();
 sg13g2_decap_8 FILLER_42_564 ();
 sg13g2_decap_8 FILLER_42_571 ();
 sg13g2_decap_8 FILLER_42_578 ();
 sg13g2_decap_8 FILLER_42_585 ();
 sg13g2_decap_8 FILLER_42_592 ();
 sg13g2_decap_8 FILLER_42_599 ();
 sg13g2_decap_8 FILLER_42_606 ();
 sg13g2_decap_8 FILLER_42_613 ();
 sg13g2_decap_8 FILLER_42_620 ();
 sg13g2_decap_8 FILLER_42_627 ();
 sg13g2_decap_8 FILLER_42_634 ();
 sg13g2_decap_8 FILLER_42_641 ();
 sg13g2_decap_8 FILLER_42_648 ();
 sg13g2_decap_8 FILLER_42_655 ();
 sg13g2_decap_8 FILLER_42_662 ();
 sg13g2_decap_8 FILLER_42_669 ();
 sg13g2_decap_8 FILLER_42_676 ();
 sg13g2_decap_8 FILLER_42_683 ();
 sg13g2_decap_8 FILLER_42_690 ();
 sg13g2_decap_8 FILLER_42_697 ();
 sg13g2_decap_8 FILLER_42_704 ();
 sg13g2_decap_8 FILLER_42_711 ();
 sg13g2_decap_8 FILLER_42_718 ();
 sg13g2_decap_8 FILLER_42_725 ();
 sg13g2_decap_8 FILLER_42_732 ();
 sg13g2_decap_8 FILLER_42_739 ();
 sg13g2_decap_8 FILLER_42_746 ();
 sg13g2_decap_8 FILLER_42_753 ();
 sg13g2_decap_8 FILLER_42_760 ();
 sg13g2_decap_8 FILLER_42_767 ();
 sg13g2_decap_8 FILLER_42_774 ();
 sg13g2_decap_8 FILLER_42_781 ();
 sg13g2_decap_8 FILLER_42_788 ();
 sg13g2_decap_8 FILLER_42_795 ();
 sg13g2_decap_8 FILLER_42_802 ();
 sg13g2_decap_8 FILLER_42_809 ();
 sg13g2_decap_8 FILLER_42_816 ();
 sg13g2_decap_8 FILLER_42_823 ();
 sg13g2_decap_8 FILLER_42_830 ();
 sg13g2_decap_8 FILLER_42_837 ();
 sg13g2_decap_8 FILLER_42_844 ();
 sg13g2_decap_8 FILLER_42_851 ();
 sg13g2_decap_8 FILLER_42_858 ();
 sg13g2_decap_8 FILLER_42_865 ();
 sg13g2_decap_8 FILLER_42_872 ();
 sg13g2_decap_8 FILLER_42_879 ();
 sg13g2_decap_8 FILLER_42_886 ();
 sg13g2_decap_8 FILLER_42_893 ();
 sg13g2_decap_8 FILLER_42_900 ();
 sg13g2_decap_8 FILLER_42_907 ();
 sg13g2_decap_8 FILLER_42_914 ();
 sg13g2_decap_8 FILLER_42_921 ();
 sg13g2_decap_8 FILLER_42_928 ();
 sg13g2_decap_8 FILLER_42_935 ();
 sg13g2_decap_8 FILLER_42_942 ();
 sg13g2_decap_8 FILLER_42_949 ();
 sg13g2_decap_8 FILLER_42_956 ();
 sg13g2_decap_8 FILLER_42_963 ();
 sg13g2_decap_8 FILLER_42_970 ();
 sg13g2_decap_8 FILLER_42_977 ();
 sg13g2_decap_8 FILLER_42_984 ();
 sg13g2_decap_8 FILLER_42_991 ();
 sg13g2_decap_8 FILLER_42_998 ();
 sg13g2_decap_8 FILLER_42_1005 ();
 sg13g2_decap_8 FILLER_42_1012 ();
 sg13g2_decap_8 FILLER_42_1019 ();
 sg13g2_fill_2 FILLER_42_1026 ();
 sg13g2_fill_1 FILLER_42_1028 ();
 sg13g2_decap_8 FILLER_43_0 ();
 sg13g2_decap_8 FILLER_43_7 ();
 sg13g2_decap_8 FILLER_43_14 ();
 sg13g2_decap_8 FILLER_43_21 ();
 sg13g2_decap_8 FILLER_43_28 ();
 sg13g2_decap_8 FILLER_43_35 ();
 sg13g2_decap_8 FILLER_43_42 ();
 sg13g2_decap_8 FILLER_43_49 ();
 sg13g2_decap_8 FILLER_43_56 ();
 sg13g2_decap_8 FILLER_43_63 ();
 sg13g2_decap_8 FILLER_43_70 ();
 sg13g2_decap_8 FILLER_43_77 ();
 sg13g2_decap_8 FILLER_43_84 ();
 sg13g2_decap_8 FILLER_43_91 ();
 sg13g2_decap_8 FILLER_43_98 ();
 sg13g2_decap_8 FILLER_43_105 ();
 sg13g2_decap_8 FILLER_43_112 ();
 sg13g2_decap_8 FILLER_43_119 ();
 sg13g2_decap_8 FILLER_43_126 ();
 sg13g2_decap_8 FILLER_43_133 ();
 sg13g2_decap_8 FILLER_43_140 ();
 sg13g2_decap_8 FILLER_43_147 ();
 sg13g2_decap_8 FILLER_43_154 ();
 sg13g2_decap_8 FILLER_43_161 ();
 sg13g2_decap_8 FILLER_43_168 ();
 sg13g2_decap_8 FILLER_43_175 ();
 sg13g2_decap_8 FILLER_43_182 ();
 sg13g2_decap_8 FILLER_43_189 ();
 sg13g2_decap_8 FILLER_43_196 ();
 sg13g2_decap_8 FILLER_43_203 ();
 sg13g2_decap_8 FILLER_43_210 ();
 sg13g2_decap_8 FILLER_43_217 ();
 sg13g2_decap_8 FILLER_43_224 ();
 sg13g2_decap_8 FILLER_43_231 ();
 sg13g2_decap_8 FILLER_43_238 ();
 sg13g2_decap_8 FILLER_43_245 ();
 sg13g2_decap_8 FILLER_43_252 ();
 sg13g2_decap_8 FILLER_43_259 ();
 sg13g2_decap_8 FILLER_43_266 ();
 sg13g2_decap_8 FILLER_43_273 ();
 sg13g2_decap_8 FILLER_43_280 ();
 sg13g2_decap_8 FILLER_43_287 ();
 sg13g2_decap_8 FILLER_43_294 ();
 sg13g2_decap_8 FILLER_43_301 ();
 sg13g2_decap_8 FILLER_43_308 ();
 sg13g2_decap_8 FILLER_43_315 ();
 sg13g2_decap_8 FILLER_43_322 ();
 sg13g2_decap_8 FILLER_43_329 ();
 sg13g2_decap_8 FILLER_43_336 ();
 sg13g2_decap_8 FILLER_43_343 ();
 sg13g2_decap_8 FILLER_43_350 ();
 sg13g2_decap_8 FILLER_43_357 ();
 sg13g2_decap_8 FILLER_43_364 ();
 sg13g2_decap_8 FILLER_43_371 ();
 sg13g2_decap_8 FILLER_43_378 ();
 sg13g2_decap_8 FILLER_43_385 ();
 sg13g2_decap_8 FILLER_43_392 ();
 sg13g2_decap_8 FILLER_43_399 ();
 sg13g2_decap_8 FILLER_43_406 ();
 sg13g2_decap_8 FILLER_43_413 ();
 sg13g2_decap_8 FILLER_43_420 ();
 sg13g2_decap_8 FILLER_43_427 ();
 sg13g2_decap_8 FILLER_43_434 ();
 sg13g2_decap_8 FILLER_43_441 ();
 sg13g2_decap_8 FILLER_43_448 ();
 sg13g2_decap_8 FILLER_43_455 ();
 sg13g2_decap_8 FILLER_43_462 ();
 sg13g2_decap_8 FILLER_43_469 ();
 sg13g2_decap_8 FILLER_43_476 ();
 sg13g2_decap_8 FILLER_43_483 ();
 sg13g2_decap_8 FILLER_43_490 ();
 sg13g2_decap_8 FILLER_43_497 ();
 sg13g2_decap_8 FILLER_43_504 ();
 sg13g2_decap_8 FILLER_43_511 ();
 sg13g2_decap_8 FILLER_43_518 ();
 sg13g2_decap_8 FILLER_43_525 ();
 sg13g2_decap_8 FILLER_43_532 ();
 sg13g2_decap_8 FILLER_43_539 ();
 sg13g2_decap_8 FILLER_43_546 ();
 sg13g2_decap_8 FILLER_43_553 ();
 sg13g2_decap_8 FILLER_43_560 ();
 sg13g2_decap_8 FILLER_43_567 ();
 sg13g2_decap_8 FILLER_43_574 ();
 sg13g2_decap_8 FILLER_43_581 ();
 sg13g2_decap_8 FILLER_43_588 ();
 sg13g2_decap_8 FILLER_43_595 ();
 sg13g2_decap_8 FILLER_43_602 ();
 sg13g2_decap_8 FILLER_43_609 ();
 sg13g2_decap_8 FILLER_43_616 ();
 sg13g2_decap_8 FILLER_43_623 ();
 sg13g2_decap_8 FILLER_43_630 ();
 sg13g2_decap_8 FILLER_43_637 ();
 sg13g2_decap_8 FILLER_43_644 ();
 sg13g2_decap_8 FILLER_43_651 ();
 sg13g2_decap_8 FILLER_43_658 ();
 sg13g2_decap_8 FILLER_43_665 ();
 sg13g2_decap_8 FILLER_43_672 ();
 sg13g2_decap_8 FILLER_43_679 ();
 sg13g2_decap_8 FILLER_43_686 ();
 sg13g2_decap_8 FILLER_43_693 ();
 sg13g2_decap_8 FILLER_43_700 ();
 sg13g2_decap_8 FILLER_43_707 ();
 sg13g2_decap_8 FILLER_43_714 ();
 sg13g2_decap_8 FILLER_43_721 ();
 sg13g2_decap_8 FILLER_43_728 ();
 sg13g2_decap_8 FILLER_43_735 ();
 sg13g2_decap_8 FILLER_43_742 ();
 sg13g2_decap_8 FILLER_43_749 ();
 sg13g2_decap_8 FILLER_43_756 ();
 sg13g2_decap_8 FILLER_43_763 ();
 sg13g2_decap_8 FILLER_43_770 ();
 sg13g2_decap_8 FILLER_43_777 ();
 sg13g2_decap_8 FILLER_43_784 ();
 sg13g2_decap_8 FILLER_43_791 ();
 sg13g2_decap_8 FILLER_43_798 ();
 sg13g2_decap_8 FILLER_43_805 ();
 sg13g2_decap_8 FILLER_43_812 ();
 sg13g2_decap_8 FILLER_43_819 ();
 sg13g2_decap_8 FILLER_43_826 ();
 sg13g2_decap_8 FILLER_43_833 ();
 sg13g2_decap_8 FILLER_43_840 ();
 sg13g2_decap_8 FILLER_43_847 ();
 sg13g2_decap_8 FILLER_43_854 ();
 sg13g2_decap_8 FILLER_43_861 ();
 sg13g2_decap_8 FILLER_43_868 ();
 sg13g2_decap_8 FILLER_43_875 ();
 sg13g2_decap_8 FILLER_43_882 ();
 sg13g2_decap_8 FILLER_43_889 ();
 sg13g2_decap_8 FILLER_43_896 ();
 sg13g2_decap_8 FILLER_43_903 ();
 sg13g2_decap_8 FILLER_43_910 ();
 sg13g2_decap_8 FILLER_43_917 ();
 sg13g2_decap_8 FILLER_43_924 ();
 sg13g2_decap_8 FILLER_43_931 ();
 sg13g2_decap_8 FILLER_43_938 ();
 sg13g2_decap_8 FILLER_43_945 ();
 sg13g2_decap_8 FILLER_43_952 ();
 sg13g2_decap_8 FILLER_43_959 ();
 sg13g2_decap_8 FILLER_43_966 ();
 sg13g2_decap_8 FILLER_43_973 ();
 sg13g2_decap_8 FILLER_43_980 ();
 sg13g2_decap_8 FILLER_43_987 ();
 sg13g2_decap_8 FILLER_43_994 ();
 sg13g2_decap_8 FILLER_43_1001 ();
 sg13g2_decap_8 FILLER_43_1008 ();
 sg13g2_decap_8 FILLER_43_1015 ();
 sg13g2_decap_8 FILLER_43_1022 ();
 sg13g2_decap_8 FILLER_44_4 ();
 sg13g2_decap_8 FILLER_44_11 ();
 sg13g2_decap_8 FILLER_44_18 ();
 sg13g2_decap_8 FILLER_44_25 ();
 sg13g2_decap_8 FILLER_44_32 ();
 sg13g2_decap_8 FILLER_44_39 ();
 sg13g2_decap_8 FILLER_44_46 ();
 sg13g2_decap_8 FILLER_44_53 ();
 sg13g2_decap_8 FILLER_44_60 ();
 sg13g2_decap_8 FILLER_44_67 ();
 sg13g2_decap_8 FILLER_44_74 ();
 sg13g2_decap_8 FILLER_44_81 ();
 sg13g2_decap_8 FILLER_44_88 ();
 sg13g2_decap_8 FILLER_44_95 ();
 sg13g2_decap_8 FILLER_44_102 ();
 sg13g2_decap_8 FILLER_44_109 ();
 sg13g2_decap_8 FILLER_44_116 ();
 sg13g2_decap_8 FILLER_44_123 ();
 sg13g2_decap_8 FILLER_44_130 ();
 sg13g2_decap_8 FILLER_44_137 ();
 sg13g2_decap_8 FILLER_44_144 ();
 sg13g2_decap_8 FILLER_44_151 ();
 sg13g2_decap_8 FILLER_44_158 ();
 sg13g2_decap_8 FILLER_44_165 ();
 sg13g2_decap_8 FILLER_44_172 ();
 sg13g2_decap_8 FILLER_44_179 ();
 sg13g2_decap_8 FILLER_44_186 ();
 sg13g2_decap_8 FILLER_44_193 ();
 sg13g2_decap_8 FILLER_44_200 ();
 sg13g2_decap_8 FILLER_44_207 ();
 sg13g2_decap_8 FILLER_44_214 ();
 sg13g2_decap_8 FILLER_44_221 ();
 sg13g2_decap_8 FILLER_44_228 ();
 sg13g2_decap_8 FILLER_44_235 ();
 sg13g2_decap_8 FILLER_44_242 ();
 sg13g2_decap_8 FILLER_44_249 ();
 sg13g2_decap_8 FILLER_44_256 ();
 sg13g2_decap_8 FILLER_44_263 ();
 sg13g2_decap_8 FILLER_44_270 ();
 sg13g2_decap_8 FILLER_44_277 ();
 sg13g2_decap_8 FILLER_44_284 ();
 sg13g2_decap_8 FILLER_44_291 ();
 sg13g2_decap_8 FILLER_44_298 ();
 sg13g2_decap_8 FILLER_44_305 ();
 sg13g2_decap_8 FILLER_44_312 ();
 sg13g2_decap_8 FILLER_44_319 ();
 sg13g2_decap_8 FILLER_44_326 ();
 sg13g2_decap_8 FILLER_44_333 ();
 sg13g2_decap_8 FILLER_44_340 ();
 sg13g2_decap_8 FILLER_44_347 ();
 sg13g2_decap_8 FILLER_44_354 ();
 sg13g2_decap_8 FILLER_44_361 ();
 sg13g2_decap_8 FILLER_44_368 ();
 sg13g2_decap_8 FILLER_44_375 ();
 sg13g2_decap_8 FILLER_44_382 ();
 sg13g2_decap_8 FILLER_44_389 ();
 sg13g2_decap_8 FILLER_44_396 ();
 sg13g2_decap_8 FILLER_44_403 ();
 sg13g2_decap_8 FILLER_44_410 ();
 sg13g2_decap_8 FILLER_44_417 ();
 sg13g2_decap_8 FILLER_44_424 ();
 sg13g2_decap_8 FILLER_44_431 ();
 sg13g2_decap_8 FILLER_44_438 ();
 sg13g2_decap_8 FILLER_44_445 ();
 sg13g2_decap_8 FILLER_44_452 ();
 sg13g2_decap_8 FILLER_44_459 ();
 sg13g2_decap_8 FILLER_44_466 ();
 sg13g2_decap_8 FILLER_44_473 ();
 sg13g2_decap_8 FILLER_44_480 ();
 sg13g2_decap_8 FILLER_44_487 ();
 sg13g2_decap_8 FILLER_44_494 ();
 sg13g2_decap_8 FILLER_44_501 ();
 sg13g2_decap_8 FILLER_44_508 ();
 sg13g2_decap_8 FILLER_44_515 ();
 sg13g2_decap_8 FILLER_44_522 ();
 sg13g2_decap_8 FILLER_44_529 ();
 sg13g2_decap_8 FILLER_44_536 ();
 sg13g2_decap_8 FILLER_44_543 ();
 sg13g2_decap_8 FILLER_44_550 ();
 sg13g2_decap_8 FILLER_44_557 ();
 sg13g2_decap_8 FILLER_44_564 ();
 sg13g2_decap_8 FILLER_44_571 ();
 sg13g2_decap_8 FILLER_44_578 ();
 sg13g2_decap_8 FILLER_44_585 ();
 sg13g2_decap_8 FILLER_44_592 ();
 sg13g2_decap_8 FILLER_44_599 ();
 sg13g2_decap_8 FILLER_44_606 ();
 sg13g2_decap_8 FILLER_44_613 ();
 sg13g2_decap_8 FILLER_44_620 ();
 sg13g2_decap_8 FILLER_44_627 ();
 sg13g2_decap_8 FILLER_44_634 ();
 sg13g2_decap_8 FILLER_44_641 ();
 sg13g2_decap_8 FILLER_44_648 ();
 sg13g2_decap_8 FILLER_44_655 ();
 sg13g2_decap_8 FILLER_44_662 ();
 sg13g2_decap_8 FILLER_44_669 ();
 sg13g2_decap_8 FILLER_44_676 ();
 sg13g2_decap_8 FILLER_44_683 ();
 sg13g2_decap_8 FILLER_44_690 ();
 sg13g2_decap_8 FILLER_44_697 ();
 sg13g2_decap_8 FILLER_44_704 ();
 sg13g2_decap_8 FILLER_44_711 ();
 sg13g2_decap_8 FILLER_44_718 ();
 sg13g2_decap_8 FILLER_44_725 ();
 sg13g2_decap_8 FILLER_44_732 ();
 sg13g2_decap_8 FILLER_44_739 ();
 sg13g2_decap_8 FILLER_44_746 ();
 sg13g2_decap_8 FILLER_44_753 ();
 sg13g2_decap_8 FILLER_44_760 ();
 sg13g2_decap_8 FILLER_44_767 ();
 sg13g2_decap_8 FILLER_44_774 ();
 sg13g2_decap_8 FILLER_44_781 ();
 sg13g2_decap_8 FILLER_44_788 ();
 sg13g2_decap_8 FILLER_44_795 ();
 sg13g2_decap_8 FILLER_44_802 ();
 sg13g2_decap_8 FILLER_44_809 ();
 sg13g2_decap_8 FILLER_44_816 ();
 sg13g2_decap_8 FILLER_44_823 ();
 sg13g2_decap_8 FILLER_44_830 ();
 sg13g2_decap_8 FILLER_44_837 ();
 sg13g2_decap_8 FILLER_44_844 ();
 sg13g2_decap_8 FILLER_44_851 ();
 sg13g2_decap_8 FILLER_44_858 ();
 sg13g2_decap_8 FILLER_44_865 ();
 sg13g2_decap_8 FILLER_44_872 ();
 sg13g2_decap_8 FILLER_44_879 ();
 sg13g2_decap_8 FILLER_44_886 ();
 sg13g2_decap_8 FILLER_44_893 ();
 sg13g2_decap_8 FILLER_44_900 ();
 sg13g2_decap_8 FILLER_44_907 ();
 sg13g2_decap_8 FILLER_44_914 ();
 sg13g2_decap_8 FILLER_44_921 ();
 sg13g2_decap_8 FILLER_44_928 ();
 sg13g2_decap_8 FILLER_44_935 ();
 sg13g2_decap_8 FILLER_44_942 ();
 sg13g2_decap_8 FILLER_44_949 ();
 sg13g2_decap_8 FILLER_44_956 ();
 sg13g2_decap_8 FILLER_44_963 ();
 sg13g2_decap_8 FILLER_44_970 ();
 sg13g2_decap_8 FILLER_44_977 ();
 sg13g2_decap_8 FILLER_44_984 ();
 sg13g2_decap_8 FILLER_44_991 ();
 sg13g2_decap_8 FILLER_44_998 ();
 sg13g2_decap_8 FILLER_44_1005 ();
 sg13g2_decap_8 FILLER_44_1012 ();
 sg13g2_decap_8 FILLER_44_1019 ();
 sg13g2_fill_2 FILLER_44_1026 ();
 sg13g2_fill_1 FILLER_44_1028 ();
 sg13g2_decap_8 FILLER_45_0 ();
 sg13g2_decap_8 FILLER_45_7 ();
 sg13g2_decap_8 FILLER_45_14 ();
 sg13g2_decap_8 FILLER_45_21 ();
 sg13g2_decap_8 FILLER_45_28 ();
 sg13g2_decap_8 FILLER_45_35 ();
 sg13g2_decap_8 FILLER_45_42 ();
 sg13g2_decap_8 FILLER_45_49 ();
 sg13g2_decap_8 FILLER_45_56 ();
 sg13g2_decap_8 FILLER_45_63 ();
 sg13g2_decap_8 FILLER_45_70 ();
 sg13g2_decap_8 FILLER_45_77 ();
 sg13g2_decap_8 FILLER_45_84 ();
 sg13g2_decap_8 FILLER_45_91 ();
 sg13g2_decap_8 FILLER_45_98 ();
 sg13g2_decap_8 FILLER_45_105 ();
 sg13g2_decap_8 FILLER_45_112 ();
 sg13g2_decap_8 FILLER_45_119 ();
 sg13g2_decap_8 FILLER_45_126 ();
 sg13g2_decap_8 FILLER_45_133 ();
 sg13g2_decap_8 FILLER_45_140 ();
 sg13g2_decap_8 FILLER_45_147 ();
 sg13g2_decap_8 FILLER_45_154 ();
 sg13g2_decap_8 FILLER_45_161 ();
 sg13g2_decap_8 FILLER_45_168 ();
 sg13g2_decap_8 FILLER_45_175 ();
 sg13g2_decap_8 FILLER_45_182 ();
 sg13g2_decap_8 FILLER_45_189 ();
 sg13g2_decap_8 FILLER_45_196 ();
 sg13g2_decap_8 FILLER_45_203 ();
 sg13g2_decap_8 FILLER_45_210 ();
 sg13g2_decap_8 FILLER_45_217 ();
 sg13g2_decap_8 FILLER_45_224 ();
 sg13g2_decap_8 FILLER_45_231 ();
 sg13g2_decap_8 FILLER_45_238 ();
 sg13g2_decap_8 FILLER_45_245 ();
 sg13g2_decap_8 FILLER_45_252 ();
 sg13g2_decap_8 FILLER_45_259 ();
 sg13g2_decap_8 FILLER_45_266 ();
 sg13g2_decap_8 FILLER_45_273 ();
 sg13g2_decap_8 FILLER_45_280 ();
 sg13g2_decap_8 FILLER_45_287 ();
 sg13g2_decap_8 FILLER_45_294 ();
 sg13g2_decap_8 FILLER_45_301 ();
 sg13g2_decap_8 FILLER_45_308 ();
 sg13g2_decap_8 FILLER_45_315 ();
 sg13g2_decap_8 FILLER_45_322 ();
 sg13g2_decap_8 FILLER_45_329 ();
 sg13g2_decap_8 FILLER_45_336 ();
 sg13g2_decap_8 FILLER_45_343 ();
 sg13g2_decap_8 FILLER_45_350 ();
 sg13g2_decap_8 FILLER_45_357 ();
 sg13g2_decap_8 FILLER_45_364 ();
 sg13g2_decap_8 FILLER_45_371 ();
 sg13g2_decap_8 FILLER_45_378 ();
 sg13g2_decap_8 FILLER_45_385 ();
 sg13g2_decap_8 FILLER_45_392 ();
 sg13g2_decap_8 FILLER_45_399 ();
 sg13g2_decap_8 FILLER_45_406 ();
 sg13g2_decap_8 FILLER_45_413 ();
 sg13g2_decap_8 FILLER_45_420 ();
 sg13g2_decap_8 FILLER_45_427 ();
 sg13g2_decap_8 FILLER_45_434 ();
 sg13g2_decap_8 FILLER_45_441 ();
 sg13g2_decap_8 FILLER_45_448 ();
 sg13g2_decap_8 FILLER_45_455 ();
 sg13g2_decap_8 FILLER_45_462 ();
 sg13g2_decap_8 FILLER_45_469 ();
 sg13g2_decap_8 FILLER_45_476 ();
 sg13g2_decap_8 FILLER_45_483 ();
 sg13g2_decap_8 FILLER_45_490 ();
 sg13g2_decap_8 FILLER_45_497 ();
 sg13g2_decap_8 FILLER_45_504 ();
 sg13g2_decap_8 FILLER_45_511 ();
 sg13g2_decap_8 FILLER_45_518 ();
 sg13g2_decap_8 FILLER_45_525 ();
 sg13g2_decap_8 FILLER_45_532 ();
 sg13g2_decap_8 FILLER_45_539 ();
 sg13g2_decap_8 FILLER_45_546 ();
 sg13g2_decap_8 FILLER_45_553 ();
 sg13g2_decap_8 FILLER_45_560 ();
 sg13g2_decap_8 FILLER_45_567 ();
 sg13g2_decap_8 FILLER_45_574 ();
 sg13g2_decap_8 FILLER_45_581 ();
 sg13g2_decap_8 FILLER_45_588 ();
 sg13g2_decap_8 FILLER_45_595 ();
 sg13g2_decap_8 FILLER_45_602 ();
 sg13g2_decap_8 FILLER_45_609 ();
 sg13g2_decap_8 FILLER_45_616 ();
 sg13g2_decap_8 FILLER_45_623 ();
 sg13g2_decap_8 FILLER_45_630 ();
 sg13g2_decap_8 FILLER_45_637 ();
 sg13g2_decap_8 FILLER_45_644 ();
 sg13g2_decap_8 FILLER_45_651 ();
 sg13g2_decap_8 FILLER_45_658 ();
 sg13g2_decap_8 FILLER_45_665 ();
 sg13g2_decap_8 FILLER_45_672 ();
 sg13g2_decap_8 FILLER_45_679 ();
 sg13g2_decap_8 FILLER_45_686 ();
 sg13g2_decap_8 FILLER_45_693 ();
 sg13g2_decap_8 FILLER_45_700 ();
 sg13g2_decap_8 FILLER_45_707 ();
 sg13g2_decap_8 FILLER_45_714 ();
 sg13g2_decap_8 FILLER_45_721 ();
 sg13g2_decap_8 FILLER_45_728 ();
 sg13g2_decap_8 FILLER_45_735 ();
 sg13g2_decap_8 FILLER_45_742 ();
 sg13g2_decap_8 FILLER_45_749 ();
 sg13g2_decap_8 FILLER_45_756 ();
 sg13g2_decap_8 FILLER_45_763 ();
 sg13g2_decap_8 FILLER_45_770 ();
 sg13g2_decap_8 FILLER_45_777 ();
 sg13g2_decap_8 FILLER_45_784 ();
 sg13g2_decap_8 FILLER_45_791 ();
 sg13g2_decap_8 FILLER_45_798 ();
 sg13g2_decap_8 FILLER_45_805 ();
 sg13g2_decap_8 FILLER_45_812 ();
 sg13g2_decap_8 FILLER_45_819 ();
 sg13g2_decap_8 FILLER_45_826 ();
 sg13g2_decap_8 FILLER_45_833 ();
 sg13g2_decap_8 FILLER_45_840 ();
 sg13g2_decap_8 FILLER_45_847 ();
 sg13g2_decap_8 FILLER_45_854 ();
 sg13g2_decap_8 FILLER_45_861 ();
 sg13g2_decap_8 FILLER_45_868 ();
 sg13g2_decap_8 FILLER_45_875 ();
 sg13g2_decap_8 FILLER_45_882 ();
 sg13g2_decap_8 FILLER_45_889 ();
 sg13g2_decap_8 FILLER_45_896 ();
 sg13g2_decap_8 FILLER_45_903 ();
 sg13g2_decap_8 FILLER_45_910 ();
 sg13g2_decap_8 FILLER_45_917 ();
 sg13g2_decap_8 FILLER_45_924 ();
 sg13g2_decap_8 FILLER_45_931 ();
 sg13g2_decap_8 FILLER_45_938 ();
 sg13g2_decap_8 FILLER_45_945 ();
 sg13g2_decap_8 FILLER_45_952 ();
 sg13g2_decap_8 FILLER_45_959 ();
 sg13g2_decap_8 FILLER_45_966 ();
 sg13g2_decap_8 FILLER_45_973 ();
 sg13g2_decap_8 FILLER_45_980 ();
 sg13g2_decap_8 FILLER_45_987 ();
 sg13g2_decap_8 FILLER_45_994 ();
 sg13g2_decap_8 FILLER_45_1001 ();
 sg13g2_decap_8 FILLER_45_1008 ();
 sg13g2_decap_8 FILLER_45_1015 ();
 sg13g2_decap_8 FILLER_45_1022 ();
 sg13g2_decap_8 FILLER_46_4 ();
 sg13g2_decap_8 FILLER_46_11 ();
 sg13g2_decap_8 FILLER_46_18 ();
 sg13g2_decap_8 FILLER_46_25 ();
 sg13g2_decap_8 FILLER_46_32 ();
 sg13g2_decap_8 FILLER_46_39 ();
 sg13g2_decap_8 FILLER_46_46 ();
 sg13g2_decap_8 FILLER_46_53 ();
 sg13g2_decap_8 FILLER_46_60 ();
 sg13g2_decap_8 FILLER_46_67 ();
 sg13g2_decap_8 FILLER_46_74 ();
 sg13g2_decap_8 FILLER_46_81 ();
 sg13g2_decap_8 FILLER_46_88 ();
 sg13g2_decap_8 FILLER_46_95 ();
 sg13g2_decap_8 FILLER_46_102 ();
 sg13g2_decap_8 FILLER_46_109 ();
 sg13g2_decap_8 FILLER_46_116 ();
 sg13g2_decap_8 FILLER_46_123 ();
 sg13g2_decap_8 FILLER_46_130 ();
 sg13g2_decap_8 FILLER_46_137 ();
 sg13g2_decap_8 FILLER_46_144 ();
 sg13g2_decap_8 FILLER_46_151 ();
 sg13g2_decap_8 FILLER_46_158 ();
 sg13g2_decap_8 FILLER_46_165 ();
 sg13g2_decap_8 FILLER_46_172 ();
 sg13g2_decap_8 FILLER_46_179 ();
 sg13g2_decap_8 FILLER_46_186 ();
 sg13g2_decap_8 FILLER_46_193 ();
 sg13g2_decap_8 FILLER_46_200 ();
 sg13g2_decap_8 FILLER_46_207 ();
 sg13g2_decap_8 FILLER_46_214 ();
 sg13g2_decap_8 FILLER_46_221 ();
 sg13g2_decap_8 FILLER_46_228 ();
 sg13g2_decap_8 FILLER_46_235 ();
 sg13g2_decap_8 FILLER_46_242 ();
 sg13g2_decap_8 FILLER_46_249 ();
 sg13g2_decap_8 FILLER_46_256 ();
 sg13g2_decap_8 FILLER_46_263 ();
 sg13g2_decap_8 FILLER_46_270 ();
 sg13g2_decap_8 FILLER_46_277 ();
 sg13g2_decap_8 FILLER_46_284 ();
 sg13g2_decap_8 FILLER_46_291 ();
 sg13g2_decap_8 FILLER_46_298 ();
 sg13g2_decap_8 FILLER_46_305 ();
 sg13g2_decap_8 FILLER_46_312 ();
 sg13g2_decap_8 FILLER_46_319 ();
 sg13g2_decap_8 FILLER_46_326 ();
 sg13g2_decap_8 FILLER_46_333 ();
 sg13g2_decap_8 FILLER_46_340 ();
 sg13g2_decap_8 FILLER_46_347 ();
 sg13g2_decap_8 FILLER_46_354 ();
 sg13g2_decap_8 FILLER_46_361 ();
 sg13g2_decap_8 FILLER_46_368 ();
 sg13g2_decap_8 FILLER_46_375 ();
 sg13g2_decap_8 FILLER_46_382 ();
 sg13g2_decap_8 FILLER_46_389 ();
 sg13g2_decap_8 FILLER_46_396 ();
 sg13g2_decap_8 FILLER_46_403 ();
 sg13g2_decap_8 FILLER_46_410 ();
 sg13g2_decap_8 FILLER_46_417 ();
 sg13g2_decap_8 FILLER_46_424 ();
 sg13g2_decap_8 FILLER_46_431 ();
 sg13g2_decap_8 FILLER_46_438 ();
 sg13g2_decap_8 FILLER_46_445 ();
 sg13g2_decap_8 FILLER_46_452 ();
 sg13g2_decap_8 FILLER_46_459 ();
 sg13g2_decap_8 FILLER_46_466 ();
 sg13g2_decap_8 FILLER_46_473 ();
 sg13g2_decap_8 FILLER_46_480 ();
 sg13g2_decap_8 FILLER_46_487 ();
 sg13g2_decap_8 FILLER_46_494 ();
 sg13g2_decap_8 FILLER_46_501 ();
 sg13g2_decap_8 FILLER_46_508 ();
 sg13g2_decap_8 FILLER_46_515 ();
 sg13g2_decap_8 FILLER_46_522 ();
 sg13g2_decap_8 FILLER_46_529 ();
 sg13g2_decap_8 FILLER_46_536 ();
 sg13g2_decap_8 FILLER_46_543 ();
 sg13g2_decap_8 FILLER_46_550 ();
 sg13g2_decap_8 FILLER_46_557 ();
 sg13g2_decap_8 FILLER_46_564 ();
 sg13g2_decap_8 FILLER_46_571 ();
 sg13g2_decap_8 FILLER_46_578 ();
 sg13g2_decap_8 FILLER_46_585 ();
 sg13g2_decap_8 FILLER_46_592 ();
 sg13g2_decap_8 FILLER_46_599 ();
 sg13g2_decap_8 FILLER_46_606 ();
 sg13g2_decap_8 FILLER_46_613 ();
 sg13g2_decap_8 FILLER_46_620 ();
 sg13g2_decap_8 FILLER_46_627 ();
 sg13g2_decap_8 FILLER_46_634 ();
 sg13g2_decap_8 FILLER_46_641 ();
 sg13g2_decap_8 FILLER_46_648 ();
 sg13g2_decap_8 FILLER_46_655 ();
 sg13g2_decap_8 FILLER_46_662 ();
 sg13g2_decap_8 FILLER_46_669 ();
 sg13g2_decap_8 FILLER_46_676 ();
 sg13g2_decap_8 FILLER_46_683 ();
 sg13g2_decap_8 FILLER_46_690 ();
 sg13g2_decap_8 FILLER_46_697 ();
 sg13g2_decap_8 FILLER_46_704 ();
 sg13g2_decap_8 FILLER_46_711 ();
 sg13g2_decap_8 FILLER_46_718 ();
 sg13g2_decap_8 FILLER_46_725 ();
 sg13g2_decap_8 FILLER_46_732 ();
 sg13g2_decap_8 FILLER_46_739 ();
 sg13g2_decap_8 FILLER_46_746 ();
 sg13g2_decap_8 FILLER_46_753 ();
 sg13g2_decap_8 FILLER_46_760 ();
 sg13g2_decap_8 FILLER_46_767 ();
 sg13g2_decap_8 FILLER_46_774 ();
 sg13g2_decap_8 FILLER_46_781 ();
 sg13g2_decap_8 FILLER_46_788 ();
 sg13g2_decap_8 FILLER_46_795 ();
 sg13g2_decap_8 FILLER_46_802 ();
 sg13g2_decap_8 FILLER_46_809 ();
 sg13g2_decap_8 FILLER_46_816 ();
 sg13g2_decap_8 FILLER_46_823 ();
 sg13g2_decap_8 FILLER_46_830 ();
 sg13g2_decap_8 FILLER_46_837 ();
 sg13g2_decap_8 FILLER_46_844 ();
 sg13g2_decap_8 FILLER_46_851 ();
 sg13g2_decap_8 FILLER_46_858 ();
 sg13g2_decap_8 FILLER_46_865 ();
 sg13g2_decap_8 FILLER_46_872 ();
 sg13g2_decap_8 FILLER_46_879 ();
 sg13g2_decap_8 FILLER_46_886 ();
 sg13g2_decap_8 FILLER_46_893 ();
 sg13g2_decap_8 FILLER_46_900 ();
 sg13g2_decap_8 FILLER_46_907 ();
 sg13g2_decap_8 FILLER_46_914 ();
 sg13g2_decap_8 FILLER_46_921 ();
 sg13g2_decap_8 FILLER_46_928 ();
 sg13g2_decap_8 FILLER_46_935 ();
 sg13g2_decap_8 FILLER_46_942 ();
 sg13g2_decap_8 FILLER_46_949 ();
 sg13g2_decap_8 FILLER_46_956 ();
 sg13g2_decap_8 FILLER_46_963 ();
 sg13g2_decap_8 FILLER_46_970 ();
 sg13g2_decap_8 FILLER_46_977 ();
 sg13g2_decap_8 FILLER_46_984 ();
 sg13g2_decap_8 FILLER_46_991 ();
 sg13g2_decap_8 FILLER_46_998 ();
 sg13g2_decap_8 FILLER_46_1005 ();
 sg13g2_decap_8 FILLER_46_1012 ();
 sg13g2_decap_8 FILLER_46_1019 ();
 sg13g2_fill_2 FILLER_46_1026 ();
 sg13g2_fill_1 FILLER_46_1028 ();
 sg13g2_decap_8 FILLER_47_0 ();
 sg13g2_decap_8 FILLER_47_7 ();
 sg13g2_decap_8 FILLER_47_14 ();
 sg13g2_decap_8 FILLER_47_21 ();
 sg13g2_decap_8 FILLER_47_28 ();
 sg13g2_decap_8 FILLER_47_35 ();
 sg13g2_decap_8 FILLER_47_42 ();
 sg13g2_decap_8 FILLER_47_49 ();
 sg13g2_decap_8 FILLER_47_56 ();
 sg13g2_decap_8 FILLER_47_63 ();
 sg13g2_decap_8 FILLER_47_70 ();
 sg13g2_decap_8 FILLER_47_77 ();
 sg13g2_decap_8 FILLER_47_84 ();
 sg13g2_decap_8 FILLER_47_91 ();
 sg13g2_decap_8 FILLER_47_98 ();
 sg13g2_decap_8 FILLER_47_105 ();
 sg13g2_decap_8 FILLER_47_112 ();
 sg13g2_decap_8 FILLER_47_119 ();
 sg13g2_decap_8 FILLER_47_126 ();
 sg13g2_decap_8 FILLER_47_133 ();
 sg13g2_decap_8 FILLER_47_140 ();
 sg13g2_decap_8 FILLER_47_147 ();
 sg13g2_decap_8 FILLER_47_154 ();
 sg13g2_decap_8 FILLER_47_161 ();
 sg13g2_decap_8 FILLER_47_168 ();
 sg13g2_decap_8 FILLER_47_175 ();
 sg13g2_decap_8 FILLER_47_182 ();
 sg13g2_decap_8 FILLER_47_189 ();
 sg13g2_decap_8 FILLER_47_196 ();
 sg13g2_decap_8 FILLER_47_203 ();
 sg13g2_decap_8 FILLER_47_210 ();
 sg13g2_decap_8 FILLER_47_217 ();
 sg13g2_decap_8 FILLER_47_224 ();
 sg13g2_decap_8 FILLER_47_231 ();
 sg13g2_decap_8 FILLER_47_238 ();
 sg13g2_decap_8 FILLER_47_245 ();
 sg13g2_decap_8 FILLER_47_252 ();
 sg13g2_decap_8 FILLER_47_259 ();
 sg13g2_decap_8 FILLER_47_266 ();
 sg13g2_decap_8 FILLER_47_273 ();
 sg13g2_decap_8 FILLER_47_280 ();
 sg13g2_decap_8 FILLER_47_287 ();
 sg13g2_decap_8 FILLER_47_294 ();
 sg13g2_decap_8 FILLER_47_301 ();
 sg13g2_decap_8 FILLER_47_308 ();
 sg13g2_decap_8 FILLER_47_315 ();
 sg13g2_decap_8 FILLER_47_322 ();
 sg13g2_decap_8 FILLER_47_329 ();
 sg13g2_decap_8 FILLER_47_336 ();
 sg13g2_decap_8 FILLER_47_343 ();
 sg13g2_decap_8 FILLER_47_350 ();
 sg13g2_decap_8 FILLER_47_357 ();
 sg13g2_decap_8 FILLER_47_364 ();
 sg13g2_decap_8 FILLER_47_371 ();
 sg13g2_decap_8 FILLER_47_378 ();
 sg13g2_decap_8 FILLER_47_385 ();
 sg13g2_decap_8 FILLER_47_392 ();
 sg13g2_decap_8 FILLER_47_399 ();
 sg13g2_decap_8 FILLER_47_406 ();
 sg13g2_decap_8 FILLER_47_413 ();
 sg13g2_decap_8 FILLER_47_420 ();
 sg13g2_decap_8 FILLER_47_427 ();
 sg13g2_decap_8 FILLER_47_434 ();
 sg13g2_decap_8 FILLER_47_441 ();
 sg13g2_decap_8 FILLER_47_448 ();
 sg13g2_decap_8 FILLER_47_455 ();
 sg13g2_decap_8 FILLER_47_462 ();
 sg13g2_decap_8 FILLER_47_469 ();
 sg13g2_decap_8 FILLER_47_476 ();
 sg13g2_decap_8 FILLER_47_483 ();
 sg13g2_decap_8 FILLER_47_490 ();
 sg13g2_decap_8 FILLER_47_497 ();
 sg13g2_decap_8 FILLER_47_504 ();
 sg13g2_decap_8 FILLER_47_511 ();
 sg13g2_decap_8 FILLER_47_518 ();
 sg13g2_decap_8 FILLER_47_525 ();
 sg13g2_decap_8 FILLER_47_532 ();
 sg13g2_decap_8 FILLER_47_539 ();
 sg13g2_decap_8 FILLER_47_546 ();
 sg13g2_decap_8 FILLER_47_553 ();
 sg13g2_decap_8 FILLER_47_560 ();
 sg13g2_decap_8 FILLER_47_567 ();
 sg13g2_decap_8 FILLER_47_574 ();
 sg13g2_decap_8 FILLER_47_581 ();
 sg13g2_decap_8 FILLER_47_588 ();
 sg13g2_decap_8 FILLER_47_595 ();
 sg13g2_decap_8 FILLER_47_602 ();
 sg13g2_decap_8 FILLER_47_609 ();
 sg13g2_decap_8 FILLER_47_616 ();
 sg13g2_decap_8 FILLER_47_623 ();
 sg13g2_decap_8 FILLER_47_630 ();
 sg13g2_decap_8 FILLER_47_637 ();
 sg13g2_decap_8 FILLER_47_644 ();
 sg13g2_decap_8 FILLER_47_651 ();
 sg13g2_decap_8 FILLER_47_658 ();
 sg13g2_decap_8 FILLER_47_665 ();
 sg13g2_decap_8 FILLER_47_672 ();
 sg13g2_decap_8 FILLER_47_679 ();
 sg13g2_decap_8 FILLER_47_686 ();
 sg13g2_decap_8 FILLER_47_693 ();
 sg13g2_decap_8 FILLER_47_700 ();
 sg13g2_decap_8 FILLER_47_707 ();
 sg13g2_decap_8 FILLER_47_714 ();
 sg13g2_decap_8 FILLER_47_721 ();
 sg13g2_decap_8 FILLER_47_728 ();
 sg13g2_decap_8 FILLER_47_735 ();
 sg13g2_decap_8 FILLER_47_742 ();
 sg13g2_decap_8 FILLER_47_749 ();
 sg13g2_decap_8 FILLER_47_756 ();
 sg13g2_decap_8 FILLER_47_763 ();
 sg13g2_decap_8 FILLER_47_770 ();
 sg13g2_decap_8 FILLER_47_777 ();
 sg13g2_decap_8 FILLER_47_784 ();
 sg13g2_decap_8 FILLER_47_791 ();
 sg13g2_decap_8 FILLER_47_798 ();
 sg13g2_decap_8 FILLER_47_805 ();
 sg13g2_decap_8 FILLER_47_812 ();
 sg13g2_decap_8 FILLER_47_819 ();
 sg13g2_decap_8 FILLER_47_826 ();
 sg13g2_decap_8 FILLER_47_833 ();
 sg13g2_decap_8 FILLER_47_840 ();
 sg13g2_decap_8 FILLER_47_847 ();
 sg13g2_decap_8 FILLER_47_854 ();
 sg13g2_decap_8 FILLER_47_861 ();
 sg13g2_decap_8 FILLER_47_868 ();
 sg13g2_decap_8 FILLER_47_875 ();
 sg13g2_decap_8 FILLER_47_882 ();
 sg13g2_decap_8 FILLER_47_889 ();
 sg13g2_decap_8 FILLER_47_896 ();
 sg13g2_decap_8 FILLER_47_903 ();
 sg13g2_decap_8 FILLER_47_910 ();
 sg13g2_decap_8 FILLER_47_917 ();
 sg13g2_decap_8 FILLER_47_924 ();
 sg13g2_decap_8 FILLER_47_931 ();
 sg13g2_decap_8 FILLER_47_938 ();
 sg13g2_decap_8 FILLER_47_945 ();
 sg13g2_decap_8 FILLER_47_952 ();
 sg13g2_decap_8 FILLER_47_959 ();
 sg13g2_decap_8 FILLER_47_966 ();
 sg13g2_decap_8 FILLER_47_973 ();
 sg13g2_decap_8 FILLER_47_980 ();
 sg13g2_decap_8 FILLER_47_987 ();
 sg13g2_decap_8 FILLER_47_994 ();
 sg13g2_decap_8 FILLER_47_1001 ();
 sg13g2_decap_8 FILLER_47_1008 ();
 sg13g2_decap_8 FILLER_47_1015 ();
 sg13g2_decap_8 FILLER_47_1022 ();
 sg13g2_decap_8 FILLER_48_0 ();
 sg13g2_decap_8 FILLER_48_7 ();
 sg13g2_decap_8 FILLER_48_14 ();
 sg13g2_decap_8 FILLER_48_21 ();
 sg13g2_decap_8 FILLER_48_28 ();
 sg13g2_decap_8 FILLER_48_35 ();
 sg13g2_decap_8 FILLER_48_42 ();
 sg13g2_decap_8 FILLER_48_49 ();
 sg13g2_decap_8 FILLER_48_56 ();
 sg13g2_decap_8 FILLER_48_63 ();
 sg13g2_decap_8 FILLER_48_70 ();
 sg13g2_decap_8 FILLER_48_77 ();
 sg13g2_decap_8 FILLER_48_84 ();
 sg13g2_decap_8 FILLER_48_91 ();
 sg13g2_decap_8 FILLER_48_98 ();
 sg13g2_decap_8 FILLER_48_105 ();
 sg13g2_decap_8 FILLER_48_112 ();
 sg13g2_decap_8 FILLER_48_119 ();
 sg13g2_decap_8 FILLER_48_126 ();
 sg13g2_decap_8 FILLER_48_133 ();
 sg13g2_decap_8 FILLER_48_140 ();
 sg13g2_decap_8 FILLER_48_147 ();
 sg13g2_decap_8 FILLER_48_154 ();
 sg13g2_decap_8 FILLER_48_161 ();
 sg13g2_decap_8 FILLER_48_168 ();
 sg13g2_decap_8 FILLER_48_175 ();
 sg13g2_decap_8 FILLER_48_182 ();
 sg13g2_decap_8 FILLER_48_189 ();
 sg13g2_decap_8 FILLER_48_196 ();
 sg13g2_decap_8 FILLER_48_203 ();
 sg13g2_decap_8 FILLER_48_210 ();
 sg13g2_decap_8 FILLER_48_217 ();
 sg13g2_decap_8 FILLER_48_224 ();
 sg13g2_decap_8 FILLER_48_231 ();
 sg13g2_decap_8 FILLER_48_238 ();
 sg13g2_decap_8 FILLER_48_245 ();
 sg13g2_decap_8 FILLER_48_252 ();
 sg13g2_decap_8 FILLER_48_259 ();
 sg13g2_decap_8 FILLER_48_266 ();
 sg13g2_decap_8 FILLER_48_273 ();
 sg13g2_decap_8 FILLER_48_280 ();
 sg13g2_decap_8 FILLER_48_287 ();
 sg13g2_decap_8 FILLER_48_294 ();
 sg13g2_decap_8 FILLER_48_301 ();
 sg13g2_decap_8 FILLER_48_308 ();
 sg13g2_decap_8 FILLER_48_315 ();
 sg13g2_decap_8 FILLER_48_322 ();
 sg13g2_decap_8 FILLER_48_329 ();
 sg13g2_decap_8 FILLER_48_336 ();
 sg13g2_decap_8 FILLER_48_343 ();
 sg13g2_decap_8 FILLER_48_350 ();
 sg13g2_decap_8 FILLER_48_357 ();
 sg13g2_decap_8 FILLER_48_364 ();
 sg13g2_decap_8 FILLER_48_371 ();
 sg13g2_decap_8 FILLER_48_378 ();
 sg13g2_decap_8 FILLER_48_385 ();
 sg13g2_decap_8 FILLER_48_392 ();
 sg13g2_decap_8 FILLER_48_399 ();
 sg13g2_decap_8 FILLER_48_406 ();
 sg13g2_decap_8 FILLER_48_413 ();
 sg13g2_decap_8 FILLER_48_420 ();
 sg13g2_decap_8 FILLER_48_427 ();
 sg13g2_decap_8 FILLER_48_434 ();
 sg13g2_decap_8 FILLER_48_441 ();
 sg13g2_decap_8 FILLER_48_448 ();
 sg13g2_decap_8 FILLER_48_455 ();
 sg13g2_decap_8 FILLER_48_462 ();
 sg13g2_decap_8 FILLER_48_469 ();
 sg13g2_decap_8 FILLER_48_476 ();
 sg13g2_decap_8 FILLER_48_483 ();
 sg13g2_decap_8 FILLER_48_490 ();
 sg13g2_decap_8 FILLER_48_497 ();
 sg13g2_decap_8 FILLER_48_504 ();
 sg13g2_decap_8 FILLER_48_511 ();
 sg13g2_decap_8 FILLER_48_518 ();
 sg13g2_decap_8 FILLER_48_525 ();
 sg13g2_decap_8 FILLER_48_532 ();
 sg13g2_decap_8 FILLER_48_539 ();
 sg13g2_decap_8 FILLER_48_546 ();
 sg13g2_decap_8 FILLER_48_553 ();
 sg13g2_decap_8 FILLER_48_560 ();
 sg13g2_decap_8 FILLER_48_567 ();
 sg13g2_decap_8 FILLER_48_574 ();
 sg13g2_decap_8 FILLER_48_581 ();
 sg13g2_decap_8 FILLER_48_588 ();
 sg13g2_decap_8 FILLER_48_595 ();
 sg13g2_decap_8 FILLER_48_602 ();
 sg13g2_decap_8 FILLER_48_609 ();
 sg13g2_decap_8 FILLER_48_616 ();
 sg13g2_decap_8 FILLER_48_623 ();
 sg13g2_decap_8 FILLER_48_630 ();
 sg13g2_decap_8 FILLER_48_637 ();
 sg13g2_decap_8 FILLER_48_644 ();
 sg13g2_decap_8 FILLER_48_651 ();
 sg13g2_decap_8 FILLER_48_658 ();
 sg13g2_decap_8 FILLER_48_665 ();
 sg13g2_decap_8 FILLER_48_672 ();
 sg13g2_decap_8 FILLER_48_679 ();
 sg13g2_decap_8 FILLER_48_686 ();
 sg13g2_decap_8 FILLER_48_693 ();
 sg13g2_decap_8 FILLER_48_700 ();
 sg13g2_decap_8 FILLER_48_707 ();
 sg13g2_decap_8 FILLER_48_714 ();
 sg13g2_decap_8 FILLER_48_721 ();
 sg13g2_decap_8 FILLER_48_728 ();
 sg13g2_decap_8 FILLER_48_735 ();
 sg13g2_decap_8 FILLER_48_742 ();
 sg13g2_decap_8 FILLER_48_749 ();
 sg13g2_decap_8 FILLER_48_756 ();
 sg13g2_decap_8 FILLER_48_763 ();
 sg13g2_decap_8 FILLER_48_770 ();
 sg13g2_decap_8 FILLER_48_777 ();
 sg13g2_decap_8 FILLER_48_784 ();
 sg13g2_decap_8 FILLER_48_791 ();
 sg13g2_decap_8 FILLER_48_798 ();
 sg13g2_decap_8 FILLER_48_805 ();
 sg13g2_decap_8 FILLER_48_812 ();
 sg13g2_decap_8 FILLER_48_819 ();
 sg13g2_decap_8 FILLER_48_826 ();
 sg13g2_decap_8 FILLER_48_833 ();
 sg13g2_decap_8 FILLER_48_840 ();
 sg13g2_decap_8 FILLER_48_847 ();
 sg13g2_decap_8 FILLER_48_854 ();
 sg13g2_decap_8 FILLER_48_861 ();
 sg13g2_decap_8 FILLER_48_868 ();
 sg13g2_decap_8 FILLER_48_875 ();
 sg13g2_decap_8 FILLER_48_882 ();
 sg13g2_decap_8 FILLER_48_889 ();
 sg13g2_decap_8 FILLER_48_896 ();
 sg13g2_decap_8 FILLER_48_903 ();
 sg13g2_decap_8 FILLER_48_910 ();
 sg13g2_decap_8 FILLER_48_917 ();
 sg13g2_decap_8 FILLER_48_924 ();
 sg13g2_decap_8 FILLER_48_931 ();
 sg13g2_decap_8 FILLER_48_938 ();
 sg13g2_decap_8 FILLER_48_945 ();
 sg13g2_decap_8 FILLER_48_952 ();
 sg13g2_decap_8 FILLER_48_959 ();
 sg13g2_decap_8 FILLER_48_966 ();
 sg13g2_decap_8 FILLER_48_973 ();
 sg13g2_decap_8 FILLER_48_980 ();
 sg13g2_decap_8 FILLER_48_987 ();
 sg13g2_decap_8 FILLER_48_994 ();
 sg13g2_decap_8 FILLER_48_1001 ();
 sg13g2_decap_8 FILLER_48_1008 ();
 sg13g2_decap_8 FILLER_48_1015 ();
 sg13g2_decap_8 FILLER_48_1022 ();
 sg13g2_decap_8 FILLER_49_4 ();
 sg13g2_decap_8 FILLER_49_11 ();
 sg13g2_decap_8 FILLER_49_18 ();
 sg13g2_decap_8 FILLER_49_25 ();
 sg13g2_decap_8 FILLER_49_32 ();
 sg13g2_decap_8 FILLER_49_39 ();
 sg13g2_decap_8 FILLER_49_46 ();
 sg13g2_decap_8 FILLER_49_53 ();
 sg13g2_decap_8 FILLER_49_60 ();
 sg13g2_decap_8 FILLER_49_67 ();
 sg13g2_decap_8 FILLER_49_74 ();
 sg13g2_decap_8 FILLER_49_81 ();
 sg13g2_decap_8 FILLER_49_88 ();
 sg13g2_decap_8 FILLER_49_95 ();
 sg13g2_decap_8 FILLER_49_102 ();
 sg13g2_decap_8 FILLER_49_109 ();
 sg13g2_decap_8 FILLER_49_116 ();
 sg13g2_decap_8 FILLER_49_123 ();
 sg13g2_decap_8 FILLER_49_130 ();
 sg13g2_decap_8 FILLER_49_137 ();
 sg13g2_decap_8 FILLER_49_144 ();
 sg13g2_decap_8 FILLER_49_151 ();
 sg13g2_decap_8 FILLER_49_158 ();
 sg13g2_decap_8 FILLER_49_165 ();
 sg13g2_decap_8 FILLER_49_172 ();
 sg13g2_decap_8 FILLER_49_179 ();
 sg13g2_decap_8 FILLER_49_186 ();
 sg13g2_decap_8 FILLER_49_193 ();
 sg13g2_decap_8 FILLER_49_200 ();
 sg13g2_decap_8 FILLER_49_207 ();
 sg13g2_decap_8 FILLER_49_214 ();
 sg13g2_decap_8 FILLER_49_221 ();
 sg13g2_decap_8 FILLER_49_228 ();
 sg13g2_decap_8 FILLER_49_235 ();
 sg13g2_decap_8 FILLER_49_242 ();
 sg13g2_decap_8 FILLER_49_249 ();
 sg13g2_decap_8 FILLER_49_256 ();
 sg13g2_decap_8 FILLER_49_263 ();
 sg13g2_decap_8 FILLER_49_270 ();
 sg13g2_decap_8 FILLER_49_277 ();
 sg13g2_decap_8 FILLER_49_284 ();
 sg13g2_decap_8 FILLER_49_291 ();
 sg13g2_decap_8 FILLER_49_298 ();
 sg13g2_decap_8 FILLER_49_305 ();
 sg13g2_decap_8 FILLER_49_312 ();
 sg13g2_decap_8 FILLER_49_319 ();
 sg13g2_decap_8 FILLER_49_326 ();
 sg13g2_decap_8 FILLER_49_333 ();
 sg13g2_decap_8 FILLER_49_340 ();
 sg13g2_decap_8 FILLER_49_347 ();
 sg13g2_decap_8 FILLER_49_354 ();
 sg13g2_decap_8 FILLER_49_361 ();
 sg13g2_decap_8 FILLER_49_368 ();
 sg13g2_decap_8 FILLER_49_375 ();
 sg13g2_decap_8 FILLER_49_382 ();
 sg13g2_decap_8 FILLER_49_389 ();
 sg13g2_decap_8 FILLER_49_396 ();
 sg13g2_decap_8 FILLER_49_403 ();
 sg13g2_decap_8 FILLER_49_410 ();
 sg13g2_decap_8 FILLER_49_417 ();
 sg13g2_decap_8 FILLER_49_424 ();
 sg13g2_decap_8 FILLER_49_431 ();
 sg13g2_decap_8 FILLER_49_438 ();
 sg13g2_decap_8 FILLER_49_445 ();
 sg13g2_decap_8 FILLER_49_452 ();
 sg13g2_decap_8 FILLER_49_459 ();
 sg13g2_decap_8 FILLER_49_466 ();
 sg13g2_decap_8 FILLER_49_473 ();
 sg13g2_decap_8 FILLER_49_480 ();
 sg13g2_decap_8 FILLER_49_487 ();
 sg13g2_decap_8 FILLER_49_494 ();
 sg13g2_decap_8 FILLER_49_501 ();
 sg13g2_decap_8 FILLER_49_508 ();
 sg13g2_decap_8 FILLER_49_515 ();
 sg13g2_decap_8 FILLER_49_522 ();
 sg13g2_decap_8 FILLER_49_529 ();
 sg13g2_decap_8 FILLER_49_536 ();
 sg13g2_decap_8 FILLER_49_543 ();
 sg13g2_decap_8 FILLER_49_550 ();
 sg13g2_decap_8 FILLER_49_557 ();
 sg13g2_decap_8 FILLER_49_564 ();
 sg13g2_decap_8 FILLER_49_571 ();
 sg13g2_decap_8 FILLER_49_578 ();
 sg13g2_decap_8 FILLER_49_585 ();
 sg13g2_decap_8 FILLER_49_592 ();
 sg13g2_decap_8 FILLER_49_599 ();
 sg13g2_decap_8 FILLER_49_606 ();
 sg13g2_decap_8 FILLER_49_613 ();
 sg13g2_decap_8 FILLER_49_620 ();
 sg13g2_decap_8 FILLER_49_627 ();
 sg13g2_decap_8 FILLER_49_634 ();
 sg13g2_decap_8 FILLER_49_641 ();
 sg13g2_decap_8 FILLER_49_648 ();
 sg13g2_decap_8 FILLER_49_655 ();
 sg13g2_decap_8 FILLER_49_662 ();
 sg13g2_decap_8 FILLER_49_669 ();
 sg13g2_decap_8 FILLER_49_676 ();
 sg13g2_decap_8 FILLER_49_683 ();
 sg13g2_decap_8 FILLER_49_690 ();
 sg13g2_decap_8 FILLER_49_697 ();
 sg13g2_decap_8 FILLER_49_704 ();
 sg13g2_decap_8 FILLER_49_711 ();
 sg13g2_decap_8 FILLER_49_718 ();
 sg13g2_decap_8 FILLER_49_725 ();
 sg13g2_decap_8 FILLER_49_732 ();
 sg13g2_decap_8 FILLER_49_739 ();
 sg13g2_decap_8 FILLER_49_746 ();
 sg13g2_decap_8 FILLER_49_753 ();
 sg13g2_decap_8 FILLER_49_760 ();
 sg13g2_decap_8 FILLER_49_767 ();
 sg13g2_decap_8 FILLER_49_774 ();
 sg13g2_decap_8 FILLER_49_781 ();
 sg13g2_decap_8 FILLER_49_788 ();
 sg13g2_decap_8 FILLER_49_795 ();
 sg13g2_decap_8 FILLER_49_802 ();
 sg13g2_decap_8 FILLER_49_809 ();
 sg13g2_decap_8 FILLER_49_816 ();
 sg13g2_decap_8 FILLER_49_823 ();
 sg13g2_decap_8 FILLER_49_830 ();
 sg13g2_decap_8 FILLER_49_837 ();
 sg13g2_decap_8 FILLER_49_844 ();
 sg13g2_decap_8 FILLER_49_851 ();
 sg13g2_decap_8 FILLER_49_858 ();
 sg13g2_decap_8 FILLER_49_865 ();
 sg13g2_decap_8 FILLER_49_872 ();
 sg13g2_decap_8 FILLER_49_879 ();
 sg13g2_decap_8 FILLER_49_886 ();
 sg13g2_decap_8 FILLER_49_893 ();
 sg13g2_decap_8 FILLER_49_900 ();
 sg13g2_decap_8 FILLER_49_907 ();
 sg13g2_decap_8 FILLER_49_914 ();
 sg13g2_decap_8 FILLER_49_921 ();
 sg13g2_decap_8 FILLER_49_928 ();
 sg13g2_decap_8 FILLER_49_935 ();
 sg13g2_decap_8 FILLER_49_942 ();
 sg13g2_decap_8 FILLER_49_949 ();
 sg13g2_decap_8 FILLER_49_956 ();
 sg13g2_decap_8 FILLER_49_963 ();
 sg13g2_decap_8 FILLER_49_970 ();
 sg13g2_decap_8 FILLER_49_977 ();
 sg13g2_decap_8 FILLER_49_984 ();
 sg13g2_decap_8 FILLER_49_991 ();
 sg13g2_decap_8 FILLER_49_998 ();
 sg13g2_decap_8 FILLER_49_1005 ();
 sg13g2_decap_8 FILLER_49_1012 ();
 sg13g2_decap_8 FILLER_49_1019 ();
 sg13g2_fill_2 FILLER_49_1026 ();
 sg13g2_fill_1 FILLER_49_1028 ();
 sg13g2_decap_8 FILLER_50_0 ();
 sg13g2_decap_8 FILLER_50_7 ();
 sg13g2_decap_8 FILLER_50_14 ();
 sg13g2_decap_8 FILLER_50_21 ();
 sg13g2_decap_8 FILLER_50_28 ();
 sg13g2_decap_8 FILLER_50_35 ();
 sg13g2_decap_8 FILLER_50_42 ();
 sg13g2_decap_8 FILLER_50_49 ();
 sg13g2_decap_8 FILLER_50_56 ();
 sg13g2_decap_8 FILLER_50_63 ();
 sg13g2_decap_8 FILLER_50_70 ();
 sg13g2_decap_8 FILLER_50_77 ();
 sg13g2_decap_8 FILLER_50_84 ();
 sg13g2_decap_8 FILLER_50_91 ();
 sg13g2_decap_8 FILLER_50_98 ();
 sg13g2_decap_8 FILLER_50_105 ();
 sg13g2_decap_8 FILLER_50_112 ();
 sg13g2_decap_8 FILLER_50_119 ();
 sg13g2_decap_8 FILLER_50_126 ();
 sg13g2_decap_8 FILLER_50_133 ();
 sg13g2_decap_8 FILLER_50_140 ();
 sg13g2_decap_8 FILLER_50_147 ();
 sg13g2_decap_8 FILLER_50_154 ();
 sg13g2_decap_8 FILLER_50_161 ();
 sg13g2_decap_8 FILLER_50_168 ();
 sg13g2_decap_8 FILLER_50_175 ();
 sg13g2_decap_8 FILLER_50_182 ();
 sg13g2_decap_8 FILLER_50_189 ();
 sg13g2_decap_8 FILLER_50_196 ();
 sg13g2_decap_8 FILLER_50_203 ();
 sg13g2_decap_8 FILLER_50_210 ();
 sg13g2_decap_8 FILLER_50_217 ();
 sg13g2_decap_8 FILLER_50_224 ();
 sg13g2_decap_8 FILLER_50_231 ();
 sg13g2_decap_8 FILLER_50_238 ();
 sg13g2_decap_8 FILLER_50_245 ();
 sg13g2_decap_8 FILLER_50_252 ();
 sg13g2_decap_8 FILLER_50_259 ();
 sg13g2_decap_8 FILLER_50_266 ();
 sg13g2_decap_8 FILLER_50_273 ();
 sg13g2_decap_8 FILLER_50_280 ();
 sg13g2_decap_8 FILLER_50_287 ();
 sg13g2_decap_8 FILLER_50_294 ();
 sg13g2_decap_8 FILLER_50_301 ();
 sg13g2_decap_8 FILLER_50_308 ();
 sg13g2_decap_8 FILLER_50_315 ();
 sg13g2_decap_8 FILLER_50_322 ();
 sg13g2_decap_8 FILLER_50_329 ();
 sg13g2_decap_8 FILLER_50_336 ();
 sg13g2_decap_8 FILLER_50_343 ();
 sg13g2_decap_8 FILLER_50_350 ();
 sg13g2_decap_8 FILLER_50_357 ();
 sg13g2_decap_8 FILLER_50_364 ();
 sg13g2_decap_8 FILLER_50_371 ();
 sg13g2_decap_8 FILLER_50_378 ();
 sg13g2_decap_8 FILLER_50_385 ();
 sg13g2_decap_8 FILLER_50_392 ();
 sg13g2_decap_8 FILLER_50_399 ();
 sg13g2_decap_8 FILLER_50_406 ();
 sg13g2_decap_8 FILLER_50_413 ();
 sg13g2_decap_8 FILLER_50_420 ();
 sg13g2_decap_8 FILLER_50_427 ();
 sg13g2_decap_8 FILLER_50_434 ();
 sg13g2_decap_8 FILLER_50_441 ();
 sg13g2_decap_8 FILLER_50_448 ();
 sg13g2_decap_8 FILLER_50_455 ();
 sg13g2_decap_8 FILLER_50_462 ();
 sg13g2_decap_8 FILLER_50_469 ();
 sg13g2_decap_8 FILLER_50_476 ();
 sg13g2_decap_8 FILLER_50_483 ();
 sg13g2_decap_8 FILLER_50_490 ();
 sg13g2_decap_8 FILLER_50_497 ();
 sg13g2_decap_8 FILLER_50_504 ();
 sg13g2_decap_8 FILLER_50_511 ();
 sg13g2_decap_8 FILLER_50_518 ();
 sg13g2_decap_8 FILLER_50_525 ();
 sg13g2_decap_8 FILLER_50_532 ();
 sg13g2_decap_8 FILLER_50_539 ();
 sg13g2_decap_8 FILLER_50_546 ();
 sg13g2_decap_8 FILLER_50_553 ();
 sg13g2_decap_8 FILLER_50_560 ();
 sg13g2_decap_8 FILLER_50_567 ();
 sg13g2_decap_8 FILLER_50_574 ();
 sg13g2_decap_8 FILLER_50_581 ();
 sg13g2_decap_8 FILLER_50_588 ();
 sg13g2_decap_8 FILLER_50_595 ();
 sg13g2_decap_8 FILLER_50_602 ();
 sg13g2_decap_8 FILLER_50_609 ();
 sg13g2_decap_8 FILLER_50_616 ();
 sg13g2_decap_8 FILLER_50_623 ();
 sg13g2_decap_8 FILLER_50_630 ();
 sg13g2_decap_8 FILLER_50_637 ();
 sg13g2_decap_8 FILLER_50_644 ();
 sg13g2_decap_8 FILLER_50_651 ();
 sg13g2_decap_8 FILLER_50_658 ();
 sg13g2_decap_8 FILLER_50_665 ();
 sg13g2_decap_8 FILLER_50_672 ();
 sg13g2_decap_8 FILLER_50_679 ();
 sg13g2_decap_8 FILLER_50_686 ();
 sg13g2_decap_8 FILLER_50_693 ();
 sg13g2_decap_8 FILLER_50_700 ();
 sg13g2_decap_8 FILLER_50_707 ();
 sg13g2_decap_8 FILLER_50_714 ();
 sg13g2_decap_8 FILLER_50_721 ();
 sg13g2_decap_8 FILLER_50_728 ();
 sg13g2_decap_8 FILLER_50_735 ();
 sg13g2_decap_8 FILLER_50_742 ();
 sg13g2_decap_8 FILLER_50_749 ();
 sg13g2_decap_8 FILLER_50_756 ();
 sg13g2_decap_8 FILLER_50_763 ();
 sg13g2_decap_8 FILLER_50_770 ();
 sg13g2_decap_8 FILLER_50_777 ();
 sg13g2_decap_8 FILLER_50_784 ();
 sg13g2_decap_8 FILLER_50_791 ();
 sg13g2_decap_8 FILLER_50_798 ();
 sg13g2_decap_8 FILLER_50_805 ();
 sg13g2_decap_8 FILLER_50_812 ();
 sg13g2_decap_8 FILLER_50_819 ();
 sg13g2_decap_8 FILLER_50_826 ();
 sg13g2_decap_8 FILLER_50_833 ();
 sg13g2_decap_8 FILLER_50_840 ();
 sg13g2_decap_8 FILLER_50_847 ();
 sg13g2_decap_8 FILLER_50_854 ();
 sg13g2_decap_8 FILLER_50_861 ();
 sg13g2_decap_8 FILLER_50_868 ();
 sg13g2_decap_8 FILLER_50_875 ();
 sg13g2_decap_8 FILLER_50_882 ();
 sg13g2_decap_8 FILLER_50_889 ();
 sg13g2_decap_8 FILLER_50_896 ();
 sg13g2_decap_8 FILLER_50_903 ();
 sg13g2_decap_8 FILLER_50_910 ();
 sg13g2_decap_8 FILLER_50_917 ();
 sg13g2_decap_8 FILLER_50_924 ();
 sg13g2_decap_8 FILLER_50_931 ();
 sg13g2_decap_8 FILLER_50_938 ();
 sg13g2_decap_8 FILLER_50_945 ();
 sg13g2_decap_8 FILLER_50_952 ();
 sg13g2_decap_8 FILLER_50_959 ();
 sg13g2_decap_8 FILLER_50_966 ();
 sg13g2_decap_8 FILLER_50_973 ();
 sg13g2_decap_8 FILLER_50_980 ();
 sg13g2_decap_8 FILLER_50_987 ();
 sg13g2_decap_8 FILLER_50_994 ();
 sg13g2_decap_8 FILLER_50_1001 ();
 sg13g2_decap_8 FILLER_50_1008 ();
 sg13g2_decap_8 FILLER_50_1015 ();
 sg13g2_decap_8 FILLER_50_1022 ();
 sg13g2_decap_8 FILLER_51_4 ();
 sg13g2_decap_8 FILLER_51_11 ();
 sg13g2_decap_8 FILLER_51_18 ();
 sg13g2_decap_8 FILLER_51_25 ();
 sg13g2_decap_8 FILLER_51_32 ();
 sg13g2_decap_8 FILLER_51_39 ();
 sg13g2_decap_8 FILLER_51_46 ();
 sg13g2_decap_8 FILLER_51_53 ();
 sg13g2_decap_8 FILLER_51_60 ();
 sg13g2_decap_8 FILLER_51_67 ();
 sg13g2_decap_8 FILLER_51_74 ();
 sg13g2_decap_8 FILLER_51_81 ();
 sg13g2_decap_8 FILLER_51_88 ();
 sg13g2_decap_8 FILLER_51_95 ();
 sg13g2_decap_8 FILLER_51_102 ();
 sg13g2_decap_8 FILLER_51_109 ();
 sg13g2_decap_8 FILLER_51_116 ();
 sg13g2_decap_8 FILLER_51_123 ();
 sg13g2_decap_8 FILLER_51_130 ();
 sg13g2_decap_8 FILLER_51_137 ();
 sg13g2_decap_8 FILLER_51_144 ();
 sg13g2_decap_8 FILLER_51_151 ();
 sg13g2_decap_8 FILLER_51_158 ();
 sg13g2_decap_8 FILLER_51_165 ();
 sg13g2_decap_8 FILLER_51_172 ();
 sg13g2_decap_8 FILLER_51_179 ();
 sg13g2_decap_8 FILLER_51_186 ();
 sg13g2_decap_8 FILLER_51_193 ();
 sg13g2_decap_8 FILLER_51_200 ();
 sg13g2_decap_8 FILLER_51_207 ();
 sg13g2_decap_8 FILLER_51_214 ();
 sg13g2_decap_8 FILLER_51_221 ();
 sg13g2_decap_8 FILLER_51_228 ();
 sg13g2_decap_8 FILLER_51_235 ();
 sg13g2_decap_8 FILLER_51_242 ();
 sg13g2_decap_8 FILLER_51_249 ();
 sg13g2_decap_8 FILLER_51_256 ();
 sg13g2_decap_8 FILLER_51_263 ();
 sg13g2_decap_8 FILLER_51_270 ();
 sg13g2_decap_8 FILLER_51_277 ();
 sg13g2_decap_8 FILLER_51_284 ();
 sg13g2_decap_8 FILLER_51_291 ();
 sg13g2_decap_8 FILLER_51_298 ();
 sg13g2_decap_8 FILLER_51_305 ();
 sg13g2_decap_8 FILLER_51_312 ();
 sg13g2_decap_8 FILLER_51_319 ();
 sg13g2_decap_8 FILLER_51_326 ();
 sg13g2_decap_8 FILLER_51_333 ();
 sg13g2_decap_8 FILLER_51_340 ();
 sg13g2_decap_8 FILLER_51_347 ();
 sg13g2_decap_8 FILLER_51_354 ();
 sg13g2_decap_8 FILLER_51_361 ();
 sg13g2_decap_8 FILLER_51_368 ();
 sg13g2_decap_8 FILLER_51_375 ();
 sg13g2_decap_8 FILLER_51_382 ();
 sg13g2_decap_8 FILLER_51_389 ();
 sg13g2_decap_8 FILLER_51_396 ();
 sg13g2_decap_8 FILLER_51_403 ();
 sg13g2_decap_8 FILLER_51_410 ();
 sg13g2_decap_8 FILLER_51_417 ();
 sg13g2_decap_8 FILLER_51_424 ();
 sg13g2_decap_8 FILLER_51_431 ();
 sg13g2_decap_8 FILLER_51_438 ();
 sg13g2_decap_8 FILLER_51_445 ();
 sg13g2_decap_8 FILLER_51_452 ();
 sg13g2_decap_8 FILLER_51_459 ();
 sg13g2_decap_8 FILLER_51_466 ();
 sg13g2_decap_8 FILLER_51_473 ();
 sg13g2_decap_8 FILLER_51_480 ();
 sg13g2_decap_8 FILLER_51_487 ();
 sg13g2_decap_8 FILLER_51_494 ();
 sg13g2_decap_8 FILLER_51_501 ();
 sg13g2_decap_8 FILLER_51_508 ();
 sg13g2_decap_8 FILLER_51_515 ();
 sg13g2_decap_8 FILLER_51_522 ();
 sg13g2_decap_8 FILLER_51_529 ();
 sg13g2_decap_8 FILLER_51_536 ();
 sg13g2_decap_8 FILLER_51_543 ();
 sg13g2_decap_8 FILLER_51_550 ();
 sg13g2_decap_8 FILLER_51_557 ();
 sg13g2_decap_8 FILLER_51_564 ();
 sg13g2_decap_8 FILLER_51_571 ();
 sg13g2_decap_8 FILLER_51_578 ();
 sg13g2_decap_8 FILLER_51_585 ();
 sg13g2_decap_8 FILLER_51_592 ();
 sg13g2_decap_8 FILLER_51_599 ();
 sg13g2_decap_8 FILLER_51_606 ();
 sg13g2_decap_8 FILLER_51_613 ();
 sg13g2_decap_8 FILLER_51_620 ();
 sg13g2_decap_8 FILLER_51_627 ();
 sg13g2_decap_8 FILLER_51_634 ();
 sg13g2_decap_8 FILLER_51_641 ();
 sg13g2_decap_8 FILLER_51_648 ();
 sg13g2_decap_8 FILLER_51_655 ();
 sg13g2_decap_8 FILLER_51_662 ();
 sg13g2_decap_8 FILLER_51_669 ();
 sg13g2_decap_8 FILLER_51_676 ();
 sg13g2_decap_8 FILLER_51_683 ();
 sg13g2_decap_8 FILLER_51_690 ();
 sg13g2_decap_8 FILLER_51_697 ();
 sg13g2_decap_8 FILLER_51_704 ();
 sg13g2_decap_8 FILLER_51_711 ();
 sg13g2_decap_8 FILLER_51_718 ();
 sg13g2_decap_8 FILLER_51_725 ();
 sg13g2_decap_8 FILLER_51_732 ();
 sg13g2_decap_8 FILLER_51_739 ();
 sg13g2_decap_8 FILLER_51_746 ();
 sg13g2_decap_8 FILLER_51_753 ();
 sg13g2_decap_8 FILLER_51_760 ();
 sg13g2_decap_8 FILLER_51_767 ();
 sg13g2_decap_8 FILLER_51_774 ();
 sg13g2_decap_8 FILLER_51_781 ();
 sg13g2_decap_8 FILLER_51_788 ();
 sg13g2_decap_8 FILLER_51_795 ();
 sg13g2_decap_8 FILLER_51_802 ();
 sg13g2_decap_8 FILLER_51_809 ();
 sg13g2_decap_8 FILLER_51_816 ();
 sg13g2_decap_8 FILLER_51_823 ();
 sg13g2_decap_8 FILLER_51_830 ();
 sg13g2_decap_8 FILLER_51_837 ();
 sg13g2_decap_8 FILLER_51_844 ();
 sg13g2_decap_8 FILLER_51_851 ();
 sg13g2_decap_8 FILLER_51_858 ();
 sg13g2_decap_8 FILLER_51_865 ();
 sg13g2_decap_8 FILLER_51_872 ();
 sg13g2_decap_8 FILLER_51_879 ();
 sg13g2_decap_8 FILLER_51_886 ();
 sg13g2_decap_8 FILLER_51_893 ();
 sg13g2_decap_8 FILLER_51_900 ();
 sg13g2_decap_8 FILLER_51_907 ();
 sg13g2_decap_8 FILLER_51_914 ();
 sg13g2_decap_8 FILLER_51_921 ();
 sg13g2_decap_8 FILLER_51_928 ();
 sg13g2_decap_8 FILLER_51_935 ();
 sg13g2_decap_8 FILLER_51_942 ();
 sg13g2_decap_8 FILLER_51_949 ();
 sg13g2_decap_8 FILLER_51_956 ();
 sg13g2_decap_8 FILLER_51_963 ();
 sg13g2_decap_8 FILLER_51_970 ();
 sg13g2_decap_8 FILLER_51_977 ();
 sg13g2_decap_8 FILLER_51_984 ();
 sg13g2_decap_8 FILLER_51_991 ();
 sg13g2_decap_8 FILLER_51_998 ();
 sg13g2_decap_8 FILLER_51_1005 ();
 sg13g2_decap_8 FILLER_51_1012 ();
 sg13g2_decap_8 FILLER_51_1019 ();
 sg13g2_fill_2 FILLER_51_1026 ();
 sg13g2_fill_1 FILLER_51_1028 ();
 sg13g2_decap_8 FILLER_52_0 ();
 sg13g2_decap_8 FILLER_52_7 ();
 sg13g2_decap_8 FILLER_52_14 ();
 sg13g2_decap_8 FILLER_52_21 ();
 sg13g2_decap_8 FILLER_52_28 ();
 sg13g2_decap_8 FILLER_52_35 ();
 sg13g2_decap_8 FILLER_52_42 ();
 sg13g2_decap_8 FILLER_52_49 ();
 sg13g2_decap_8 FILLER_52_56 ();
 sg13g2_decap_8 FILLER_52_63 ();
 sg13g2_decap_8 FILLER_52_70 ();
 sg13g2_decap_8 FILLER_52_77 ();
 sg13g2_decap_8 FILLER_52_84 ();
 sg13g2_decap_8 FILLER_52_91 ();
 sg13g2_decap_8 FILLER_52_98 ();
 sg13g2_decap_8 FILLER_52_105 ();
 sg13g2_decap_8 FILLER_52_112 ();
 sg13g2_decap_8 FILLER_52_119 ();
 sg13g2_decap_8 FILLER_52_126 ();
 sg13g2_decap_8 FILLER_52_133 ();
 sg13g2_decap_8 FILLER_52_140 ();
 sg13g2_decap_8 FILLER_52_147 ();
 sg13g2_decap_8 FILLER_52_154 ();
 sg13g2_decap_8 FILLER_52_161 ();
 sg13g2_decap_8 FILLER_52_168 ();
 sg13g2_decap_8 FILLER_52_175 ();
 sg13g2_decap_8 FILLER_52_182 ();
 sg13g2_decap_8 FILLER_52_189 ();
 sg13g2_decap_8 FILLER_52_196 ();
 sg13g2_decap_8 FILLER_52_203 ();
 sg13g2_decap_8 FILLER_52_210 ();
 sg13g2_decap_8 FILLER_52_217 ();
 sg13g2_decap_8 FILLER_52_224 ();
 sg13g2_decap_8 FILLER_52_231 ();
 sg13g2_decap_8 FILLER_52_238 ();
 sg13g2_decap_8 FILLER_52_245 ();
 sg13g2_decap_8 FILLER_52_252 ();
 sg13g2_decap_8 FILLER_52_259 ();
 sg13g2_decap_8 FILLER_52_266 ();
 sg13g2_decap_8 FILLER_52_273 ();
 sg13g2_decap_8 FILLER_52_280 ();
 sg13g2_decap_8 FILLER_52_287 ();
 sg13g2_decap_8 FILLER_52_294 ();
 sg13g2_decap_8 FILLER_52_301 ();
 sg13g2_decap_8 FILLER_52_308 ();
 sg13g2_decap_8 FILLER_52_315 ();
 sg13g2_decap_8 FILLER_52_322 ();
 sg13g2_decap_8 FILLER_52_329 ();
 sg13g2_decap_8 FILLER_52_336 ();
 sg13g2_decap_8 FILLER_52_343 ();
 sg13g2_decap_8 FILLER_52_350 ();
 sg13g2_decap_8 FILLER_52_357 ();
 sg13g2_decap_8 FILLER_52_364 ();
 sg13g2_decap_8 FILLER_52_371 ();
 sg13g2_decap_8 FILLER_52_378 ();
 sg13g2_decap_8 FILLER_52_385 ();
 sg13g2_decap_8 FILLER_52_392 ();
 sg13g2_decap_8 FILLER_52_399 ();
 sg13g2_decap_8 FILLER_52_406 ();
 sg13g2_decap_8 FILLER_52_413 ();
 sg13g2_decap_8 FILLER_52_420 ();
 sg13g2_decap_8 FILLER_52_427 ();
 sg13g2_decap_8 FILLER_52_434 ();
 sg13g2_decap_8 FILLER_52_441 ();
 sg13g2_decap_8 FILLER_52_448 ();
 sg13g2_decap_8 FILLER_52_455 ();
 sg13g2_decap_8 FILLER_52_462 ();
 sg13g2_decap_8 FILLER_52_469 ();
 sg13g2_decap_8 FILLER_52_476 ();
 sg13g2_decap_8 FILLER_52_483 ();
 sg13g2_decap_8 FILLER_52_490 ();
 sg13g2_decap_8 FILLER_52_497 ();
 sg13g2_decap_8 FILLER_52_504 ();
 sg13g2_decap_8 FILLER_52_511 ();
 sg13g2_decap_8 FILLER_52_518 ();
 sg13g2_decap_8 FILLER_52_525 ();
 sg13g2_decap_8 FILLER_52_532 ();
 sg13g2_decap_8 FILLER_52_539 ();
 sg13g2_decap_8 FILLER_52_546 ();
 sg13g2_decap_8 FILLER_52_553 ();
 sg13g2_decap_8 FILLER_52_560 ();
 sg13g2_decap_8 FILLER_52_567 ();
 sg13g2_decap_8 FILLER_52_574 ();
 sg13g2_decap_8 FILLER_52_581 ();
 sg13g2_decap_8 FILLER_52_588 ();
 sg13g2_decap_8 FILLER_52_595 ();
 sg13g2_decap_8 FILLER_52_602 ();
 sg13g2_decap_8 FILLER_52_609 ();
 sg13g2_decap_8 FILLER_52_616 ();
 sg13g2_decap_8 FILLER_52_623 ();
 sg13g2_decap_8 FILLER_52_630 ();
 sg13g2_decap_8 FILLER_52_637 ();
 sg13g2_decap_8 FILLER_52_644 ();
 sg13g2_decap_8 FILLER_52_651 ();
 sg13g2_decap_8 FILLER_52_658 ();
 sg13g2_decap_8 FILLER_52_665 ();
 sg13g2_decap_8 FILLER_52_672 ();
 sg13g2_decap_8 FILLER_52_679 ();
 sg13g2_decap_8 FILLER_52_686 ();
 sg13g2_decap_8 FILLER_52_693 ();
 sg13g2_decap_8 FILLER_52_700 ();
 sg13g2_decap_8 FILLER_52_707 ();
 sg13g2_decap_8 FILLER_52_714 ();
 sg13g2_decap_8 FILLER_52_721 ();
 sg13g2_decap_8 FILLER_52_728 ();
 sg13g2_decap_8 FILLER_52_735 ();
 sg13g2_decap_8 FILLER_52_742 ();
 sg13g2_decap_8 FILLER_52_749 ();
 sg13g2_decap_8 FILLER_52_756 ();
 sg13g2_decap_8 FILLER_52_763 ();
 sg13g2_decap_8 FILLER_52_770 ();
 sg13g2_decap_8 FILLER_52_777 ();
 sg13g2_decap_8 FILLER_52_784 ();
 sg13g2_decap_8 FILLER_52_791 ();
 sg13g2_decap_8 FILLER_52_798 ();
 sg13g2_decap_8 FILLER_52_805 ();
 sg13g2_decap_8 FILLER_52_812 ();
 sg13g2_decap_8 FILLER_52_819 ();
 sg13g2_decap_8 FILLER_52_826 ();
 sg13g2_decap_8 FILLER_52_833 ();
 sg13g2_decap_8 FILLER_52_840 ();
 sg13g2_decap_8 FILLER_52_847 ();
 sg13g2_decap_8 FILLER_52_854 ();
 sg13g2_decap_8 FILLER_52_861 ();
 sg13g2_decap_8 FILLER_52_868 ();
 sg13g2_decap_8 FILLER_52_875 ();
 sg13g2_decap_8 FILLER_52_882 ();
 sg13g2_decap_8 FILLER_52_889 ();
 sg13g2_decap_8 FILLER_52_896 ();
 sg13g2_decap_8 FILLER_52_903 ();
 sg13g2_decap_8 FILLER_52_910 ();
 sg13g2_decap_8 FILLER_52_917 ();
 sg13g2_decap_8 FILLER_52_924 ();
 sg13g2_decap_8 FILLER_52_931 ();
 sg13g2_decap_8 FILLER_52_938 ();
 sg13g2_decap_8 FILLER_52_945 ();
 sg13g2_decap_8 FILLER_52_952 ();
 sg13g2_decap_8 FILLER_52_959 ();
 sg13g2_decap_8 FILLER_52_966 ();
 sg13g2_decap_8 FILLER_52_973 ();
 sg13g2_decap_8 FILLER_52_980 ();
 sg13g2_decap_8 FILLER_52_987 ();
 sg13g2_decap_8 FILLER_52_994 ();
 sg13g2_decap_8 FILLER_52_1001 ();
 sg13g2_decap_8 FILLER_52_1008 ();
 sg13g2_decap_8 FILLER_52_1015 ();
 sg13g2_decap_8 FILLER_52_1022 ();
 sg13g2_decap_8 FILLER_53_0 ();
 sg13g2_decap_8 FILLER_53_7 ();
 sg13g2_decap_8 FILLER_53_14 ();
 sg13g2_decap_8 FILLER_53_21 ();
 sg13g2_decap_8 FILLER_53_28 ();
 sg13g2_decap_8 FILLER_53_35 ();
 sg13g2_decap_8 FILLER_53_42 ();
 sg13g2_decap_8 FILLER_53_49 ();
 sg13g2_decap_8 FILLER_53_56 ();
 sg13g2_decap_8 FILLER_53_63 ();
 sg13g2_decap_8 FILLER_53_70 ();
 sg13g2_decap_8 FILLER_53_77 ();
 sg13g2_decap_8 FILLER_53_84 ();
 sg13g2_decap_8 FILLER_53_91 ();
 sg13g2_decap_8 FILLER_53_98 ();
 sg13g2_decap_8 FILLER_53_105 ();
 sg13g2_decap_8 FILLER_53_112 ();
 sg13g2_decap_8 FILLER_53_119 ();
 sg13g2_decap_8 FILLER_53_126 ();
 sg13g2_decap_8 FILLER_53_133 ();
 sg13g2_decap_8 FILLER_53_140 ();
 sg13g2_decap_8 FILLER_53_147 ();
 sg13g2_decap_8 FILLER_53_154 ();
 sg13g2_decap_8 FILLER_53_161 ();
 sg13g2_decap_8 FILLER_53_168 ();
 sg13g2_decap_8 FILLER_53_175 ();
 sg13g2_decap_8 FILLER_53_182 ();
 sg13g2_decap_8 FILLER_53_189 ();
 sg13g2_decap_8 FILLER_53_196 ();
 sg13g2_decap_8 FILLER_53_203 ();
 sg13g2_decap_8 FILLER_53_210 ();
 sg13g2_decap_8 FILLER_53_217 ();
 sg13g2_decap_8 FILLER_53_224 ();
 sg13g2_decap_8 FILLER_53_231 ();
 sg13g2_decap_8 FILLER_53_238 ();
 sg13g2_decap_8 FILLER_53_245 ();
 sg13g2_decap_8 FILLER_53_252 ();
 sg13g2_decap_8 FILLER_53_259 ();
 sg13g2_decap_8 FILLER_53_266 ();
 sg13g2_decap_8 FILLER_53_273 ();
 sg13g2_decap_8 FILLER_53_280 ();
 sg13g2_decap_8 FILLER_53_287 ();
 sg13g2_decap_8 FILLER_53_294 ();
 sg13g2_decap_8 FILLER_53_301 ();
 sg13g2_decap_8 FILLER_53_308 ();
 sg13g2_decap_8 FILLER_53_315 ();
 sg13g2_decap_8 FILLER_53_322 ();
 sg13g2_decap_8 FILLER_53_329 ();
 sg13g2_decap_8 FILLER_53_336 ();
 sg13g2_decap_8 FILLER_53_343 ();
 sg13g2_decap_8 FILLER_53_350 ();
 sg13g2_decap_8 FILLER_53_357 ();
 sg13g2_decap_8 FILLER_53_364 ();
 sg13g2_decap_8 FILLER_53_371 ();
 sg13g2_decap_8 FILLER_53_378 ();
 sg13g2_decap_8 FILLER_53_385 ();
 sg13g2_decap_8 FILLER_53_392 ();
 sg13g2_decap_8 FILLER_53_399 ();
 sg13g2_decap_8 FILLER_53_406 ();
 sg13g2_decap_8 FILLER_53_413 ();
 sg13g2_decap_8 FILLER_53_420 ();
 sg13g2_decap_8 FILLER_53_427 ();
 sg13g2_decap_8 FILLER_53_434 ();
 sg13g2_decap_8 FILLER_53_441 ();
 sg13g2_decap_8 FILLER_53_448 ();
 sg13g2_decap_8 FILLER_53_455 ();
 sg13g2_decap_8 FILLER_53_462 ();
 sg13g2_decap_8 FILLER_53_469 ();
 sg13g2_decap_8 FILLER_53_476 ();
 sg13g2_decap_8 FILLER_53_483 ();
 sg13g2_decap_8 FILLER_53_490 ();
 sg13g2_decap_8 FILLER_53_497 ();
 sg13g2_decap_8 FILLER_53_504 ();
 sg13g2_decap_8 FILLER_53_511 ();
 sg13g2_decap_8 FILLER_53_518 ();
 sg13g2_decap_8 FILLER_53_525 ();
 sg13g2_decap_8 FILLER_53_532 ();
 sg13g2_decap_8 FILLER_53_539 ();
 sg13g2_decap_8 FILLER_53_546 ();
 sg13g2_decap_8 FILLER_53_553 ();
 sg13g2_decap_8 FILLER_53_560 ();
 sg13g2_decap_8 FILLER_53_567 ();
 sg13g2_decap_8 FILLER_53_574 ();
 sg13g2_decap_8 FILLER_53_581 ();
 sg13g2_decap_8 FILLER_53_588 ();
 sg13g2_decap_8 FILLER_53_595 ();
 sg13g2_decap_8 FILLER_53_602 ();
 sg13g2_decap_8 FILLER_53_609 ();
 sg13g2_decap_8 FILLER_53_616 ();
 sg13g2_decap_8 FILLER_53_623 ();
 sg13g2_decap_8 FILLER_53_630 ();
 sg13g2_decap_8 FILLER_53_637 ();
 sg13g2_decap_8 FILLER_53_644 ();
 sg13g2_decap_8 FILLER_53_651 ();
 sg13g2_decap_8 FILLER_53_658 ();
 sg13g2_decap_8 FILLER_53_665 ();
 sg13g2_decap_8 FILLER_53_672 ();
 sg13g2_decap_8 FILLER_53_679 ();
 sg13g2_decap_8 FILLER_53_686 ();
 sg13g2_decap_8 FILLER_53_693 ();
 sg13g2_decap_8 FILLER_53_700 ();
 sg13g2_decap_8 FILLER_53_707 ();
 sg13g2_decap_8 FILLER_53_714 ();
 sg13g2_decap_8 FILLER_53_721 ();
 sg13g2_decap_8 FILLER_53_728 ();
 sg13g2_decap_8 FILLER_53_735 ();
 sg13g2_decap_8 FILLER_53_742 ();
 sg13g2_decap_8 FILLER_53_749 ();
 sg13g2_decap_8 FILLER_53_756 ();
 sg13g2_decap_8 FILLER_53_763 ();
 sg13g2_decap_8 FILLER_53_770 ();
 sg13g2_decap_8 FILLER_53_777 ();
 sg13g2_decap_8 FILLER_53_784 ();
 sg13g2_decap_8 FILLER_53_791 ();
 sg13g2_decap_8 FILLER_53_798 ();
 sg13g2_decap_8 FILLER_53_805 ();
 sg13g2_decap_8 FILLER_53_812 ();
 sg13g2_decap_8 FILLER_53_819 ();
 sg13g2_decap_8 FILLER_53_826 ();
 sg13g2_decap_8 FILLER_53_833 ();
 sg13g2_decap_8 FILLER_53_840 ();
 sg13g2_decap_8 FILLER_53_847 ();
 sg13g2_decap_8 FILLER_53_854 ();
 sg13g2_decap_8 FILLER_53_861 ();
 sg13g2_decap_8 FILLER_53_868 ();
 sg13g2_decap_8 FILLER_53_875 ();
 sg13g2_decap_8 FILLER_53_882 ();
 sg13g2_decap_8 FILLER_53_889 ();
 sg13g2_decap_8 FILLER_53_896 ();
 sg13g2_decap_8 FILLER_53_903 ();
 sg13g2_decap_8 FILLER_53_910 ();
 sg13g2_decap_8 FILLER_53_917 ();
 sg13g2_decap_8 FILLER_53_924 ();
 sg13g2_decap_8 FILLER_53_931 ();
 sg13g2_decap_8 FILLER_53_938 ();
 sg13g2_decap_8 FILLER_53_945 ();
 sg13g2_decap_8 FILLER_53_952 ();
 sg13g2_decap_8 FILLER_53_959 ();
 sg13g2_decap_8 FILLER_53_966 ();
 sg13g2_decap_8 FILLER_53_973 ();
 sg13g2_decap_8 FILLER_53_980 ();
 sg13g2_decap_8 FILLER_53_987 ();
 sg13g2_decap_8 FILLER_53_994 ();
 sg13g2_decap_8 FILLER_53_1001 ();
 sg13g2_decap_8 FILLER_53_1008 ();
 sg13g2_decap_8 FILLER_53_1015 ();
 sg13g2_decap_8 FILLER_53_1022 ();
 sg13g2_decap_8 FILLER_54_4 ();
 sg13g2_decap_8 FILLER_54_11 ();
 sg13g2_decap_8 FILLER_54_18 ();
 sg13g2_decap_8 FILLER_54_25 ();
 sg13g2_decap_8 FILLER_54_32 ();
 sg13g2_decap_8 FILLER_54_39 ();
 sg13g2_decap_8 FILLER_54_46 ();
 sg13g2_decap_8 FILLER_54_53 ();
 sg13g2_decap_8 FILLER_54_60 ();
 sg13g2_decap_8 FILLER_54_67 ();
 sg13g2_decap_8 FILLER_54_74 ();
 sg13g2_decap_8 FILLER_54_81 ();
 sg13g2_decap_8 FILLER_54_88 ();
 sg13g2_decap_8 FILLER_54_95 ();
 sg13g2_decap_8 FILLER_54_102 ();
 sg13g2_decap_8 FILLER_54_109 ();
 sg13g2_decap_8 FILLER_54_116 ();
 sg13g2_decap_8 FILLER_54_123 ();
 sg13g2_decap_8 FILLER_54_130 ();
 sg13g2_decap_8 FILLER_54_137 ();
 sg13g2_decap_8 FILLER_54_144 ();
 sg13g2_decap_8 FILLER_54_151 ();
 sg13g2_decap_8 FILLER_54_158 ();
 sg13g2_decap_8 FILLER_54_165 ();
 sg13g2_decap_8 FILLER_54_172 ();
 sg13g2_decap_8 FILLER_54_179 ();
 sg13g2_decap_8 FILLER_54_186 ();
 sg13g2_decap_8 FILLER_54_193 ();
 sg13g2_decap_8 FILLER_54_200 ();
 sg13g2_decap_8 FILLER_54_207 ();
 sg13g2_decap_8 FILLER_54_214 ();
 sg13g2_decap_8 FILLER_54_221 ();
 sg13g2_decap_8 FILLER_54_228 ();
 sg13g2_decap_8 FILLER_54_235 ();
 sg13g2_decap_8 FILLER_54_242 ();
 sg13g2_decap_8 FILLER_54_249 ();
 sg13g2_decap_8 FILLER_54_256 ();
 sg13g2_decap_8 FILLER_54_263 ();
 sg13g2_decap_8 FILLER_54_270 ();
 sg13g2_decap_8 FILLER_54_277 ();
 sg13g2_decap_8 FILLER_54_284 ();
 sg13g2_decap_8 FILLER_54_291 ();
 sg13g2_decap_8 FILLER_54_298 ();
 sg13g2_decap_8 FILLER_54_305 ();
 sg13g2_decap_8 FILLER_54_312 ();
 sg13g2_decap_8 FILLER_54_319 ();
 sg13g2_decap_8 FILLER_54_326 ();
 sg13g2_decap_8 FILLER_54_333 ();
 sg13g2_decap_8 FILLER_54_340 ();
 sg13g2_decap_8 FILLER_54_347 ();
 sg13g2_decap_8 FILLER_54_354 ();
 sg13g2_decap_8 FILLER_54_361 ();
 sg13g2_decap_8 FILLER_54_368 ();
 sg13g2_decap_8 FILLER_54_375 ();
 sg13g2_decap_8 FILLER_54_382 ();
 sg13g2_decap_8 FILLER_54_389 ();
 sg13g2_decap_8 FILLER_54_396 ();
 sg13g2_decap_8 FILLER_54_403 ();
 sg13g2_decap_8 FILLER_54_410 ();
 sg13g2_decap_8 FILLER_54_417 ();
 sg13g2_decap_8 FILLER_54_424 ();
 sg13g2_decap_8 FILLER_54_431 ();
 sg13g2_decap_8 FILLER_54_438 ();
 sg13g2_decap_8 FILLER_54_445 ();
 sg13g2_decap_8 FILLER_54_452 ();
 sg13g2_decap_8 FILLER_54_459 ();
 sg13g2_decap_8 FILLER_54_466 ();
 sg13g2_decap_8 FILLER_54_473 ();
 sg13g2_decap_8 FILLER_54_480 ();
 sg13g2_decap_8 FILLER_54_487 ();
 sg13g2_decap_8 FILLER_54_494 ();
 sg13g2_decap_8 FILLER_54_501 ();
 sg13g2_decap_8 FILLER_54_508 ();
 sg13g2_decap_8 FILLER_54_515 ();
 sg13g2_decap_8 FILLER_54_522 ();
 sg13g2_decap_8 FILLER_54_529 ();
 sg13g2_decap_8 FILLER_54_536 ();
 sg13g2_decap_8 FILLER_54_543 ();
 sg13g2_decap_8 FILLER_54_550 ();
 sg13g2_decap_8 FILLER_54_557 ();
 sg13g2_decap_8 FILLER_54_564 ();
 sg13g2_decap_8 FILLER_54_571 ();
 sg13g2_decap_8 FILLER_54_578 ();
 sg13g2_decap_8 FILLER_54_585 ();
 sg13g2_decap_8 FILLER_54_592 ();
 sg13g2_decap_8 FILLER_54_599 ();
 sg13g2_decap_8 FILLER_54_606 ();
 sg13g2_decap_8 FILLER_54_613 ();
 sg13g2_decap_8 FILLER_54_620 ();
 sg13g2_decap_8 FILLER_54_627 ();
 sg13g2_decap_8 FILLER_54_634 ();
 sg13g2_decap_8 FILLER_54_641 ();
 sg13g2_decap_8 FILLER_54_648 ();
 sg13g2_decap_8 FILLER_54_655 ();
 sg13g2_decap_8 FILLER_54_662 ();
 sg13g2_decap_8 FILLER_54_669 ();
 sg13g2_decap_8 FILLER_54_676 ();
 sg13g2_decap_8 FILLER_54_683 ();
 sg13g2_decap_8 FILLER_54_690 ();
 sg13g2_decap_8 FILLER_54_697 ();
 sg13g2_decap_8 FILLER_54_704 ();
 sg13g2_decap_8 FILLER_54_711 ();
 sg13g2_decap_8 FILLER_54_718 ();
 sg13g2_decap_8 FILLER_54_725 ();
 sg13g2_decap_8 FILLER_54_732 ();
 sg13g2_decap_8 FILLER_54_739 ();
 sg13g2_decap_8 FILLER_54_746 ();
 sg13g2_decap_8 FILLER_54_753 ();
 sg13g2_decap_8 FILLER_54_760 ();
 sg13g2_decap_8 FILLER_54_767 ();
 sg13g2_decap_8 FILLER_54_774 ();
 sg13g2_decap_8 FILLER_54_781 ();
 sg13g2_decap_8 FILLER_54_788 ();
 sg13g2_decap_8 FILLER_54_795 ();
 sg13g2_decap_8 FILLER_54_802 ();
 sg13g2_decap_8 FILLER_54_809 ();
 sg13g2_decap_8 FILLER_54_816 ();
 sg13g2_decap_8 FILLER_54_823 ();
 sg13g2_decap_8 FILLER_54_830 ();
 sg13g2_decap_8 FILLER_54_837 ();
 sg13g2_decap_8 FILLER_54_844 ();
 sg13g2_decap_8 FILLER_54_851 ();
 sg13g2_decap_8 FILLER_54_858 ();
 sg13g2_decap_8 FILLER_54_865 ();
 sg13g2_decap_8 FILLER_54_872 ();
 sg13g2_decap_8 FILLER_54_879 ();
 sg13g2_decap_8 FILLER_54_886 ();
 sg13g2_decap_8 FILLER_54_893 ();
 sg13g2_decap_8 FILLER_54_900 ();
 sg13g2_decap_8 FILLER_54_907 ();
 sg13g2_decap_8 FILLER_54_914 ();
 sg13g2_decap_8 FILLER_54_921 ();
 sg13g2_decap_8 FILLER_54_928 ();
 sg13g2_decap_8 FILLER_54_935 ();
 sg13g2_decap_8 FILLER_54_942 ();
 sg13g2_decap_8 FILLER_54_949 ();
 sg13g2_decap_8 FILLER_54_956 ();
 sg13g2_decap_8 FILLER_54_963 ();
 sg13g2_decap_8 FILLER_54_970 ();
 sg13g2_decap_8 FILLER_54_977 ();
 sg13g2_decap_8 FILLER_54_984 ();
 sg13g2_decap_8 FILLER_54_991 ();
 sg13g2_decap_8 FILLER_54_998 ();
 sg13g2_decap_8 FILLER_54_1005 ();
 sg13g2_decap_8 FILLER_54_1012 ();
 sg13g2_decap_8 FILLER_54_1019 ();
 sg13g2_fill_2 FILLER_54_1026 ();
 sg13g2_fill_1 FILLER_54_1028 ();
 sg13g2_decap_8 FILLER_55_0 ();
 sg13g2_decap_8 FILLER_55_7 ();
 sg13g2_decap_8 FILLER_55_14 ();
 sg13g2_decap_8 FILLER_55_21 ();
 sg13g2_decap_8 FILLER_55_28 ();
 sg13g2_decap_8 FILLER_55_35 ();
 sg13g2_decap_8 FILLER_55_42 ();
 sg13g2_decap_8 FILLER_55_49 ();
 sg13g2_decap_8 FILLER_55_56 ();
 sg13g2_decap_8 FILLER_55_63 ();
 sg13g2_decap_8 FILLER_55_70 ();
 sg13g2_decap_8 FILLER_55_77 ();
 sg13g2_decap_8 FILLER_55_84 ();
 sg13g2_decap_8 FILLER_55_91 ();
 sg13g2_decap_8 FILLER_55_98 ();
 sg13g2_decap_8 FILLER_55_105 ();
 sg13g2_decap_8 FILLER_55_112 ();
 sg13g2_decap_8 FILLER_55_119 ();
 sg13g2_decap_8 FILLER_55_126 ();
 sg13g2_decap_8 FILLER_55_133 ();
 sg13g2_decap_8 FILLER_55_140 ();
 sg13g2_decap_8 FILLER_55_147 ();
 sg13g2_decap_8 FILLER_55_154 ();
 sg13g2_decap_8 FILLER_55_161 ();
 sg13g2_decap_8 FILLER_55_168 ();
 sg13g2_decap_8 FILLER_55_175 ();
 sg13g2_decap_8 FILLER_55_182 ();
 sg13g2_decap_8 FILLER_55_189 ();
 sg13g2_decap_8 FILLER_55_196 ();
 sg13g2_decap_8 FILLER_55_203 ();
 sg13g2_decap_8 FILLER_55_210 ();
 sg13g2_decap_8 FILLER_55_217 ();
 sg13g2_decap_8 FILLER_55_224 ();
 sg13g2_decap_8 FILLER_55_231 ();
 sg13g2_decap_8 FILLER_55_238 ();
 sg13g2_decap_8 FILLER_55_245 ();
 sg13g2_decap_8 FILLER_55_252 ();
 sg13g2_decap_8 FILLER_55_259 ();
 sg13g2_decap_8 FILLER_55_266 ();
 sg13g2_decap_8 FILLER_55_273 ();
 sg13g2_decap_8 FILLER_55_280 ();
 sg13g2_decap_8 FILLER_55_287 ();
 sg13g2_decap_8 FILLER_55_294 ();
 sg13g2_decap_8 FILLER_55_301 ();
 sg13g2_decap_8 FILLER_55_308 ();
 sg13g2_decap_8 FILLER_55_315 ();
 sg13g2_decap_8 FILLER_55_322 ();
 sg13g2_decap_8 FILLER_55_329 ();
 sg13g2_decap_8 FILLER_55_336 ();
 sg13g2_decap_8 FILLER_55_343 ();
 sg13g2_decap_8 FILLER_55_350 ();
 sg13g2_decap_8 FILLER_55_357 ();
 sg13g2_decap_8 FILLER_55_364 ();
 sg13g2_decap_8 FILLER_55_371 ();
 sg13g2_decap_8 FILLER_55_378 ();
 sg13g2_decap_8 FILLER_55_385 ();
 sg13g2_decap_8 FILLER_55_392 ();
 sg13g2_decap_8 FILLER_55_399 ();
 sg13g2_decap_8 FILLER_55_406 ();
 sg13g2_decap_8 FILLER_55_413 ();
 sg13g2_decap_8 FILLER_55_420 ();
 sg13g2_decap_8 FILLER_55_427 ();
 sg13g2_decap_8 FILLER_55_434 ();
 sg13g2_decap_8 FILLER_55_441 ();
 sg13g2_decap_8 FILLER_55_448 ();
 sg13g2_decap_8 FILLER_55_455 ();
 sg13g2_decap_8 FILLER_55_462 ();
 sg13g2_decap_8 FILLER_55_469 ();
 sg13g2_decap_8 FILLER_55_476 ();
 sg13g2_decap_8 FILLER_55_483 ();
 sg13g2_decap_8 FILLER_55_490 ();
 sg13g2_decap_8 FILLER_55_497 ();
 sg13g2_decap_8 FILLER_55_504 ();
 sg13g2_decap_8 FILLER_55_511 ();
 sg13g2_decap_8 FILLER_55_518 ();
 sg13g2_decap_8 FILLER_55_525 ();
 sg13g2_decap_8 FILLER_55_532 ();
 sg13g2_decap_8 FILLER_55_539 ();
 sg13g2_decap_8 FILLER_55_546 ();
 sg13g2_decap_8 FILLER_55_553 ();
 sg13g2_decap_8 FILLER_55_560 ();
 sg13g2_decap_8 FILLER_55_567 ();
 sg13g2_decap_8 FILLER_55_574 ();
 sg13g2_decap_8 FILLER_55_581 ();
 sg13g2_decap_8 FILLER_55_588 ();
 sg13g2_decap_8 FILLER_55_595 ();
 sg13g2_decap_8 FILLER_55_602 ();
 sg13g2_decap_8 FILLER_55_609 ();
 sg13g2_decap_8 FILLER_55_616 ();
 sg13g2_decap_8 FILLER_55_623 ();
 sg13g2_decap_8 FILLER_55_630 ();
 sg13g2_decap_8 FILLER_55_637 ();
 sg13g2_decap_8 FILLER_55_644 ();
 sg13g2_decap_8 FILLER_55_651 ();
 sg13g2_decap_8 FILLER_55_658 ();
 sg13g2_decap_8 FILLER_55_665 ();
 sg13g2_decap_8 FILLER_55_672 ();
 sg13g2_decap_8 FILLER_55_679 ();
 sg13g2_decap_8 FILLER_55_686 ();
 sg13g2_decap_8 FILLER_55_693 ();
 sg13g2_decap_8 FILLER_55_700 ();
 sg13g2_decap_8 FILLER_55_707 ();
 sg13g2_decap_8 FILLER_55_714 ();
 sg13g2_decap_8 FILLER_55_721 ();
 sg13g2_decap_8 FILLER_55_728 ();
 sg13g2_decap_8 FILLER_55_735 ();
 sg13g2_decap_8 FILLER_55_742 ();
 sg13g2_decap_8 FILLER_55_749 ();
 sg13g2_decap_8 FILLER_55_756 ();
 sg13g2_decap_8 FILLER_55_763 ();
 sg13g2_decap_8 FILLER_55_770 ();
 sg13g2_decap_8 FILLER_55_777 ();
 sg13g2_decap_8 FILLER_55_784 ();
 sg13g2_decap_8 FILLER_55_791 ();
 sg13g2_decap_8 FILLER_55_798 ();
 sg13g2_decap_8 FILLER_55_805 ();
 sg13g2_decap_8 FILLER_55_812 ();
 sg13g2_decap_8 FILLER_55_819 ();
 sg13g2_decap_8 FILLER_55_826 ();
 sg13g2_decap_8 FILLER_55_833 ();
 sg13g2_decap_8 FILLER_55_840 ();
 sg13g2_decap_8 FILLER_55_847 ();
 sg13g2_decap_8 FILLER_55_854 ();
 sg13g2_decap_8 FILLER_55_861 ();
 sg13g2_decap_8 FILLER_55_868 ();
 sg13g2_decap_8 FILLER_55_875 ();
 sg13g2_decap_8 FILLER_55_882 ();
 sg13g2_decap_8 FILLER_55_889 ();
 sg13g2_decap_8 FILLER_55_896 ();
 sg13g2_decap_8 FILLER_55_903 ();
 sg13g2_decap_8 FILLER_55_910 ();
 sg13g2_decap_8 FILLER_55_917 ();
 sg13g2_decap_8 FILLER_55_924 ();
 sg13g2_decap_8 FILLER_55_931 ();
 sg13g2_decap_8 FILLER_55_938 ();
 sg13g2_decap_8 FILLER_55_945 ();
 sg13g2_decap_8 FILLER_55_952 ();
 sg13g2_decap_8 FILLER_55_959 ();
 sg13g2_decap_8 FILLER_55_966 ();
 sg13g2_decap_8 FILLER_55_973 ();
 sg13g2_decap_8 FILLER_55_980 ();
 sg13g2_decap_8 FILLER_55_987 ();
 sg13g2_decap_8 FILLER_55_994 ();
 sg13g2_decap_8 FILLER_55_1001 ();
 sg13g2_decap_8 FILLER_55_1008 ();
 sg13g2_decap_8 FILLER_55_1015 ();
 sg13g2_decap_8 FILLER_55_1022 ();
 sg13g2_decap_8 FILLER_56_4 ();
 sg13g2_decap_8 FILLER_56_11 ();
 sg13g2_decap_8 FILLER_56_18 ();
 sg13g2_decap_8 FILLER_56_25 ();
 sg13g2_decap_8 FILLER_56_32 ();
 sg13g2_decap_8 FILLER_56_39 ();
 sg13g2_decap_8 FILLER_56_46 ();
 sg13g2_decap_8 FILLER_56_53 ();
 sg13g2_decap_8 FILLER_56_60 ();
 sg13g2_decap_8 FILLER_56_67 ();
 sg13g2_decap_8 FILLER_56_74 ();
 sg13g2_decap_8 FILLER_56_81 ();
 sg13g2_decap_8 FILLER_56_88 ();
 sg13g2_decap_8 FILLER_56_95 ();
 sg13g2_decap_8 FILLER_56_102 ();
 sg13g2_decap_8 FILLER_56_109 ();
 sg13g2_decap_8 FILLER_56_116 ();
 sg13g2_decap_8 FILLER_56_123 ();
 sg13g2_decap_8 FILLER_56_130 ();
 sg13g2_decap_8 FILLER_56_137 ();
 sg13g2_decap_8 FILLER_56_144 ();
 sg13g2_decap_8 FILLER_56_151 ();
 sg13g2_decap_8 FILLER_56_158 ();
 sg13g2_decap_8 FILLER_56_165 ();
 sg13g2_decap_8 FILLER_56_172 ();
 sg13g2_decap_8 FILLER_56_179 ();
 sg13g2_decap_8 FILLER_56_186 ();
 sg13g2_decap_8 FILLER_56_193 ();
 sg13g2_decap_8 FILLER_56_200 ();
 sg13g2_decap_8 FILLER_56_207 ();
 sg13g2_decap_8 FILLER_56_214 ();
 sg13g2_decap_8 FILLER_56_221 ();
 sg13g2_decap_8 FILLER_56_228 ();
 sg13g2_decap_8 FILLER_56_235 ();
 sg13g2_decap_8 FILLER_56_242 ();
 sg13g2_decap_8 FILLER_56_249 ();
 sg13g2_decap_8 FILLER_56_256 ();
 sg13g2_decap_8 FILLER_56_263 ();
 sg13g2_decap_8 FILLER_56_270 ();
 sg13g2_decap_8 FILLER_56_277 ();
 sg13g2_decap_8 FILLER_56_284 ();
 sg13g2_decap_8 FILLER_56_291 ();
 sg13g2_decap_8 FILLER_56_298 ();
 sg13g2_decap_8 FILLER_56_305 ();
 sg13g2_decap_8 FILLER_56_312 ();
 sg13g2_decap_8 FILLER_56_319 ();
 sg13g2_decap_8 FILLER_56_326 ();
 sg13g2_decap_8 FILLER_56_333 ();
 sg13g2_decap_8 FILLER_56_340 ();
 sg13g2_decap_8 FILLER_56_347 ();
 sg13g2_decap_8 FILLER_56_354 ();
 sg13g2_decap_8 FILLER_56_361 ();
 sg13g2_decap_8 FILLER_56_368 ();
 sg13g2_decap_8 FILLER_56_375 ();
 sg13g2_decap_8 FILLER_56_382 ();
 sg13g2_decap_8 FILLER_56_389 ();
 sg13g2_decap_8 FILLER_56_396 ();
 sg13g2_decap_8 FILLER_56_403 ();
 sg13g2_decap_8 FILLER_56_410 ();
 sg13g2_decap_8 FILLER_56_417 ();
 sg13g2_decap_8 FILLER_56_424 ();
 sg13g2_decap_8 FILLER_56_431 ();
 sg13g2_decap_8 FILLER_56_438 ();
 sg13g2_decap_8 FILLER_56_445 ();
 sg13g2_decap_8 FILLER_56_452 ();
 sg13g2_decap_8 FILLER_56_459 ();
 sg13g2_decap_8 FILLER_56_466 ();
 sg13g2_decap_8 FILLER_56_473 ();
 sg13g2_decap_8 FILLER_56_480 ();
 sg13g2_decap_8 FILLER_56_487 ();
 sg13g2_decap_8 FILLER_56_494 ();
 sg13g2_decap_8 FILLER_56_501 ();
 sg13g2_decap_8 FILLER_56_508 ();
 sg13g2_decap_8 FILLER_56_515 ();
 sg13g2_decap_8 FILLER_56_522 ();
 sg13g2_decap_8 FILLER_56_529 ();
 sg13g2_decap_8 FILLER_56_536 ();
 sg13g2_decap_8 FILLER_56_543 ();
 sg13g2_decap_8 FILLER_56_550 ();
 sg13g2_decap_8 FILLER_56_557 ();
 sg13g2_decap_8 FILLER_56_564 ();
 sg13g2_decap_8 FILLER_56_571 ();
 sg13g2_decap_8 FILLER_56_578 ();
 sg13g2_decap_8 FILLER_56_585 ();
 sg13g2_decap_8 FILLER_56_592 ();
 sg13g2_decap_8 FILLER_56_599 ();
 sg13g2_decap_8 FILLER_56_606 ();
 sg13g2_decap_8 FILLER_56_613 ();
 sg13g2_decap_8 FILLER_56_620 ();
 sg13g2_decap_8 FILLER_56_627 ();
 sg13g2_decap_8 FILLER_56_634 ();
 sg13g2_decap_8 FILLER_56_641 ();
 sg13g2_decap_8 FILLER_56_648 ();
 sg13g2_decap_8 FILLER_56_655 ();
 sg13g2_decap_8 FILLER_56_662 ();
 sg13g2_decap_8 FILLER_56_669 ();
 sg13g2_decap_8 FILLER_56_676 ();
 sg13g2_decap_8 FILLER_56_683 ();
 sg13g2_decap_8 FILLER_56_690 ();
 sg13g2_decap_8 FILLER_56_697 ();
 sg13g2_decap_8 FILLER_56_704 ();
 sg13g2_decap_8 FILLER_56_711 ();
 sg13g2_decap_8 FILLER_56_718 ();
 sg13g2_decap_8 FILLER_56_725 ();
 sg13g2_decap_8 FILLER_56_732 ();
 sg13g2_decap_8 FILLER_56_739 ();
 sg13g2_decap_8 FILLER_56_746 ();
 sg13g2_decap_8 FILLER_56_753 ();
 sg13g2_decap_8 FILLER_56_760 ();
 sg13g2_decap_8 FILLER_56_767 ();
 sg13g2_decap_8 FILLER_56_774 ();
 sg13g2_decap_8 FILLER_56_781 ();
 sg13g2_decap_8 FILLER_56_788 ();
 sg13g2_decap_8 FILLER_56_795 ();
 sg13g2_decap_8 FILLER_56_802 ();
 sg13g2_decap_8 FILLER_56_809 ();
 sg13g2_decap_8 FILLER_56_816 ();
 sg13g2_decap_8 FILLER_56_823 ();
 sg13g2_decap_8 FILLER_56_830 ();
 sg13g2_decap_8 FILLER_56_837 ();
 sg13g2_decap_8 FILLER_56_844 ();
 sg13g2_decap_8 FILLER_56_851 ();
 sg13g2_decap_8 FILLER_56_858 ();
 sg13g2_decap_8 FILLER_56_865 ();
 sg13g2_decap_8 FILLER_56_872 ();
 sg13g2_decap_8 FILLER_56_879 ();
 sg13g2_decap_8 FILLER_56_886 ();
 sg13g2_decap_8 FILLER_56_893 ();
 sg13g2_decap_8 FILLER_56_900 ();
 sg13g2_decap_8 FILLER_56_907 ();
 sg13g2_decap_8 FILLER_56_914 ();
 sg13g2_decap_8 FILLER_56_921 ();
 sg13g2_decap_8 FILLER_56_928 ();
 sg13g2_decap_8 FILLER_56_935 ();
 sg13g2_decap_8 FILLER_56_942 ();
 sg13g2_decap_8 FILLER_56_949 ();
 sg13g2_decap_8 FILLER_56_956 ();
 sg13g2_decap_8 FILLER_56_963 ();
 sg13g2_decap_8 FILLER_56_970 ();
 sg13g2_decap_8 FILLER_56_977 ();
 sg13g2_decap_8 FILLER_56_984 ();
 sg13g2_decap_8 FILLER_56_991 ();
 sg13g2_decap_8 FILLER_56_998 ();
 sg13g2_decap_8 FILLER_56_1005 ();
 sg13g2_decap_8 FILLER_56_1012 ();
 sg13g2_decap_8 FILLER_56_1019 ();
 sg13g2_fill_2 FILLER_56_1026 ();
 sg13g2_fill_1 FILLER_56_1028 ();
 sg13g2_decap_8 FILLER_57_0 ();
 sg13g2_decap_8 FILLER_57_7 ();
 sg13g2_decap_8 FILLER_57_14 ();
 sg13g2_decap_8 FILLER_57_21 ();
 sg13g2_decap_8 FILLER_57_28 ();
 sg13g2_decap_8 FILLER_57_35 ();
 sg13g2_decap_8 FILLER_57_42 ();
 sg13g2_decap_8 FILLER_57_49 ();
 sg13g2_decap_8 FILLER_57_56 ();
 sg13g2_decap_8 FILLER_57_63 ();
 sg13g2_decap_8 FILLER_57_70 ();
 sg13g2_decap_8 FILLER_57_77 ();
 sg13g2_decap_8 FILLER_57_84 ();
 sg13g2_decap_8 FILLER_57_91 ();
 sg13g2_decap_8 FILLER_57_98 ();
 sg13g2_decap_8 FILLER_57_105 ();
 sg13g2_decap_8 FILLER_57_112 ();
 sg13g2_decap_8 FILLER_57_119 ();
 sg13g2_decap_8 FILLER_57_126 ();
 sg13g2_decap_8 FILLER_57_133 ();
 sg13g2_decap_8 FILLER_57_140 ();
 sg13g2_decap_8 FILLER_57_147 ();
 sg13g2_decap_8 FILLER_57_154 ();
 sg13g2_decap_8 FILLER_57_161 ();
 sg13g2_decap_8 FILLER_57_168 ();
 sg13g2_decap_8 FILLER_57_175 ();
 sg13g2_decap_8 FILLER_57_182 ();
 sg13g2_decap_8 FILLER_57_189 ();
 sg13g2_decap_8 FILLER_57_196 ();
 sg13g2_decap_8 FILLER_57_203 ();
 sg13g2_decap_8 FILLER_57_210 ();
 sg13g2_decap_8 FILLER_57_217 ();
 sg13g2_decap_8 FILLER_57_224 ();
 sg13g2_decap_8 FILLER_57_231 ();
 sg13g2_decap_8 FILLER_57_238 ();
 sg13g2_decap_8 FILLER_57_245 ();
 sg13g2_decap_8 FILLER_57_252 ();
 sg13g2_decap_8 FILLER_57_259 ();
 sg13g2_decap_8 FILLER_57_266 ();
 sg13g2_decap_8 FILLER_57_273 ();
 sg13g2_decap_8 FILLER_57_280 ();
 sg13g2_decap_8 FILLER_57_287 ();
 sg13g2_decap_8 FILLER_57_294 ();
 sg13g2_decap_8 FILLER_57_301 ();
 sg13g2_decap_8 FILLER_57_308 ();
 sg13g2_decap_8 FILLER_57_315 ();
 sg13g2_decap_8 FILLER_57_322 ();
 sg13g2_decap_8 FILLER_57_329 ();
 sg13g2_decap_8 FILLER_57_336 ();
 sg13g2_decap_8 FILLER_57_343 ();
 sg13g2_decap_8 FILLER_57_350 ();
 sg13g2_decap_8 FILLER_57_357 ();
 sg13g2_decap_8 FILLER_57_364 ();
 sg13g2_decap_8 FILLER_57_371 ();
 sg13g2_decap_8 FILLER_57_378 ();
 sg13g2_decap_8 FILLER_57_385 ();
 sg13g2_decap_8 FILLER_57_392 ();
 sg13g2_decap_8 FILLER_57_399 ();
 sg13g2_decap_8 FILLER_57_406 ();
 sg13g2_decap_8 FILLER_57_413 ();
 sg13g2_decap_8 FILLER_57_420 ();
 sg13g2_decap_8 FILLER_57_427 ();
 sg13g2_decap_8 FILLER_57_434 ();
 sg13g2_decap_8 FILLER_57_441 ();
 sg13g2_decap_8 FILLER_57_448 ();
 sg13g2_decap_8 FILLER_57_455 ();
 sg13g2_decap_8 FILLER_57_462 ();
 sg13g2_decap_8 FILLER_57_469 ();
 sg13g2_decap_8 FILLER_57_476 ();
 sg13g2_decap_8 FILLER_57_483 ();
 sg13g2_decap_8 FILLER_57_490 ();
 sg13g2_decap_8 FILLER_57_497 ();
 sg13g2_decap_8 FILLER_57_504 ();
 sg13g2_decap_8 FILLER_57_511 ();
 sg13g2_decap_8 FILLER_57_518 ();
 sg13g2_decap_8 FILLER_57_525 ();
 sg13g2_decap_8 FILLER_57_532 ();
 sg13g2_decap_8 FILLER_57_539 ();
 sg13g2_decap_8 FILLER_57_546 ();
 sg13g2_decap_8 FILLER_57_553 ();
 sg13g2_decap_8 FILLER_57_560 ();
 sg13g2_decap_8 FILLER_57_567 ();
 sg13g2_decap_8 FILLER_57_574 ();
 sg13g2_decap_8 FILLER_57_581 ();
 sg13g2_decap_8 FILLER_57_588 ();
 sg13g2_decap_8 FILLER_57_595 ();
 sg13g2_decap_8 FILLER_57_602 ();
 sg13g2_decap_8 FILLER_57_609 ();
 sg13g2_decap_8 FILLER_57_616 ();
 sg13g2_decap_8 FILLER_57_623 ();
 sg13g2_decap_8 FILLER_57_630 ();
 sg13g2_decap_8 FILLER_57_637 ();
 sg13g2_decap_8 FILLER_57_644 ();
 sg13g2_decap_8 FILLER_57_651 ();
 sg13g2_decap_8 FILLER_57_658 ();
 sg13g2_decap_8 FILLER_57_665 ();
 sg13g2_decap_8 FILLER_57_672 ();
 sg13g2_decap_8 FILLER_57_679 ();
 sg13g2_decap_8 FILLER_57_686 ();
 sg13g2_decap_8 FILLER_57_693 ();
 sg13g2_decap_8 FILLER_57_700 ();
 sg13g2_decap_8 FILLER_57_707 ();
 sg13g2_decap_8 FILLER_57_714 ();
 sg13g2_decap_8 FILLER_57_721 ();
 sg13g2_decap_8 FILLER_57_728 ();
 sg13g2_decap_8 FILLER_57_735 ();
 sg13g2_decap_8 FILLER_57_742 ();
 sg13g2_decap_8 FILLER_57_749 ();
 sg13g2_decap_8 FILLER_57_756 ();
 sg13g2_decap_8 FILLER_57_763 ();
 sg13g2_decap_8 FILLER_57_770 ();
 sg13g2_decap_8 FILLER_57_777 ();
 sg13g2_decap_8 FILLER_57_784 ();
 sg13g2_decap_8 FILLER_57_791 ();
 sg13g2_decap_8 FILLER_57_798 ();
 sg13g2_decap_8 FILLER_57_805 ();
 sg13g2_decap_8 FILLER_57_812 ();
 sg13g2_decap_8 FILLER_57_819 ();
 sg13g2_decap_8 FILLER_57_826 ();
 sg13g2_decap_8 FILLER_57_833 ();
 sg13g2_decap_8 FILLER_57_840 ();
 sg13g2_decap_8 FILLER_57_847 ();
 sg13g2_decap_8 FILLER_57_854 ();
 sg13g2_decap_8 FILLER_57_861 ();
 sg13g2_decap_8 FILLER_57_868 ();
 sg13g2_decap_8 FILLER_57_875 ();
 sg13g2_decap_8 FILLER_57_882 ();
 sg13g2_decap_8 FILLER_57_889 ();
 sg13g2_decap_8 FILLER_57_896 ();
 sg13g2_decap_8 FILLER_57_903 ();
 sg13g2_decap_8 FILLER_57_910 ();
 sg13g2_decap_8 FILLER_57_917 ();
 sg13g2_decap_8 FILLER_57_924 ();
 sg13g2_decap_8 FILLER_57_931 ();
 sg13g2_decap_8 FILLER_57_938 ();
 sg13g2_decap_8 FILLER_57_945 ();
 sg13g2_decap_8 FILLER_57_952 ();
 sg13g2_decap_8 FILLER_57_959 ();
 sg13g2_decap_8 FILLER_57_966 ();
 sg13g2_decap_8 FILLER_57_973 ();
 sg13g2_decap_8 FILLER_57_980 ();
 sg13g2_decap_8 FILLER_57_987 ();
 sg13g2_decap_8 FILLER_57_994 ();
 sg13g2_decap_8 FILLER_57_1001 ();
 sg13g2_decap_8 FILLER_57_1008 ();
 sg13g2_decap_8 FILLER_57_1015 ();
 sg13g2_decap_8 FILLER_57_1022 ();
 sg13g2_decap_8 FILLER_58_0 ();
 sg13g2_decap_8 FILLER_58_7 ();
 sg13g2_decap_8 FILLER_58_14 ();
 sg13g2_decap_8 FILLER_58_21 ();
 sg13g2_decap_8 FILLER_58_28 ();
 sg13g2_decap_8 FILLER_58_35 ();
 sg13g2_decap_8 FILLER_58_42 ();
 sg13g2_decap_8 FILLER_58_49 ();
 sg13g2_decap_8 FILLER_58_56 ();
 sg13g2_decap_8 FILLER_58_63 ();
 sg13g2_decap_8 FILLER_58_70 ();
 sg13g2_decap_8 FILLER_58_77 ();
 sg13g2_decap_8 FILLER_58_84 ();
 sg13g2_decap_8 FILLER_58_91 ();
 sg13g2_decap_8 FILLER_58_98 ();
 sg13g2_decap_8 FILLER_58_105 ();
 sg13g2_decap_8 FILLER_58_112 ();
 sg13g2_decap_8 FILLER_58_119 ();
 sg13g2_decap_8 FILLER_58_126 ();
 sg13g2_decap_4 FILLER_58_133 ();
 sg13g2_fill_2 FILLER_58_137 ();
 sg13g2_decap_8 FILLER_58_147 ();
 sg13g2_decap_8 FILLER_58_154 ();
 sg13g2_decap_8 FILLER_58_161 ();
 sg13g2_decap_8 FILLER_58_168 ();
 sg13g2_decap_8 FILLER_58_175 ();
 sg13g2_decap_8 FILLER_58_182 ();
 sg13g2_decap_8 FILLER_58_189 ();
 sg13g2_decap_8 FILLER_58_196 ();
 sg13g2_decap_8 FILLER_58_203 ();
 sg13g2_decap_8 FILLER_58_210 ();
 sg13g2_decap_8 FILLER_58_217 ();
 sg13g2_decap_8 FILLER_58_224 ();
 sg13g2_decap_8 FILLER_58_231 ();
 sg13g2_decap_8 FILLER_58_238 ();
 sg13g2_decap_8 FILLER_58_245 ();
 sg13g2_decap_8 FILLER_58_252 ();
 sg13g2_decap_8 FILLER_58_259 ();
 sg13g2_decap_8 FILLER_58_266 ();
 sg13g2_decap_8 FILLER_58_273 ();
 sg13g2_decap_8 FILLER_58_280 ();
 sg13g2_decap_8 FILLER_58_287 ();
 sg13g2_decap_8 FILLER_58_294 ();
 sg13g2_decap_8 FILLER_58_301 ();
 sg13g2_decap_8 FILLER_58_308 ();
 sg13g2_decap_8 FILLER_58_315 ();
 sg13g2_decap_8 FILLER_58_322 ();
 sg13g2_decap_8 FILLER_58_329 ();
 sg13g2_decap_8 FILLER_58_336 ();
 sg13g2_decap_8 FILLER_58_343 ();
 sg13g2_decap_8 FILLER_58_350 ();
 sg13g2_decap_8 FILLER_58_357 ();
 sg13g2_decap_8 FILLER_58_364 ();
 sg13g2_decap_8 FILLER_58_371 ();
 sg13g2_decap_8 FILLER_58_378 ();
 sg13g2_decap_8 FILLER_58_385 ();
 sg13g2_decap_8 FILLER_58_392 ();
 sg13g2_decap_8 FILLER_58_399 ();
 sg13g2_decap_8 FILLER_58_406 ();
 sg13g2_decap_8 FILLER_58_413 ();
 sg13g2_decap_8 FILLER_58_420 ();
 sg13g2_decap_8 FILLER_58_427 ();
 sg13g2_decap_8 FILLER_58_434 ();
 sg13g2_decap_8 FILLER_58_441 ();
 sg13g2_decap_8 FILLER_58_448 ();
 sg13g2_decap_8 FILLER_58_455 ();
 sg13g2_decap_8 FILLER_58_462 ();
 sg13g2_decap_8 FILLER_58_469 ();
 sg13g2_decap_8 FILLER_58_476 ();
 sg13g2_decap_8 FILLER_58_483 ();
 sg13g2_decap_8 FILLER_58_490 ();
 sg13g2_decap_8 FILLER_58_497 ();
 sg13g2_decap_8 FILLER_58_504 ();
 sg13g2_decap_8 FILLER_58_511 ();
 sg13g2_decap_8 FILLER_58_518 ();
 sg13g2_decap_8 FILLER_58_525 ();
 sg13g2_decap_8 FILLER_58_532 ();
 sg13g2_decap_8 FILLER_58_539 ();
 sg13g2_decap_8 FILLER_58_546 ();
 sg13g2_decap_8 FILLER_58_553 ();
 sg13g2_decap_8 FILLER_58_560 ();
 sg13g2_decap_8 FILLER_58_567 ();
 sg13g2_decap_8 FILLER_58_574 ();
 sg13g2_decap_8 FILLER_58_581 ();
 sg13g2_decap_8 FILLER_58_588 ();
 sg13g2_decap_8 FILLER_58_595 ();
 sg13g2_decap_8 FILLER_58_602 ();
 sg13g2_decap_8 FILLER_58_609 ();
 sg13g2_decap_8 FILLER_58_616 ();
 sg13g2_decap_8 FILLER_58_623 ();
 sg13g2_decap_8 FILLER_58_630 ();
 sg13g2_decap_8 FILLER_58_637 ();
 sg13g2_decap_8 FILLER_58_644 ();
 sg13g2_decap_8 FILLER_58_651 ();
 sg13g2_decap_8 FILLER_58_658 ();
 sg13g2_decap_8 FILLER_58_665 ();
 sg13g2_decap_8 FILLER_58_672 ();
 sg13g2_decap_8 FILLER_58_679 ();
 sg13g2_decap_8 FILLER_58_686 ();
 sg13g2_decap_8 FILLER_58_693 ();
 sg13g2_decap_8 FILLER_58_700 ();
 sg13g2_decap_8 FILLER_58_707 ();
 sg13g2_decap_8 FILLER_58_714 ();
 sg13g2_decap_8 FILLER_58_721 ();
 sg13g2_decap_8 FILLER_58_728 ();
 sg13g2_decap_8 FILLER_58_735 ();
 sg13g2_decap_8 FILLER_58_742 ();
 sg13g2_decap_8 FILLER_58_749 ();
 sg13g2_decap_8 FILLER_58_756 ();
 sg13g2_decap_8 FILLER_58_763 ();
 sg13g2_decap_8 FILLER_58_770 ();
 sg13g2_decap_8 FILLER_58_777 ();
 sg13g2_decap_8 FILLER_58_784 ();
 sg13g2_decap_8 FILLER_58_791 ();
 sg13g2_decap_8 FILLER_58_798 ();
 sg13g2_decap_8 FILLER_58_805 ();
 sg13g2_decap_8 FILLER_58_812 ();
 sg13g2_decap_8 FILLER_58_819 ();
 sg13g2_decap_8 FILLER_58_826 ();
 sg13g2_decap_8 FILLER_58_833 ();
 sg13g2_decap_8 FILLER_58_840 ();
 sg13g2_decap_8 FILLER_58_847 ();
 sg13g2_decap_8 FILLER_58_854 ();
 sg13g2_decap_8 FILLER_58_861 ();
 sg13g2_decap_8 FILLER_58_868 ();
 sg13g2_decap_8 FILLER_58_875 ();
 sg13g2_decap_8 FILLER_58_882 ();
 sg13g2_decap_8 FILLER_58_889 ();
 sg13g2_decap_8 FILLER_58_896 ();
 sg13g2_decap_8 FILLER_58_903 ();
 sg13g2_decap_8 FILLER_58_910 ();
 sg13g2_decap_8 FILLER_58_917 ();
 sg13g2_decap_8 FILLER_58_924 ();
 sg13g2_decap_8 FILLER_58_931 ();
 sg13g2_decap_8 FILLER_58_938 ();
 sg13g2_decap_8 FILLER_58_945 ();
 sg13g2_decap_8 FILLER_58_952 ();
 sg13g2_decap_8 FILLER_58_959 ();
 sg13g2_decap_8 FILLER_58_966 ();
 sg13g2_decap_8 FILLER_58_973 ();
 sg13g2_decap_8 FILLER_58_980 ();
 sg13g2_decap_8 FILLER_58_987 ();
 sg13g2_decap_8 FILLER_58_994 ();
 sg13g2_decap_8 FILLER_58_1001 ();
 sg13g2_decap_8 FILLER_58_1008 ();
 sg13g2_decap_8 FILLER_58_1015 ();
 sg13g2_decap_8 FILLER_58_1022 ();
 sg13g2_decap_8 FILLER_59_4 ();
 sg13g2_decap_8 FILLER_59_11 ();
 sg13g2_decap_8 FILLER_59_18 ();
 sg13g2_decap_8 FILLER_59_25 ();
 sg13g2_decap_8 FILLER_59_32 ();
 sg13g2_decap_8 FILLER_59_39 ();
 sg13g2_decap_8 FILLER_59_46 ();
 sg13g2_decap_8 FILLER_59_53 ();
 sg13g2_decap_8 FILLER_59_60 ();
 sg13g2_decap_4 FILLER_59_67 ();
 sg13g2_fill_1 FILLER_59_71 ();
 sg13g2_decap_8 FILLER_59_85 ();
 sg13g2_decap_8 FILLER_59_92 ();
 sg13g2_decap_8 FILLER_59_99 ();
 sg13g2_decap_8 FILLER_59_106 ();
 sg13g2_decap_8 FILLER_59_113 ();
 sg13g2_decap_8 FILLER_59_120 ();
 sg13g2_decap_8 FILLER_59_127 ();
 sg13g2_decap_4 FILLER_59_134 ();
 sg13g2_fill_2 FILLER_59_138 ();
 sg13g2_decap_8 FILLER_59_145 ();
 sg13g2_decap_8 FILLER_59_152 ();
 sg13g2_decap_8 FILLER_59_159 ();
 sg13g2_decap_8 FILLER_59_166 ();
 sg13g2_decap_8 FILLER_59_173 ();
 sg13g2_decap_8 FILLER_59_180 ();
 sg13g2_decap_8 FILLER_59_187 ();
 sg13g2_decap_8 FILLER_59_194 ();
 sg13g2_decap_8 FILLER_59_201 ();
 sg13g2_decap_8 FILLER_59_208 ();
 sg13g2_decap_8 FILLER_59_215 ();
 sg13g2_decap_8 FILLER_59_222 ();
 sg13g2_decap_8 FILLER_59_229 ();
 sg13g2_decap_8 FILLER_59_236 ();
 sg13g2_decap_8 FILLER_59_243 ();
 sg13g2_decap_8 FILLER_59_250 ();
 sg13g2_decap_8 FILLER_59_257 ();
 sg13g2_decap_8 FILLER_59_264 ();
 sg13g2_decap_8 FILLER_59_271 ();
 sg13g2_decap_8 FILLER_59_278 ();
 sg13g2_decap_8 FILLER_59_285 ();
 sg13g2_decap_8 FILLER_59_292 ();
 sg13g2_decap_8 FILLER_59_299 ();
 sg13g2_decap_8 FILLER_59_306 ();
 sg13g2_decap_8 FILLER_59_313 ();
 sg13g2_decap_8 FILLER_59_320 ();
 sg13g2_decap_8 FILLER_59_327 ();
 sg13g2_decap_8 FILLER_59_334 ();
 sg13g2_decap_8 FILLER_59_341 ();
 sg13g2_decap_8 FILLER_59_348 ();
 sg13g2_decap_8 FILLER_59_355 ();
 sg13g2_decap_8 FILLER_59_362 ();
 sg13g2_decap_8 FILLER_59_369 ();
 sg13g2_decap_8 FILLER_59_376 ();
 sg13g2_decap_8 FILLER_59_383 ();
 sg13g2_decap_8 FILLER_59_390 ();
 sg13g2_decap_8 FILLER_59_397 ();
 sg13g2_decap_8 FILLER_59_404 ();
 sg13g2_decap_8 FILLER_59_411 ();
 sg13g2_decap_8 FILLER_59_418 ();
 sg13g2_decap_8 FILLER_59_425 ();
 sg13g2_decap_8 FILLER_59_432 ();
 sg13g2_decap_8 FILLER_59_439 ();
 sg13g2_decap_8 FILLER_59_446 ();
 sg13g2_decap_8 FILLER_59_453 ();
 sg13g2_decap_8 FILLER_59_460 ();
 sg13g2_decap_8 FILLER_59_467 ();
 sg13g2_decap_8 FILLER_59_474 ();
 sg13g2_decap_8 FILLER_59_481 ();
 sg13g2_decap_8 FILLER_59_488 ();
 sg13g2_decap_8 FILLER_59_495 ();
 sg13g2_decap_8 FILLER_59_502 ();
 sg13g2_decap_8 FILLER_59_509 ();
 sg13g2_decap_8 FILLER_59_516 ();
 sg13g2_decap_8 FILLER_59_523 ();
 sg13g2_decap_8 FILLER_59_530 ();
 sg13g2_decap_8 FILLER_59_537 ();
 sg13g2_decap_8 FILLER_59_544 ();
 sg13g2_decap_8 FILLER_59_551 ();
 sg13g2_decap_8 FILLER_59_558 ();
 sg13g2_decap_8 FILLER_59_565 ();
 sg13g2_decap_8 FILLER_59_572 ();
 sg13g2_decap_8 FILLER_59_579 ();
 sg13g2_decap_8 FILLER_59_586 ();
 sg13g2_decap_8 FILLER_59_593 ();
 sg13g2_decap_8 FILLER_59_600 ();
 sg13g2_decap_8 FILLER_59_607 ();
 sg13g2_decap_8 FILLER_59_614 ();
 sg13g2_decap_8 FILLER_59_621 ();
 sg13g2_decap_8 FILLER_59_628 ();
 sg13g2_decap_8 FILLER_59_635 ();
 sg13g2_decap_8 FILLER_59_642 ();
 sg13g2_decap_8 FILLER_59_649 ();
 sg13g2_decap_8 FILLER_59_656 ();
 sg13g2_decap_8 FILLER_59_663 ();
 sg13g2_decap_8 FILLER_59_670 ();
 sg13g2_decap_8 FILLER_59_677 ();
 sg13g2_decap_8 FILLER_59_684 ();
 sg13g2_decap_8 FILLER_59_691 ();
 sg13g2_decap_8 FILLER_59_698 ();
 sg13g2_decap_8 FILLER_59_705 ();
 sg13g2_decap_8 FILLER_59_712 ();
 sg13g2_decap_8 FILLER_59_719 ();
 sg13g2_decap_8 FILLER_59_726 ();
 sg13g2_decap_8 FILLER_59_733 ();
 sg13g2_decap_8 FILLER_59_740 ();
 sg13g2_decap_8 FILLER_59_747 ();
 sg13g2_decap_8 FILLER_59_754 ();
 sg13g2_decap_8 FILLER_59_761 ();
 sg13g2_decap_8 FILLER_59_768 ();
 sg13g2_decap_8 FILLER_59_775 ();
 sg13g2_decap_8 FILLER_59_782 ();
 sg13g2_decap_8 FILLER_59_789 ();
 sg13g2_decap_8 FILLER_59_796 ();
 sg13g2_decap_8 FILLER_59_803 ();
 sg13g2_decap_8 FILLER_59_810 ();
 sg13g2_decap_8 FILLER_59_817 ();
 sg13g2_decap_8 FILLER_59_824 ();
 sg13g2_decap_8 FILLER_59_831 ();
 sg13g2_decap_8 FILLER_59_838 ();
 sg13g2_decap_8 FILLER_59_845 ();
 sg13g2_decap_8 FILLER_59_852 ();
 sg13g2_decap_8 FILLER_59_859 ();
 sg13g2_decap_8 FILLER_59_866 ();
 sg13g2_decap_8 FILLER_59_873 ();
 sg13g2_decap_8 FILLER_59_880 ();
 sg13g2_decap_8 FILLER_59_887 ();
 sg13g2_decap_8 FILLER_59_894 ();
 sg13g2_decap_8 FILLER_59_901 ();
 sg13g2_decap_8 FILLER_59_908 ();
 sg13g2_decap_8 FILLER_59_915 ();
 sg13g2_decap_8 FILLER_59_922 ();
 sg13g2_decap_8 FILLER_59_929 ();
 sg13g2_decap_8 FILLER_59_936 ();
 sg13g2_decap_8 FILLER_59_943 ();
 sg13g2_decap_8 FILLER_59_950 ();
 sg13g2_decap_8 FILLER_59_957 ();
 sg13g2_decap_8 FILLER_59_964 ();
 sg13g2_decap_8 FILLER_59_971 ();
 sg13g2_decap_8 FILLER_59_978 ();
 sg13g2_decap_8 FILLER_59_985 ();
 sg13g2_decap_8 FILLER_59_992 ();
 sg13g2_decap_8 FILLER_59_999 ();
 sg13g2_decap_8 FILLER_59_1006 ();
 sg13g2_decap_8 FILLER_59_1013 ();
 sg13g2_decap_8 FILLER_59_1020 ();
 sg13g2_fill_2 FILLER_59_1027 ();
 sg13g2_decap_8 FILLER_60_0 ();
 sg13g2_decap_8 FILLER_60_7 ();
 sg13g2_decap_4 FILLER_60_14 ();
 sg13g2_fill_2 FILLER_60_18 ();
 sg13g2_decap_8 FILLER_60_25 ();
 sg13g2_decap_8 FILLER_60_32 ();
 sg13g2_decap_8 FILLER_60_39 ();
 sg13g2_decap_8 FILLER_60_46 ();
 sg13g2_decap_8 FILLER_60_53 ();
 sg13g2_decap_8 FILLER_60_60 ();
 sg13g2_decap_8 FILLER_60_67 ();
 sg13g2_decap_8 FILLER_60_74 ();
 sg13g2_decap_8 FILLER_60_81 ();
 sg13g2_decap_8 FILLER_60_88 ();
 sg13g2_decap_8 FILLER_60_95 ();
 sg13g2_decap_8 FILLER_60_102 ();
 sg13g2_decap_8 FILLER_60_109 ();
 sg13g2_decap_8 FILLER_60_116 ();
 sg13g2_decap_8 FILLER_60_123 ();
 sg13g2_decap_4 FILLER_60_130 ();
 sg13g2_fill_2 FILLER_60_134 ();
 sg13g2_decap_8 FILLER_60_144 ();
 sg13g2_decap_8 FILLER_60_151 ();
 sg13g2_decap_8 FILLER_60_158 ();
 sg13g2_decap_8 FILLER_60_165 ();
 sg13g2_decap_8 FILLER_60_172 ();
 sg13g2_decap_8 FILLER_60_179 ();
 sg13g2_decap_8 FILLER_60_186 ();
 sg13g2_decap_8 FILLER_60_193 ();
 sg13g2_decap_8 FILLER_60_200 ();
 sg13g2_decap_8 FILLER_60_207 ();
 sg13g2_decap_8 FILLER_60_214 ();
 sg13g2_decap_8 FILLER_60_221 ();
 sg13g2_decap_8 FILLER_60_228 ();
 sg13g2_decap_8 FILLER_60_235 ();
 sg13g2_decap_8 FILLER_60_242 ();
 sg13g2_decap_8 FILLER_60_249 ();
 sg13g2_decap_8 FILLER_60_256 ();
 sg13g2_decap_8 FILLER_60_263 ();
 sg13g2_decap_8 FILLER_60_270 ();
 sg13g2_decap_8 FILLER_60_277 ();
 sg13g2_decap_8 FILLER_60_284 ();
 sg13g2_decap_8 FILLER_60_291 ();
 sg13g2_decap_8 FILLER_60_298 ();
 sg13g2_decap_8 FILLER_60_305 ();
 sg13g2_decap_8 FILLER_60_312 ();
 sg13g2_decap_8 FILLER_60_319 ();
 sg13g2_decap_8 FILLER_60_326 ();
 sg13g2_decap_8 FILLER_60_333 ();
 sg13g2_decap_8 FILLER_60_340 ();
 sg13g2_decap_8 FILLER_60_347 ();
 sg13g2_decap_8 FILLER_60_354 ();
 sg13g2_decap_8 FILLER_60_361 ();
 sg13g2_decap_8 FILLER_60_368 ();
 sg13g2_decap_8 FILLER_60_375 ();
 sg13g2_decap_8 FILLER_60_382 ();
 sg13g2_decap_8 FILLER_60_389 ();
 sg13g2_decap_8 FILLER_60_396 ();
 sg13g2_decap_8 FILLER_60_403 ();
 sg13g2_decap_8 FILLER_60_410 ();
 sg13g2_decap_8 FILLER_60_417 ();
 sg13g2_decap_8 FILLER_60_424 ();
 sg13g2_decap_8 FILLER_60_431 ();
 sg13g2_decap_8 FILLER_60_438 ();
 sg13g2_decap_8 FILLER_60_445 ();
 sg13g2_decap_8 FILLER_60_452 ();
 sg13g2_decap_8 FILLER_60_459 ();
 sg13g2_decap_8 FILLER_60_466 ();
 sg13g2_decap_8 FILLER_60_473 ();
 sg13g2_decap_8 FILLER_60_480 ();
 sg13g2_decap_8 FILLER_60_487 ();
 sg13g2_decap_8 FILLER_60_494 ();
 sg13g2_decap_8 FILLER_60_501 ();
 sg13g2_decap_8 FILLER_60_508 ();
 sg13g2_decap_8 FILLER_60_515 ();
 sg13g2_decap_8 FILLER_60_522 ();
 sg13g2_decap_8 FILLER_60_529 ();
 sg13g2_decap_8 FILLER_60_536 ();
 sg13g2_decap_8 FILLER_60_543 ();
 sg13g2_decap_8 FILLER_60_550 ();
 sg13g2_decap_8 FILLER_60_557 ();
 sg13g2_decap_8 FILLER_60_564 ();
 sg13g2_decap_8 FILLER_60_571 ();
 sg13g2_decap_8 FILLER_60_578 ();
 sg13g2_decap_8 FILLER_60_585 ();
 sg13g2_decap_8 FILLER_60_592 ();
 sg13g2_decap_8 FILLER_60_599 ();
 sg13g2_decap_8 FILLER_60_606 ();
 sg13g2_decap_8 FILLER_60_613 ();
 sg13g2_decap_8 FILLER_60_620 ();
 sg13g2_decap_8 FILLER_60_627 ();
 sg13g2_decap_8 FILLER_60_634 ();
 sg13g2_decap_8 FILLER_60_641 ();
 sg13g2_decap_8 FILLER_60_648 ();
 sg13g2_decap_8 FILLER_60_655 ();
 sg13g2_decap_8 FILLER_60_662 ();
 sg13g2_decap_8 FILLER_60_669 ();
 sg13g2_decap_8 FILLER_60_676 ();
 sg13g2_decap_8 FILLER_60_683 ();
 sg13g2_decap_8 FILLER_60_690 ();
 sg13g2_decap_8 FILLER_60_697 ();
 sg13g2_decap_8 FILLER_60_704 ();
 sg13g2_decap_8 FILLER_60_711 ();
 sg13g2_decap_8 FILLER_60_718 ();
 sg13g2_decap_8 FILLER_60_725 ();
 sg13g2_decap_8 FILLER_60_732 ();
 sg13g2_decap_8 FILLER_60_739 ();
 sg13g2_decap_8 FILLER_60_746 ();
 sg13g2_decap_8 FILLER_60_753 ();
 sg13g2_decap_8 FILLER_60_760 ();
 sg13g2_decap_8 FILLER_60_767 ();
 sg13g2_decap_8 FILLER_60_774 ();
 sg13g2_decap_8 FILLER_60_781 ();
 sg13g2_decap_8 FILLER_60_788 ();
 sg13g2_decap_8 FILLER_60_795 ();
 sg13g2_decap_8 FILLER_60_802 ();
 sg13g2_decap_8 FILLER_60_809 ();
 sg13g2_decap_8 FILLER_60_816 ();
 sg13g2_decap_8 FILLER_60_823 ();
 sg13g2_decap_8 FILLER_60_830 ();
 sg13g2_decap_8 FILLER_60_837 ();
 sg13g2_decap_8 FILLER_60_844 ();
 sg13g2_decap_8 FILLER_60_851 ();
 sg13g2_decap_8 FILLER_60_858 ();
 sg13g2_decap_8 FILLER_60_865 ();
 sg13g2_decap_8 FILLER_60_872 ();
 sg13g2_decap_8 FILLER_60_879 ();
 sg13g2_decap_8 FILLER_60_886 ();
 sg13g2_decap_8 FILLER_60_893 ();
 sg13g2_decap_8 FILLER_60_900 ();
 sg13g2_decap_8 FILLER_60_907 ();
 sg13g2_decap_8 FILLER_60_914 ();
 sg13g2_decap_8 FILLER_60_921 ();
 sg13g2_decap_8 FILLER_60_928 ();
 sg13g2_decap_8 FILLER_60_935 ();
 sg13g2_decap_8 FILLER_60_942 ();
 sg13g2_decap_8 FILLER_60_949 ();
 sg13g2_decap_8 FILLER_60_956 ();
 sg13g2_decap_8 FILLER_60_963 ();
 sg13g2_decap_8 FILLER_60_970 ();
 sg13g2_decap_8 FILLER_60_977 ();
 sg13g2_decap_8 FILLER_60_984 ();
 sg13g2_decap_8 FILLER_60_991 ();
 sg13g2_decap_8 FILLER_60_998 ();
 sg13g2_decap_8 FILLER_60_1005 ();
 sg13g2_decap_8 FILLER_60_1012 ();
 sg13g2_decap_8 FILLER_60_1019 ();
 sg13g2_fill_2 FILLER_60_1026 ();
 sg13g2_fill_1 FILLER_60_1028 ();
 sg13g2_decap_8 FILLER_61_4 ();
 sg13g2_fill_2 FILLER_61_11 ();
 sg13g2_fill_1 FILLER_61_13 ();
 sg13g2_decap_4 FILLER_61_27 ();
 sg13g2_fill_1 FILLER_61_31 ();
 sg13g2_decap_8 FILLER_61_37 ();
 sg13g2_decap_8 FILLER_61_44 ();
 sg13g2_fill_2 FILLER_61_68 ();
 sg13g2_decap_8 FILLER_61_74 ();
 sg13g2_decap_8 FILLER_61_81 ();
 sg13g2_decap_8 FILLER_61_88 ();
 sg13g2_decap_8 FILLER_61_95 ();
 sg13g2_decap_8 FILLER_61_102 ();
 sg13g2_decap_8 FILLER_61_109 ();
 sg13g2_decap_8 FILLER_61_116 ();
 sg13g2_decap_8 FILLER_61_123 ();
 sg13g2_decap_8 FILLER_61_151 ();
 sg13g2_decap_8 FILLER_61_158 ();
 sg13g2_decap_8 FILLER_61_165 ();
 sg13g2_decap_8 FILLER_61_172 ();
 sg13g2_decap_8 FILLER_61_179 ();
 sg13g2_decap_8 FILLER_61_186 ();
 sg13g2_decap_8 FILLER_61_193 ();
 sg13g2_decap_8 FILLER_61_200 ();
 sg13g2_decap_8 FILLER_61_207 ();
 sg13g2_decap_8 FILLER_61_214 ();
 sg13g2_decap_8 FILLER_61_221 ();
 sg13g2_decap_8 FILLER_61_228 ();
 sg13g2_decap_8 FILLER_61_235 ();
 sg13g2_decap_8 FILLER_61_242 ();
 sg13g2_decap_8 FILLER_61_249 ();
 sg13g2_decap_8 FILLER_61_256 ();
 sg13g2_decap_8 FILLER_61_263 ();
 sg13g2_decap_8 FILLER_61_270 ();
 sg13g2_decap_8 FILLER_61_277 ();
 sg13g2_decap_8 FILLER_61_284 ();
 sg13g2_decap_8 FILLER_61_291 ();
 sg13g2_decap_8 FILLER_61_298 ();
 sg13g2_decap_8 FILLER_61_305 ();
 sg13g2_decap_8 FILLER_61_312 ();
 sg13g2_decap_8 FILLER_61_319 ();
 sg13g2_decap_8 FILLER_61_326 ();
 sg13g2_decap_8 FILLER_61_333 ();
 sg13g2_decap_8 FILLER_61_340 ();
 sg13g2_decap_8 FILLER_61_347 ();
 sg13g2_decap_8 FILLER_61_354 ();
 sg13g2_decap_8 FILLER_61_361 ();
 sg13g2_decap_8 FILLER_61_368 ();
 sg13g2_decap_8 FILLER_61_375 ();
 sg13g2_decap_8 FILLER_61_382 ();
 sg13g2_decap_8 FILLER_61_389 ();
 sg13g2_decap_8 FILLER_61_396 ();
 sg13g2_decap_8 FILLER_61_403 ();
 sg13g2_decap_8 FILLER_61_410 ();
 sg13g2_decap_8 FILLER_61_417 ();
 sg13g2_decap_8 FILLER_61_424 ();
 sg13g2_decap_8 FILLER_61_431 ();
 sg13g2_decap_8 FILLER_61_438 ();
 sg13g2_decap_8 FILLER_61_445 ();
 sg13g2_decap_8 FILLER_61_452 ();
 sg13g2_decap_8 FILLER_61_459 ();
 sg13g2_decap_8 FILLER_61_466 ();
 sg13g2_decap_8 FILLER_61_473 ();
 sg13g2_decap_8 FILLER_61_480 ();
 sg13g2_decap_8 FILLER_61_487 ();
 sg13g2_decap_8 FILLER_61_494 ();
 sg13g2_decap_8 FILLER_61_501 ();
 sg13g2_decap_8 FILLER_61_508 ();
 sg13g2_decap_8 FILLER_61_515 ();
 sg13g2_decap_8 FILLER_61_522 ();
 sg13g2_decap_8 FILLER_61_529 ();
 sg13g2_decap_8 FILLER_61_536 ();
 sg13g2_decap_8 FILLER_61_543 ();
 sg13g2_decap_8 FILLER_61_550 ();
 sg13g2_decap_8 FILLER_61_557 ();
 sg13g2_decap_8 FILLER_61_564 ();
 sg13g2_decap_8 FILLER_61_571 ();
 sg13g2_decap_8 FILLER_61_578 ();
 sg13g2_decap_8 FILLER_61_585 ();
 sg13g2_decap_8 FILLER_61_592 ();
 sg13g2_decap_8 FILLER_61_599 ();
 sg13g2_decap_8 FILLER_61_606 ();
 sg13g2_decap_8 FILLER_61_613 ();
 sg13g2_decap_8 FILLER_61_620 ();
 sg13g2_decap_8 FILLER_61_627 ();
 sg13g2_decap_8 FILLER_61_634 ();
 sg13g2_decap_8 FILLER_61_641 ();
 sg13g2_decap_8 FILLER_61_648 ();
 sg13g2_decap_8 FILLER_61_655 ();
 sg13g2_decap_8 FILLER_61_662 ();
 sg13g2_decap_8 FILLER_61_669 ();
 sg13g2_decap_8 FILLER_61_676 ();
 sg13g2_decap_8 FILLER_61_683 ();
 sg13g2_decap_8 FILLER_61_690 ();
 sg13g2_decap_8 FILLER_61_697 ();
 sg13g2_decap_8 FILLER_61_704 ();
 sg13g2_decap_8 FILLER_61_711 ();
 sg13g2_decap_8 FILLER_61_718 ();
 sg13g2_decap_8 FILLER_61_725 ();
 sg13g2_decap_8 FILLER_61_732 ();
 sg13g2_decap_8 FILLER_61_739 ();
 sg13g2_decap_8 FILLER_61_746 ();
 sg13g2_decap_8 FILLER_61_753 ();
 sg13g2_decap_8 FILLER_61_760 ();
 sg13g2_decap_8 FILLER_61_767 ();
 sg13g2_decap_8 FILLER_61_774 ();
 sg13g2_decap_8 FILLER_61_781 ();
 sg13g2_decap_8 FILLER_61_788 ();
 sg13g2_decap_8 FILLER_61_795 ();
 sg13g2_decap_8 FILLER_61_802 ();
 sg13g2_decap_8 FILLER_61_809 ();
 sg13g2_decap_8 FILLER_61_816 ();
 sg13g2_decap_8 FILLER_61_823 ();
 sg13g2_decap_8 FILLER_61_830 ();
 sg13g2_decap_8 FILLER_61_837 ();
 sg13g2_decap_8 FILLER_61_844 ();
 sg13g2_decap_8 FILLER_61_851 ();
 sg13g2_decap_8 FILLER_61_858 ();
 sg13g2_decap_8 FILLER_61_865 ();
 sg13g2_decap_8 FILLER_61_872 ();
 sg13g2_decap_8 FILLER_61_879 ();
 sg13g2_decap_8 FILLER_61_886 ();
 sg13g2_decap_8 FILLER_61_893 ();
 sg13g2_decap_8 FILLER_61_900 ();
 sg13g2_decap_8 FILLER_61_907 ();
 sg13g2_decap_8 FILLER_61_914 ();
 sg13g2_decap_8 FILLER_61_921 ();
 sg13g2_decap_8 FILLER_61_928 ();
 sg13g2_decap_8 FILLER_61_935 ();
 sg13g2_decap_8 FILLER_61_942 ();
 sg13g2_decap_8 FILLER_61_949 ();
 sg13g2_decap_8 FILLER_61_956 ();
 sg13g2_decap_8 FILLER_61_963 ();
 sg13g2_decap_8 FILLER_61_970 ();
 sg13g2_decap_8 FILLER_61_977 ();
 sg13g2_decap_8 FILLER_61_984 ();
 sg13g2_decap_8 FILLER_61_991 ();
 sg13g2_decap_8 FILLER_61_998 ();
 sg13g2_decap_8 FILLER_61_1005 ();
 sg13g2_decap_8 FILLER_61_1012 ();
 sg13g2_decap_8 FILLER_61_1019 ();
 sg13g2_fill_2 FILLER_61_1026 ();
 sg13g2_fill_1 FILLER_61_1028 ();
 sg13g2_decap_8 FILLER_62_0 ();
 sg13g2_decap_8 FILLER_62_7 ();
 sg13g2_decap_8 FILLER_62_14 ();
 sg13g2_decap_8 FILLER_62_21 ();
 sg13g2_decap_8 FILLER_62_28 ();
 sg13g2_decap_8 FILLER_62_35 ();
 sg13g2_decap_8 FILLER_62_42 ();
 sg13g2_decap_8 FILLER_62_49 ();
 sg13g2_fill_1 FILLER_62_56 ();
 sg13g2_decap_8 FILLER_62_62 ();
 sg13g2_decap_8 FILLER_62_69 ();
 sg13g2_decap_8 FILLER_62_76 ();
 sg13g2_decap_8 FILLER_62_83 ();
 sg13g2_decap_8 FILLER_62_98 ();
 sg13g2_decap_8 FILLER_62_105 ();
 sg13g2_decap_8 FILLER_62_112 ();
 sg13g2_decap_8 FILLER_62_119 ();
 sg13g2_decap_8 FILLER_62_126 ();
 sg13g2_decap_8 FILLER_62_133 ();
 sg13g2_decap_8 FILLER_62_140 ();
 sg13g2_decap_8 FILLER_62_147 ();
 sg13g2_decap_8 FILLER_62_154 ();
 sg13g2_decap_8 FILLER_62_161 ();
 sg13g2_decap_8 FILLER_62_168 ();
 sg13g2_decap_8 FILLER_62_175 ();
 sg13g2_decap_8 FILLER_62_182 ();
 sg13g2_decap_8 FILLER_62_189 ();
 sg13g2_decap_8 FILLER_62_196 ();
 sg13g2_decap_8 FILLER_62_203 ();
 sg13g2_decap_8 FILLER_62_210 ();
 sg13g2_decap_8 FILLER_62_217 ();
 sg13g2_decap_8 FILLER_62_224 ();
 sg13g2_decap_8 FILLER_62_231 ();
 sg13g2_decap_8 FILLER_62_238 ();
 sg13g2_decap_8 FILLER_62_245 ();
 sg13g2_decap_8 FILLER_62_252 ();
 sg13g2_decap_8 FILLER_62_259 ();
 sg13g2_decap_8 FILLER_62_266 ();
 sg13g2_decap_8 FILLER_62_273 ();
 sg13g2_decap_8 FILLER_62_280 ();
 sg13g2_decap_8 FILLER_62_287 ();
 sg13g2_decap_8 FILLER_62_294 ();
 sg13g2_decap_8 FILLER_62_301 ();
 sg13g2_decap_8 FILLER_62_308 ();
 sg13g2_decap_8 FILLER_62_315 ();
 sg13g2_decap_8 FILLER_62_322 ();
 sg13g2_decap_8 FILLER_62_329 ();
 sg13g2_decap_8 FILLER_62_336 ();
 sg13g2_decap_8 FILLER_62_343 ();
 sg13g2_decap_8 FILLER_62_350 ();
 sg13g2_decap_8 FILLER_62_357 ();
 sg13g2_decap_8 FILLER_62_364 ();
 sg13g2_decap_8 FILLER_62_371 ();
 sg13g2_decap_8 FILLER_62_378 ();
 sg13g2_decap_8 FILLER_62_385 ();
 sg13g2_decap_8 FILLER_62_392 ();
 sg13g2_decap_8 FILLER_62_399 ();
 sg13g2_decap_8 FILLER_62_406 ();
 sg13g2_decap_8 FILLER_62_413 ();
 sg13g2_decap_8 FILLER_62_420 ();
 sg13g2_decap_8 FILLER_62_427 ();
 sg13g2_decap_8 FILLER_62_434 ();
 sg13g2_decap_8 FILLER_62_441 ();
 sg13g2_decap_8 FILLER_62_448 ();
 sg13g2_decap_8 FILLER_62_455 ();
 sg13g2_decap_8 FILLER_62_462 ();
 sg13g2_decap_8 FILLER_62_469 ();
 sg13g2_decap_8 FILLER_62_476 ();
 sg13g2_decap_8 FILLER_62_483 ();
 sg13g2_decap_8 FILLER_62_490 ();
 sg13g2_decap_8 FILLER_62_497 ();
 sg13g2_decap_8 FILLER_62_504 ();
 sg13g2_decap_8 FILLER_62_511 ();
 sg13g2_decap_8 FILLER_62_518 ();
 sg13g2_decap_8 FILLER_62_525 ();
 sg13g2_decap_8 FILLER_62_532 ();
 sg13g2_decap_8 FILLER_62_539 ();
 sg13g2_decap_8 FILLER_62_546 ();
 sg13g2_decap_8 FILLER_62_553 ();
 sg13g2_decap_8 FILLER_62_560 ();
 sg13g2_decap_8 FILLER_62_567 ();
 sg13g2_decap_8 FILLER_62_574 ();
 sg13g2_decap_8 FILLER_62_581 ();
 sg13g2_decap_8 FILLER_62_588 ();
 sg13g2_decap_8 FILLER_62_595 ();
 sg13g2_decap_8 FILLER_62_602 ();
 sg13g2_decap_8 FILLER_62_609 ();
 sg13g2_decap_8 FILLER_62_616 ();
 sg13g2_decap_8 FILLER_62_623 ();
 sg13g2_decap_8 FILLER_62_630 ();
 sg13g2_decap_8 FILLER_62_637 ();
 sg13g2_decap_8 FILLER_62_644 ();
 sg13g2_decap_8 FILLER_62_651 ();
 sg13g2_decap_8 FILLER_62_658 ();
 sg13g2_decap_8 FILLER_62_665 ();
 sg13g2_decap_8 FILLER_62_672 ();
 sg13g2_decap_8 FILLER_62_679 ();
 sg13g2_decap_8 FILLER_62_686 ();
 sg13g2_decap_8 FILLER_62_693 ();
 sg13g2_decap_8 FILLER_62_700 ();
 sg13g2_decap_8 FILLER_62_707 ();
 sg13g2_decap_8 FILLER_62_714 ();
 sg13g2_decap_8 FILLER_62_721 ();
 sg13g2_decap_8 FILLER_62_728 ();
 sg13g2_decap_8 FILLER_62_735 ();
 sg13g2_decap_8 FILLER_62_742 ();
 sg13g2_decap_8 FILLER_62_749 ();
 sg13g2_decap_8 FILLER_62_756 ();
 sg13g2_decap_8 FILLER_62_763 ();
 sg13g2_decap_8 FILLER_62_770 ();
 sg13g2_decap_8 FILLER_62_777 ();
 sg13g2_decap_8 FILLER_62_784 ();
 sg13g2_decap_8 FILLER_62_791 ();
 sg13g2_decap_8 FILLER_62_798 ();
 sg13g2_decap_8 FILLER_62_805 ();
 sg13g2_decap_8 FILLER_62_812 ();
 sg13g2_decap_8 FILLER_62_819 ();
 sg13g2_decap_8 FILLER_62_826 ();
 sg13g2_decap_8 FILLER_62_833 ();
 sg13g2_decap_8 FILLER_62_840 ();
 sg13g2_decap_8 FILLER_62_847 ();
 sg13g2_decap_8 FILLER_62_854 ();
 sg13g2_decap_8 FILLER_62_861 ();
 sg13g2_decap_8 FILLER_62_868 ();
 sg13g2_decap_8 FILLER_62_875 ();
 sg13g2_decap_8 FILLER_62_882 ();
 sg13g2_decap_8 FILLER_62_889 ();
 sg13g2_decap_8 FILLER_62_896 ();
 sg13g2_decap_8 FILLER_62_903 ();
 sg13g2_decap_8 FILLER_62_910 ();
 sg13g2_decap_8 FILLER_62_917 ();
 sg13g2_decap_8 FILLER_62_924 ();
 sg13g2_decap_8 FILLER_62_931 ();
 sg13g2_decap_8 FILLER_62_938 ();
 sg13g2_decap_8 FILLER_62_945 ();
 sg13g2_decap_8 FILLER_62_952 ();
 sg13g2_decap_8 FILLER_62_959 ();
 sg13g2_decap_8 FILLER_62_966 ();
 sg13g2_decap_8 FILLER_62_973 ();
 sg13g2_decap_8 FILLER_62_980 ();
 sg13g2_decap_8 FILLER_62_987 ();
 sg13g2_decap_8 FILLER_62_994 ();
 sg13g2_decap_8 FILLER_62_1001 ();
 sg13g2_decap_8 FILLER_62_1008 ();
 sg13g2_decap_8 FILLER_62_1015 ();
 sg13g2_decap_8 FILLER_62_1022 ();
 sg13g2_decap_8 FILLER_63_0 ();
 sg13g2_decap_8 FILLER_63_7 ();
 sg13g2_decap_8 FILLER_63_14 ();
 sg13g2_decap_8 FILLER_63_21 ();
 sg13g2_decap_8 FILLER_63_28 ();
 sg13g2_decap_8 FILLER_63_35 ();
 sg13g2_decap_8 FILLER_63_42 ();
 sg13g2_decap_8 FILLER_63_49 ();
 sg13g2_decap_8 FILLER_63_56 ();
 sg13g2_decap_8 FILLER_63_63 ();
 sg13g2_decap_8 FILLER_63_70 ();
 sg13g2_decap_8 FILLER_63_77 ();
 sg13g2_decap_8 FILLER_63_84 ();
 sg13g2_decap_8 FILLER_63_91 ();
 sg13g2_decap_8 FILLER_63_98 ();
 sg13g2_decap_8 FILLER_63_105 ();
 sg13g2_decap_8 FILLER_63_112 ();
 sg13g2_decap_8 FILLER_63_119 ();
 sg13g2_decap_8 FILLER_63_126 ();
 sg13g2_decap_8 FILLER_63_133 ();
 sg13g2_decap_8 FILLER_63_140 ();
 sg13g2_decap_8 FILLER_63_147 ();
 sg13g2_decap_8 FILLER_63_154 ();
 sg13g2_decap_8 FILLER_63_161 ();
 sg13g2_decap_8 FILLER_63_168 ();
 sg13g2_decap_8 FILLER_63_175 ();
 sg13g2_decap_8 FILLER_63_182 ();
 sg13g2_decap_8 FILLER_63_189 ();
 sg13g2_decap_8 FILLER_63_196 ();
 sg13g2_decap_8 FILLER_63_203 ();
 sg13g2_decap_8 FILLER_63_210 ();
 sg13g2_decap_8 FILLER_63_217 ();
 sg13g2_decap_8 FILLER_63_224 ();
 sg13g2_decap_8 FILLER_63_231 ();
 sg13g2_decap_8 FILLER_63_238 ();
 sg13g2_decap_8 FILLER_63_245 ();
 sg13g2_decap_8 FILLER_63_252 ();
 sg13g2_decap_8 FILLER_63_259 ();
 sg13g2_decap_8 FILLER_63_266 ();
 sg13g2_decap_8 FILLER_63_273 ();
 sg13g2_decap_8 FILLER_63_280 ();
 sg13g2_decap_8 FILLER_63_287 ();
 sg13g2_decap_8 FILLER_63_294 ();
 sg13g2_decap_8 FILLER_63_301 ();
 sg13g2_decap_8 FILLER_63_308 ();
 sg13g2_decap_8 FILLER_63_315 ();
 sg13g2_decap_8 FILLER_63_322 ();
 sg13g2_decap_8 FILLER_63_329 ();
 sg13g2_decap_8 FILLER_63_336 ();
 sg13g2_decap_8 FILLER_63_343 ();
 sg13g2_decap_8 FILLER_63_350 ();
 sg13g2_decap_8 FILLER_63_357 ();
 sg13g2_decap_8 FILLER_63_364 ();
 sg13g2_decap_8 FILLER_63_371 ();
 sg13g2_decap_8 FILLER_63_378 ();
 sg13g2_decap_8 FILLER_63_385 ();
 sg13g2_decap_8 FILLER_63_392 ();
 sg13g2_decap_8 FILLER_63_399 ();
 sg13g2_decap_8 FILLER_63_406 ();
 sg13g2_decap_8 FILLER_63_413 ();
 sg13g2_decap_8 FILLER_63_420 ();
 sg13g2_decap_8 FILLER_63_427 ();
 sg13g2_decap_8 FILLER_63_434 ();
 sg13g2_decap_8 FILLER_63_441 ();
 sg13g2_decap_8 FILLER_63_448 ();
 sg13g2_decap_8 FILLER_63_455 ();
 sg13g2_decap_8 FILLER_63_462 ();
 sg13g2_decap_8 FILLER_63_469 ();
 sg13g2_decap_8 FILLER_63_476 ();
 sg13g2_decap_8 FILLER_63_483 ();
 sg13g2_decap_8 FILLER_63_490 ();
 sg13g2_decap_8 FILLER_63_497 ();
 sg13g2_decap_8 FILLER_63_504 ();
 sg13g2_decap_8 FILLER_63_511 ();
 sg13g2_decap_8 FILLER_63_518 ();
 sg13g2_decap_8 FILLER_63_525 ();
 sg13g2_decap_8 FILLER_63_532 ();
 sg13g2_decap_8 FILLER_63_539 ();
 sg13g2_decap_8 FILLER_63_546 ();
 sg13g2_decap_8 FILLER_63_553 ();
 sg13g2_decap_8 FILLER_63_560 ();
 sg13g2_decap_8 FILLER_63_567 ();
 sg13g2_decap_8 FILLER_63_574 ();
 sg13g2_decap_8 FILLER_63_581 ();
 sg13g2_decap_8 FILLER_63_588 ();
 sg13g2_decap_8 FILLER_63_595 ();
 sg13g2_decap_8 FILLER_63_602 ();
 sg13g2_decap_8 FILLER_63_609 ();
 sg13g2_decap_8 FILLER_63_616 ();
 sg13g2_decap_8 FILLER_63_623 ();
 sg13g2_decap_8 FILLER_63_630 ();
 sg13g2_decap_8 FILLER_63_637 ();
 sg13g2_decap_8 FILLER_63_644 ();
 sg13g2_decap_8 FILLER_63_651 ();
 sg13g2_decap_8 FILLER_63_658 ();
 sg13g2_decap_8 FILLER_63_665 ();
 sg13g2_decap_8 FILLER_63_672 ();
 sg13g2_decap_8 FILLER_63_679 ();
 sg13g2_decap_8 FILLER_63_686 ();
 sg13g2_decap_8 FILLER_63_693 ();
 sg13g2_decap_8 FILLER_63_700 ();
 sg13g2_decap_8 FILLER_63_707 ();
 sg13g2_decap_8 FILLER_63_714 ();
 sg13g2_decap_8 FILLER_63_721 ();
 sg13g2_decap_8 FILLER_63_728 ();
 sg13g2_decap_8 FILLER_63_735 ();
 sg13g2_decap_8 FILLER_63_742 ();
 sg13g2_decap_8 FILLER_63_749 ();
 sg13g2_decap_8 FILLER_63_756 ();
 sg13g2_decap_8 FILLER_63_763 ();
 sg13g2_decap_8 FILLER_63_770 ();
 sg13g2_decap_8 FILLER_63_777 ();
 sg13g2_decap_8 FILLER_63_784 ();
 sg13g2_decap_8 FILLER_63_791 ();
 sg13g2_decap_8 FILLER_63_798 ();
 sg13g2_decap_8 FILLER_63_805 ();
 sg13g2_decap_8 FILLER_63_812 ();
 sg13g2_decap_8 FILLER_63_819 ();
 sg13g2_decap_8 FILLER_63_826 ();
 sg13g2_decap_8 FILLER_63_833 ();
 sg13g2_decap_8 FILLER_63_840 ();
 sg13g2_decap_8 FILLER_63_847 ();
 sg13g2_decap_8 FILLER_63_854 ();
 sg13g2_decap_8 FILLER_63_861 ();
 sg13g2_decap_8 FILLER_63_868 ();
 sg13g2_decap_8 FILLER_63_875 ();
 sg13g2_decap_8 FILLER_63_882 ();
 sg13g2_decap_8 FILLER_63_889 ();
 sg13g2_decap_8 FILLER_63_896 ();
 sg13g2_decap_8 FILLER_63_903 ();
 sg13g2_decap_8 FILLER_63_910 ();
 sg13g2_decap_8 FILLER_63_917 ();
 sg13g2_decap_8 FILLER_63_924 ();
 sg13g2_decap_8 FILLER_63_931 ();
 sg13g2_decap_8 FILLER_63_938 ();
 sg13g2_decap_8 FILLER_63_945 ();
 sg13g2_decap_8 FILLER_63_952 ();
 sg13g2_decap_8 FILLER_63_959 ();
 sg13g2_decap_8 FILLER_63_966 ();
 sg13g2_decap_8 FILLER_63_973 ();
 sg13g2_decap_8 FILLER_63_980 ();
 sg13g2_decap_8 FILLER_63_987 ();
 sg13g2_decap_8 FILLER_63_994 ();
 sg13g2_decap_8 FILLER_63_1001 ();
 sg13g2_decap_8 FILLER_63_1008 ();
 sg13g2_decap_8 FILLER_63_1015 ();
 sg13g2_decap_8 FILLER_63_1022 ();
 sg13g2_decap_8 FILLER_64_4 ();
 sg13g2_decap_8 FILLER_64_11 ();
 sg13g2_decap_8 FILLER_64_18 ();
 sg13g2_decap_8 FILLER_64_25 ();
 sg13g2_decap_8 FILLER_64_32 ();
 sg13g2_decap_8 FILLER_64_39 ();
 sg13g2_decap_8 FILLER_64_46 ();
 sg13g2_decap_8 FILLER_64_53 ();
 sg13g2_decap_8 FILLER_64_60 ();
 sg13g2_decap_8 FILLER_64_67 ();
 sg13g2_decap_8 FILLER_64_74 ();
 sg13g2_decap_8 FILLER_64_81 ();
 sg13g2_decap_8 FILLER_64_88 ();
 sg13g2_decap_8 FILLER_64_95 ();
 sg13g2_decap_8 FILLER_64_102 ();
 sg13g2_decap_8 FILLER_64_109 ();
 sg13g2_decap_8 FILLER_64_116 ();
 sg13g2_decap_8 FILLER_64_123 ();
 sg13g2_decap_8 FILLER_64_130 ();
 sg13g2_decap_8 FILLER_64_137 ();
 sg13g2_decap_8 FILLER_64_144 ();
 sg13g2_decap_8 FILLER_64_151 ();
 sg13g2_decap_8 FILLER_64_158 ();
 sg13g2_decap_8 FILLER_64_165 ();
 sg13g2_decap_8 FILLER_64_172 ();
 sg13g2_decap_8 FILLER_64_179 ();
 sg13g2_decap_8 FILLER_64_186 ();
 sg13g2_decap_8 FILLER_64_193 ();
 sg13g2_decap_8 FILLER_64_200 ();
 sg13g2_decap_8 FILLER_64_207 ();
 sg13g2_decap_8 FILLER_64_214 ();
 sg13g2_decap_8 FILLER_64_221 ();
 sg13g2_decap_8 FILLER_64_228 ();
 sg13g2_decap_8 FILLER_64_235 ();
 sg13g2_decap_8 FILLER_64_242 ();
 sg13g2_decap_8 FILLER_64_249 ();
 sg13g2_decap_8 FILLER_64_256 ();
 sg13g2_decap_8 FILLER_64_263 ();
 sg13g2_decap_8 FILLER_64_270 ();
 sg13g2_decap_8 FILLER_64_277 ();
 sg13g2_decap_8 FILLER_64_284 ();
 sg13g2_decap_8 FILLER_64_291 ();
 sg13g2_decap_8 FILLER_64_298 ();
 sg13g2_decap_8 FILLER_64_305 ();
 sg13g2_decap_8 FILLER_64_312 ();
 sg13g2_decap_8 FILLER_64_319 ();
 sg13g2_decap_8 FILLER_64_326 ();
 sg13g2_decap_8 FILLER_64_333 ();
 sg13g2_decap_8 FILLER_64_340 ();
 sg13g2_decap_8 FILLER_64_347 ();
 sg13g2_decap_8 FILLER_64_354 ();
 sg13g2_decap_8 FILLER_64_361 ();
 sg13g2_decap_8 FILLER_64_368 ();
 sg13g2_decap_8 FILLER_64_375 ();
 sg13g2_decap_8 FILLER_64_382 ();
 sg13g2_decap_8 FILLER_64_389 ();
 sg13g2_decap_8 FILLER_64_396 ();
 sg13g2_decap_8 FILLER_64_403 ();
 sg13g2_decap_8 FILLER_64_410 ();
 sg13g2_decap_8 FILLER_64_417 ();
 sg13g2_decap_8 FILLER_64_424 ();
 sg13g2_decap_8 FILLER_64_431 ();
 sg13g2_decap_8 FILLER_64_438 ();
 sg13g2_decap_8 FILLER_64_445 ();
 sg13g2_decap_8 FILLER_64_452 ();
 sg13g2_decap_8 FILLER_64_459 ();
 sg13g2_decap_8 FILLER_64_466 ();
 sg13g2_decap_8 FILLER_64_473 ();
 sg13g2_decap_8 FILLER_64_480 ();
 sg13g2_decap_8 FILLER_64_487 ();
 sg13g2_decap_8 FILLER_64_494 ();
 sg13g2_decap_8 FILLER_64_501 ();
 sg13g2_decap_8 FILLER_64_508 ();
 sg13g2_decap_8 FILLER_64_515 ();
 sg13g2_decap_8 FILLER_64_522 ();
 sg13g2_decap_8 FILLER_64_529 ();
 sg13g2_decap_8 FILLER_64_536 ();
 sg13g2_decap_8 FILLER_64_543 ();
 sg13g2_decap_8 FILLER_64_550 ();
 sg13g2_decap_8 FILLER_64_557 ();
 sg13g2_decap_8 FILLER_64_564 ();
 sg13g2_decap_8 FILLER_64_571 ();
 sg13g2_decap_8 FILLER_64_578 ();
 sg13g2_decap_8 FILLER_64_585 ();
 sg13g2_decap_8 FILLER_64_592 ();
 sg13g2_decap_8 FILLER_64_599 ();
 sg13g2_decap_8 FILLER_64_606 ();
 sg13g2_decap_8 FILLER_64_613 ();
 sg13g2_decap_8 FILLER_64_620 ();
 sg13g2_decap_8 FILLER_64_627 ();
 sg13g2_decap_8 FILLER_64_634 ();
 sg13g2_decap_8 FILLER_64_641 ();
 sg13g2_decap_8 FILLER_64_648 ();
 sg13g2_decap_8 FILLER_64_655 ();
 sg13g2_decap_8 FILLER_64_662 ();
 sg13g2_decap_8 FILLER_64_669 ();
 sg13g2_decap_8 FILLER_64_676 ();
 sg13g2_decap_8 FILLER_64_683 ();
 sg13g2_decap_8 FILLER_64_690 ();
 sg13g2_decap_8 FILLER_64_697 ();
 sg13g2_decap_8 FILLER_64_704 ();
 sg13g2_decap_8 FILLER_64_711 ();
 sg13g2_decap_8 FILLER_64_718 ();
 sg13g2_decap_8 FILLER_64_725 ();
 sg13g2_decap_8 FILLER_64_732 ();
 sg13g2_decap_8 FILLER_64_739 ();
 sg13g2_decap_8 FILLER_64_746 ();
 sg13g2_decap_8 FILLER_64_753 ();
 sg13g2_decap_8 FILLER_64_760 ();
 sg13g2_decap_8 FILLER_64_767 ();
 sg13g2_decap_8 FILLER_64_774 ();
 sg13g2_decap_8 FILLER_64_781 ();
 sg13g2_decap_8 FILLER_64_788 ();
 sg13g2_decap_8 FILLER_64_795 ();
 sg13g2_decap_8 FILLER_64_802 ();
 sg13g2_decap_8 FILLER_64_809 ();
 sg13g2_decap_8 FILLER_64_816 ();
 sg13g2_decap_8 FILLER_64_823 ();
 sg13g2_decap_8 FILLER_64_830 ();
 sg13g2_decap_8 FILLER_64_837 ();
 sg13g2_decap_8 FILLER_64_844 ();
 sg13g2_decap_8 FILLER_64_851 ();
 sg13g2_decap_8 FILLER_64_858 ();
 sg13g2_decap_8 FILLER_64_865 ();
 sg13g2_decap_8 FILLER_64_872 ();
 sg13g2_decap_8 FILLER_64_879 ();
 sg13g2_decap_8 FILLER_64_886 ();
 sg13g2_decap_8 FILLER_64_893 ();
 sg13g2_decap_8 FILLER_64_900 ();
 sg13g2_decap_8 FILLER_64_907 ();
 sg13g2_decap_8 FILLER_64_914 ();
 sg13g2_decap_8 FILLER_64_921 ();
 sg13g2_decap_8 FILLER_64_928 ();
 sg13g2_decap_8 FILLER_64_935 ();
 sg13g2_decap_8 FILLER_64_942 ();
 sg13g2_decap_8 FILLER_64_949 ();
 sg13g2_decap_8 FILLER_64_956 ();
 sg13g2_decap_8 FILLER_64_963 ();
 sg13g2_decap_8 FILLER_64_970 ();
 sg13g2_decap_8 FILLER_64_977 ();
 sg13g2_decap_8 FILLER_64_984 ();
 sg13g2_decap_8 FILLER_64_991 ();
 sg13g2_decap_8 FILLER_64_998 ();
 sg13g2_decap_8 FILLER_64_1005 ();
 sg13g2_decap_8 FILLER_64_1012 ();
 sg13g2_decap_8 FILLER_64_1019 ();
 sg13g2_fill_2 FILLER_64_1026 ();
 sg13g2_fill_1 FILLER_64_1028 ();
 sg13g2_decap_8 FILLER_65_0 ();
 sg13g2_decap_8 FILLER_65_7 ();
 sg13g2_decap_8 FILLER_65_14 ();
 sg13g2_decap_8 FILLER_65_21 ();
 sg13g2_decap_8 FILLER_65_28 ();
 sg13g2_decap_8 FILLER_65_35 ();
 sg13g2_decap_8 FILLER_65_42 ();
 sg13g2_decap_8 FILLER_65_49 ();
 sg13g2_decap_8 FILLER_65_56 ();
 sg13g2_decap_8 FILLER_65_63 ();
 sg13g2_decap_8 FILLER_65_70 ();
 sg13g2_decap_8 FILLER_65_77 ();
 sg13g2_decap_8 FILLER_65_84 ();
 sg13g2_decap_8 FILLER_65_91 ();
 sg13g2_decap_8 FILLER_65_98 ();
 sg13g2_decap_8 FILLER_65_105 ();
 sg13g2_decap_8 FILLER_65_112 ();
 sg13g2_decap_8 FILLER_65_119 ();
 sg13g2_decap_8 FILLER_65_126 ();
 sg13g2_decap_8 FILLER_65_133 ();
 sg13g2_decap_8 FILLER_65_140 ();
 sg13g2_decap_8 FILLER_65_147 ();
 sg13g2_decap_8 FILLER_65_154 ();
 sg13g2_decap_8 FILLER_65_161 ();
 sg13g2_decap_8 FILLER_65_168 ();
 sg13g2_decap_8 FILLER_65_175 ();
 sg13g2_decap_8 FILLER_65_182 ();
 sg13g2_decap_8 FILLER_65_189 ();
 sg13g2_decap_8 FILLER_65_196 ();
 sg13g2_decap_8 FILLER_65_203 ();
 sg13g2_decap_8 FILLER_65_210 ();
 sg13g2_decap_8 FILLER_65_217 ();
 sg13g2_decap_8 FILLER_65_224 ();
 sg13g2_decap_8 FILLER_65_231 ();
 sg13g2_decap_8 FILLER_65_238 ();
 sg13g2_decap_8 FILLER_65_245 ();
 sg13g2_decap_8 FILLER_65_252 ();
 sg13g2_decap_8 FILLER_65_259 ();
 sg13g2_decap_8 FILLER_65_266 ();
 sg13g2_decap_8 FILLER_65_273 ();
 sg13g2_decap_8 FILLER_65_280 ();
 sg13g2_decap_8 FILLER_65_287 ();
 sg13g2_decap_8 FILLER_65_294 ();
 sg13g2_decap_8 FILLER_65_301 ();
 sg13g2_decap_8 FILLER_65_308 ();
 sg13g2_decap_8 FILLER_65_315 ();
 sg13g2_decap_8 FILLER_65_322 ();
 sg13g2_decap_8 FILLER_65_329 ();
 sg13g2_decap_8 FILLER_65_336 ();
 sg13g2_decap_8 FILLER_65_343 ();
 sg13g2_decap_8 FILLER_65_350 ();
 sg13g2_decap_8 FILLER_65_357 ();
 sg13g2_decap_8 FILLER_65_364 ();
 sg13g2_decap_8 FILLER_65_371 ();
 sg13g2_decap_8 FILLER_65_378 ();
 sg13g2_decap_8 FILLER_65_385 ();
 sg13g2_decap_8 FILLER_65_392 ();
 sg13g2_decap_8 FILLER_65_399 ();
 sg13g2_decap_8 FILLER_65_406 ();
 sg13g2_decap_8 FILLER_65_413 ();
 sg13g2_decap_8 FILLER_65_420 ();
 sg13g2_decap_8 FILLER_65_427 ();
 sg13g2_decap_8 FILLER_65_434 ();
 sg13g2_decap_8 FILLER_65_441 ();
 sg13g2_decap_8 FILLER_65_448 ();
 sg13g2_decap_8 FILLER_65_455 ();
 sg13g2_decap_8 FILLER_65_462 ();
 sg13g2_decap_8 FILLER_65_469 ();
 sg13g2_decap_8 FILLER_65_476 ();
 sg13g2_decap_8 FILLER_65_483 ();
 sg13g2_decap_8 FILLER_65_490 ();
 sg13g2_decap_8 FILLER_65_497 ();
 sg13g2_decap_8 FILLER_65_504 ();
 sg13g2_decap_8 FILLER_65_511 ();
 sg13g2_decap_8 FILLER_65_518 ();
 sg13g2_decap_8 FILLER_65_525 ();
 sg13g2_decap_8 FILLER_65_532 ();
 sg13g2_decap_8 FILLER_65_539 ();
 sg13g2_decap_8 FILLER_65_546 ();
 sg13g2_decap_8 FILLER_65_553 ();
 sg13g2_decap_8 FILLER_65_560 ();
 sg13g2_decap_8 FILLER_65_567 ();
 sg13g2_decap_8 FILLER_65_574 ();
 sg13g2_decap_8 FILLER_65_581 ();
 sg13g2_decap_8 FILLER_65_588 ();
 sg13g2_decap_8 FILLER_65_595 ();
 sg13g2_decap_8 FILLER_65_602 ();
 sg13g2_decap_8 FILLER_65_609 ();
 sg13g2_decap_8 FILLER_65_616 ();
 sg13g2_decap_8 FILLER_65_623 ();
 sg13g2_decap_8 FILLER_65_630 ();
 sg13g2_decap_8 FILLER_65_637 ();
 sg13g2_decap_8 FILLER_65_644 ();
 sg13g2_decap_8 FILLER_65_651 ();
 sg13g2_decap_8 FILLER_65_658 ();
 sg13g2_decap_8 FILLER_65_665 ();
 sg13g2_decap_8 FILLER_65_672 ();
 sg13g2_decap_8 FILLER_65_679 ();
 sg13g2_decap_8 FILLER_65_686 ();
 sg13g2_decap_8 FILLER_65_693 ();
 sg13g2_decap_8 FILLER_65_700 ();
 sg13g2_decap_8 FILLER_65_707 ();
 sg13g2_decap_8 FILLER_65_714 ();
 sg13g2_decap_8 FILLER_65_721 ();
 sg13g2_decap_8 FILLER_65_728 ();
 sg13g2_decap_8 FILLER_65_735 ();
 sg13g2_decap_8 FILLER_65_742 ();
 sg13g2_decap_8 FILLER_65_749 ();
 sg13g2_decap_8 FILLER_65_756 ();
 sg13g2_decap_8 FILLER_65_763 ();
 sg13g2_decap_8 FILLER_65_770 ();
 sg13g2_decap_8 FILLER_65_777 ();
 sg13g2_decap_8 FILLER_65_784 ();
 sg13g2_decap_8 FILLER_65_791 ();
 sg13g2_decap_8 FILLER_65_798 ();
 sg13g2_decap_8 FILLER_65_805 ();
 sg13g2_decap_8 FILLER_65_812 ();
 sg13g2_decap_8 FILLER_65_819 ();
 sg13g2_decap_8 FILLER_65_826 ();
 sg13g2_decap_8 FILLER_65_833 ();
 sg13g2_decap_8 FILLER_65_840 ();
 sg13g2_decap_8 FILLER_65_847 ();
 sg13g2_decap_8 FILLER_65_854 ();
 sg13g2_decap_8 FILLER_65_861 ();
 sg13g2_decap_8 FILLER_65_868 ();
 sg13g2_decap_8 FILLER_65_875 ();
 sg13g2_decap_8 FILLER_65_882 ();
 sg13g2_decap_8 FILLER_65_889 ();
 sg13g2_decap_8 FILLER_65_896 ();
 sg13g2_decap_8 FILLER_65_903 ();
 sg13g2_decap_8 FILLER_65_910 ();
 sg13g2_decap_8 FILLER_65_917 ();
 sg13g2_decap_8 FILLER_65_924 ();
 sg13g2_decap_8 FILLER_65_931 ();
 sg13g2_decap_8 FILLER_65_938 ();
 sg13g2_decap_8 FILLER_65_945 ();
 sg13g2_decap_8 FILLER_65_952 ();
 sg13g2_decap_8 FILLER_65_959 ();
 sg13g2_decap_8 FILLER_65_966 ();
 sg13g2_decap_8 FILLER_65_973 ();
 sg13g2_decap_8 FILLER_65_980 ();
 sg13g2_decap_8 FILLER_65_987 ();
 sg13g2_decap_8 FILLER_65_994 ();
 sg13g2_decap_8 FILLER_65_1001 ();
 sg13g2_decap_8 FILLER_65_1008 ();
 sg13g2_decap_8 FILLER_65_1015 ();
 sg13g2_decap_8 FILLER_65_1022 ();
 sg13g2_decap_8 FILLER_66_4 ();
 sg13g2_decap_8 FILLER_66_11 ();
 sg13g2_fill_1 FILLER_66_18 ();
 sg13g2_decap_8 FILLER_66_27 ();
 sg13g2_decap_8 FILLER_66_34 ();
 sg13g2_decap_8 FILLER_66_41 ();
 sg13g2_decap_8 FILLER_66_48 ();
 sg13g2_decap_8 FILLER_66_55 ();
 sg13g2_decap_8 FILLER_66_62 ();
 sg13g2_decap_8 FILLER_66_69 ();
 sg13g2_decap_8 FILLER_66_76 ();
 sg13g2_decap_8 FILLER_66_83 ();
 sg13g2_decap_8 FILLER_66_90 ();
 sg13g2_decap_8 FILLER_66_97 ();
 sg13g2_decap_8 FILLER_66_104 ();
 sg13g2_decap_8 FILLER_66_111 ();
 sg13g2_decap_8 FILLER_66_118 ();
 sg13g2_decap_8 FILLER_66_125 ();
 sg13g2_decap_8 FILLER_66_132 ();
 sg13g2_decap_8 FILLER_66_139 ();
 sg13g2_decap_8 FILLER_66_146 ();
 sg13g2_decap_8 FILLER_66_153 ();
 sg13g2_decap_8 FILLER_66_160 ();
 sg13g2_decap_8 FILLER_66_167 ();
 sg13g2_decap_8 FILLER_66_174 ();
 sg13g2_decap_8 FILLER_66_181 ();
 sg13g2_decap_8 FILLER_66_188 ();
 sg13g2_decap_8 FILLER_66_195 ();
 sg13g2_decap_8 FILLER_66_202 ();
 sg13g2_decap_8 FILLER_66_209 ();
 sg13g2_decap_8 FILLER_66_216 ();
 sg13g2_decap_8 FILLER_66_223 ();
 sg13g2_decap_8 FILLER_66_230 ();
 sg13g2_decap_8 FILLER_66_237 ();
 sg13g2_decap_8 FILLER_66_244 ();
 sg13g2_decap_8 FILLER_66_251 ();
 sg13g2_decap_8 FILLER_66_258 ();
 sg13g2_decap_8 FILLER_66_265 ();
 sg13g2_decap_8 FILLER_66_272 ();
 sg13g2_decap_8 FILLER_66_279 ();
 sg13g2_decap_8 FILLER_66_286 ();
 sg13g2_decap_8 FILLER_66_293 ();
 sg13g2_decap_8 FILLER_66_300 ();
 sg13g2_decap_8 FILLER_66_307 ();
 sg13g2_decap_8 FILLER_66_314 ();
 sg13g2_decap_8 FILLER_66_321 ();
 sg13g2_decap_8 FILLER_66_328 ();
 sg13g2_decap_8 FILLER_66_335 ();
 sg13g2_decap_8 FILLER_66_342 ();
 sg13g2_decap_8 FILLER_66_349 ();
 sg13g2_decap_8 FILLER_66_356 ();
 sg13g2_decap_8 FILLER_66_363 ();
 sg13g2_decap_8 FILLER_66_370 ();
 sg13g2_decap_8 FILLER_66_377 ();
 sg13g2_decap_8 FILLER_66_384 ();
 sg13g2_decap_8 FILLER_66_391 ();
 sg13g2_decap_8 FILLER_66_398 ();
 sg13g2_decap_8 FILLER_66_405 ();
 sg13g2_decap_8 FILLER_66_412 ();
 sg13g2_decap_8 FILLER_66_419 ();
 sg13g2_decap_8 FILLER_66_426 ();
 sg13g2_decap_8 FILLER_66_433 ();
 sg13g2_decap_8 FILLER_66_440 ();
 sg13g2_decap_8 FILLER_66_447 ();
 sg13g2_decap_8 FILLER_66_454 ();
 sg13g2_decap_8 FILLER_66_461 ();
 sg13g2_decap_8 FILLER_66_468 ();
 sg13g2_decap_8 FILLER_66_475 ();
 sg13g2_decap_8 FILLER_66_482 ();
 sg13g2_decap_8 FILLER_66_489 ();
 sg13g2_decap_8 FILLER_66_496 ();
 sg13g2_decap_8 FILLER_66_503 ();
 sg13g2_decap_8 FILLER_66_510 ();
 sg13g2_decap_8 FILLER_66_517 ();
 sg13g2_decap_8 FILLER_66_524 ();
 sg13g2_decap_8 FILLER_66_531 ();
 sg13g2_decap_8 FILLER_66_538 ();
 sg13g2_decap_8 FILLER_66_545 ();
 sg13g2_decap_8 FILLER_66_552 ();
 sg13g2_decap_8 FILLER_66_559 ();
 sg13g2_decap_8 FILLER_66_566 ();
 sg13g2_decap_8 FILLER_66_573 ();
 sg13g2_decap_8 FILLER_66_580 ();
 sg13g2_decap_8 FILLER_66_587 ();
 sg13g2_decap_8 FILLER_66_594 ();
 sg13g2_decap_8 FILLER_66_601 ();
 sg13g2_decap_8 FILLER_66_608 ();
 sg13g2_decap_8 FILLER_66_615 ();
 sg13g2_decap_8 FILLER_66_622 ();
 sg13g2_decap_8 FILLER_66_629 ();
 sg13g2_decap_8 FILLER_66_636 ();
 sg13g2_decap_8 FILLER_66_643 ();
 sg13g2_decap_8 FILLER_66_650 ();
 sg13g2_decap_8 FILLER_66_657 ();
 sg13g2_decap_8 FILLER_66_664 ();
 sg13g2_decap_8 FILLER_66_671 ();
 sg13g2_decap_8 FILLER_66_678 ();
 sg13g2_decap_8 FILLER_66_685 ();
 sg13g2_decap_8 FILLER_66_692 ();
 sg13g2_decap_8 FILLER_66_699 ();
 sg13g2_decap_8 FILLER_66_706 ();
 sg13g2_decap_8 FILLER_66_713 ();
 sg13g2_decap_8 FILLER_66_720 ();
 sg13g2_decap_8 FILLER_66_727 ();
 sg13g2_decap_8 FILLER_66_734 ();
 sg13g2_decap_8 FILLER_66_741 ();
 sg13g2_decap_8 FILLER_66_748 ();
 sg13g2_decap_8 FILLER_66_755 ();
 sg13g2_decap_8 FILLER_66_762 ();
 sg13g2_decap_8 FILLER_66_769 ();
 sg13g2_decap_8 FILLER_66_776 ();
 sg13g2_decap_8 FILLER_66_783 ();
 sg13g2_decap_8 FILLER_66_790 ();
 sg13g2_decap_8 FILLER_66_797 ();
 sg13g2_decap_8 FILLER_66_804 ();
 sg13g2_decap_8 FILLER_66_811 ();
 sg13g2_decap_8 FILLER_66_818 ();
 sg13g2_decap_8 FILLER_66_825 ();
 sg13g2_decap_8 FILLER_66_832 ();
 sg13g2_decap_8 FILLER_66_839 ();
 sg13g2_decap_8 FILLER_66_846 ();
 sg13g2_decap_8 FILLER_66_853 ();
 sg13g2_decap_8 FILLER_66_860 ();
 sg13g2_decap_8 FILLER_66_867 ();
 sg13g2_decap_8 FILLER_66_874 ();
 sg13g2_decap_8 FILLER_66_881 ();
 sg13g2_decap_8 FILLER_66_888 ();
 sg13g2_decap_8 FILLER_66_895 ();
 sg13g2_decap_8 FILLER_66_902 ();
 sg13g2_decap_8 FILLER_66_909 ();
 sg13g2_decap_8 FILLER_66_916 ();
 sg13g2_decap_8 FILLER_66_923 ();
 sg13g2_decap_8 FILLER_66_930 ();
 sg13g2_decap_8 FILLER_66_937 ();
 sg13g2_decap_8 FILLER_66_944 ();
 sg13g2_decap_8 FILLER_66_951 ();
 sg13g2_decap_8 FILLER_66_958 ();
 sg13g2_decap_8 FILLER_66_965 ();
 sg13g2_decap_8 FILLER_66_972 ();
 sg13g2_decap_8 FILLER_66_979 ();
 sg13g2_decap_8 FILLER_66_986 ();
 sg13g2_decap_8 FILLER_66_993 ();
 sg13g2_decap_8 FILLER_66_1000 ();
 sg13g2_decap_8 FILLER_66_1007 ();
 sg13g2_decap_8 FILLER_66_1014 ();
 sg13g2_decap_8 FILLER_66_1021 ();
 sg13g2_fill_1 FILLER_66_1028 ();
 sg13g2_decap_8 FILLER_67_0 ();
 sg13g2_decap_8 FILLER_67_7 ();
 sg13g2_fill_1 FILLER_67_14 ();
 sg13g2_fill_2 FILLER_67_31 ();
 sg13g2_fill_1 FILLER_67_33 ();
 sg13g2_decap_8 FILLER_67_38 ();
 sg13g2_fill_2 FILLER_67_45 ();
 sg13g2_fill_1 FILLER_67_47 ();
 sg13g2_fill_2 FILLER_67_55 ();
 sg13g2_fill_1 FILLER_67_57 ();
 sg13g2_decap_8 FILLER_67_70 ();
 sg13g2_decap_8 FILLER_67_77 ();
 sg13g2_decap_8 FILLER_67_84 ();
 sg13g2_decap_8 FILLER_67_91 ();
 sg13g2_decap_8 FILLER_67_98 ();
 sg13g2_decap_8 FILLER_67_105 ();
 sg13g2_decap_8 FILLER_67_112 ();
 sg13g2_decap_8 FILLER_67_119 ();
 sg13g2_decap_8 FILLER_67_126 ();
 sg13g2_decap_8 FILLER_67_133 ();
 sg13g2_decap_8 FILLER_67_140 ();
 sg13g2_decap_8 FILLER_67_147 ();
 sg13g2_decap_8 FILLER_67_154 ();
 sg13g2_decap_8 FILLER_67_161 ();
 sg13g2_decap_8 FILLER_67_168 ();
 sg13g2_decap_8 FILLER_67_175 ();
 sg13g2_decap_8 FILLER_67_182 ();
 sg13g2_decap_8 FILLER_67_189 ();
 sg13g2_decap_8 FILLER_67_196 ();
 sg13g2_decap_8 FILLER_67_203 ();
 sg13g2_decap_8 FILLER_67_210 ();
 sg13g2_decap_8 FILLER_67_217 ();
 sg13g2_decap_8 FILLER_67_224 ();
 sg13g2_decap_8 FILLER_67_231 ();
 sg13g2_decap_8 FILLER_67_238 ();
 sg13g2_decap_8 FILLER_67_245 ();
 sg13g2_decap_8 FILLER_67_252 ();
 sg13g2_decap_8 FILLER_67_259 ();
 sg13g2_decap_8 FILLER_67_266 ();
 sg13g2_decap_8 FILLER_67_273 ();
 sg13g2_decap_8 FILLER_67_280 ();
 sg13g2_decap_8 FILLER_67_287 ();
 sg13g2_decap_8 FILLER_67_294 ();
 sg13g2_decap_8 FILLER_67_301 ();
 sg13g2_decap_8 FILLER_67_308 ();
 sg13g2_decap_8 FILLER_67_315 ();
 sg13g2_decap_8 FILLER_67_322 ();
 sg13g2_decap_8 FILLER_67_329 ();
 sg13g2_decap_8 FILLER_67_336 ();
 sg13g2_decap_8 FILLER_67_343 ();
 sg13g2_decap_8 FILLER_67_350 ();
 sg13g2_decap_8 FILLER_67_357 ();
 sg13g2_decap_8 FILLER_67_364 ();
 sg13g2_decap_8 FILLER_67_371 ();
 sg13g2_decap_8 FILLER_67_378 ();
 sg13g2_decap_8 FILLER_67_385 ();
 sg13g2_decap_8 FILLER_67_392 ();
 sg13g2_decap_8 FILLER_67_399 ();
 sg13g2_decap_8 FILLER_67_406 ();
 sg13g2_decap_8 FILLER_67_413 ();
 sg13g2_decap_8 FILLER_67_420 ();
 sg13g2_decap_8 FILLER_67_427 ();
 sg13g2_decap_8 FILLER_67_434 ();
 sg13g2_decap_8 FILLER_67_441 ();
 sg13g2_decap_8 FILLER_67_448 ();
 sg13g2_decap_8 FILLER_67_455 ();
 sg13g2_decap_8 FILLER_67_462 ();
 sg13g2_decap_8 FILLER_67_469 ();
 sg13g2_decap_8 FILLER_67_476 ();
 sg13g2_decap_8 FILLER_67_483 ();
 sg13g2_decap_8 FILLER_67_490 ();
 sg13g2_decap_8 FILLER_67_497 ();
 sg13g2_decap_8 FILLER_67_504 ();
 sg13g2_decap_8 FILLER_67_511 ();
 sg13g2_decap_8 FILLER_67_518 ();
 sg13g2_decap_8 FILLER_67_525 ();
 sg13g2_decap_8 FILLER_67_532 ();
 sg13g2_decap_8 FILLER_67_539 ();
 sg13g2_decap_8 FILLER_67_546 ();
 sg13g2_decap_8 FILLER_67_553 ();
 sg13g2_decap_8 FILLER_67_560 ();
 sg13g2_decap_8 FILLER_67_567 ();
 sg13g2_decap_8 FILLER_67_574 ();
 sg13g2_decap_8 FILLER_67_581 ();
 sg13g2_decap_8 FILLER_67_588 ();
 sg13g2_decap_8 FILLER_67_595 ();
 sg13g2_decap_8 FILLER_67_602 ();
 sg13g2_decap_8 FILLER_67_609 ();
 sg13g2_decap_8 FILLER_67_616 ();
 sg13g2_decap_8 FILLER_67_623 ();
 sg13g2_decap_8 FILLER_67_630 ();
 sg13g2_decap_8 FILLER_67_637 ();
 sg13g2_decap_8 FILLER_67_644 ();
 sg13g2_decap_8 FILLER_67_651 ();
 sg13g2_decap_8 FILLER_67_658 ();
 sg13g2_decap_8 FILLER_67_665 ();
 sg13g2_decap_8 FILLER_67_672 ();
 sg13g2_decap_8 FILLER_67_679 ();
 sg13g2_decap_8 FILLER_67_686 ();
 sg13g2_decap_8 FILLER_67_693 ();
 sg13g2_decap_8 FILLER_67_700 ();
 sg13g2_decap_8 FILLER_67_707 ();
 sg13g2_decap_8 FILLER_67_714 ();
 sg13g2_decap_8 FILLER_67_721 ();
 sg13g2_decap_8 FILLER_67_728 ();
 sg13g2_decap_8 FILLER_67_735 ();
 sg13g2_decap_8 FILLER_67_742 ();
 sg13g2_decap_8 FILLER_67_749 ();
 sg13g2_decap_8 FILLER_67_756 ();
 sg13g2_decap_8 FILLER_67_763 ();
 sg13g2_decap_8 FILLER_67_770 ();
 sg13g2_decap_8 FILLER_67_777 ();
 sg13g2_decap_8 FILLER_67_784 ();
 sg13g2_decap_8 FILLER_67_791 ();
 sg13g2_decap_8 FILLER_67_798 ();
 sg13g2_decap_8 FILLER_67_805 ();
 sg13g2_decap_8 FILLER_67_812 ();
 sg13g2_decap_8 FILLER_67_819 ();
 sg13g2_decap_8 FILLER_67_826 ();
 sg13g2_decap_8 FILLER_67_833 ();
 sg13g2_decap_8 FILLER_67_840 ();
 sg13g2_decap_8 FILLER_67_847 ();
 sg13g2_decap_8 FILLER_67_854 ();
 sg13g2_decap_8 FILLER_67_861 ();
 sg13g2_decap_8 FILLER_67_868 ();
 sg13g2_decap_8 FILLER_67_875 ();
 sg13g2_decap_8 FILLER_67_882 ();
 sg13g2_decap_8 FILLER_67_889 ();
 sg13g2_decap_8 FILLER_67_896 ();
 sg13g2_decap_8 FILLER_67_903 ();
 sg13g2_decap_8 FILLER_67_910 ();
 sg13g2_decap_8 FILLER_67_917 ();
 sg13g2_decap_8 FILLER_67_924 ();
 sg13g2_decap_8 FILLER_67_931 ();
 sg13g2_decap_8 FILLER_67_938 ();
 sg13g2_decap_8 FILLER_67_945 ();
 sg13g2_decap_8 FILLER_67_952 ();
 sg13g2_decap_8 FILLER_67_959 ();
 sg13g2_decap_8 FILLER_67_966 ();
 sg13g2_decap_8 FILLER_67_973 ();
 sg13g2_decap_8 FILLER_67_980 ();
 sg13g2_decap_8 FILLER_67_987 ();
 sg13g2_decap_8 FILLER_67_994 ();
 sg13g2_decap_8 FILLER_67_1001 ();
 sg13g2_decap_8 FILLER_67_1008 ();
 sg13g2_decap_8 FILLER_67_1015 ();
 sg13g2_decap_8 FILLER_67_1022 ();
 sg13g2_decap_8 FILLER_68_4 ();
 sg13g2_decap_8 FILLER_68_11 ();
 sg13g2_decap_8 FILLER_68_18 ();
 sg13g2_decap_8 FILLER_68_25 ();
 sg13g2_decap_8 FILLER_68_32 ();
 sg13g2_decap_8 FILLER_68_39 ();
 sg13g2_decap_4 FILLER_68_46 ();
 sg13g2_fill_2 FILLER_68_50 ();
 sg13g2_decap_8 FILLER_68_68 ();
 sg13g2_decap_8 FILLER_68_75 ();
 sg13g2_decap_8 FILLER_68_82 ();
 sg13g2_decap_8 FILLER_68_89 ();
 sg13g2_decap_8 FILLER_68_96 ();
 sg13g2_decap_8 FILLER_68_103 ();
 sg13g2_decap_8 FILLER_68_110 ();
 sg13g2_decap_8 FILLER_68_117 ();
 sg13g2_decap_8 FILLER_68_124 ();
 sg13g2_decap_8 FILLER_68_131 ();
 sg13g2_decap_8 FILLER_68_138 ();
 sg13g2_decap_8 FILLER_68_145 ();
 sg13g2_decap_8 FILLER_68_152 ();
 sg13g2_decap_8 FILLER_68_159 ();
 sg13g2_decap_8 FILLER_68_166 ();
 sg13g2_decap_8 FILLER_68_173 ();
 sg13g2_decap_8 FILLER_68_180 ();
 sg13g2_decap_8 FILLER_68_187 ();
 sg13g2_decap_8 FILLER_68_194 ();
 sg13g2_decap_8 FILLER_68_201 ();
 sg13g2_decap_8 FILLER_68_208 ();
 sg13g2_decap_8 FILLER_68_215 ();
 sg13g2_decap_8 FILLER_68_222 ();
 sg13g2_decap_8 FILLER_68_229 ();
 sg13g2_decap_8 FILLER_68_236 ();
 sg13g2_decap_8 FILLER_68_243 ();
 sg13g2_decap_8 FILLER_68_250 ();
 sg13g2_decap_8 FILLER_68_257 ();
 sg13g2_decap_8 FILLER_68_264 ();
 sg13g2_decap_8 FILLER_68_271 ();
 sg13g2_decap_8 FILLER_68_278 ();
 sg13g2_decap_8 FILLER_68_285 ();
 sg13g2_decap_8 FILLER_68_292 ();
 sg13g2_decap_8 FILLER_68_299 ();
 sg13g2_decap_8 FILLER_68_306 ();
 sg13g2_decap_8 FILLER_68_313 ();
 sg13g2_decap_8 FILLER_68_320 ();
 sg13g2_decap_8 FILLER_68_327 ();
 sg13g2_decap_8 FILLER_68_334 ();
 sg13g2_decap_8 FILLER_68_341 ();
 sg13g2_decap_8 FILLER_68_348 ();
 sg13g2_decap_8 FILLER_68_355 ();
 sg13g2_decap_8 FILLER_68_362 ();
 sg13g2_decap_8 FILLER_68_369 ();
 sg13g2_decap_8 FILLER_68_376 ();
 sg13g2_decap_8 FILLER_68_383 ();
 sg13g2_decap_8 FILLER_68_390 ();
 sg13g2_decap_8 FILLER_68_397 ();
 sg13g2_decap_8 FILLER_68_404 ();
 sg13g2_decap_8 FILLER_68_411 ();
 sg13g2_decap_8 FILLER_68_418 ();
 sg13g2_decap_8 FILLER_68_425 ();
 sg13g2_decap_8 FILLER_68_432 ();
 sg13g2_decap_8 FILLER_68_439 ();
 sg13g2_decap_8 FILLER_68_446 ();
 sg13g2_decap_8 FILLER_68_453 ();
 sg13g2_decap_8 FILLER_68_460 ();
 sg13g2_decap_8 FILLER_68_467 ();
 sg13g2_decap_8 FILLER_68_474 ();
 sg13g2_decap_8 FILLER_68_481 ();
 sg13g2_decap_8 FILLER_68_488 ();
 sg13g2_decap_8 FILLER_68_495 ();
 sg13g2_decap_8 FILLER_68_502 ();
 sg13g2_decap_8 FILLER_68_509 ();
 sg13g2_decap_8 FILLER_68_516 ();
 sg13g2_decap_8 FILLER_68_523 ();
 sg13g2_decap_8 FILLER_68_530 ();
 sg13g2_decap_8 FILLER_68_537 ();
 sg13g2_decap_8 FILLER_68_544 ();
 sg13g2_decap_8 FILLER_68_551 ();
 sg13g2_decap_8 FILLER_68_558 ();
 sg13g2_decap_8 FILLER_68_565 ();
 sg13g2_decap_8 FILLER_68_572 ();
 sg13g2_decap_8 FILLER_68_579 ();
 sg13g2_decap_8 FILLER_68_586 ();
 sg13g2_decap_8 FILLER_68_593 ();
 sg13g2_decap_8 FILLER_68_600 ();
 sg13g2_decap_8 FILLER_68_607 ();
 sg13g2_decap_8 FILLER_68_614 ();
 sg13g2_decap_8 FILLER_68_621 ();
 sg13g2_decap_8 FILLER_68_628 ();
 sg13g2_decap_8 FILLER_68_635 ();
 sg13g2_decap_8 FILLER_68_642 ();
 sg13g2_decap_8 FILLER_68_649 ();
 sg13g2_decap_8 FILLER_68_656 ();
 sg13g2_decap_8 FILLER_68_663 ();
 sg13g2_decap_8 FILLER_68_670 ();
 sg13g2_decap_8 FILLER_68_677 ();
 sg13g2_decap_8 FILLER_68_684 ();
 sg13g2_decap_8 FILLER_68_691 ();
 sg13g2_decap_8 FILLER_68_698 ();
 sg13g2_decap_8 FILLER_68_705 ();
 sg13g2_decap_8 FILLER_68_712 ();
 sg13g2_decap_8 FILLER_68_719 ();
 sg13g2_decap_8 FILLER_68_726 ();
 sg13g2_decap_8 FILLER_68_733 ();
 sg13g2_decap_8 FILLER_68_740 ();
 sg13g2_decap_8 FILLER_68_747 ();
 sg13g2_decap_8 FILLER_68_754 ();
 sg13g2_decap_8 FILLER_68_761 ();
 sg13g2_decap_8 FILLER_68_768 ();
 sg13g2_decap_8 FILLER_68_775 ();
 sg13g2_decap_8 FILLER_68_782 ();
 sg13g2_decap_8 FILLER_68_789 ();
 sg13g2_decap_8 FILLER_68_796 ();
 sg13g2_decap_8 FILLER_68_803 ();
 sg13g2_decap_8 FILLER_68_810 ();
 sg13g2_decap_8 FILLER_68_817 ();
 sg13g2_decap_8 FILLER_68_824 ();
 sg13g2_decap_8 FILLER_68_831 ();
 sg13g2_decap_8 FILLER_68_838 ();
 sg13g2_decap_8 FILLER_68_845 ();
 sg13g2_decap_8 FILLER_68_852 ();
 sg13g2_decap_8 FILLER_68_859 ();
 sg13g2_decap_8 FILLER_68_866 ();
 sg13g2_decap_8 FILLER_68_873 ();
 sg13g2_decap_8 FILLER_68_880 ();
 sg13g2_decap_8 FILLER_68_887 ();
 sg13g2_decap_8 FILLER_68_894 ();
 sg13g2_decap_8 FILLER_68_901 ();
 sg13g2_decap_8 FILLER_68_908 ();
 sg13g2_decap_8 FILLER_68_915 ();
 sg13g2_decap_8 FILLER_68_922 ();
 sg13g2_decap_8 FILLER_68_929 ();
 sg13g2_decap_8 FILLER_68_936 ();
 sg13g2_decap_8 FILLER_68_943 ();
 sg13g2_decap_8 FILLER_68_950 ();
 sg13g2_decap_8 FILLER_68_957 ();
 sg13g2_decap_8 FILLER_68_964 ();
 sg13g2_decap_8 FILLER_68_971 ();
 sg13g2_decap_8 FILLER_68_978 ();
 sg13g2_decap_8 FILLER_68_985 ();
 sg13g2_decap_8 FILLER_68_992 ();
 sg13g2_decap_8 FILLER_68_999 ();
 sg13g2_decap_8 FILLER_68_1006 ();
 sg13g2_decap_8 FILLER_68_1013 ();
 sg13g2_decap_8 FILLER_68_1020 ();
 sg13g2_fill_2 FILLER_68_1027 ();
 sg13g2_decap_8 FILLER_69_0 ();
 sg13g2_decap_8 FILLER_69_7 ();
 sg13g2_decap_8 FILLER_69_14 ();
 sg13g2_decap_8 FILLER_69_21 ();
 sg13g2_decap_8 FILLER_69_28 ();
 sg13g2_decap_8 FILLER_69_35 ();
 sg13g2_decap_8 FILLER_69_42 ();
 sg13g2_decap_8 FILLER_69_49 ();
 sg13g2_decap_4 FILLER_69_56 ();
 sg13g2_decap_8 FILLER_69_64 ();
 sg13g2_decap_8 FILLER_69_71 ();
 sg13g2_decap_8 FILLER_69_78 ();
 sg13g2_decap_8 FILLER_69_85 ();
 sg13g2_decap_8 FILLER_69_92 ();
 sg13g2_decap_8 FILLER_69_99 ();
 sg13g2_decap_8 FILLER_69_106 ();
 sg13g2_decap_8 FILLER_69_113 ();
 sg13g2_decap_8 FILLER_69_120 ();
 sg13g2_decap_8 FILLER_69_127 ();
 sg13g2_decap_8 FILLER_69_134 ();
 sg13g2_decap_8 FILLER_69_141 ();
 sg13g2_decap_8 FILLER_69_148 ();
 sg13g2_decap_8 FILLER_69_155 ();
 sg13g2_decap_8 FILLER_69_162 ();
 sg13g2_decap_8 FILLER_69_169 ();
 sg13g2_decap_8 FILLER_69_176 ();
 sg13g2_decap_8 FILLER_69_183 ();
 sg13g2_decap_8 FILLER_69_190 ();
 sg13g2_decap_8 FILLER_69_197 ();
 sg13g2_decap_8 FILLER_69_204 ();
 sg13g2_decap_8 FILLER_69_211 ();
 sg13g2_decap_8 FILLER_69_218 ();
 sg13g2_decap_8 FILLER_69_225 ();
 sg13g2_decap_8 FILLER_69_232 ();
 sg13g2_decap_8 FILLER_69_239 ();
 sg13g2_decap_8 FILLER_69_246 ();
 sg13g2_decap_8 FILLER_69_253 ();
 sg13g2_decap_8 FILLER_69_260 ();
 sg13g2_decap_8 FILLER_69_267 ();
 sg13g2_decap_8 FILLER_69_274 ();
 sg13g2_decap_8 FILLER_69_281 ();
 sg13g2_decap_8 FILLER_69_288 ();
 sg13g2_decap_8 FILLER_69_295 ();
 sg13g2_decap_8 FILLER_69_302 ();
 sg13g2_decap_8 FILLER_69_309 ();
 sg13g2_decap_8 FILLER_69_316 ();
 sg13g2_decap_8 FILLER_69_323 ();
 sg13g2_decap_8 FILLER_69_330 ();
 sg13g2_decap_8 FILLER_69_337 ();
 sg13g2_decap_8 FILLER_69_344 ();
 sg13g2_decap_8 FILLER_69_351 ();
 sg13g2_decap_8 FILLER_69_358 ();
 sg13g2_decap_8 FILLER_69_365 ();
 sg13g2_decap_8 FILLER_69_372 ();
 sg13g2_decap_8 FILLER_69_379 ();
 sg13g2_decap_8 FILLER_69_386 ();
 sg13g2_decap_8 FILLER_69_393 ();
 sg13g2_decap_8 FILLER_69_400 ();
 sg13g2_decap_8 FILLER_69_407 ();
 sg13g2_decap_8 FILLER_69_414 ();
 sg13g2_decap_8 FILLER_69_421 ();
 sg13g2_decap_8 FILLER_69_428 ();
 sg13g2_decap_8 FILLER_69_435 ();
 sg13g2_decap_8 FILLER_69_442 ();
 sg13g2_decap_8 FILLER_69_449 ();
 sg13g2_decap_8 FILLER_69_456 ();
 sg13g2_decap_8 FILLER_69_463 ();
 sg13g2_decap_8 FILLER_69_470 ();
 sg13g2_decap_8 FILLER_69_477 ();
 sg13g2_decap_8 FILLER_69_484 ();
 sg13g2_decap_8 FILLER_69_491 ();
 sg13g2_decap_8 FILLER_69_498 ();
 sg13g2_decap_8 FILLER_69_505 ();
 sg13g2_decap_8 FILLER_69_512 ();
 sg13g2_decap_8 FILLER_69_519 ();
 sg13g2_decap_8 FILLER_69_526 ();
 sg13g2_decap_8 FILLER_69_533 ();
 sg13g2_decap_8 FILLER_69_540 ();
 sg13g2_decap_8 FILLER_69_547 ();
 sg13g2_decap_8 FILLER_69_554 ();
 sg13g2_decap_8 FILLER_69_561 ();
 sg13g2_decap_8 FILLER_69_568 ();
 sg13g2_decap_8 FILLER_69_575 ();
 sg13g2_decap_8 FILLER_69_582 ();
 sg13g2_decap_8 FILLER_69_589 ();
 sg13g2_decap_8 FILLER_69_596 ();
 sg13g2_decap_8 FILLER_69_603 ();
 sg13g2_decap_8 FILLER_69_610 ();
 sg13g2_decap_8 FILLER_69_617 ();
 sg13g2_decap_8 FILLER_69_624 ();
 sg13g2_decap_8 FILLER_69_631 ();
 sg13g2_decap_8 FILLER_69_638 ();
 sg13g2_decap_8 FILLER_69_645 ();
 sg13g2_decap_8 FILLER_69_652 ();
 sg13g2_decap_8 FILLER_69_659 ();
 sg13g2_decap_8 FILLER_69_666 ();
 sg13g2_decap_8 FILLER_69_673 ();
 sg13g2_decap_8 FILLER_69_680 ();
 sg13g2_decap_8 FILLER_69_687 ();
 sg13g2_decap_8 FILLER_69_694 ();
 sg13g2_decap_8 FILLER_69_701 ();
 sg13g2_decap_8 FILLER_69_708 ();
 sg13g2_decap_8 FILLER_69_715 ();
 sg13g2_decap_8 FILLER_69_722 ();
 sg13g2_decap_8 FILLER_69_729 ();
 sg13g2_decap_8 FILLER_69_736 ();
 sg13g2_decap_8 FILLER_69_743 ();
 sg13g2_decap_8 FILLER_69_750 ();
 sg13g2_decap_8 FILLER_69_757 ();
 sg13g2_decap_8 FILLER_69_764 ();
 sg13g2_decap_8 FILLER_69_771 ();
 sg13g2_decap_8 FILLER_69_778 ();
 sg13g2_decap_8 FILLER_69_785 ();
 sg13g2_decap_8 FILLER_69_792 ();
 sg13g2_decap_8 FILLER_69_799 ();
 sg13g2_decap_8 FILLER_69_806 ();
 sg13g2_decap_8 FILLER_69_813 ();
 sg13g2_decap_8 FILLER_69_820 ();
 sg13g2_decap_8 FILLER_69_827 ();
 sg13g2_decap_8 FILLER_69_834 ();
 sg13g2_decap_8 FILLER_69_841 ();
 sg13g2_decap_8 FILLER_69_848 ();
 sg13g2_decap_8 FILLER_69_855 ();
 sg13g2_decap_8 FILLER_69_862 ();
 sg13g2_decap_8 FILLER_69_869 ();
 sg13g2_decap_8 FILLER_69_876 ();
 sg13g2_decap_8 FILLER_69_883 ();
 sg13g2_decap_8 FILLER_69_890 ();
 sg13g2_decap_8 FILLER_69_897 ();
 sg13g2_decap_8 FILLER_69_904 ();
 sg13g2_decap_8 FILLER_69_911 ();
 sg13g2_decap_8 FILLER_69_918 ();
 sg13g2_decap_8 FILLER_69_925 ();
 sg13g2_decap_8 FILLER_69_932 ();
 sg13g2_decap_8 FILLER_69_939 ();
 sg13g2_decap_8 FILLER_69_946 ();
 sg13g2_decap_8 FILLER_69_953 ();
 sg13g2_decap_8 FILLER_69_960 ();
 sg13g2_decap_8 FILLER_69_967 ();
 sg13g2_decap_8 FILLER_69_974 ();
 sg13g2_decap_8 FILLER_69_981 ();
 sg13g2_decap_8 FILLER_69_988 ();
 sg13g2_decap_8 FILLER_69_995 ();
 sg13g2_decap_8 FILLER_69_1002 ();
 sg13g2_decap_8 FILLER_69_1009 ();
 sg13g2_decap_8 FILLER_69_1016 ();
 sg13g2_decap_4 FILLER_69_1023 ();
 sg13g2_fill_2 FILLER_69_1027 ();
 sg13g2_decap_8 FILLER_70_0 ();
 sg13g2_decap_8 FILLER_70_7 ();
 sg13g2_decap_8 FILLER_70_14 ();
 sg13g2_decap_8 FILLER_70_21 ();
 sg13g2_decap_8 FILLER_70_28 ();
 sg13g2_decap_8 FILLER_70_35 ();
 sg13g2_decap_8 FILLER_70_42 ();
 sg13g2_decap_8 FILLER_70_49 ();
 sg13g2_decap_8 FILLER_70_56 ();
 sg13g2_decap_8 FILLER_70_63 ();
 sg13g2_decap_8 FILLER_70_70 ();
 sg13g2_decap_8 FILLER_70_77 ();
 sg13g2_decap_8 FILLER_70_84 ();
 sg13g2_decap_8 FILLER_70_91 ();
 sg13g2_decap_8 FILLER_70_98 ();
 sg13g2_decap_8 FILLER_70_105 ();
 sg13g2_decap_8 FILLER_70_112 ();
 sg13g2_decap_8 FILLER_70_119 ();
 sg13g2_decap_8 FILLER_70_126 ();
 sg13g2_decap_8 FILLER_70_133 ();
 sg13g2_decap_8 FILLER_70_140 ();
 sg13g2_decap_8 FILLER_70_147 ();
 sg13g2_decap_8 FILLER_70_154 ();
 sg13g2_decap_8 FILLER_70_161 ();
 sg13g2_decap_8 FILLER_70_168 ();
 sg13g2_decap_8 FILLER_70_175 ();
 sg13g2_decap_8 FILLER_70_182 ();
 sg13g2_decap_8 FILLER_70_189 ();
 sg13g2_decap_8 FILLER_70_196 ();
 sg13g2_decap_8 FILLER_70_203 ();
 sg13g2_decap_8 FILLER_70_210 ();
 sg13g2_decap_8 FILLER_70_217 ();
 sg13g2_decap_8 FILLER_70_224 ();
 sg13g2_decap_8 FILLER_70_231 ();
 sg13g2_decap_8 FILLER_70_238 ();
 sg13g2_decap_8 FILLER_70_245 ();
 sg13g2_decap_8 FILLER_70_252 ();
 sg13g2_decap_8 FILLER_70_259 ();
 sg13g2_decap_8 FILLER_70_266 ();
 sg13g2_decap_8 FILLER_70_273 ();
 sg13g2_decap_8 FILLER_70_280 ();
 sg13g2_decap_8 FILLER_70_287 ();
 sg13g2_decap_8 FILLER_70_294 ();
 sg13g2_decap_8 FILLER_70_301 ();
 sg13g2_decap_8 FILLER_70_308 ();
 sg13g2_decap_8 FILLER_70_315 ();
 sg13g2_decap_8 FILLER_70_322 ();
 sg13g2_decap_8 FILLER_70_329 ();
 sg13g2_decap_8 FILLER_70_336 ();
 sg13g2_decap_8 FILLER_70_343 ();
 sg13g2_decap_8 FILLER_70_350 ();
 sg13g2_decap_8 FILLER_70_357 ();
 sg13g2_decap_8 FILLER_70_364 ();
 sg13g2_decap_8 FILLER_70_371 ();
 sg13g2_decap_8 FILLER_70_378 ();
 sg13g2_decap_8 FILLER_70_385 ();
 sg13g2_decap_8 FILLER_70_392 ();
 sg13g2_decap_8 FILLER_70_399 ();
 sg13g2_decap_8 FILLER_70_406 ();
 sg13g2_decap_8 FILLER_70_413 ();
 sg13g2_decap_8 FILLER_70_420 ();
 sg13g2_decap_8 FILLER_70_427 ();
 sg13g2_decap_8 FILLER_70_434 ();
 sg13g2_decap_8 FILLER_70_441 ();
 sg13g2_decap_8 FILLER_70_448 ();
 sg13g2_decap_8 FILLER_70_455 ();
 sg13g2_decap_8 FILLER_70_462 ();
 sg13g2_decap_8 FILLER_70_469 ();
 sg13g2_decap_8 FILLER_70_476 ();
 sg13g2_decap_8 FILLER_70_483 ();
 sg13g2_decap_8 FILLER_70_490 ();
 sg13g2_decap_8 FILLER_70_497 ();
 sg13g2_decap_8 FILLER_70_504 ();
 sg13g2_decap_8 FILLER_70_511 ();
 sg13g2_decap_8 FILLER_70_518 ();
 sg13g2_decap_8 FILLER_70_525 ();
 sg13g2_decap_8 FILLER_70_532 ();
 sg13g2_decap_8 FILLER_70_539 ();
 sg13g2_decap_8 FILLER_70_546 ();
 sg13g2_decap_8 FILLER_70_553 ();
 sg13g2_decap_8 FILLER_70_560 ();
 sg13g2_decap_8 FILLER_70_567 ();
 sg13g2_decap_8 FILLER_70_574 ();
 sg13g2_decap_8 FILLER_70_581 ();
 sg13g2_decap_8 FILLER_70_588 ();
 sg13g2_decap_8 FILLER_70_595 ();
 sg13g2_decap_8 FILLER_70_602 ();
 sg13g2_decap_8 FILLER_70_609 ();
 sg13g2_decap_8 FILLER_70_616 ();
 sg13g2_decap_8 FILLER_70_623 ();
 sg13g2_decap_8 FILLER_70_630 ();
 sg13g2_decap_8 FILLER_70_637 ();
 sg13g2_decap_8 FILLER_70_644 ();
 sg13g2_decap_8 FILLER_70_651 ();
 sg13g2_decap_8 FILLER_70_658 ();
 sg13g2_decap_8 FILLER_70_665 ();
 sg13g2_decap_8 FILLER_70_672 ();
 sg13g2_decap_8 FILLER_70_679 ();
 sg13g2_decap_8 FILLER_70_686 ();
 sg13g2_decap_8 FILLER_70_693 ();
 sg13g2_decap_8 FILLER_70_700 ();
 sg13g2_decap_8 FILLER_70_707 ();
 sg13g2_decap_8 FILLER_70_714 ();
 sg13g2_decap_8 FILLER_70_721 ();
 sg13g2_decap_8 FILLER_70_728 ();
 sg13g2_decap_8 FILLER_70_735 ();
 sg13g2_decap_8 FILLER_70_742 ();
 sg13g2_decap_8 FILLER_70_749 ();
 sg13g2_decap_8 FILLER_70_756 ();
 sg13g2_decap_8 FILLER_70_763 ();
 sg13g2_decap_8 FILLER_70_770 ();
 sg13g2_decap_8 FILLER_70_777 ();
 sg13g2_decap_8 FILLER_70_784 ();
 sg13g2_decap_8 FILLER_70_791 ();
 sg13g2_decap_8 FILLER_70_798 ();
 sg13g2_decap_8 FILLER_70_805 ();
 sg13g2_decap_8 FILLER_70_812 ();
 sg13g2_decap_8 FILLER_70_819 ();
 sg13g2_decap_8 FILLER_70_826 ();
 sg13g2_decap_8 FILLER_70_833 ();
 sg13g2_decap_8 FILLER_70_840 ();
 sg13g2_decap_8 FILLER_70_847 ();
 sg13g2_decap_8 FILLER_70_854 ();
 sg13g2_decap_8 FILLER_70_861 ();
 sg13g2_decap_8 FILLER_70_868 ();
 sg13g2_decap_8 FILLER_70_875 ();
 sg13g2_decap_8 FILLER_70_882 ();
 sg13g2_decap_8 FILLER_70_889 ();
 sg13g2_decap_8 FILLER_70_896 ();
 sg13g2_decap_8 FILLER_70_903 ();
 sg13g2_decap_8 FILLER_70_910 ();
 sg13g2_decap_8 FILLER_70_917 ();
 sg13g2_decap_8 FILLER_70_924 ();
 sg13g2_decap_8 FILLER_70_931 ();
 sg13g2_decap_8 FILLER_70_938 ();
 sg13g2_decap_8 FILLER_70_945 ();
 sg13g2_decap_8 FILLER_70_952 ();
 sg13g2_decap_8 FILLER_70_959 ();
 sg13g2_decap_8 FILLER_70_966 ();
 sg13g2_decap_8 FILLER_70_973 ();
 sg13g2_decap_8 FILLER_70_980 ();
 sg13g2_decap_8 FILLER_70_987 ();
 sg13g2_decap_8 FILLER_70_994 ();
 sg13g2_decap_8 FILLER_70_1001 ();
 sg13g2_decap_8 FILLER_70_1008 ();
 sg13g2_decap_8 FILLER_70_1015 ();
 sg13g2_decap_8 FILLER_70_1022 ();
 sg13g2_decap_8 FILLER_71_4 ();
 sg13g2_decap_8 FILLER_71_11 ();
 sg13g2_decap_8 FILLER_71_18 ();
 sg13g2_decap_8 FILLER_71_25 ();
 sg13g2_decap_8 FILLER_71_32 ();
 sg13g2_decap_8 FILLER_71_39 ();
 sg13g2_decap_8 FILLER_71_46 ();
 sg13g2_decap_8 FILLER_71_53 ();
 sg13g2_decap_8 FILLER_71_60 ();
 sg13g2_decap_8 FILLER_71_67 ();
 sg13g2_decap_8 FILLER_71_74 ();
 sg13g2_decap_8 FILLER_71_81 ();
 sg13g2_decap_8 FILLER_71_88 ();
 sg13g2_decap_8 FILLER_71_95 ();
 sg13g2_decap_8 FILLER_71_102 ();
 sg13g2_decap_8 FILLER_71_109 ();
 sg13g2_decap_8 FILLER_71_116 ();
 sg13g2_decap_8 FILLER_71_123 ();
 sg13g2_decap_8 FILLER_71_130 ();
 sg13g2_decap_8 FILLER_71_137 ();
 sg13g2_decap_8 FILLER_71_144 ();
 sg13g2_decap_8 FILLER_71_151 ();
 sg13g2_decap_8 FILLER_71_158 ();
 sg13g2_decap_8 FILLER_71_165 ();
 sg13g2_decap_8 FILLER_71_172 ();
 sg13g2_decap_8 FILLER_71_179 ();
 sg13g2_decap_8 FILLER_71_186 ();
 sg13g2_decap_8 FILLER_71_193 ();
 sg13g2_decap_8 FILLER_71_200 ();
 sg13g2_decap_8 FILLER_71_207 ();
 sg13g2_decap_8 FILLER_71_214 ();
 sg13g2_decap_8 FILLER_71_221 ();
 sg13g2_decap_8 FILLER_71_228 ();
 sg13g2_decap_8 FILLER_71_235 ();
 sg13g2_decap_8 FILLER_71_242 ();
 sg13g2_decap_8 FILLER_71_249 ();
 sg13g2_decap_8 FILLER_71_256 ();
 sg13g2_decap_8 FILLER_71_263 ();
 sg13g2_decap_8 FILLER_71_270 ();
 sg13g2_decap_8 FILLER_71_277 ();
 sg13g2_decap_8 FILLER_71_284 ();
 sg13g2_decap_8 FILLER_71_291 ();
 sg13g2_decap_8 FILLER_71_298 ();
 sg13g2_decap_8 FILLER_71_305 ();
 sg13g2_decap_8 FILLER_71_312 ();
 sg13g2_decap_8 FILLER_71_319 ();
 sg13g2_decap_8 FILLER_71_326 ();
 sg13g2_decap_8 FILLER_71_333 ();
 sg13g2_decap_8 FILLER_71_340 ();
 sg13g2_decap_8 FILLER_71_347 ();
 sg13g2_decap_8 FILLER_71_354 ();
 sg13g2_decap_8 FILLER_71_361 ();
 sg13g2_decap_8 FILLER_71_368 ();
 sg13g2_decap_8 FILLER_71_375 ();
 sg13g2_decap_8 FILLER_71_382 ();
 sg13g2_decap_8 FILLER_71_389 ();
 sg13g2_decap_8 FILLER_71_396 ();
 sg13g2_decap_8 FILLER_71_403 ();
 sg13g2_decap_8 FILLER_71_410 ();
 sg13g2_decap_8 FILLER_71_417 ();
 sg13g2_decap_8 FILLER_71_424 ();
 sg13g2_decap_8 FILLER_71_431 ();
 sg13g2_decap_8 FILLER_71_438 ();
 sg13g2_decap_8 FILLER_71_445 ();
 sg13g2_decap_8 FILLER_71_452 ();
 sg13g2_decap_8 FILLER_71_459 ();
 sg13g2_decap_8 FILLER_71_466 ();
 sg13g2_decap_8 FILLER_71_473 ();
 sg13g2_decap_8 FILLER_71_480 ();
 sg13g2_decap_8 FILLER_71_487 ();
 sg13g2_decap_8 FILLER_71_494 ();
 sg13g2_decap_8 FILLER_71_501 ();
 sg13g2_decap_8 FILLER_71_508 ();
 sg13g2_decap_8 FILLER_71_515 ();
 sg13g2_decap_8 FILLER_71_522 ();
 sg13g2_decap_8 FILLER_71_529 ();
 sg13g2_decap_8 FILLER_71_536 ();
 sg13g2_decap_8 FILLER_71_543 ();
 sg13g2_decap_8 FILLER_71_550 ();
 sg13g2_decap_8 FILLER_71_557 ();
 sg13g2_decap_8 FILLER_71_564 ();
 sg13g2_decap_8 FILLER_71_571 ();
 sg13g2_decap_8 FILLER_71_578 ();
 sg13g2_decap_8 FILLER_71_585 ();
 sg13g2_decap_8 FILLER_71_592 ();
 sg13g2_decap_8 FILLER_71_599 ();
 sg13g2_decap_8 FILLER_71_606 ();
 sg13g2_decap_8 FILLER_71_613 ();
 sg13g2_decap_8 FILLER_71_620 ();
 sg13g2_decap_8 FILLER_71_627 ();
 sg13g2_decap_8 FILLER_71_634 ();
 sg13g2_decap_8 FILLER_71_641 ();
 sg13g2_decap_8 FILLER_71_648 ();
 sg13g2_decap_8 FILLER_71_655 ();
 sg13g2_decap_8 FILLER_71_662 ();
 sg13g2_decap_8 FILLER_71_669 ();
 sg13g2_decap_8 FILLER_71_676 ();
 sg13g2_decap_8 FILLER_71_683 ();
 sg13g2_decap_8 FILLER_71_690 ();
 sg13g2_decap_8 FILLER_71_697 ();
 sg13g2_decap_8 FILLER_71_704 ();
 sg13g2_decap_8 FILLER_71_711 ();
 sg13g2_decap_8 FILLER_71_718 ();
 sg13g2_decap_8 FILLER_71_725 ();
 sg13g2_decap_8 FILLER_71_732 ();
 sg13g2_decap_8 FILLER_71_739 ();
 sg13g2_decap_8 FILLER_71_746 ();
 sg13g2_decap_8 FILLER_71_753 ();
 sg13g2_decap_8 FILLER_71_760 ();
 sg13g2_decap_8 FILLER_71_767 ();
 sg13g2_decap_8 FILLER_71_774 ();
 sg13g2_decap_8 FILLER_71_781 ();
 sg13g2_decap_8 FILLER_71_788 ();
 sg13g2_decap_8 FILLER_71_795 ();
 sg13g2_decap_8 FILLER_71_802 ();
 sg13g2_decap_8 FILLER_71_809 ();
 sg13g2_decap_8 FILLER_71_816 ();
 sg13g2_decap_8 FILLER_71_823 ();
 sg13g2_decap_8 FILLER_71_830 ();
 sg13g2_decap_8 FILLER_71_837 ();
 sg13g2_decap_8 FILLER_71_844 ();
 sg13g2_decap_8 FILLER_71_851 ();
 sg13g2_decap_8 FILLER_71_858 ();
 sg13g2_decap_8 FILLER_71_865 ();
 sg13g2_decap_8 FILLER_71_872 ();
 sg13g2_decap_8 FILLER_71_879 ();
 sg13g2_decap_8 FILLER_71_886 ();
 sg13g2_decap_8 FILLER_71_893 ();
 sg13g2_decap_8 FILLER_71_900 ();
 sg13g2_decap_8 FILLER_71_907 ();
 sg13g2_decap_8 FILLER_71_914 ();
 sg13g2_decap_8 FILLER_71_921 ();
 sg13g2_decap_8 FILLER_71_928 ();
 sg13g2_decap_8 FILLER_71_935 ();
 sg13g2_decap_8 FILLER_71_942 ();
 sg13g2_decap_8 FILLER_71_949 ();
 sg13g2_decap_8 FILLER_71_956 ();
 sg13g2_decap_8 FILLER_71_963 ();
 sg13g2_decap_8 FILLER_71_970 ();
 sg13g2_decap_8 FILLER_71_977 ();
 sg13g2_decap_8 FILLER_71_984 ();
 sg13g2_decap_8 FILLER_71_991 ();
 sg13g2_decap_8 FILLER_71_998 ();
 sg13g2_decap_8 FILLER_71_1005 ();
 sg13g2_decap_8 FILLER_71_1012 ();
 sg13g2_decap_8 FILLER_71_1019 ();
 sg13g2_fill_2 FILLER_71_1026 ();
 sg13g2_fill_1 FILLER_71_1028 ();
 sg13g2_decap_8 FILLER_72_0 ();
 sg13g2_decap_8 FILLER_72_7 ();
 sg13g2_decap_8 FILLER_72_14 ();
 sg13g2_decap_8 FILLER_72_21 ();
 sg13g2_decap_8 FILLER_72_28 ();
 sg13g2_decap_8 FILLER_72_35 ();
 sg13g2_decap_8 FILLER_72_42 ();
 sg13g2_decap_8 FILLER_72_49 ();
 sg13g2_decap_8 FILLER_72_56 ();
 sg13g2_decap_8 FILLER_72_63 ();
 sg13g2_decap_8 FILLER_72_70 ();
 sg13g2_decap_8 FILLER_72_77 ();
 sg13g2_decap_8 FILLER_72_84 ();
 sg13g2_decap_8 FILLER_72_91 ();
 sg13g2_decap_8 FILLER_72_98 ();
 sg13g2_decap_8 FILLER_72_105 ();
 sg13g2_decap_8 FILLER_72_112 ();
 sg13g2_decap_8 FILLER_72_119 ();
 sg13g2_decap_8 FILLER_72_126 ();
 sg13g2_decap_8 FILLER_72_133 ();
 sg13g2_decap_8 FILLER_72_140 ();
 sg13g2_decap_8 FILLER_72_147 ();
 sg13g2_decap_8 FILLER_72_154 ();
 sg13g2_decap_8 FILLER_72_161 ();
 sg13g2_decap_8 FILLER_72_168 ();
 sg13g2_decap_8 FILLER_72_175 ();
 sg13g2_decap_8 FILLER_72_182 ();
 sg13g2_decap_8 FILLER_72_189 ();
 sg13g2_decap_8 FILLER_72_196 ();
 sg13g2_decap_8 FILLER_72_203 ();
 sg13g2_decap_8 FILLER_72_210 ();
 sg13g2_decap_8 FILLER_72_217 ();
 sg13g2_decap_8 FILLER_72_224 ();
 sg13g2_decap_8 FILLER_72_231 ();
 sg13g2_decap_8 FILLER_72_238 ();
 sg13g2_decap_8 FILLER_72_245 ();
 sg13g2_decap_8 FILLER_72_252 ();
 sg13g2_decap_8 FILLER_72_259 ();
 sg13g2_decap_8 FILLER_72_266 ();
 sg13g2_decap_8 FILLER_72_273 ();
 sg13g2_decap_8 FILLER_72_280 ();
 sg13g2_decap_8 FILLER_72_287 ();
 sg13g2_decap_8 FILLER_72_294 ();
 sg13g2_decap_8 FILLER_72_301 ();
 sg13g2_decap_8 FILLER_72_308 ();
 sg13g2_decap_8 FILLER_72_315 ();
 sg13g2_decap_8 FILLER_72_322 ();
 sg13g2_decap_8 FILLER_72_329 ();
 sg13g2_decap_8 FILLER_72_336 ();
 sg13g2_decap_8 FILLER_72_343 ();
 sg13g2_decap_8 FILLER_72_350 ();
 sg13g2_decap_8 FILLER_72_357 ();
 sg13g2_decap_8 FILLER_72_364 ();
 sg13g2_decap_8 FILLER_72_371 ();
 sg13g2_decap_8 FILLER_72_378 ();
 sg13g2_decap_8 FILLER_72_385 ();
 sg13g2_decap_8 FILLER_72_392 ();
 sg13g2_decap_8 FILLER_72_399 ();
 sg13g2_decap_8 FILLER_72_406 ();
 sg13g2_decap_8 FILLER_72_413 ();
 sg13g2_decap_8 FILLER_72_420 ();
 sg13g2_decap_8 FILLER_72_427 ();
 sg13g2_decap_8 FILLER_72_434 ();
 sg13g2_decap_8 FILLER_72_441 ();
 sg13g2_decap_8 FILLER_72_448 ();
 sg13g2_decap_8 FILLER_72_455 ();
 sg13g2_decap_8 FILLER_72_462 ();
 sg13g2_decap_8 FILLER_72_469 ();
 sg13g2_decap_8 FILLER_72_476 ();
 sg13g2_decap_8 FILLER_72_483 ();
 sg13g2_decap_8 FILLER_72_490 ();
 sg13g2_decap_8 FILLER_72_497 ();
 sg13g2_decap_8 FILLER_72_504 ();
 sg13g2_decap_8 FILLER_72_511 ();
 sg13g2_decap_8 FILLER_72_518 ();
 sg13g2_decap_8 FILLER_72_525 ();
 sg13g2_decap_8 FILLER_72_532 ();
 sg13g2_decap_8 FILLER_72_539 ();
 sg13g2_decap_8 FILLER_72_546 ();
 sg13g2_decap_8 FILLER_72_553 ();
 sg13g2_decap_8 FILLER_72_560 ();
 sg13g2_decap_8 FILLER_72_567 ();
 sg13g2_decap_8 FILLER_72_574 ();
 sg13g2_decap_8 FILLER_72_581 ();
 sg13g2_decap_8 FILLER_72_588 ();
 sg13g2_decap_8 FILLER_72_595 ();
 sg13g2_decap_8 FILLER_72_602 ();
 sg13g2_decap_8 FILLER_72_609 ();
 sg13g2_decap_8 FILLER_72_616 ();
 sg13g2_decap_8 FILLER_72_623 ();
 sg13g2_decap_8 FILLER_72_630 ();
 sg13g2_decap_8 FILLER_72_637 ();
 sg13g2_decap_8 FILLER_72_644 ();
 sg13g2_decap_8 FILLER_72_651 ();
 sg13g2_decap_8 FILLER_72_658 ();
 sg13g2_decap_8 FILLER_72_665 ();
 sg13g2_decap_8 FILLER_72_672 ();
 sg13g2_decap_8 FILLER_72_679 ();
 sg13g2_decap_8 FILLER_72_686 ();
 sg13g2_decap_8 FILLER_72_693 ();
 sg13g2_decap_8 FILLER_72_700 ();
 sg13g2_decap_8 FILLER_72_707 ();
 sg13g2_decap_8 FILLER_72_714 ();
 sg13g2_decap_8 FILLER_72_721 ();
 sg13g2_decap_8 FILLER_72_728 ();
 sg13g2_decap_8 FILLER_72_735 ();
 sg13g2_decap_8 FILLER_72_742 ();
 sg13g2_decap_8 FILLER_72_749 ();
 sg13g2_decap_8 FILLER_72_756 ();
 sg13g2_decap_8 FILLER_72_763 ();
 sg13g2_decap_8 FILLER_72_770 ();
 sg13g2_decap_8 FILLER_72_777 ();
 sg13g2_decap_8 FILLER_72_784 ();
 sg13g2_decap_8 FILLER_72_791 ();
 sg13g2_decap_8 FILLER_72_798 ();
 sg13g2_decap_8 FILLER_72_805 ();
 sg13g2_decap_8 FILLER_72_812 ();
 sg13g2_decap_8 FILLER_72_819 ();
 sg13g2_decap_8 FILLER_72_826 ();
 sg13g2_decap_8 FILLER_72_833 ();
 sg13g2_decap_8 FILLER_72_840 ();
 sg13g2_decap_8 FILLER_72_847 ();
 sg13g2_decap_8 FILLER_72_854 ();
 sg13g2_decap_8 FILLER_72_861 ();
 sg13g2_decap_8 FILLER_72_868 ();
 sg13g2_decap_8 FILLER_72_875 ();
 sg13g2_decap_8 FILLER_72_882 ();
 sg13g2_decap_8 FILLER_72_889 ();
 sg13g2_decap_8 FILLER_72_896 ();
 sg13g2_decap_8 FILLER_72_903 ();
 sg13g2_decap_8 FILLER_72_910 ();
 sg13g2_decap_8 FILLER_72_917 ();
 sg13g2_decap_8 FILLER_72_924 ();
 sg13g2_decap_8 FILLER_72_931 ();
 sg13g2_decap_8 FILLER_72_938 ();
 sg13g2_decap_8 FILLER_72_945 ();
 sg13g2_decap_8 FILLER_72_952 ();
 sg13g2_decap_8 FILLER_72_959 ();
 sg13g2_decap_8 FILLER_72_966 ();
 sg13g2_decap_8 FILLER_72_973 ();
 sg13g2_decap_8 FILLER_72_980 ();
 sg13g2_decap_8 FILLER_72_987 ();
 sg13g2_decap_8 FILLER_72_994 ();
 sg13g2_decap_8 FILLER_72_1001 ();
 sg13g2_decap_8 FILLER_72_1008 ();
 sg13g2_decap_8 FILLER_72_1015 ();
 sg13g2_decap_8 FILLER_72_1022 ();
 sg13g2_decap_8 FILLER_73_4 ();
 sg13g2_decap_8 FILLER_73_11 ();
 sg13g2_decap_8 FILLER_73_18 ();
 sg13g2_decap_8 FILLER_73_25 ();
 sg13g2_decap_8 FILLER_73_32 ();
 sg13g2_decap_8 FILLER_73_39 ();
 sg13g2_decap_8 FILLER_73_46 ();
 sg13g2_decap_4 FILLER_73_53 ();
 sg13g2_fill_2 FILLER_73_57 ();
 sg13g2_decap_8 FILLER_73_67 ();
 sg13g2_decap_8 FILLER_73_74 ();
 sg13g2_decap_8 FILLER_73_81 ();
 sg13g2_decap_8 FILLER_73_88 ();
 sg13g2_decap_8 FILLER_73_95 ();
 sg13g2_decap_8 FILLER_73_102 ();
 sg13g2_decap_8 FILLER_73_109 ();
 sg13g2_decap_8 FILLER_73_116 ();
 sg13g2_decap_8 FILLER_73_123 ();
 sg13g2_decap_8 FILLER_73_130 ();
 sg13g2_decap_8 FILLER_73_137 ();
 sg13g2_decap_8 FILLER_73_144 ();
 sg13g2_decap_8 FILLER_73_151 ();
 sg13g2_decap_8 FILLER_73_158 ();
 sg13g2_decap_8 FILLER_73_165 ();
 sg13g2_decap_8 FILLER_73_172 ();
 sg13g2_decap_8 FILLER_73_179 ();
 sg13g2_decap_8 FILLER_73_186 ();
 sg13g2_decap_8 FILLER_73_193 ();
 sg13g2_decap_8 FILLER_73_200 ();
 sg13g2_decap_8 FILLER_73_207 ();
 sg13g2_decap_8 FILLER_73_214 ();
 sg13g2_decap_8 FILLER_73_221 ();
 sg13g2_decap_8 FILLER_73_228 ();
 sg13g2_decap_8 FILLER_73_235 ();
 sg13g2_decap_8 FILLER_73_242 ();
 sg13g2_decap_8 FILLER_73_249 ();
 sg13g2_decap_8 FILLER_73_256 ();
 sg13g2_decap_8 FILLER_73_263 ();
 sg13g2_decap_8 FILLER_73_270 ();
 sg13g2_decap_8 FILLER_73_277 ();
 sg13g2_decap_8 FILLER_73_284 ();
 sg13g2_decap_8 FILLER_73_291 ();
 sg13g2_decap_8 FILLER_73_298 ();
 sg13g2_decap_8 FILLER_73_305 ();
 sg13g2_decap_8 FILLER_73_312 ();
 sg13g2_decap_8 FILLER_73_319 ();
 sg13g2_decap_8 FILLER_73_326 ();
 sg13g2_decap_8 FILLER_73_333 ();
 sg13g2_decap_8 FILLER_73_340 ();
 sg13g2_decap_8 FILLER_73_347 ();
 sg13g2_decap_8 FILLER_73_354 ();
 sg13g2_decap_8 FILLER_73_361 ();
 sg13g2_decap_8 FILLER_73_368 ();
 sg13g2_decap_8 FILLER_73_375 ();
 sg13g2_decap_8 FILLER_73_382 ();
 sg13g2_decap_8 FILLER_73_389 ();
 sg13g2_decap_8 FILLER_73_396 ();
 sg13g2_decap_8 FILLER_73_403 ();
 sg13g2_decap_8 FILLER_73_410 ();
 sg13g2_decap_8 FILLER_73_417 ();
 sg13g2_decap_8 FILLER_73_424 ();
 sg13g2_decap_8 FILLER_73_431 ();
 sg13g2_decap_8 FILLER_73_438 ();
 sg13g2_decap_8 FILLER_73_445 ();
 sg13g2_decap_8 FILLER_73_452 ();
 sg13g2_decap_8 FILLER_73_459 ();
 sg13g2_decap_8 FILLER_73_466 ();
 sg13g2_decap_8 FILLER_73_473 ();
 sg13g2_decap_8 FILLER_73_480 ();
 sg13g2_decap_8 FILLER_73_487 ();
 sg13g2_decap_8 FILLER_73_494 ();
 sg13g2_decap_8 FILLER_73_501 ();
 sg13g2_decap_8 FILLER_73_508 ();
 sg13g2_decap_8 FILLER_73_515 ();
 sg13g2_decap_8 FILLER_73_522 ();
 sg13g2_decap_8 FILLER_73_529 ();
 sg13g2_decap_8 FILLER_73_536 ();
 sg13g2_decap_8 FILLER_73_543 ();
 sg13g2_decap_8 FILLER_73_550 ();
 sg13g2_decap_8 FILLER_73_557 ();
 sg13g2_decap_8 FILLER_73_564 ();
 sg13g2_decap_8 FILLER_73_571 ();
 sg13g2_decap_8 FILLER_73_578 ();
 sg13g2_decap_8 FILLER_73_585 ();
 sg13g2_decap_8 FILLER_73_592 ();
 sg13g2_decap_8 FILLER_73_599 ();
 sg13g2_decap_8 FILLER_73_606 ();
 sg13g2_decap_8 FILLER_73_613 ();
 sg13g2_decap_8 FILLER_73_620 ();
 sg13g2_decap_8 FILLER_73_627 ();
 sg13g2_decap_8 FILLER_73_634 ();
 sg13g2_decap_8 FILLER_73_641 ();
 sg13g2_decap_8 FILLER_73_648 ();
 sg13g2_decap_8 FILLER_73_655 ();
 sg13g2_decap_8 FILLER_73_662 ();
 sg13g2_decap_8 FILLER_73_669 ();
 sg13g2_decap_8 FILLER_73_676 ();
 sg13g2_decap_8 FILLER_73_683 ();
 sg13g2_decap_8 FILLER_73_690 ();
 sg13g2_decap_8 FILLER_73_697 ();
 sg13g2_decap_8 FILLER_73_704 ();
 sg13g2_decap_8 FILLER_73_711 ();
 sg13g2_decap_8 FILLER_73_718 ();
 sg13g2_decap_8 FILLER_73_725 ();
 sg13g2_decap_8 FILLER_73_732 ();
 sg13g2_decap_8 FILLER_73_739 ();
 sg13g2_decap_8 FILLER_73_746 ();
 sg13g2_decap_8 FILLER_73_753 ();
 sg13g2_decap_8 FILLER_73_760 ();
 sg13g2_decap_8 FILLER_73_767 ();
 sg13g2_decap_8 FILLER_73_774 ();
 sg13g2_decap_8 FILLER_73_781 ();
 sg13g2_decap_8 FILLER_73_788 ();
 sg13g2_decap_8 FILLER_73_795 ();
 sg13g2_decap_8 FILLER_73_802 ();
 sg13g2_decap_8 FILLER_73_809 ();
 sg13g2_decap_8 FILLER_73_816 ();
 sg13g2_decap_8 FILLER_73_823 ();
 sg13g2_decap_8 FILLER_73_830 ();
 sg13g2_decap_8 FILLER_73_837 ();
 sg13g2_decap_8 FILLER_73_844 ();
 sg13g2_decap_8 FILLER_73_851 ();
 sg13g2_decap_8 FILLER_73_858 ();
 sg13g2_decap_8 FILLER_73_865 ();
 sg13g2_decap_8 FILLER_73_872 ();
 sg13g2_decap_8 FILLER_73_879 ();
 sg13g2_decap_8 FILLER_73_886 ();
 sg13g2_decap_8 FILLER_73_893 ();
 sg13g2_decap_8 FILLER_73_900 ();
 sg13g2_decap_8 FILLER_73_907 ();
 sg13g2_decap_8 FILLER_73_914 ();
 sg13g2_decap_8 FILLER_73_921 ();
 sg13g2_decap_8 FILLER_73_928 ();
 sg13g2_decap_8 FILLER_73_935 ();
 sg13g2_decap_8 FILLER_73_942 ();
 sg13g2_decap_8 FILLER_73_949 ();
 sg13g2_decap_8 FILLER_73_956 ();
 sg13g2_decap_8 FILLER_73_963 ();
 sg13g2_decap_8 FILLER_73_970 ();
 sg13g2_decap_8 FILLER_73_977 ();
 sg13g2_decap_8 FILLER_73_984 ();
 sg13g2_decap_8 FILLER_73_991 ();
 sg13g2_decap_8 FILLER_73_998 ();
 sg13g2_decap_8 FILLER_73_1005 ();
 sg13g2_decap_8 FILLER_73_1012 ();
 sg13g2_decap_8 FILLER_73_1019 ();
 sg13g2_fill_2 FILLER_73_1026 ();
 sg13g2_fill_1 FILLER_73_1028 ();
 sg13g2_decap_8 FILLER_74_0 ();
 sg13g2_decap_8 FILLER_74_7 ();
 sg13g2_decap_8 FILLER_74_14 ();
 sg13g2_decap_8 FILLER_74_21 ();
 sg13g2_decap_8 FILLER_74_28 ();
 sg13g2_decap_8 FILLER_74_35 ();
 sg13g2_decap_8 FILLER_74_42 ();
 sg13g2_decap_4 FILLER_74_49 ();
 sg13g2_fill_1 FILLER_74_53 ();
 sg13g2_decap_8 FILLER_74_71 ();
 sg13g2_decap_8 FILLER_74_78 ();
 sg13g2_decap_8 FILLER_74_85 ();
 sg13g2_decap_8 FILLER_74_92 ();
 sg13g2_decap_8 FILLER_74_99 ();
 sg13g2_decap_8 FILLER_74_106 ();
 sg13g2_decap_8 FILLER_74_113 ();
 sg13g2_decap_8 FILLER_74_120 ();
 sg13g2_decap_8 FILLER_74_127 ();
 sg13g2_decap_8 FILLER_74_134 ();
 sg13g2_decap_8 FILLER_74_141 ();
 sg13g2_decap_8 FILLER_74_148 ();
 sg13g2_decap_8 FILLER_74_155 ();
 sg13g2_decap_8 FILLER_74_162 ();
 sg13g2_decap_8 FILLER_74_169 ();
 sg13g2_decap_8 FILLER_74_176 ();
 sg13g2_decap_8 FILLER_74_183 ();
 sg13g2_decap_8 FILLER_74_190 ();
 sg13g2_decap_8 FILLER_74_197 ();
 sg13g2_decap_8 FILLER_74_204 ();
 sg13g2_decap_8 FILLER_74_211 ();
 sg13g2_decap_8 FILLER_74_218 ();
 sg13g2_decap_8 FILLER_74_225 ();
 sg13g2_decap_8 FILLER_74_232 ();
 sg13g2_decap_8 FILLER_74_239 ();
 sg13g2_decap_8 FILLER_74_246 ();
 sg13g2_decap_8 FILLER_74_253 ();
 sg13g2_decap_8 FILLER_74_260 ();
 sg13g2_decap_8 FILLER_74_267 ();
 sg13g2_decap_8 FILLER_74_274 ();
 sg13g2_decap_8 FILLER_74_281 ();
 sg13g2_decap_8 FILLER_74_288 ();
 sg13g2_decap_8 FILLER_74_295 ();
 sg13g2_decap_8 FILLER_74_302 ();
 sg13g2_decap_8 FILLER_74_309 ();
 sg13g2_decap_8 FILLER_74_316 ();
 sg13g2_decap_8 FILLER_74_323 ();
 sg13g2_decap_8 FILLER_74_330 ();
 sg13g2_decap_8 FILLER_74_337 ();
 sg13g2_decap_8 FILLER_74_344 ();
 sg13g2_decap_8 FILLER_74_351 ();
 sg13g2_decap_8 FILLER_74_358 ();
 sg13g2_decap_8 FILLER_74_365 ();
 sg13g2_decap_8 FILLER_74_372 ();
 sg13g2_decap_8 FILLER_74_379 ();
 sg13g2_decap_8 FILLER_74_386 ();
 sg13g2_decap_8 FILLER_74_393 ();
 sg13g2_decap_8 FILLER_74_400 ();
 sg13g2_decap_8 FILLER_74_407 ();
 sg13g2_decap_8 FILLER_74_414 ();
 sg13g2_decap_8 FILLER_74_421 ();
 sg13g2_decap_8 FILLER_74_428 ();
 sg13g2_decap_8 FILLER_74_435 ();
 sg13g2_decap_8 FILLER_74_442 ();
 sg13g2_decap_8 FILLER_74_449 ();
 sg13g2_decap_8 FILLER_74_456 ();
 sg13g2_decap_8 FILLER_74_463 ();
 sg13g2_decap_8 FILLER_74_470 ();
 sg13g2_decap_8 FILLER_74_477 ();
 sg13g2_decap_8 FILLER_74_484 ();
 sg13g2_decap_8 FILLER_74_491 ();
 sg13g2_decap_8 FILLER_74_498 ();
 sg13g2_decap_8 FILLER_74_505 ();
 sg13g2_decap_8 FILLER_74_512 ();
 sg13g2_decap_8 FILLER_74_519 ();
 sg13g2_decap_8 FILLER_74_526 ();
 sg13g2_decap_8 FILLER_74_533 ();
 sg13g2_decap_8 FILLER_74_540 ();
 sg13g2_decap_8 FILLER_74_547 ();
 sg13g2_decap_8 FILLER_74_554 ();
 sg13g2_decap_8 FILLER_74_561 ();
 sg13g2_decap_8 FILLER_74_568 ();
 sg13g2_decap_8 FILLER_74_575 ();
 sg13g2_decap_8 FILLER_74_582 ();
 sg13g2_decap_8 FILLER_74_589 ();
 sg13g2_decap_8 FILLER_74_596 ();
 sg13g2_decap_8 FILLER_74_603 ();
 sg13g2_decap_8 FILLER_74_610 ();
 sg13g2_decap_8 FILLER_74_617 ();
 sg13g2_decap_8 FILLER_74_624 ();
 sg13g2_decap_8 FILLER_74_631 ();
 sg13g2_decap_8 FILLER_74_638 ();
 sg13g2_decap_8 FILLER_74_645 ();
 sg13g2_decap_8 FILLER_74_652 ();
 sg13g2_decap_8 FILLER_74_659 ();
 sg13g2_decap_8 FILLER_74_666 ();
 sg13g2_decap_8 FILLER_74_673 ();
 sg13g2_decap_8 FILLER_74_680 ();
 sg13g2_decap_8 FILLER_74_687 ();
 sg13g2_decap_8 FILLER_74_694 ();
 sg13g2_decap_8 FILLER_74_701 ();
 sg13g2_decap_8 FILLER_74_708 ();
 sg13g2_decap_8 FILLER_74_715 ();
 sg13g2_decap_8 FILLER_74_722 ();
 sg13g2_decap_8 FILLER_74_729 ();
 sg13g2_decap_8 FILLER_74_736 ();
 sg13g2_decap_8 FILLER_74_743 ();
 sg13g2_decap_8 FILLER_74_750 ();
 sg13g2_decap_8 FILLER_74_757 ();
 sg13g2_decap_8 FILLER_74_764 ();
 sg13g2_decap_8 FILLER_74_771 ();
 sg13g2_decap_8 FILLER_74_778 ();
 sg13g2_decap_8 FILLER_74_785 ();
 sg13g2_decap_8 FILLER_74_792 ();
 sg13g2_decap_8 FILLER_74_799 ();
 sg13g2_decap_8 FILLER_74_806 ();
 sg13g2_decap_8 FILLER_74_813 ();
 sg13g2_decap_8 FILLER_74_820 ();
 sg13g2_decap_8 FILLER_74_827 ();
 sg13g2_decap_8 FILLER_74_834 ();
 sg13g2_decap_8 FILLER_74_841 ();
 sg13g2_decap_8 FILLER_74_848 ();
 sg13g2_decap_8 FILLER_74_855 ();
 sg13g2_decap_8 FILLER_74_862 ();
 sg13g2_decap_8 FILLER_74_869 ();
 sg13g2_decap_8 FILLER_74_876 ();
 sg13g2_decap_8 FILLER_74_883 ();
 sg13g2_decap_8 FILLER_74_890 ();
 sg13g2_decap_8 FILLER_74_897 ();
 sg13g2_decap_8 FILLER_74_904 ();
 sg13g2_decap_8 FILLER_74_911 ();
 sg13g2_decap_8 FILLER_74_918 ();
 sg13g2_decap_8 FILLER_74_925 ();
 sg13g2_decap_8 FILLER_74_932 ();
 sg13g2_decap_8 FILLER_74_939 ();
 sg13g2_decap_8 FILLER_74_946 ();
 sg13g2_decap_8 FILLER_74_953 ();
 sg13g2_decap_8 FILLER_74_960 ();
 sg13g2_decap_8 FILLER_74_967 ();
 sg13g2_decap_8 FILLER_74_974 ();
 sg13g2_decap_8 FILLER_74_981 ();
 sg13g2_decap_8 FILLER_74_988 ();
 sg13g2_decap_8 FILLER_74_995 ();
 sg13g2_decap_8 FILLER_74_1002 ();
 sg13g2_decap_8 FILLER_74_1009 ();
 sg13g2_decap_8 FILLER_74_1016 ();
 sg13g2_decap_4 FILLER_74_1023 ();
 sg13g2_fill_2 FILLER_74_1027 ();
 sg13g2_decap_8 FILLER_75_0 ();
 sg13g2_decap_8 FILLER_75_7 ();
 sg13g2_decap_8 FILLER_75_14 ();
 sg13g2_decap_8 FILLER_75_21 ();
 sg13g2_decap_8 FILLER_75_28 ();
 sg13g2_decap_8 FILLER_75_35 ();
 sg13g2_decap_8 FILLER_75_42 ();
 sg13g2_decap_8 FILLER_75_49 ();
 sg13g2_fill_2 FILLER_75_56 ();
 sg13g2_fill_1 FILLER_75_58 ();
 sg13g2_decap_8 FILLER_75_63 ();
 sg13g2_decap_8 FILLER_75_70 ();
 sg13g2_decap_8 FILLER_75_77 ();
 sg13g2_decap_8 FILLER_75_84 ();
 sg13g2_decap_8 FILLER_75_91 ();
 sg13g2_decap_8 FILLER_75_98 ();
 sg13g2_decap_8 FILLER_75_105 ();
 sg13g2_decap_8 FILLER_75_112 ();
 sg13g2_decap_8 FILLER_75_119 ();
 sg13g2_decap_8 FILLER_75_126 ();
 sg13g2_decap_8 FILLER_75_133 ();
 sg13g2_decap_8 FILLER_75_140 ();
 sg13g2_decap_8 FILLER_75_147 ();
 sg13g2_decap_8 FILLER_75_154 ();
 sg13g2_decap_8 FILLER_75_161 ();
 sg13g2_decap_8 FILLER_75_168 ();
 sg13g2_decap_8 FILLER_75_175 ();
 sg13g2_decap_8 FILLER_75_182 ();
 sg13g2_decap_8 FILLER_75_189 ();
 sg13g2_decap_8 FILLER_75_196 ();
 sg13g2_decap_8 FILLER_75_203 ();
 sg13g2_decap_8 FILLER_75_210 ();
 sg13g2_decap_8 FILLER_75_217 ();
 sg13g2_decap_8 FILLER_75_224 ();
 sg13g2_decap_8 FILLER_75_231 ();
 sg13g2_decap_8 FILLER_75_238 ();
 sg13g2_decap_8 FILLER_75_245 ();
 sg13g2_decap_8 FILLER_75_252 ();
 sg13g2_decap_8 FILLER_75_259 ();
 sg13g2_decap_8 FILLER_75_266 ();
 sg13g2_decap_8 FILLER_75_273 ();
 sg13g2_decap_8 FILLER_75_280 ();
 sg13g2_decap_8 FILLER_75_287 ();
 sg13g2_decap_8 FILLER_75_294 ();
 sg13g2_decap_8 FILLER_75_301 ();
 sg13g2_decap_8 FILLER_75_308 ();
 sg13g2_decap_8 FILLER_75_315 ();
 sg13g2_decap_8 FILLER_75_322 ();
 sg13g2_decap_8 FILLER_75_329 ();
 sg13g2_decap_8 FILLER_75_336 ();
 sg13g2_decap_8 FILLER_75_343 ();
 sg13g2_decap_8 FILLER_75_350 ();
 sg13g2_decap_8 FILLER_75_357 ();
 sg13g2_decap_8 FILLER_75_364 ();
 sg13g2_decap_8 FILLER_75_371 ();
 sg13g2_decap_8 FILLER_75_378 ();
 sg13g2_decap_8 FILLER_75_385 ();
 sg13g2_decap_8 FILLER_75_392 ();
 sg13g2_decap_8 FILLER_75_399 ();
 sg13g2_decap_8 FILLER_75_406 ();
 sg13g2_decap_8 FILLER_75_413 ();
 sg13g2_decap_8 FILLER_75_420 ();
 sg13g2_decap_8 FILLER_75_427 ();
 sg13g2_decap_8 FILLER_75_434 ();
 sg13g2_decap_8 FILLER_75_441 ();
 sg13g2_decap_8 FILLER_75_448 ();
 sg13g2_decap_8 FILLER_75_455 ();
 sg13g2_decap_8 FILLER_75_462 ();
 sg13g2_decap_8 FILLER_75_469 ();
 sg13g2_decap_8 FILLER_75_476 ();
 sg13g2_decap_8 FILLER_75_483 ();
 sg13g2_decap_8 FILLER_75_490 ();
 sg13g2_decap_8 FILLER_75_497 ();
 sg13g2_decap_8 FILLER_75_504 ();
 sg13g2_decap_8 FILLER_75_511 ();
 sg13g2_decap_8 FILLER_75_518 ();
 sg13g2_decap_8 FILLER_75_525 ();
 sg13g2_decap_8 FILLER_75_532 ();
 sg13g2_decap_8 FILLER_75_539 ();
 sg13g2_decap_8 FILLER_75_546 ();
 sg13g2_decap_8 FILLER_75_553 ();
 sg13g2_decap_8 FILLER_75_560 ();
 sg13g2_decap_8 FILLER_75_567 ();
 sg13g2_decap_8 FILLER_75_574 ();
 sg13g2_decap_8 FILLER_75_581 ();
 sg13g2_decap_8 FILLER_75_588 ();
 sg13g2_decap_8 FILLER_75_595 ();
 sg13g2_decap_8 FILLER_75_602 ();
 sg13g2_decap_8 FILLER_75_609 ();
 sg13g2_decap_8 FILLER_75_616 ();
 sg13g2_decap_8 FILLER_75_623 ();
 sg13g2_decap_8 FILLER_75_630 ();
 sg13g2_decap_8 FILLER_75_637 ();
 sg13g2_decap_8 FILLER_75_644 ();
 sg13g2_decap_8 FILLER_75_651 ();
 sg13g2_decap_8 FILLER_75_658 ();
 sg13g2_decap_8 FILLER_75_665 ();
 sg13g2_decap_8 FILLER_75_672 ();
 sg13g2_decap_8 FILLER_75_679 ();
 sg13g2_decap_8 FILLER_75_686 ();
 sg13g2_decap_8 FILLER_75_693 ();
 sg13g2_decap_8 FILLER_75_700 ();
 sg13g2_decap_8 FILLER_75_707 ();
 sg13g2_decap_8 FILLER_75_714 ();
 sg13g2_decap_8 FILLER_75_721 ();
 sg13g2_decap_8 FILLER_75_728 ();
 sg13g2_decap_8 FILLER_75_735 ();
 sg13g2_decap_8 FILLER_75_742 ();
 sg13g2_decap_8 FILLER_75_749 ();
 sg13g2_decap_8 FILLER_75_756 ();
 sg13g2_decap_8 FILLER_75_763 ();
 sg13g2_decap_8 FILLER_75_770 ();
 sg13g2_decap_8 FILLER_75_777 ();
 sg13g2_decap_8 FILLER_75_784 ();
 sg13g2_decap_8 FILLER_75_791 ();
 sg13g2_decap_8 FILLER_75_798 ();
 sg13g2_decap_8 FILLER_75_805 ();
 sg13g2_decap_8 FILLER_75_812 ();
 sg13g2_decap_8 FILLER_75_819 ();
 sg13g2_decap_8 FILLER_75_826 ();
 sg13g2_decap_8 FILLER_75_833 ();
 sg13g2_decap_8 FILLER_75_840 ();
 sg13g2_decap_8 FILLER_75_847 ();
 sg13g2_decap_8 FILLER_75_854 ();
 sg13g2_decap_8 FILLER_75_861 ();
 sg13g2_decap_8 FILLER_75_868 ();
 sg13g2_decap_8 FILLER_75_875 ();
 sg13g2_decap_8 FILLER_75_882 ();
 sg13g2_decap_8 FILLER_75_889 ();
 sg13g2_decap_8 FILLER_75_896 ();
 sg13g2_decap_8 FILLER_75_903 ();
 sg13g2_decap_8 FILLER_75_910 ();
 sg13g2_decap_8 FILLER_75_917 ();
 sg13g2_decap_8 FILLER_75_924 ();
 sg13g2_decap_8 FILLER_75_931 ();
 sg13g2_decap_8 FILLER_75_938 ();
 sg13g2_decap_8 FILLER_75_945 ();
 sg13g2_decap_8 FILLER_75_952 ();
 sg13g2_decap_8 FILLER_75_959 ();
 sg13g2_decap_8 FILLER_75_966 ();
 sg13g2_decap_8 FILLER_75_973 ();
 sg13g2_decap_8 FILLER_75_980 ();
 sg13g2_decap_8 FILLER_75_987 ();
 sg13g2_decap_8 FILLER_75_994 ();
 sg13g2_decap_8 FILLER_75_1001 ();
 sg13g2_decap_8 FILLER_75_1008 ();
 sg13g2_decap_8 FILLER_75_1015 ();
 sg13g2_decap_8 FILLER_75_1022 ();
 sg13g2_decap_8 FILLER_76_4 ();
 sg13g2_decap_8 FILLER_76_11 ();
 sg13g2_decap_8 FILLER_76_18 ();
 sg13g2_decap_8 FILLER_76_25 ();
 sg13g2_decap_8 FILLER_76_32 ();
 sg13g2_decap_8 FILLER_76_39 ();
 sg13g2_decap_8 FILLER_76_46 ();
 sg13g2_decap_8 FILLER_76_53 ();
 sg13g2_decap_8 FILLER_76_60 ();
 sg13g2_decap_8 FILLER_76_67 ();
 sg13g2_decap_8 FILLER_76_74 ();
 sg13g2_decap_8 FILLER_76_81 ();
 sg13g2_decap_8 FILLER_76_88 ();
 sg13g2_decap_8 FILLER_76_95 ();
 sg13g2_decap_8 FILLER_76_102 ();
 sg13g2_decap_8 FILLER_76_109 ();
 sg13g2_decap_8 FILLER_76_116 ();
 sg13g2_decap_8 FILLER_76_123 ();
 sg13g2_decap_8 FILLER_76_130 ();
 sg13g2_decap_8 FILLER_76_137 ();
 sg13g2_decap_8 FILLER_76_144 ();
 sg13g2_decap_8 FILLER_76_151 ();
 sg13g2_decap_8 FILLER_76_158 ();
 sg13g2_decap_8 FILLER_76_165 ();
 sg13g2_decap_8 FILLER_76_172 ();
 sg13g2_decap_8 FILLER_76_179 ();
 sg13g2_decap_8 FILLER_76_186 ();
 sg13g2_decap_8 FILLER_76_193 ();
 sg13g2_decap_8 FILLER_76_200 ();
 sg13g2_decap_8 FILLER_76_207 ();
 sg13g2_decap_8 FILLER_76_214 ();
 sg13g2_decap_8 FILLER_76_221 ();
 sg13g2_decap_8 FILLER_76_228 ();
 sg13g2_decap_8 FILLER_76_235 ();
 sg13g2_decap_8 FILLER_76_242 ();
 sg13g2_decap_8 FILLER_76_249 ();
 sg13g2_decap_8 FILLER_76_256 ();
 sg13g2_decap_8 FILLER_76_263 ();
 sg13g2_decap_8 FILLER_76_270 ();
 sg13g2_decap_8 FILLER_76_277 ();
 sg13g2_decap_8 FILLER_76_284 ();
 sg13g2_decap_8 FILLER_76_291 ();
 sg13g2_decap_8 FILLER_76_298 ();
 sg13g2_decap_8 FILLER_76_305 ();
 sg13g2_decap_8 FILLER_76_312 ();
 sg13g2_decap_8 FILLER_76_319 ();
 sg13g2_decap_8 FILLER_76_326 ();
 sg13g2_decap_8 FILLER_76_333 ();
 sg13g2_decap_8 FILLER_76_340 ();
 sg13g2_decap_8 FILLER_76_347 ();
 sg13g2_decap_8 FILLER_76_354 ();
 sg13g2_decap_8 FILLER_76_361 ();
 sg13g2_decap_8 FILLER_76_368 ();
 sg13g2_decap_8 FILLER_76_375 ();
 sg13g2_decap_8 FILLER_76_382 ();
 sg13g2_decap_8 FILLER_76_389 ();
 sg13g2_decap_8 FILLER_76_396 ();
 sg13g2_decap_8 FILLER_76_403 ();
 sg13g2_decap_8 FILLER_76_410 ();
 sg13g2_decap_8 FILLER_76_417 ();
 sg13g2_decap_8 FILLER_76_424 ();
 sg13g2_decap_8 FILLER_76_431 ();
 sg13g2_decap_8 FILLER_76_438 ();
 sg13g2_decap_8 FILLER_76_445 ();
 sg13g2_decap_8 FILLER_76_452 ();
 sg13g2_decap_8 FILLER_76_459 ();
 sg13g2_decap_8 FILLER_76_466 ();
 sg13g2_decap_8 FILLER_76_473 ();
 sg13g2_decap_8 FILLER_76_480 ();
 sg13g2_decap_8 FILLER_76_487 ();
 sg13g2_decap_8 FILLER_76_494 ();
 sg13g2_decap_8 FILLER_76_501 ();
 sg13g2_decap_8 FILLER_76_508 ();
 sg13g2_decap_8 FILLER_76_515 ();
 sg13g2_decap_8 FILLER_76_522 ();
 sg13g2_decap_8 FILLER_76_529 ();
 sg13g2_decap_8 FILLER_76_536 ();
 sg13g2_decap_8 FILLER_76_543 ();
 sg13g2_decap_8 FILLER_76_550 ();
 sg13g2_decap_8 FILLER_76_557 ();
 sg13g2_decap_8 FILLER_76_564 ();
 sg13g2_decap_8 FILLER_76_571 ();
 sg13g2_decap_8 FILLER_76_578 ();
 sg13g2_decap_8 FILLER_76_585 ();
 sg13g2_decap_8 FILLER_76_592 ();
 sg13g2_decap_8 FILLER_76_599 ();
 sg13g2_decap_8 FILLER_76_606 ();
 sg13g2_decap_8 FILLER_76_613 ();
 sg13g2_decap_8 FILLER_76_620 ();
 sg13g2_decap_8 FILLER_76_627 ();
 sg13g2_decap_8 FILLER_76_634 ();
 sg13g2_decap_8 FILLER_76_641 ();
 sg13g2_decap_8 FILLER_76_648 ();
 sg13g2_decap_8 FILLER_76_655 ();
 sg13g2_decap_8 FILLER_76_662 ();
 sg13g2_decap_8 FILLER_76_669 ();
 sg13g2_decap_8 FILLER_76_676 ();
 sg13g2_decap_8 FILLER_76_683 ();
 sg13g2_decap_8 FILLER_76_690 ();
 sg13g2_decap_8 FILLER_76_697 ();
 sg13g2_decap_8 FILLER_76_704 ();
 sg13g2_decap_8 FILLER_76_711 ();
 sg13g2_decap_8 FILLER_76_718 ();
 sg13g2_decap_8 FILLER_76_725 ();
 sg13g2_decap_8 FILLER_76_732 ();
 sg13g2_decap_8 FILLER_76_739 ();
 sg13g2_decap_8 FILLER_76_746 ();
 sg13g2_decap_8 FILLER_76_753 ();
 sg13g2_decap_8 FILLER_76_760 ();
 sg13g2_decap_8 FILLER_76_767 ();
 sg13g2_decap_8 FILLER_76_774 ();
 sg13g2_decap_8 FILLER_76_781 ();
 sg13g2_decap_8 FILLER_76_788 ();
 sg13g2_decap_8 FILLER_76_795 ();
 sg13g2_decap_8 FILLER_76_802 ();
 sg13g2_decap_8 FILLER_76_809 ();
 sg13g2_decap_8 FILLER_76_816 ();
 sg13g2_decap_8 FILLER_76_823 ();
 sg13g2_decap_8 FILLER_76_830 ();
 sg13g2_decap_8 FILLER_76_837 ();
 sg13g2_decap_8 FILLER_76_844 ();
 sg13g2_decap_8 FILLER_76_851 ();
 sg13g2_decap_8 FILLER_76_858 ();
 sg13g2_decap_8 FILLER_76_865 ();
 sg13g2_decap_8 FILLER_76_872 ();
 sg13g2_decap_8 FILLER_76_879 ();
 sg13g2_decap_8 FILLER_76_886 ();
 sg13g2_decap_8 FILLER_76_893 ();
 sg13g2_decap_8 FILLER_76_900 ();
 sg13g2_decap_8 FILLER_76_907 ();
 sg13g2_decap_8 FILLER_76_914 ();
 sg13g2_decap_8 FILLER_76_921 ();
 sg13g2_decap_8 FILLER_76_928 ();
 sg13g2_decap_8 FILLER_76_935 ();
 sg13g2_decap_8 FILLER_76_942 ();
 sg13g2_decap_8 FILLER_76_949 ();
 sg13g2_decap_8 FILLER_76_956 ();
 sg13g2_decap_8 FILLER_76_963 ();
 sg13g2_decap_8 FILLER_76_970 ();
 sg13g2_decap_8 FILLER_76_977 ();
 sg13g2_decap_8 FILLER_76_984 ();
 sg13g2_decap_8 FILLER_76_991 ();
 sg13g2_decap_8 FILLER_76_998 ();
 sg13g2_decap_8 FILLER_76_1005 ();
 sg13g2_decap_8 FILLER_76_1012 ();
 sg13g2_decap_8 FILLER_76_1019 ();
 sg13g2_fill_2 FILLER_76_1026 ();
 sg13g2_fill_1 FILLER_76_1028 ();
 sg13g2_decap_8 FILLER_77_0 ();
 sg13g2_decap_8 FILLER_77_7 ();
 sg13g2_decap_8 FILLER_77_14 ();
 sg13g2_decap_8 FILLER_77_21 ();
 sg13g2_decap_8 FILLER_77_28 ();
 sg13g2_decap_8 FILLER_77_35 ();
 sg13g2_decap_8 FILLER_77_42 ();
 sg13g2_decap_8 FILLER_77_49 ();
 sg13g2_decap_8 FILLER_77_56 ();
 sg13g2_decap_8 FILLER_77_63 ();
 sg13g2_decap_8 FILLER_77_70 ();
 sg13g2_decap_8 FILLER_77_77 ();
 sg13g2_decap_8 FILLER_77_84 ();
 sg13g2_decap_8 FILLER_77_91 ();
 sg13g2_decap_8 FILLER_77_98 ();
 sg13g2_decap_8 FILLER_77_105 ();
 sg13g2_decap_8 FILLER_77_112 ();
 sg13g2_decap_8 FILLER_77_119 ();
 sg13g2_decap_8 FILLER_77_126 ();
 sg13g2_decap_8 FILLER_77_133 ();
 sg13g2_decap_8 FILLER_77_140 ();
 sg13g2_decap_8 FILLER_77_147 ();
 sg13g2_decap_8 FILLER_77_154 ();
 sg13g2_decap_8 FILLER_77_161 ();
 sg13g2_decap_8 FILLER_77_168 ();
 sg13g2_decap_8 FILLER_77_175 ();
 sg13g2_decap_8 FILLER_77_182 ();
 sg13g2_decap_8 FILLER_77_189 ();
 sg13g2_decap_8 FILLER_77_196 ();
 sg13g2_decap_8 FILLER_77_203 ();
 sg13g2_decap_8 FILLER_77_210 ();
 sg13g2_decap_8 FILLER_77_217 ();
 sg13g2_decap_8 FILLER_77_224 ();
 sg13g2_decap_8 FILLER_77_231 ();
 sg13g2_decap_8 FILLER_77_238 ();
 sg13g2_decap_8 FILLER_77_245 ();
 sg13g2_decap_8 FILLER_77_252 ();
 sg13g2_decap_8 FILLER_77_259 ();
 sg13g2_decap_8 FILLER_77_266 ();
 sg13g2_decap_8 FILLER_77_273 ();
 sg13g2_decap_8 FILLER_77_280 ();
 sg13g2_decap_8 FILLER_77_287 ();
 sg13g2_decap_8 FILLER_77_294 ();
 sg13g2_decap_8 FILLER_77_301 ();
 sg13g2_decap_8 FILLER_77_308 ();
 sg13g2_decap_8 FILLER_77_315 ();
 sg13g2_decap_8 FILLER_77_322 ();
 sg13g2_decap_8 FILLER_77_329 ();
 sg13g2_decap_8 FILLER_77_336 ();
 sg13g2_decap_8 FILLER_77_343 ();
 sg13g2_decap_8 FILLER_77_350 ();
 sg13g2_decap_8 FILLER_77_357 ();
 sg13g2_decap_8 FILLER_77_364 ();
 sg13g2_decap_8 FILLER_77_371 ();
 sg13g2_decap_8 FILLER_77_378 ();
 sg13g2_decap_8 FILLER_77_385 ();
 sg13g2_decap_8 FILLER_77_392 ();
 sg13g2_decap_8 FILLER_77_399 ();
 sg13g2_decap_8 FILLER_77_406 ();
 sg13g2_decap_8 FILLER_77_413 ();
 sg13g2_decap_8 FILLER_77_420 ();
 sg13g2_decap_8 FILLER_77_427 ();
 sg13g2_decap_8 FILLER_77_434 ();
 sg13g2_decap_8 FILLER_77_441 ();
 sg13g2_decap_8 FILLER_77_448 ();
 sg13g2_decap_8 FILLER_77_455 ();
 sg13g2_decap_8 FILLER_77_462 ();
 sg13g2_decap_8 FILLER_77_469 ();
 sg13g2_decap_8 FILLER_77_476 ();
 sg13g2_decap_8 FILLER_77_483 ();
 sg13g2_decap_8 FILLER_77_490 ();
 sg13g2_decap_8 FILLER_77_497 ();
 sg13g2_decap_8 FILLER_77_504 ();
 sg13g2_decap_8 FILLER_77_511 ();
 sg13g2_decap_8 FILLER_77_518 ();
 sg13g2_decap_8 FILLER_77_525 ();
 sg13g2_decap_8 FILLER_77_532 ();
 sg13g2_decap_8 FILLER_77_539 ();
 sg13g2_decap_8 FILLER_77_546 ();
 sg13g2_decap_8 FILLER_77_553 ();
 sg13g2_decap_8 FILLER_77_560 ();
 sg13g2_decap_8 FILLER_77_567 ();
 sg13g2_decap_8 FILLER_77_574 ();
 sg13g2_decap_8 FILLER_77_581 ();
 sg13g2_decap_8 FILLER_77_588 ();
 sg13g2_decap_8 FILLER_77_595 ();
 sg13g2_decap_8 FILLER_77_602 ();
 sg13g2_decap_8 FILLER_77_609 ();
 sg13g2_decap_8 FILLER_77_616 ();
 sg13g2_decap_8 FILLER_77_623 ();
 sg13g2_decap_8 FILLER_77_630 ();
 sg13g2_decap_8 FILLER_77_637 ();
 sg13g2_decap_8 FILLER_77_644 ();
 sg13g2_decap_8 FILLER_77_651 ();
 sg13g2_decap_8 FILLER_77_658 ();
 sg13g2_decap_8 FILLER_77_665 ();
 sg13g2_decap_8 FILLER_77_672 ();
 sg13g2_decap_8 FILLER_77_679 ();
 sg13g2_decap_8 FILLER_77_686 ();
 sg13g2_decap_8 FILLER_77_693 ();
 sg13g2_decap_8 FILLER_77_700 ();
 sg13g2_decap_8 FILLER_77_707 ();
 sg13g2_decap_8 FILLER_77_714 ();
 sg13g2_decap_8 FILLER_77_721 ();
 sg13g2_decap_8 FILLER_77_728 ();
 sg13g2_decap_8 FILLER_77_735 ();
 sg13g2_decap_8 FILLER_77_742 ();
 sg13g2_decap_8 FILLER_77_749 ();
 sg13g2_decap_8 FILLER_77_756 ();
 sg13g2_decap_8 FILLER_77_763 ();
 sg13g2_decap_8 FILLER_77_770 ();
 sg13g2_decap_8 FILLER_77_777 ();
 sg13g2_decap_8 FILLER_77_784 ();
 sg13g2_decap_8 FILLER_77_791 ();
 sg13g2_decap_8 FILLER_77_798 ();
 sg13g2_decap_8 FILLER_77_805 ();
 sg13g2_decap_8 FILLER_77_812 ();
 sg13g2_decap_8 FILLER_77_819 ();
 sg13g2_decap_8 FILLER_77_826 ();
 sg13g2_decap_8 FILLER_77_833 ();
 sg13g2_decap_8 FILLER_77_840 ();
 sg13g2_decap_8 FILLER_77_847 ();
 sg13g2_decap_8 FILLER_77_854 ();
 sg13g2_decap_8 FILLER_77_861 ();
 sg13g2_decap_8 FILLER_77_868 ();
 sg13g2_decap_8 FILLER_77_875 ();
 sg13g2_decap_8 FILLER_77_882 ();
 sg13g2_decap_8 FILLER_77_889 ();
 sg13g2_decap_8 FILLER_77_896 ();
 sg13g2_decap_8 FILLER_77_903 ();
 sg13g2_decap_8 FILLER_77_910 ();
 sg13g2_decap_8 FILLER_77_917 ();
 sg13g2_decap_8 FILLER_77_924 ();
 sg13g2_decap_8 FILLER_77_931 ();
 sg13g2_decap_8 FILLER_77_938 ();
 sg13g2_decap_8 FILLER_77_945 ();
 sg13g2_decap_8 FILLER_77_952 ();
 sg13g2_decap_8 FILLER_77_959 ();
 sg13g2_decap_8 FILLER_77_966 ();
 sg13g2_decap_8 FILLER_77_973 ();
 sg13g2_decap_8 FILLER_77_980 ();
 sg13g2_decap_8 FILLER_77_987 ();
 sg13g2_decap_8 FILLER_77_994 ();
 sg13g2_decap_8 FILLER_77_1001 ();
 sg13g2_decap_8 FILLER_77_1008 ();
 sg13g2_decap_8 FILLER_77_1015 ();
 sg13g2_decap_8 FILLER_77_1022 ();
 sg13g2_decap_8 FILLER_78_4 ();
 sg13g2_decap_8 FILLER_78_11 ();
 sg13g2_decap_8 FILLER_78_18 ();
 sg13g2_decap_8 FILLER_78_25 ();
 sg13g2_decap_8 FILLER_78_32 ();
 sg13g2_decap_8 FILLER_78_39 ();
 sg13g2_decap_8 FILLER_78_46 ();
 sg13g2_decap_8 FILLER_78_53 ();
 sg13g2_fill_1 FILLER_78_60 ();
 sg13g2_decap_8 FILLER_78_69 ();
 sg13g2_decap_8 FILLER_78_76 ();
 sg13g2_decap_8 FILLER_78_83 ();
 sg13g2_decap_8 FILLER_78_90 ();
 sg13g2_decap_8 FILLER_78_97 ();
 sg13g2_decap_8 FILLER_78_104 ();
 sg13g2_decap_8 FILLER_78_111 ();
 sg13g2_decap_8 FILLER_78_118 ();
 sg13g2_decap_8 FILLER_78_125 ();
 sg13g2_decap_8 FILLER_78_132 ();
 sg13g2_decap_8 FILLER_78_139 ();
 sg13g2_decap_8 FILLER_78_146 ();
 sg13g2_decap_8 FILLER_78_153 ();
 sg13g2_decap_8 FILLER_78_160 ();
 sg13g2_decap_8 FILLER_78_167 ();
 sg13g2_decap_8 FILLER_78_174 ();
 sg13g2_decap_8 FILLER_78_181 ();
 sg13g2_decap_8 FILLER_78_188 ();
 sg13g2_decap_8 FILLER_78_195 ();
 sg13g2_decap_8 FILLER_78_202 ();
 sg13g2_decap_8 FILLER_78_209 ();
 sg13g2_decap_8 FILLER_78_216 ();
 sg13g2_decap_8 FILLER_78_223 ();
 sg13g2_decap_8 FILLER_78_230 ();
 sg13g2_decap_8 FILLER_78_237 ();
 sg13g2_decap_8 FILLER_78_244 ();
 sg13g2_decap_8 FILLER_78_251 ();
 sg13g2_decap_8 FILLER_78_258 ();
 sg13g2_decap_8 FILLER_78_265 ();
 sg13g2_decap_8 FILLER_78_272 ();
 sg13g2_decap_8 FILLER_78_279 ();
 sg13g2_decap_8 FILLER_78_286 ();
 sg13g2_decap_8 FILLER_78_293 ();
 sg13g2_decap_8 FILLER_78_300 ();
 sg13g2_decap_8 FILLER_78_307 ();
 sg13g2_decap_8 FILLER_78_314 ();
 sg13g2_decap_8 FILLER_78_321 ();
 sg13g2_decap_8 FILLER_78_328 ();
 sg13g2_decap_8 FILLER_78_335 ();
 sg13g2_decap_8 FILLER_78_342 ();
 sg13g2_decap_8 FILLER_78_349 ();
 sg13g2_decap_8 FILLER_78_356 ();
 sg13g2_decap_8 FILLER_78_363 ();
 sg13g2_decap_8 FILLER_78_370 ();
 sg13g2_decap_8 FILLER_78_377 ();
 sg13g2_decap_8 FILLER_78_384 ();
 sg13g2_decap_8 FILLER_78_391 ();
 sg13g2_decap_8 FILLER_78_398 ();
 sg13g2_decap_8 FILLER_78_405 ();
 sg13g2_decap_8 FILLER_78_412 ();
 sg13g2_decap_8 FILLER_78_419 ();
 sg13g2_decap_8 FILLER_78_426 ();
 sg13g2_decap_8 FILLER_78_433 ();
 sg13g2_decap_8 FILLER_78_440 ();
 sg13g2_decap_8 FILLER_78_447 ();
 sg13g2_decap_8 FILLER_78_454 ();
 sg13g2_decap_8 FILLER_78_461 ();
 sg13g2_decap_8 FILLER_78_468 ();
 sg13g2_decap_8 FILLER_78_475 ();
 sg13g2_decap_8 FILLER_78_482 ();
 sg13g2_decap_8 FILLER_78_489 ();
 sg13g2_decap_8 FILLER_78_496 ();
 sg13g2_decap_8 FILLER_78_503 ();
 sg13g2_decap_8 FILLER_78_510 ();
 sg13g2_decap_8 FILLER_78_517 ();
 sg13g2_decap_8 FILLER_78_524 ();
 sg13g2_decap_8 FILLER_78_531 ();
 sg13g2_decap_8 FILLER_78_538 ();
 sg13g2_decap_8 FILLER_78_545 ();
 sg13g2_decap_8 FILLER_78_552 ();
 sg13g2_decap_8 FILLER_78_559 ();
 sg13g2_decap_8 FILLER_78_566 ();
 sg13g2_decap_8 FILLER_78_573 ();
 sg13g2_decap_8 FILLER_78_580 ();
 sg13g2_decap_8 FILLER_78_587 ();
 sg13g2_decap_8 FILLER_78_594 ();
 sg13g2_decap_8 FILLER_78_601 ();
 sg13g2_decap_8 FILLER_78_608 ();
 sg13g2_decap_8 FILLER_78_615 ();
 sg13g2_decap_8 FILLER_78_622 ();
 sg13g2_decap_8 FILLER_78_629 ();
 sg13g2_decap_8 FILLER_78_636 ();
 sg13g2_decap_8 FILLER_78_643 ();
 sg13g2_decap_8 FILLER_78_650 ();
 sg13g2_decap_8 FILLER_78_657 ();
 sg13g2_decap_8 FILLER_78_664 ();
 sg13g2_decap_8 FILLER_78_671 ();
 sg13g2_decap_8 FILLER_78_678 ();
 sg13g2_decap_8 FILLER_78_685 ();
 sg13g2_decap_8 FILLER_78_692 ();
 sg13g2_decap_8 FILLER_78_699 ();
 sg13g2_decap_8 FILLER_78_706 ();
 sg13g2_decap_8 FILLER_78_713 ();
 sg13g2_decap_8 FILLER_78_720 ();
 sg13g2_decap_8 FILLER_78_727 ();
 sg13g2_decap_8 FILLER_78_734 ();
 sg13g2_decap_8 FILLER_78_741 ();
 sg13g2_decap_8 FILLER_78_748 ();
 sg13g2_decap_8 FILLER_78_755 ();
 sg13g2_decap_8 FILLER_78_762 ();
 sg13g2_decap_8 FILLER_78_769 ();
 sg13g2_decap_8 FILLER_78_776 ();
 sg13g2_decap_8 FILLER_78_783 ();
 sg13g2_decap_8 FILLER_78_790 ();
 sg13g2_decap_8 FILLER_78_797 ();
 sg13g2_decap_8 FILLER_78_804 ();
 sg13g2_decap_8 FILLER_78_811 ();
 sg13g2_decap_8 FILLER_78_818 ();
 sg13g2_decap_8 FILLER_78_825 ();
 sg13g2_decap_8 FILLER_78_832 ();
 sg13g2_decap_8 FILLER_78_839 ();
 sg13g2_decap_8 FILLER_78_846 ();
 sg13g2_decap_8 FILLER_78_853 ();
 sg13g2_decap_8 FILLER_78_860 ();
 sg13g2_decap_8 FILLER_78_867 ();
 sg13g2_decap_8 FILLER_78_874 ();
 sg13g2_decap_8 FILLER_78_881 ();
 sg13g2_decap_8 FILLER_78_888 ();
 sg13g2_decap_8 FILLER_78_895 ();
 sg13g2_decap_8 FILLER_78_902 ();
 sg13g2_decap_8 FILLER_78_909 ();
 sg13g2_decap_8 FILLER_78_916 ();
 sg13g2_decap_8 FILLER_78_923 ();
 sg13g2_decap_8 FILLER_78_930 ();
 sg13g2_decap_8 FILLER_78_937 ();
 sg13g2_decap_8 FILLER_78_944 ();
 sg13g2_decap_8 FILLER_78_951 ();
 sg13g2_decap_8 FILLER_78_958 ();
 sg13g2_decap_8 FILLER_78_965 ();
 sg13g2_decap_8 FILLER_78_972 ();
 sg13g2_decap_8 FILLER_78_979 ();
 sg13g2_decap_8 FILLER_78_986 ();
 sg13g2_decap_8 FILLER_78_993 ();
 sg13g2_decap_8 FILLER_78_1000 ();
 sg13g2_decap_8 FILLER_78_1007 ();
 sg13g2_decap_8 FILLER_78_1014 ();
 sg13g2_decap_8 FILLER_78_1021 ();
 sg13g2_fill_1 FILLER_78_1028 ();
 sg13g2_decap_8 FILLER_79_0 ();
 sg13g2_decap_8 FILLER_79_7 ();
 sg13g2_decap_8 FILLER_79_14 ();
 sg13g2_decap_8 FILLER_79_21 ();
 sg13g2_decap_8 FILLER_79_28 ();
 sg13g2_decap_8 FILLER_79_35 ();
 sg13g2_decap_8 FILLER_79_42 ();
 sg13g2_decap_8 FILLER_79_49 ();
 sg13g2_fill_2 FILLER_79_56 ();
 sg13g2_fill_1 FILLER_79_58 ();
 sg13g2_decap_8 FILLER_79_67 ();
 sg13g2_decap_8 FILLER_79_74 ();
 sg13g2_decap_8 FILLER_79_81 ();
 sg13g2_decap_8 FILLER_79_88 ();
 sg13g2_decap_8 FILLER_79_95 ();
 sg13g2_decap_8 FILLER_79_102 ();
 sg13g2_decap_8 FILLER_79_109 ();
 sg13g2_decap_8 FILLER_79_116 ();
 sg13g2_decap_8 FILLER_79_123 ();
 sg13g2_decap_8 FILLER_79_130 ();
 sg13g2_decap_8 FILLER_79_137 ();
 sg13g2_decap_8 FILLER_79_144 ();
 sg13g2_decap_8 FILLER_79_151 ();
 sg13g2_decap_8 FILLER_79_158 ();
 sg13g2_decap_8 FILLER_79_165 ();
 sg13g2_decap_8 FILLER_79_172 ();
 sg13g2_decap_8 FILLER_79_179 ();
 sg13g2_decap_8 FILLER_79_186 ();
 sg13g2_decap_8 FILLER_79_193 ();
 sg13g2_decap_8 FILLER_79_200 ();
 sg13g2_decap_8 FILLER_79_207 ();
 sg13g2_decap_8 FILLER_79_214 ();
 sg13g2_decap_8 FILLER_79_221 ();
 sg13g2_decap_8 FILLER_79_228 ();
 sg13g2_decap_8 FILLER_79_235 ();
 sg13g2_decap_8 FILLER_79_242 ();
 sg13g2_decap_8 FILLER_79_249 ();
 sg13g2_decap_8 FILLER_79_256 ();
 sg13g2_decap_8 FILLER_79_263 ();
 sg13g2_decap_8 FILLER_79_270 ();
 sg13g2_decap_8 FILLER_79_277 ();
 sg13g2_decap_8 FILLER_79_284 ();
 sg13g2_decap_8 FILLER_79_291 ();
 sg13g2_decap_8 FILLER_79_298 ();
 sg13g2_decap_8 FILLER_79_305 ();
 sg13g2_decap_8 FILLER_79_312 ();
 sg13g2_decap_8 FILLER_79_319 ();
 sg13g2_decap_8 FILLER_79_326 ();
 sg13g2_decap_8 FILLER_79_333 ();
 sg13g2_decap_8 FILLER_79_340 ();
 sg13g2_decap_8 FILLER_79_347 ();
 sg13g2_decap_8 FILLER_79_354 ();
 sg13g2_decap_8 FILLER_79_361 ();
 sg13g2_decap_8 FILLER_79_368 ();
 sg13g2_decap_8 FILLER_79_375 ();
 sg13g2_decap_8 FILLER_79_382 ();
 sg13g2_decap_8 FILLER_79_389 ();
 sg13g2_decap_8 FILLER_79_396 ();
 sg13g2_decap_8 FILLER_79_403 ();
 sg13g2_decap_8 FILLER_79_410 ();
 sg13g2_decap_8 FILLER_79_417 ();
 sg13g2_decap_8 FILLER_79_424 ();
 sg13g2_decap_8 FILLER_79_431 ();
 sg13g2_decap_8 FILLER_79_438 ();
 sg13g2_decap_8 FILLER_79_445 ();
 sg13g2_decap_8 FILLER_79_452 ();
 sg13g2_decap_8 FILLER_79_459 ();
 sg13g2_decap_8 FILLER_79_466 ();
 sg13g2_decap_8 FILLER_79_473 ();
 sg13g2_decap_8 FILLER_79_480 ();
 sg13g2_decap_8 FILLER_79_487 ();
 sg13g2_decap_8 FILLER_79_494 ();
 sg13g2_decap_8 FILLER_79_501 ();
 sg13g2_decap_8 FILLER_79_508 ();
 sg13g2_decap_8 FILLER_79_515 ();
 sg13g2_decap_8 FILLER_79_522 ();
 sg13g2_decap_8 FILLER_79_529 ();
 sg13g2_decap_8 FILLER_79_536 ();
 sg13g2_decap_8 FILLER_79_543 ();
 sg13g2_decap_8 FILLER_79_550 ();
 sg13g2_decap_8 FILLER_79_557 ();
 sg13g2_decap_8 FILLER_79_564 ();
 sg13g2_decap_8 FILLER_79_571 ();
 sg13g2_decap_8 FILLER_79_578 ();
 sg13g2_decap_8 FILLER_79_585 ();
 sg13g2_decap_8 FILLER_79_592 ();
 sg13g2_decap_8 FILLER_79_599 ();
 sg13g2_decap_8 FILLER_79_606 ();
 sg13g2_decap_8 FILLER_79_613 ();
 sg13g2_decap_8 FILLER_79_620 ();
 sg13g2_decap_8 FILLER_79_627 ();
 sg13g2_decap_8 FILLER_79_634 ();
 sg13g2_decap_8 FILLER_79_641 ();
 sg13g2_decap_8 FILLER_79_648 ();
 sg13g2_decap_8 FILLER_79_655 ();
 sg13g2_decap_8 FILLER_79_662 ();
 sg13g2_decap_8 FILLER_79_669 ();
 sg13g2_decap_8 FILLER_79_676 ();
 sg13g2_decap_8 FILLER_79_683 ();
 sg13g2_decap_8 FILLER_79_690 ();
 sg13g2_decap_8 FILLER_79_697 ();
 sg13g2_decap_8 FILLER_79_704 ();
 sg13g2_decap_8 FILLER_79_711 ();
 sg13g2_decap_8 FILLER_79_718 ();
 sg13g2_decap_8 FILLER_79_725 ();
 sg13g2_decap_8 FILLER_79_732 ();
 sg13g2_decap_8 FILLER_79_739 ();
 sg13g2_decap_8 FILLER_79_746 ();
 sg13g2_decap_8 FILLER_79_753 ();
 sg13g2_decap_8 FILLER_79_760 ();
 sg13g2_decap_8 FILLER_79_767 ();
 sg13g2_decap_8 FILLER_79_774 ();
 sg13g2_decap_8 FILLER_79_781 ();
 sg13g2_decap_8 FILLER_79_788 ();
 sg13g2_decap_8 FILLER_79_795 ();
 sg13g2_decap_8 FILLER_79_802 ();
 sg13g2_decap_8 FILLER_79_809 ();
 sg13g2_decap_8 FILLER_79_816 ();
 sg13g2_decap_8 FILLER_79_823 ();
 sg13g2_decap_8 FILLER_79_830 ();
 sg13g2_decap_8 FILLER_79_837 ();
 sg13g2_decap_8 FILLER_79_844 ();
 sg13g2_decap_8 FILLER_79_851 ();
 sg13g2_decap_8 FILLER_79_858 ();
 sg13g2_decap_8 FILLER_79_865 ();
 sg13g2_decap_8 FILLER_79_872 ();
 sg13g2_decap_8 FILLER_79_879 ();
 sg13g2_decap_8 FILLER_79_886 ();
 sg13g2_decap_8 FILLER_79_893 ();
 sg13g2_decap_8 FILLER_79_900 ();
 sg13g2_decap_8 FILLER_79_907 ();
 sg13g2_decap_8 FILLER_79_914 ();
 sg13g2_decap_8 FILLER_79_921 ();
 sg13g2_decap_8 FILLER_79_928 ();
 sg13g2_decap_8 FILLER_79_935 ();
 sg13g2_decap_8 FILLER_79_942 ();
 sg13g2_decap_8 FILLER_79_949 ();
 sg13g2_decap_8 FILLER_79_956 ();
 sg13g2_decap_8 FILLER_79_963 ();
 sg13g2_decap_8 FILLER_79_970 ();
 sg13g2_decap_8 FILLER_79_977 ();
 sg13g2_decap_8 FILLER_79_984 ();
 sg13g2_decap_8 FILLER_79_991 ();
 sg13g2_decap_8 FILLER_79_998 ();
 sg13g2_decap_8 FILLER_79_1005 ();
 sg13g2_decap_8 FILLER_79_1012 ();
 sg13g2_decap_8 FILLER_79_1019 ();
 sg13g2_fill_2 FILLER_79_1026 ();
 sg13g2_fill_1 FILLER_79_1028 ();
 sg13g2_decap_8 FILLER_80_0 ();
 sg13g2_decap_8 FILLER_80_7 ();
 sg13g2_decap_8 FILLER_80_14 ();
 sg13g2_decap_8 FILLER_80_21 ();
 sg13g2_decap_8 FILLER_80_28 ();
 sg13g2_decap_8 FILLER_80_35 ();
 sg13g2_decap_8 FILLER_80_42 ();
 sg13g2_decap_8 FILLER_80_49 ();
 sg13g2_decap_8 FILLER_80_56 ();
 sg13g2_decap_8 FILLER_80_63 ();
 sg13g2_decap_8 FILLER_80_70 ();
 sg13g2_decap_8 FILLER_80_77 ();
 sg13g2_decap_8 FILLER_80_84 ();
 sg13g2_decap_8 FILLER_80_91 ();
 sg13g2_decap_8 FILLER_80_98 ();
 sg13g2_decap_8 FILLER_80_105 ();
 sg13g2_decap_8 FILLER_80_112 ();
 sg13g2_decap_8 FILLER_80_119 ();
 sg13g2_decap_8 FILLER_80_126 ();
 sg13g2_decap_8 FILLER_80_133 ();
 sg13g2_decap_8 FILLER_80_140 ();
 sg13g2_decap_8 FILLER_80_147 ();
 sg13g2_decap_8 FILLER_80_154 ();
 sg13g2_decap_8 FILLER_80_161 ();
 sg13g2_decap_8 FILLER_80_168 ();
 sg13g2_decap_8 FILLER_80_175 ();
 sg13g2_decap_8 FILLER_80_182 ();
 sg13g2_decap_8 FILLER_80_189 ();
 sg13g2_decap_8 FILLER_80_196 ();
 sg13g2_decap_8 FILLER_80_203 ();
 sg13g2_decap_8 FILLER_80_210 ();
 sg13g2_decap_8 FILLER_80_217 ();
 sg13g2_decap_8 FILLER_80_224 ();
 sg13g2_decap_8 FILLER_80_231 ();
 sg13g2_decap_8 FILLER_80_238 ();
 sg13g2_decap_8 FILLER_80_245 ();
 sg13g2_decap_8 FILLER_80_252 ();
 sg13g2_decap_8 FILLER_80_259 ();
 sg13g2_decap_8 FILLER_80_266 ();
 sg13g2_decap_8 FILLER_80_273 ();
 sg13g2_decap_8 FILLER_80_280 ();
 sg13g2_decap_8 FILLER_80_287 ();
 sg13g2_decap_8 FILLER_80_294 ();
 sg13g2_decap_8 FILLER_80_301 ();
 sg13g2_decap_8 FILLER_80_308 ();
 sg13g2_decap_8 FILLER_80_315 ();
 sg13g2_decap_8 FILLER_80_322 ();
 sg13g2_decap_8 FILLER_80_329 ();
 sg13g2_decap_8 FILLER_80_336 ();
 sg13g2_decap_8 FILLER_80_343 ();
 sg13g2_decap_8 FILLER_80_350 ();
 sg13g2_decap_8 FILLER_80_357 ();
 sg13g2_decap_8 FILLER_80_364 ();
 sg13g2_decap_8 FILLER_80_371 ();
 sg13g2_decap_8 FILLER_80_378 ();
 sg13g2_decap_8 FILLER_80_385 ();
 sg13g2_decap_8 FILLER_80_392 ();
 sg13g2_decap_8 FILLER_80_399 ();
 sg13g2_decap_8 FILLER_80_406 ();
 sg13g2_decap_8 FILLER_80_413 ();
 sg13g2_decap_8 FILLER_80_420 ();
 sg13g2_decap_8 FILLER_80_427 ();
 sg13g2_decap_8 FILLER_80_434 ();
 sg13g2_decap_8 FILLER_80_441 ();
 sg13g2_decap_8 FILLER_80_448 ();
 sg13g2_decap_8 FILLER_80_455 ();
 sg13g2_decap_8 FILLER_80_462 ();
 sg13g2_decap_8 FILLER_80_469 ();
 sg13g2_decap_8 FILLER_80_476 ();
 sg13g2_decap_8 FILLER_80_483 ();
 sg13g2_decap_8 FILLER_80_490 ();
 sg13g2_decap_8 FILLER_80_497 ();
 sg13g2_decap_8 FILLER_80_504 ();
 sg13g2_decap_8 FILLER_80_511 ();
 sg13g2_decap_8 FILLER_80_518 ();
 sg13g2_decap_8 FILLER_80_525 ();
 sg13g2_decap_8 FILLER_80_532 ();
 sg13g2_decap_8 FILLER_80_539 ();
 sg13g2_decap_8 FILLER_80_546 ();
 sg13g2_decap_8 FILLER_80_553 ();
 sg13g2_decap_8 FILLER_80_560 ();
 sg13g2_decap_8 FILLER_80_567 ();
 sg13g2_decap_8 FILLER_80_574 ();
 sg13g2_decap_8 FILLER_80_581 ();
 sg13g2_decap_8 FILLER_80_588 ();
 sg13g2_decap_8 FILLER_80_595 ();
 sg13g2_decap_8 FILLER_80_602 ();
 sg13g2_decap_8 FILLER_80_609 ();
 sg13g2_decap_8 FILLER_80_616 ();
 sg13g2_decap_8 FILLER_80_623 ();
 sg13g2_decap_8 FILLER_80_630 ();
 sg13g2_decap_8 FILLER_80_637 ();
 sg13g2_decap_8 FILLER_80_644 ();
 sg13g2_decap_8 FILLER_80_651 ();
 sg13g2_decap_8 FILLER_80_658 ();
 sg13g2_decap_8 FILLER_80_665 ();
 sg13g2_decap_8 FILLER_80_672 ();
 sg13g2_decap_8 FILLER_80_679 ();
 sg13g2_decap_8 FILLER_80_686 ();
 sg13g2_decap_8 FILLER_80_693 ();
 sg13g2_decap_8 FILLER_80_700 ();
 sg13g2_decap_8 FILLER_80_707 ();
 sg13g2_decap_8 FILLER_80_714 ();
 sg13g2_decap_8 FILLER_80_721 ();
 sg13g2_decap_8 FILLER_80_728 ();
 sg13g2_decap_8 FILLER_80_735 ();
 sg13g2_decap_8 FILLER_80_742 ();
 sg13g2_decap_8 FILLER_80_749 ();
 sg13g2_decap_8 FILLER_80_756 ();
 sg13g2_decap_8 FILLER_80_763 ();
 sg13g2_decap_8 FILLER_80_770 ();
 sg13g2_decap_8 FILLER_80_777 ();
 sg13g2_decap_8 FILLER_80_784 ();
 sg13g2_decap_8 FILLER_80_791 ();
 sg13g2_decap_8 FILLER_80_798 ();
 sg13g2_decap_8 FILLER_80_805 ();
 sg13g2_decap_8 FILLER_80_812 ();
 sg13g2_decap_8 FILLER_80_819 ();
 sg13g2_decap_8 FILLER_80_826 ();
 sg13g2_decap_8 FILLER_80_833 ();
 sg13g2_decap_8 FILLER_80_840 ();
 sg13g2_decap_8 FILLER_80_847 ();
 sg13g2_decap_8 FILLER_80_854 ();
 sg13g2_decap_8 FILLER_80_861 ();
 sg13g2_decap_8 FILLER_80_868 ();
 sg13g2_decap_8 FILLER_80_875 ();
 sg13g2_decap_8 FILLER_80_882 ();
 sg13g2_decap_8 FILLER_80_889 ();
 sg13g2_decap_8 FILLER_80_896 ();
 sg13g2_decap_8 FILLER_80_903 ();
 sg13g2_decap_8 FILLER_80_910 ();
 sg13g2_decap_8 FILLER_80_917 ();
 sg13g2_decap_8 FILLER_80_924 ();
 sg13g2_decap_8 FILLER_80_931 ();
 sg13g2_decap_8 FILLER_80_938 ();
 sg13g2_decap_8 FILLER_80_945 ();
 sg13g2_decap_8 FILLER_80_952 ();
 sg13g2_decap_8 FILLER_80_959 ();
 sg13g2_decap_8 FILLER_80_966 ();
 sg13g2_decap_8 FILLER_80_973 ();
 sg13g2_decap_8 FILLER_80_980 ();
 sg13g2_decap_8 FILLER_80_987 ();
 sg13g2_decap_8 FILLER_80_994 ();
 sg13g2_decap_8 FILLER_80_1001 ();
 sg13g2_decap_8 FILLER_80_1008 ();
 sg13g2_decap_8 FILLER_80_1015 ();
 sg13g2_decap_8 FILLER_80_1022 ();
 sg13g2_decap_8 FILLER_81_4 ();
 sg13g2_decap_8 FILLER_81_11 ();
 sg13g2_decap_8 FILLER_81_18 ();
 sg13g2_decap_8 FILLER_81_25 ();
 sg13g2_decap_8 FILLER_81_32 ();
 sg13g2_decap_8 FILLER_81_39 ();
 sg13g2_decap_8 FILLER_81_46 ();
 sg13g2_decap_8 FILLER_81_53 ();
 sg13g2_decap_8 FILLER_81_60 ();
 sg13g2_decap_8 FILLER_81_67 ();
 sg13g2_decap_8 FILLER_81_74 ();
 sg13g2_decap_8 FILLER_81_81 ();
 sg13g2_decap_8 FILLER_81_88 ();
 sg13g2_decap_8 FILLER_81_95 ();
 sg13g2_decap_8 FILLER_81_102 ();
 sg13g2_decap_8 FILLER_81_109 ();
 sg13g2_decap_8 FILLER_81_116 ();
 sg13g2_decap_8 FILLER_81_123 ();
 sg13g2_decap_8 FILLER_81_130 ();
 sg13g2_decap_8 FILLER_81_137 ();
 sg13g2_decap_8 FILLER_81_144 ();
 sg13g2_decap_8 FILLER_81_151 ();
 sg13g2_decap_8 FILLER_81_158 ();
 sg13g2_decap_8 FILLER_81_165 ();
 sg13g2_decap_8 FILLER_81_172 ();
 sg13g2_decap_8 FILLER_81_179 ();
 sg13g2_decap_8 FILLER_81_186 ();
 sg13g2_decap_8 FILLER_81_193 ();
 sg13g2_decap_8 FILLER_81_200 ();
 sg13g2_decap_8 FILLER_81_207 ();
 sg13g2_decap_8 FILLER_81_214 ();
 sg13g2_decap_8 FILLER_81_221 ();
 sg13g2_decap_8 FILLER_81_228 ();
 sg13g2_decap_8 FILLER_81_235 ();
 sg13g2_decap_8 FILLER_81_242 ();
 sg13g2_decap_8 FILLER_81_249 ();
 sg13g2_decap_8 FILLER_81_256 ();
 sg13g2_decap_8 FILLER_81_263 ();
 sg13g2_decap_8 FILLER_81_270 ();
 sg13g2_decap_8 FILLER_81_277 ();
 sg13g2_decap_8 FILLER_81_284 ();
 sg13g2_decap_8 FILLER_81_291 ();
 sg13g2_decap_8 FILLER_81_298 ();
 sg13g2_decap_8 FILLER_81_305 ();
 sg13g2_decap_8 FILLER_81_312 ();
 sg13g2_decap_8 FILLER_81_319 ();
 sg13g2_decap_8 FILLER_81_326 ();
 sg13g2_decap_8 FILLER_81_333 ();
 sg13g2_decap_8 FILLER_81_340 ();
 sg13g2_decap_8 FILLER_81_347 ();
 sg13g2_decap_8 FILLER_81_354 ();
 sg13g2_decap_8 FILLER_81_361 ();
 sg13g2_decap_8 FILLER_81_368 ();
 sg13g2_decap_8 FILLER_81_375 ();
 sg13g2_decap_8 FILLER_81_382 ();
 sg13g2_decap_8 FILLER_81_389 ();
 sg13g2_decap_8 FILLER_81_396 ();
 sg13g2_decap_8 FILLER_81_403 ();
 sg13g2_decap_8 FILLER_81_410 ();
 sg13g2_decap_8 FILLER_81_417 ();
 sg13g2_decap_8 FILLER_81_424 ();
 sg13g2_decap_8 FILLER_81_431 ();
 sg13g2_decap_8 FILLER_81_438 ();
 sg13g2_decap_8 FILLER_81_445 ();
 sg13g2_decap_8 FILLER_81_452 ();
 sg13g2_decap_8 FILLER_81_459 ();
 sg13g2_decap_8 FILLER_81_466 ();
 sg13g2_decap_8 FILLER_81_473 ();
 sg13g2_decap_8 FILLER_81_480 ();
 sg13g2_decap_8 FILLER_81_487 ();
 sg13g2_decap_8 FILLER_81_494 ();
 sg13g2_decap_8 FILLER_81_501 ();
 sg13g2_decap_8 FILLER_81_508 ();
 sg13g2_decap_8 FILLER_81_515 ();
 sg13g2_decap_8 FILLER_81_522 ();
 sg13g2_decap_8 FILLER_81_529 ();
 sg13g2_decap_8 FILLER_81_536 ();
 sg13g2_decap_8 FILLER_81_543 ();
 sg13g2_decap_8 FILLER_81_550 ();
 sg13g2_decap_8 FILLER_81_557 ();
 sg13g2_decap_8 FILLER_81_564 ();
 sg13g2_decap_8 FILLER_81_571 ();
 sg13g2_decap_8 FILLER_81_578 ();
 sg13g2_decap_8 FILLER_81_585 ();
 sg13g2_decap_8 FILLER_81_592 ();
 sg13g2_decap_8 FILLER_81_599 ();
 sg13g2_decap_8 FILLER_81_606 ();
 sg13g2_decap_8 FILLER_81_613 ();
 sg13g2_decap_8 FILLER_81_620 ();
 sg13g2_decap_8 FILLER_81_627 ();
 sg13g2_decap_8 FILLER_81_634 ();
 sg13g2_decap_8 FILLER_81_641 ();
 sg13g2_decap_8 FILLER_81_648 ();
 sg13g2_decap_8 FILLER_81_655 ();
 sg13g2_decap_8 FILLER_81_662 ();
 sg13g2_decap_8 FILLER_81_669 ();
 sg13g2_decap_8 FILLER_81_676 ();
 sg13g2_decap_8 FILLER_81_683 ();
 sg13g2_decap_8 FILLER_81_690 ();
 sg13g2_decap_8 FILLER_81_697 ();
 sg13g2_decap_8 FILLER_81_704 ();
 sg13g2_decap_8 FILLER_81_711 ();
 sg13g2_decap_8 FILLER_81_718 ();
 sg13g2_decap_8 FILLER_81_725 ();
 sg13g2_decap_8 FILLER_81_732 ();
 sg13g2_decap_8 FILLER_81_739 ();
 sg13g2_decap_8 FILLER_81_746 ();
 sg13g2_decap_8 FILLER_81_753 ();
 sg13g2_decap_8 FILLER_81_760 ();
 sg13g2_decap_8 FILLER_81_767 ();
 sg13g2_decap_8 FILLER_81_774 ();
 sg13g2_decap_8 FILLER_81_781 ();
 sg13g2_decap_8 FILLER_81_788 ();
 sg13g2_decap_8 FILLER_81_795 ();
 sg13g2_decap_8 FILLER_81_802 ();
 sg13g2_decap_8 FILLER_81_809 ();
 sg13g2_decap_8 FILLER_81_816 ();
 sg13g2_decap_8 FILLER_81_823 ();
 sg13g2_decap_8 FILLER_81_830 ();
 sg13g2_decap_8 FILLER_81_837 ();
 sg13g2_decap_8 FILLER_81_844 ();
 sg13g2_decap_8 FILLER_81_851 ();
 sg13g2_decap_8 FILLER_81_858 ();
 sg13g2_decap_8 FILLER_81_865 ();
 sg13g2_decap_8 FILLER_81_872 ();
 sg13g2_decap_8 FILLER_81_879 ();
 sg13g2_decap_8 FILLER_81_886 ();
 sg13g2_decap_8 FILLER_81_893 ();
 sg13g2_decap_8 FILLER_81_900 ();
 sg13g2_decap_8 FILLER_81_907 ();
 sg13g2_decap_8 FILLER_81_914 ();
 sg13g2_decap_8 FILLER_81_921 ();
 sg13g2_decap_8 FILLER_81_928 ();
 sg13g2_decap_8 FILLER_81_935 ();
 sg13g2_decap_8 FILLER_81_942 ();
 sg13g2_decap_8 FILLER_81_949 ();
 sg13g2_decap_8 FILLER_81_956 ();
 sg13g2_decap_8 FILLER_81_963 ();
 sg13g2_decap_8 FILLER_81_970 ();
 sg13g2_decap_8 FILLER_81_977 ();
 sg13g2_decap_8 FILLER_81_984 ();
 sg13g2_decap_8 FILLER_81_991 ();
 sg13g2_decap_8 FILLER_81_998 ();
 sg13g2_decap_8 FILLER_81_1005 ();
 sg13g2_decap_8 FILLER_81_1012 ();
 sg13g2_decap_8 FILLER_81_1019 ();
 sg13g2_fill_2 FILLER_81_1026 ();
 sg13g2_fill_1 FILLER_81_1028 ();
 sg13g2_decap_8 FILLER_82_0 ();
 sg13g2_decap_8 FILLER_82_7 ();
 sg13g2_decap_8 FILLER_82_14 ();
 sg13g2_decap_8 FILLER_82_21 ();
 sg13g2_decap_8 FILLER_82_28 ();
 sg13g2_decap_8 FILLER_82_35 ();
 sg13g2_decap_8 FILLER_82_42 ();
 sg13g2_decap_8 FILLER_82_49 ();
 sg13g2_decap_8 FILLER_82_56 ();
 sg13g2_decap_8 FILLER_82_63 ();
 sg13g2_decap_8 FILLER_82_70 ();
 sg13g2_decap_8 FILLER_82_77 ();
 sg13g2_decap_8 FILLER_82_84 ();
 sg13g2_decap_8 FILLER_82_91 ();
 sg13g2_decap_8 FILLER_82_98 ();
 sg13g2_decap_8 FILLER_82_105 ();
 sg13g2_decap_8 FILLER_82_112 ();
 sg13g2_decap_8 FILLER_82_119 ();
 sg13g2_decap_8 FILLER_82_126 ();
 sg13g2_decap_8 FILLER_82_133 ();
 sg13g2_decap_8 FILLER_82_140 ();
 sg13g2_decap_8 FILLER_82_147 ();
 sg13g2_decap_8 FILLER_82_154 ();
 sg13g2_decap_8 FILLER_82_161 ();
 sg13g2_decap_8 FILLER_82_168 ();
 sg13g2_decap_8 FILLER_82_175 ();
 sg13g2_decap_8 FILLER_82_182 ();
 sg13g2_decap_8 FILLER_82_189 ();
 sg13g2_decap_8 FILLER_82_196 ();
 sg13g2_decap_8 FILLER_82_203 ();
 sg13g2_decap_8 FILLER_82_210 ();
 sg13g2_decap_8 FILLER_82_217 ();
 sg13g2_decap_8 FILLER_82_224 ();
 sg13g2_decap_8 FILLER_82_231 ();
 sg13g2_decap_8 FILLER_82_238 ();
 sg13g2_decap_8 FILLER_82_245 ();
 sg13g2_decap_8 FILLER_82_252 ();
 sg13g2_decap_8 FILLER_82_259 ();
 sg13g2_decap_8 FILLER_82_266 ();
 sg13g2_decap_8 FILLER_82_273 ();
 sg13g2_decap_8 FILLER_82_280 ();
 sg13g2_decap_8 FILLER_82_287 ();
 sg13g2_decap_8 FILLER_82_294 ();
 sg13g2_decap_8 FILLER_82_301 ();
 sg13g2_decap_8 FILLER_82_308 ();
 sg13g2_decap_8 FILLER_82_315 ();
 sg13g2_decap_8 FILLER_82_322 ();
 sg13g2_decap_8 FILLER_82_329 ();
 sg13g2_decap_8 FILLER_82_336 ();
 sg13g2_decap_8 FILLER_82_343 ();
 sg13g2_decap_8 FILLER_82_350 ();
 sg13g2_decap_8 FILLER_82_357 ();
 sg13g2_decap_8 FILLER_82_364 ();
 sg13g2_decap_8 FILLER_82_371 ();
 sg13g2_decap_8 FILLER_82_378 ();
 sg13g2_decap_8 FILLER_82_385 ();
 sg13g2_decap_8 FILLER_82_392 ();
 sg13g2_decap_8 FILLER_82_399 ();
 sg13g2_decap_8 FILLER_82_406 ();
 sg13g2_decap_8 FILLER_82_413 ();
 sg13g2_decap_8 FILLER_82_420 ();
 sg13g2_decap_8 FILLER_82_427 ();
 sg13g2_decap_8 FILLER_82_434 ();
 sg13g2_decap_8 FILLER_82_441 ();
 sg13g2_decap_8 FILLER_82_448 ();
 sg13g2_decap_8 FILLER_82_455 ();
 sg13g2_decap_8 FILLER_82_462 ();
 sg13g2_decap_8 FILLER_82_469 ();
 sg13g2_decap_8 FILLER_82_476 ();
 sg13g2_decap_8 FILLER_82_483 ();
 sg13g2_decap_8 FILLER_82_490 ();
 sg13g2_decap_8 FILLER_82_497 ();
 sg13g2_decap_8 FILLER_82_504 ();
 sg13g2_decap_8 FILLER_82_511 ();
 sg13g2_decap_8 FILLER_82_518 ();
 sg13g2_decap_8 FILLER_82_525 ();
 sg13g2_decap_8 FILLER_82_532 ();
 sg13g2_decap_8 FILLER_82_539 ();
 sg13g2_decap_8 FILLER_82_546 ();
 sg13g2_decap_8 FILLER_82_553 ();
 sg13g2_decap_8 FILLER_82_560 ();
 sg13g2_decap_8 FILLER_82_567 ();
 sg13g2_decap_8 FILLER_82_574 ();
 sg13g2_decap_8 FILLER_82_581 ();
 sg13g2_decap_8 FILLER_82_588 ();
 sg13g2_decap_8 FILLER_82_595 ();
 sg13g2_decap_8 FILLER_82_602 ();
 sg13g2_decap_8 FILLER_82_609 ();
 sg13g2_decap_8 FILLER_82_616 ();
 sg13g2_decap_8 FILLER_82_623 ();
 sg13g2_decap_8 FILLER_82_630 ();
 sg13g2_decap_8 FILLER_82_637 ();
 sg13g2_decap_8 FILLER_82_644 ();
 sg13g2_decap_8 FILLER_82_651 ();
 sg13g2_decap_8 FILLER_82_658 ();
 sg13g2_decap_8 FILLER_82_665 ();
 sg13g2_decap_8 FILLER_82_672 ();
 sg13g2_decap_8 FILLER_82_679 ();
 sg13g2_decap_8 FILLER_82_686 ();
 sg13g2_decap_8 FILLER_82_693 ();
 sg13g2_decap_8 FILLER_82_700 ();
 sg13g2_decap_8 FILLER_82_707 ();
 sg13g2_decap_8 FILLER_82_714 ();
 sg13g2_decap_8 FILLER_82_721 ();
 sg13g2_decap_8 FILLER_82_728 ();
 sg13g2_decap_8 FILLER_82_735 ();
 sg13g2_decap_8 FILLER_82_742 ();
 sg13g2_decap_8 FILLER_82_749 ();
 sg13g2_decap_8 FILLER_82_756 ();
 sg13g2_decap_8 FILLER_82_763 ();
 sg13g2_decap_8 FILLER_82_770 ();
 sg13g2_decap_8 FILLER_82_777 ();
 sg13g2_decap_8 FILLER_82_784 ();
 sg13g2_decap_8 FILLER_82_791 ();
 sg13g2_decap_8 FILLER_82_798 ();
 sg13g2_decap_8 FILLER_82_805 ();
 sg13g2_decap_8 FILLER_82_812 ();
 sg13g2_decap_8 FILLER_82_819 ();
 sg13g2_decap_8 FILLER_82_826 ();
 sg13g2_decap_8 FILLER_82_833 ();
 sg13g2_decap_8 FILLER_82_840 ();
 sg13g2_decap_8 FILLER_82_847 ();
 sg13g2_decap_8 FILLER_82_854 ();
 sg13g2_decap_8 FILLER_82_861 ();
 sg13g2_decap_8 FILLER_82_868 ();
 sg13g2_decap_8 FILLER_82_875 ();
 sg13g2_decap_8 FILLER_82_882 ();
 sg13g2_decap_8 FILLER_82_889 ();
 sg13g2_decap_8 FILLER_82_896 ();
 sg13g2_decap_8 FILLER_82_903 ();
 sg13g2_decap_8 FILLER_82_910 ();
 sg13g2_decap_8 FILLER_82_917 ();
 sg13g2_decap_8 FILLER_82_924 ();
 sg13g2_decap_8 FILLER_82_931 ();
 sg13g2_decap_8 FILLER_82_938 ();
 sg13g2_decap_8 FILLER_82_945 ();
 sg13g2_decap_8 FILLER_82_952 ();
 sg13g2_decap_8 FILLER_82_959 ();
 sg13g2_decap_8 FILLER_82_966 ();
 sg13g2_decap_8 FILLER_82_973 ();
 sg13g2_decap_8 FILLER_82_980 ();
 sg13g2_decap_8 FILLER_82_987 ();
 sg13g2_decap_8 FILLER_82_994 ();
 sg13g2_decap_8 FILLER_82_1001 ();
 sg13g2_decap_8 FILLER_82_1008 ();
 sg13g2_decap_8 FILLER_82_1015 ();
 sg13g2_decap_8 FILLER_82_1022 ();
 sg13g2_decap_8 FILLER_83_4 ();
 sg13g2_decap_8 FILLER_83_11 ();
 sg13g2_decap_8 FILLER_83_18 ();
 sg13g2_decap_8 FILLER_83_25 ();
 sg13g2_decap_8 FILLER_83_32 ();
 sg13g2_decap_8 FILLER_83_39 ();
 sg13g2_decap_8 FILLER_83_46 ();
 sg13g2_decap_8 FILLER_83_53 ();
 sg13g2_decap_8 FILLER_83_60 ();
 sg13g2_decap_8 FILLER_83_67 ();
 sg13g2_decap_8 FILLER_83_74 ();
 sg13g2_decap_8 FILLER_83_81 ();
 sg13g2_decap_8 FILLER_83_88 ();
 sg13g2_decap_8 FILLER_83_95 ();
 sg13g2_decap_8 FILLER_83_102 ();
 sg13g2_decap_8 FILLER_83_109 ();
 sg13g2_decap_8 FILLER_83_116 ();
 sg13g2_decap_8 FILLER_83_123 ();
 sg13g2_decap_8 FILLER_83_130 ();
 sg13g2_decap_8 FILLER_83_137 ();
 sg13g2_decap_8 FILLER_83_144 ();
 sg13g2_decap_8 FILLER_83_151 ();
 sg13g2_decap_8 FILLER_83_158 ();
 sg13g2_decap_8 FILLER_83_165 ();
 sg13g2_decap_8 FILLER_83_172 ();
 sg13g2_decap_8 FILLER_83_179 ();
 sg13g2_decap_8 FILLER_83_186 ();
 sg13g2_decap_8 FILLER_83_193 ();
 sg13g2_decap_8 FILLER_83_200 ();
 sg13g2_decap_8 FILLER_83_207 ();
 sg13g2_decap_8 FILLER_83_214 ();
 sg13g2_decap_8 FILLER_83_221 ();
 sg13g2_decap_8 FILLER_83_228 ();
 sg13g2_decap_8 FILLER_83_235 ();
 sg13g2_decap_8 FILLER_83_242 ();
 sg13g2_decap_8 FILLER_83_249 ();
 sg13g2_decap_8 FILLER_83_256 ();
 sg13g2_decap_8 FILLER_83_263 ();
 sg13g2_decap_8 FILLER_83_270 ();
 sg13g2_decap_8 FILLER_83_277 ();
 sg13g2_decap_8 FILLER_83_284 ();
 sg13g2_decap_8 FILLER_83_291 ();
 sg13g2_decap_8 FILLER_83_298 ();
 sg13g2_decap_8 FILLER_83_305 ();
 sg13g2_decap_8 FILLER_83_312 ();
 sg13g2_decap_8 FILLER_83_319 ();
 sg13g2_decap_8 FILLER_83_326 ();
 sg13g2_decap_8 FILLER_83_333 ();
 sg13g2_decap_8 FILLER_83_340 ();
 sg13g2_decap_8 FILLER_83_347 ();
 sg13g2_decap_8 FILLER_83_354 ();
 sg13g2_decap_8 FILLER_83_361 ();
 sg13g2_decap_8 FILLER_83_368 ();
 sg13g2_decap_8 FILLER_83_375 ();
 sg13g2_decap_8 FILLER_83_382 ();
 sg13g2_decap_8 FILLER_83_389 ();
 sg13g2_decap_8 FILLER_83_396 ();
 sg13g2_decap_8 FILLER_83_403 ();
 sg13g2_decap_8 FILLER_83_410 ();
 sg13g2_decap_8 FILLER_83_417 ();
 sg13g2_decap_8 FILLER_83_424 ();
 sg13g2_decap_8 FILLER_83_431 ();
 sg13g2_decap_8 FILLER_83_438 ();
 sg13g2_decap_8 FILLER_83_445 ();
 sg13g2_decap_8 FILLER_83_452 ();
 sg13g2_decap_8 FILLER_83_459 ();
 sg13g2_decap_8 FILLER_83_466 ();
 sg13g2_decap_8 FILLER_83_473 ();
 sg13g2_decap_8 FILLER_83_480 ();
 sg13g2_decap_8 FILLER_83_487 ();
 sg13g2_decap_8 FILLER_83_494 ();
 sg13g2_decap_8 FILLER_83_501 ();
 sg13g2_decap_8 FILLER_83_508 ();
 sg13g2_decap_8 FILLER_83_515 ();
 sg13g2_decap_8 FILLER_83_522 ();
 sg13g2_decap_8 FILLER_83_529 ();
 sg13g2_decap_8 FILLER_83_536 ();
 sg13g2_decap_8 FILLER_83_543 ();
 sg13g2_decap_8 FILLER_83_550 ();
 sg13g2_decap_8 FILLER_83_557 ();
 sg13g2_decap_8 FILLER_83_564 ();
 sg13g2_decap_8 FILLER_83_571 ();
 sg13g2_decap_8 FILLER_83_578 ();
 sg13g2_decap_8 FILLER_83_585 ();
 sg13g2_decap_8 FILLER_83_592 ();
 sg13g2_decap_8 FILLER_83_599 ();
 sg13g2_decap_8 FILLER_83_606 ();
 sg13g2_decap_8 FILLER_83_613 ();
 sg13g2_decap_8 FILLER_83_620 ();
 sg13g2_decap_8 FILLER_83_627 ();
 sg13g2_decap_8 FILLER_83_634 ();
 sg13g2_decap_8 FILLER_83_641 ();
 sg13g2_decap_8 FILLER_83_648 ();
 sg13g2_decap_8 FILLER_83_655 ();
 sg13g2_decap_8 FILLER_83_662 ();
 sg13g2_decap_8 FILLER_83_669 ();
 sg13g2_decap_8 FILLER_83_676 ();
 sg13g2_decap_8 FILLER_83_683 ();
 sg13g2_decap_8 FILLER_83_690 ();
 sg13g2_decap_8 FILLER_83_697 ();
 sg13g2_decap_8 FILLER_83_704 ();
 sg13g2_decap_8 FILLER_83_711 ();
 sg13g2_decap_8 FILLER_83_718 ();
 sg13g2_decap_8 FILLER_83_725 ();
 sg13g2_decap_8 FILLER_83_732 ();
 sg13g2_decap_8 FILLER_83_739 ();
 sg13g2_decap_8 FILLER_83_746 ();
 sg13g2_decap_8 FILLER_83_753 ();
 sg13g2_decap_8 FILLER_83_760 ();
 sg13g2_decap_8 FILLER_83_767 ();
 sg13g2_decap_8 FILLER_83_774 ();
 sg13g2_decap_8 FILLER_83_781 ();
 sg13g2_decap_8 FILLER_83_788 ();
 sg13g2_decap_8 FILLER_83_795 ();
 sg13g2_decap_8 FILLER_83_802 ();
 sg13g2_decap_8 FILLER_83_809 ();
 sg13g2_decap_8 FILLER_83_816 ();
 sg13g2_decap_8 FILLER_83_823 ();
 sg13g2_decap_8 FILLER_83_830 ();
 sg13g2_decap_8 FILLER_83_837 ();
 sg13g2_decap_8 FILLER_83_844 ();
 sg13g2_decap_8 FILLER_83_851 ();
 sg13g2_decap_8 FILLER_83_858 ();
 sg13g2_decap_8 FILLER_83_865 ();
 sg13g2_decap_8 FILLER_83_872 ();
 sg13g2_decap_8 FILLER_83_879 ();
 sg13g2_decap_8 FILLER_83_886 ();
 sg13g2_decap_8 FILLER_83_893 ();
 sg13g2_decap_8 FILLER_83_900 ();
 sg13g2_decap_8 FILLER_83_907 ();
 sg13g2_decap_8 FILLER_83_914 ();
 sg13g2_decap_8 FILLER_83_921 ();
 sg13g2_decap_8 FILLER_83_928 ();
 sg13g2_decap_8 FILLER_83_935 ();
 sg13g2_decap_8 FILLER_83_942 ();
 sg13g2_decap_8 FILLER_83_949 ();
 sg13g2_decap_8 FILLER_83_956 ();
 sg13g2_decap_8 FILLER_83_963 ();
 sg13g2_decap_8 FILLER_83_970 ();
 sg13g2_decap_8 FILLER_83_977 ();
 sg13g2_decap_8 FILLER_83_984 ();
 sg13g2_decap_8 FILLER_83_991 ();
 sg13g2_decap_8 FILLER_83_998 ();
 sg13g2_decap_8 FILLER_83_1005 ();
 sg13g2_decap_8 FILLER_83_1012 ();
 sg13g2_decap_8 FILLER_83_1019 ();
 sg13g2_fill_2 FILLER_83_1026 ();
 sg13g2_fill_1 FILLER_83_1028 ();
 sg13g2_decap_8 FILLER_84_0 ();
 sg13g2_decap_8 FILLER_84_7 ();
 sg13g2_decap_8 FILLER_84_14 ();
 sg13g2_decap_8 FILLER_84_21 ();
 sg13g2_decap_8 FILLER_84_28 ();
 sg13g2_decap_8 FILLER_84_35 ();
 sg13g2_decap_8 FILLER_84_42 ();
 sg13g2_decap_8 FILLER_84_49 ();
 sg13g2_decap_8 FILLER_84_56 ();
 sg13g2_decap_8 FILLER_84_63 ();
 sg13g2_decap_8 FILLER_84_70 ();
 sg13g2_decap_8 FILLER_84_77 ();
 sg13g2_decap_8 FILLER_84_84 ();
 sg13g2_decap_8 FILLER_84_91 ();
 sg13g2_decap_8 FILLER_84_98 ();
 sg13g2_decap_8 FILLER_84_105 ();
 sg13g2_decap_8 FILLER_84_112 ();
 sg13g2_decap_8 FILLER_84_119 ();
 sg13g2_decap_8 FILLER_84_126 ();
 sg13g2_decap_8 FILLER_84_133 ();
 sg13g2_decap_8 FILLER_84_140 ();
 sg13g2_decap_8 FILLER_84_147 ();
 sg13g2_decap_8 FILLER_84_154 ();
 sg13g2_decap_8 FILLER_84_161 ();
 sg13g2_decap_8 FILLER_84_168 ();
 sg13g2_decap_8 FILLER_84_175 ();
 sg13g2_decap_8 FILLER_84_182 ();
 sg13g2_decap_8 FILLER_84_189 ();
 sg13g2_decap_8 FILLER_84_196 ();
 sg13g2_decap_8 FILLER_84_203 ();
 sg13g2_decap_8 FILLER_84_210 ();
 sg13g2_decap_8 FILLER_84_217 ();
 sg13g2_decap_8 FILLER_84_224 ();
 sg13g2_decap_8 FILLER_84_231 ();
 sg13g2_decap_8 FILLER_84_238 ();
 sg13g2_decap_8 FILLER_84_245 ();
 sg13g2_decap_8 FILLER_84_252 ();
 sg13g2_decap_8 FILLER_84_259 ();
 sg13g2_decap_8 FILLER_84_266 ();
 sg13g2_decap_8 FILLER_84_273 ();
 sg13g2_decap_8 FILLER_84_280 ();
 sg13g2_decap_8 FILLER_84_287 ();
 sg13g2_decap_8 FILLER_84_294 ();
 sg13g2_decap_8 FILLER_84_301 ();
 sg13g2_decap_8 FILLER_84_308 ();
 sg13g2_decap_8 FILLER_84_315 ();
 sg13g2_decap_8 FILLER_84_322 ();
 sg13g2_decap_8 FILLER_84_329 ();
 sg13g2_decap_8 FILLER_84_336 ();
 sg13g2_decap_8 FILLER_84_343 ();
 sg13g2_decap_8 FILLER_84_350 ();
 sg13g2_decap_8 FILLER_84_357 ();
 sg13g2_decap_8 FILLER_84_364 ();
 sg13g2_decap_8 FILLER_84_371 ();
 sg13g2_decap_8 FILLER_84_378 ();
 sg13g2_decap_8 FILLER_84_385 ();
 sg13g2_decap_8 FILLER_84_392 ();
 sg13g2_decap_8 FILLER_84_399 ();
 sg13g2_decap_8 FILLER_84_406 ();
 sg13g2_decap_8 FILLER_84_413 ();
 sg13g2_decap_8 FILLER_84_420 ();
 sg13g2_decap_8 FILLER_84_427 ();
 sg13g2_decap_8 FILLER_84_434 ();
 sg13g2_decap_8 FILLER_84_441 ();
 sg13g2_decap_8 FILLER_84_448 ();
 sg13g2_decap_8 FILLER_84_455 ();
 sg13g2_decap_8 FILLER_84_462 ();
 sg13g2_decap_8 FILLER_84_469 ();
 sg13g2_decap_8 FILLER_84_476 ();
 sg13g2_decap_8 FILLER_84_483 ();
 sg13g2_decap_8 FILLER_84_490 ();
 sg13g2_decap_8 FILLER_84_497 ();
 sg13g2_decap_8 FILLER_84_504 ();
 sg13g2_decap_8 FILLER_84_511 ();
 sg13g2_decap_8 FILLER_84_518 ();
 sg13g2_decap_8 FILLER_84_525 ();
 sg13g2_decap_8 FILLER_84_532 ();
 sg13g2_decap_8 FILLER_84_539 ();
 sg13g2_decap_8 FILLER_84_546 ();
 sg13g2_decap_8 FILLER_84_553 ();
 sg13g2_decap_8 FILLER_84_560 ();
 sg13g2_decap_8 FILLER_84_567 ();
 sg13g2_decap_8 FILLER_84_574 ();
 sg13g2_decap_8 FILLER_84_581 ();
 sg13g2_decap_8 FILLER_84_588 ();
 sg13g2_decap_8 FILLER_84_595 ();
 sg13g2_decap_8 FILLER_84_602 ();
 sg13g2_decap_8 FILLER_84_609 ();
 sg13g2_decap_8 FILLER_84_616 ();
 sg13g2_decap_8 FILLER_84_623 ();
 sg13g2_decap_8 FILLER_84_630 ();
 sg13g2_decap_8 FILLER_84_637 ();
 sg13g2_decap_8 FILLER_84_644 ();
 sg13g2_decap_8 FILLER_84_651 ();
 sg13g2_decap_8 FILLER_84_658 ();
 sg13g2_decap_8 FILLER_84_665 ();
 sg13g2_decap_8 FILLER_84_672 ();
 sg13g2_decap_8 FILLER_84_679 ();
 sg13g2_decap_8 FILLER_84_686 ();
 sg13g2_decap_8 FILLER_84_693 ();
 sg13g2_decap_8 FILLER_84_700 ();
 sg13g2_decap_8 FILLER_84_707 ();
 sg13g2_decap_8 FILLER_84_714 ();
 sg13g2_decap_8 FILLER_84_721 ();
 sg13g2_decap_8 FILLER_84_728 ();
 sg13g2_decap_8 FILLER_84_735 ();
 sg13g2_decap_8 FILLER_84_742 ();
 sg13g2_decap_8 FILLER_84_749 ();
 sg13g2_decap_8 FILLER_84_756 ();
 sg13g2_decap_8 FILLER_84_763 ();
 sg13g2_decap_8 FILLER_84_770 ();
 sg13g2_decap_8 FILLER_84_777 ();
 sg13g2_decap_8 FILLER_84_784 ();
 sg13g2_decap_8 FILLER_84_791 ();
 sg13g2_decap_8 FILLER_84_798 ();
 sg13g2_decap_8 FILLER_84_805 ();
 sg13g2_decap_8 FILLER_84_812 ();
 sg13g2_decap_8 FILLER_84_819 ();
 sg13g2_decap_8 FILLER_84_826 ();
 sg13g2_decap_8 FILLER_84_833 ();
 sg13g2_decap_8 FILLER_84_840 ();
 sg13g2_decap_8 FILLER_84_847 ();
 sg13g2_decap_8 FILLER_84_854 ();
 sg13g2_decap_8 FILLER_84_861 ();
 sg13g2_decap_8 FILLER_84_868 ();
 sg13g2_decap_8 FILLER_84_875 ();
 sg13g2_decap_8 FILLER_84_882 ();
 sg13g2_decap_8 FILLER_84_889 ();
 sg13g2_decap_8 FILLER_84_896 ();
 sg13g2_decap_8 FILLER_84_903 ();
 sg13g2_decap_8 FILLER_84_910 ();
 sg13g2_decap_8 FILLER_84_917 ();
 sg13g2_decap_8 FILLER_84_924 ();
 sg13g2_decap_8 FILLER_84_931 ();
 sg13g2_decap_8 FILLER_84_938 ();
 sg13g2_decap_8 FILLER_84_945 ();
 sg13g2_decap_8 FILLER_84_952 ();
 sg13g2_decap_8 FILLER_84_959 ();
 sg13g2_decap_8 FILLER_84_966 ();
 sg13g2_decap_8 FILLER_84_973 ();
 sg13g2_decap_8 FILLER_84_980 ();
 sg13g2_decap_8 FILLER_84_987 ();
 sg13g2_decap_8 FILLER_84_994 ();
 sg13g2_decap_8 FILLER_84_1001 ();
 sg13g2_decap_8 FILLER_84_1008 ();
 sg13g2_decap_8 FILLER_84_1015 ();
 sg13g2_decap_8 FILLER_84_1022 ();
 sg13g2_decap_8 FILLER_85_0 ();
 sg13g2_decap_8 FILLER_85_7 ();
 sg13g2_decap_8 FILLER_85_14 ();
 sg13g2_decap_8 FILLER_85_21 ();
 sg13g2_decap_8 FILLER_85_28 ();
 sg13g2_decap_8 FILLER_85_35 ();
 sg13g2_decap_8 FILLER_85_42 ();
 sg13g2_decap_8 FILLER_85_49 ();
 sg13g2_decap_8 FILLER_85_56 ();
 sg13g2_decap_8 FILLER_85_63 ();
 sg13g2_decap_8 FILLER_85_70 ();
 sg13g2_decap_8 FILLER_85_77 ();
 sg13g2_decap_8 FILLER_85_84 ();
 sg13g2_decap_8 FILLER_85_91 ();
 sg13g2_decap_8 FILLER_85_98 ();
 sg13g2_decap_8 FILLER_85_105 ();
 sg13g2_decap_8 FILLER_85_112 ();
 sg13g2_decap_8 FILLER_85_119 ();
 sg13g2_decap_8 FILLER_85_126 ();
 sg13g2_decap_8 FILLER_85_133 ();
 sg13g2_decap_8 FILLER_85_140 ();
 sg13g2_decap_8 FILLER_85_147 ();
 sg13g2_decap_8 FILLER_85_154 ();
 sg13g2_decap_8 FILLER_85_161 ();
 sg13g2_decap_8 FILLER_85_168 ();
 sg13g2_decap_8 FILLER_85_175 ();
 sg13g2_decap_8 FILLER_85_182 ();
 sg13g2_decap_8 FILLER_85_189 ();
 sg13g2_decap_8 FILLER_85_196 ();
 sg13g2_decap_8 FILLER_85_203 ();
 sg13g2_decap_8 FILLER_85_210 ();
 sg13g2_decap_8 FILLER_85_217 ();
 sg13g2_decap_8 FILLER_85_224 ();
 sg13g2_decap_8 FILLER_85_231 ();
 sg13g2_decap_8 FILLER_85_238 ();
 sg13g2_decap_8 FILLER_85_245 ();
 sg13g2_decap_8 FILLER_85_252 ();
 sg13g2_decap_8 FILLER_85_259 ();
 sg13g2_decap_8 FILLER_85_266 ();
 sg13g2_decap_8 FILLER_85_273 ();
 sg13g2_decap_8 FILLER_85_280 ();
 sg13g2_decap_8 FILLER_85_287 ();
 sg13g2_decap_8 FILLER_85_294 ();
 sg13g2_decap_8 FILLER_85_301 ();
 sg13g2_decap_8 FILLER_85_308 ();
 sg13g2_decap_8 FILLER_85_315 ();
 sg13g2_decap_8 FILLER_85_322 ();
 sg13g2_decap_8 FILLER_85_329 ();
 sg13g2_decap_8 FILLER_85_336 ();
 sg13g2_decap_8 FILLER_85_343 ();
 sg13g2_decap_8 FILLER_85_350 ();
 sg13g2_decap_8 FILLER_85_357 ();
 sg13g2_decap_8 FILLER_85_364 ();
 sg13g2_decap_8 FILLER_85_371 ();
 sg13g2_decap_8 FILLER_85_378 ();
 sg13g2_decap_8 FILLER_85_385 ();
 sg13g2_decap_8 FILLER_85_392 ();
 sg13g2_decap_8 FILLER_85_399 ();
 sg13g2_decap_8 FILLER_85_406 ();
 sg13g2_decap_8 FILLER_85_413 ();
 sg13g2_decap_8 FILLER_85_420 ();
 sg13g2_decap_8 FILLER_85_427 ();
 sg13g2_decap_8 FILLER_85_434 ();
 sg13g2_decap_8 FILLER_85_441 ();
 sg13g2_decap_8 FILLER_85_448 ();
 sg13g2_decap_8 FILLER_85_455 ();
 sg13g2_decap_8 FILLER_85_462 ();
 sg13g2_decap_8 FILLER_85_469 ();
 sg13g2_decap_8 FILLER_85_476 ();
 sg13g2_decap_8 FILLER_85_483 ();
 sg13g2_decap_8 FILLER_85_490 ();
 sg13g2_decap_8 FILLER_85_497 ();
 sg13g2_decap_8 FILLER_85_504 ();
 sg13g2_decap_8 FILLER_85_511 ();
 sg13g2_decap_8 FILLER_85_518 ();
 sg13g2_decap_8 FILLER_85_525 ();
 sg13g2_decap_8 FILLER_85_532 ();
 sg13g2_decap_8 FILLER_85_539 ();
 sg13g2_decap_8 FILLER_85_546 ();
 sg13g2_decap_8 FILLER_85_553 ();
 sg13g2_decap_8 FILLER_85_560 ();
 sg13g2_decap_8 FILLER_85_567 ();
 sg13g2_decap_8 FILLER_85_574 ();
 sg13g2_decap_8 FILLER_85_581 ();
 sg13g2_decap_8 FILLER_85_588 ();
 sg13g2_decap_8 FILLER_85_595 ();
 sg13g2_decap_8 FILLER_85_602 ();
 sg13g2_decap_8 FILLER_85_609 ();
 sg13g2_decap_8 FILLER_85_616 ();
 sg13g2_decap_8 FILLER_85_623 ();
 sg13g2_decap_8 FILLER_85_630 ();
 sg13g2_decap_8 FILLER_85_637 ();
 sg13g2_decap_8 FILLER_85_644 ();
 sg13g2_decap_8 FILLER_85_651 ();
 sg13g2_decap_8 FILLER_85_658 ();
 sg13g2_decap_8 FILLER_85_665 ();
 sg13g2_decap_8 FILLER_85_672 ();
 sg13g2_decap_8 FILLER_85_679 ();
 sg13g2_decap_8 FILLER_85_686 ();
 sg13g2_decap_8 FILLER_85_693 ();
 sg13g2_decap_8 FILLER_85_700 ();
 sg13g2_decap_8 FILLER_85_707 ();
 sg13g2_decap_8 FILLER_85_714 ();
 sg13g2_decap_8 FILLER_85_721 ();
 sg13g2_decap_8 FILLER_85_728 ();
 sg13g2_decap_8 FILLER_85_735 ();
 sg13g2_decap_8 FILLER_85_742 ();
 sg13g2_decap_8 FILLER_85_749 ();
 sg13g2_decap_8 FILLER_85_756 ();
 sg13g2_decap_8 FILLER_85_763 ();
 sg13g2_decap_8 FILLER_85_770 ();
 sg13g2_decap_8 FILLER_85_777 ();
 sg13g2_decap_8 FILLER_85_784 ();
 sg13g2_decap_8 FILLER_85_791 ();
 sg13g2_decap_8 FILLER_85_798 ();
 sg13g2_decap_8 FILLER_85_805 ();
 sg13g2_decap_8 FILLER_85_812 ();
 sg13g2_decap_8 FILLER_85_819 ();
 sg13g2_decap_8 FILLER_85_826 ();
 sg13g2_decap_8 FILLER_85_833 ();
 sg13g2_decap_8 FILLER_85_840 ();
 sg13g2_decap_8 FILLER_85_847 ();
 sg13g2_decap_8 FILLER_85_854 ();
 sg13g2_decap_8 FILLER_85_861 ();
 sg13g2_decap_8 FILLER_85_868 ();
 sg13g2_decap_8 FILLER_85_875 ();
 sg13g2_decap_8 FILLER_85_882 ();
 sg13g2_decap_8 FILLER_85_889 ();
 sg13g2_decap_8 FILLER_85_896 ();
 sg13g2_decap_8 FILLER_85_903 ();
 sg13g2_decap_8 FILLER_85_910 ();
 sg13g2_decap_8 FILLER_85_917 ();
 sg13g2_decap_8 FILLER_85_924 ();
 sg13g2_decap_8 FILLER_85_931 ();
 sg13g2_decap_8 FILLER_85_938 ();
 sg13g2_decap_8 FILLER_85_945 ();
 sg13g2_decap_8 FILLER_85_952 ();
 sg13g2_decap_8 FILLER_85_959 ();
 sg13g2_decap_8 FILLER_85_966 ();
 sg13g2_decap_8 FILLER_85_973 ();
 sg13g2_decap_8 FILLER_85_980 ();
 sg13g2_decap_8 FILLER_85_987 ();
 sg13g2_decap_8 FILLER_85_994 ();
 sg13g2_decap_8 FILLER_85_1001 ();
 sg13g2_decap_8 FILLER_85_1008 ();
 sg13g2_decap_8 FILLER_85_1015 ();
 sg13g2_decap_8 FILLER_85_1022 ();
 sg13g2_decap_8 FILLER_86_4 ();
 sg13g2_decap_8 FILLER_86_11 ();
 sg13g2_decap_8 FILLER_86_18 ();
 sg13g2_decap_8 FILLER_86_25 ();
 sg13g2_decap_8 FILLER_86_32 ();
 sg13g2_decap_8 FILLER_86_39 ();
 sg13g2_decap_8 FILLER_86_46 ();
 sg13g2_decap_8 FILLER_86_53 ();
 sg13g2_decap_8 FILLER_86_60 ();
 sg13g2_decap_8 FILLER_86_67 ();
 sg13g2_decap_8 FILLER_86_74 ();
 sg13g2_decap_8 FILLER_86_81 ();
 sg13g2_decap_8 FILLER_86_88 ();
 sg13g2_decap_8 FILLER_86_95 ();
 sg13g2_decap_8 FILLER_86_102 ();
 sg13g2_decap_8 FILLER_86_109 ();
 sg13g2_decap_8 FILLER_86_116 ();
 sg13g2_decap_8 FILLER_86_123 ();
 sg13g2_decap_8 FILLER_86_130 ();
 sg13g2_decap_8 FILLER_86_137 ();
 sg13g2_decap_8 FILLER_86_144 ();
 sg13g2_decap_8 FILLER_86_151 ();
 sg13g2_decap_8 FILLER_86_158 ();
 sg13g2_decap_8 FILLER_86_165 ();
 sg13g2_decap_8 FILLER_86_172 ();
 sg13g2_decap_8 FILLER_86_179 ();
 sg13g2_decap_8 FILLER_86_186 ();
 sg13g2_decap_8 FILLER_86_193 ();
 sg13g2_decap_8 FILLER_86_200 ();
 sg13g2_decap_8 FILLER_86_207 ();
 sg13g2_decap_8 FILLER_86_214 ();
 sg13g2_decap_8 FILLER_86_221 ();
 sg13g2_decap_8 FILLER_86_228 ();
 sg13g2_decap_8 FILLER_86_235 ();
 sg13g2_decap_8 FILLER_86_242 ();
 sg13g2_decap_8 FILLER_86_249 ();
 sg13g2_decap_8 FILLER_86_256 ();
 sg13g2_decap_8 FILLER_86_263 ();
 sg13g2_decap_8 FILLER_86_270 ();
 sg13g2_decap_8 FILLER_86_277 ();
 sg13g2_decap_8 FILLER_86_284 ();
 sg13g2_decap_8 FILLER_86_291 ();
 sg13g2_decap_8 FILLER_86_298 ();
 sg13g2_decap_8 FILLER_86_305 ();
 sg13g2_decap_8 FILLER_86_312 ();
 sg13g2_decap_8 FILLER_86_319 ();
 sg13g2_decap_8 FILLER_86_326 ();
 sg13g2_decap_8 FILLER_86_333 ();
 sg13g2_decap_8 FILLER_86_340 ();
 sg13g2_decap_8 FILLER_86_347 ();
 sg13g2_decap_8 FILLER_86_354 ();
 sg13g2_decap_8 FILLER_86_361 ();
 sg13g2_decap_8 FILLER_86_368 ();
 sg13g2_decap_8 FILLER_86_375 ();
 sg13g2_decap_8 FILLER_86_382 ();
 sg13g2_decap_8 FILLER_86_389 ();
 sg13g2_decap_8 FILLER_86_396 ();
 sg13g2_decap_8 FILLER_86_403 ();
 sg13g2_decap_8 FILLER_86_410 ();
 sg13g2_decap_8 FILLER_86_417 ();
 sg13g2_decap_8 FILLER_86_424 ();
 sg13g2_decap_8 FILLER_86_431 ();
 sg13g2_decap_8 FILLER_86_438 ();
 sg13g2_decap_8 FILLER_86_445 ();
 sg13g2_decap_8 FILLER_86_452 ();
 sg13g2_decap_8 FILLER_86_459 ();
 sg13g2_decap_8 FILLER_86_466 ();
 sg13g2_decap_8 FILLER_86_473 ();
 sg13g2_decap_8 FILLER_86_480 ();
 sg13g2_decap_8 FILLER_86_487 ();
 sg13g2_decap_8 FILLER_86_494 ();
 sg13g2_decap_8 FILLER_86_501 ();
 sg13g2_decap_8 FILLER_86_508 ();
 sg13g2_decap_8 FILLER_86_515 ();
 sg13g2_decap_8 FILLER_86_522 ();
 sg13g2_decap_8 FILLER_86_529 ();
 sg13g2_decap_8 FILLER_86_536 ();
 sg13g2_decap_8 FILLER_86_543 ();
 sg13g2_decap_8 FILLER_86_550 ();
 sg13g2_decap_8 FILLER_86_557 ();
 sg13g2_decap_8 FILLER_86_564 ();
 sg13g2_decap_8 FILLER_86_571 ();
 sg13g2_decap_8 FILLER_86_578 ();
 sg13g2_decap_8 FILLER_86_585 ();
 sg13g2_decap_8 FILLER_86_592 ();
 sg13g2_decap_8 FILLER_86_599 ();
 sg13g2_decap_8 FILLER_86_606 ();
 sg13g2_decap_8 FILLER_86_613 ();
 sg13g2_decap_8 FILLER_86_620 ();
 sg13g2_decap_8 FILLER_86_627 ();
 sg13g2_decap_8 FILLER_86_634 ();
 sg13g2_decap_8 FILLER_86_641 ();
 sg13g2_decap_8 FILLER_86_648 ();
 sg13g2_decap_8 FILLER_86_655 ();
 sg13g2_decap_8 FILLER_86_662 ();
 sg13g2_decap_8 FILLER_86_669 ();
 sg13g2_decap_8 FILLER_86_676 ();
 sg13g2_decap_8 FILLER_86_683 ();
 sg13g2_decap_8 FILLER_86_690 ();
 sg13g2_decap_8 FILLER_86_697 ();
 sg13g2_decap_8 FILLER_86_704 ();
 sg13g2_decap_8 FILLER_86_711 ();
 sg13g2_decap_8 FILLER_86_718 ();
 sg13g2_decap_8 FILLER_86_725 ();
 sg13g2_decap_8 FILLER_86_732 ();
 sg13g2_decap_8 FILLER_86_739 ();
 sg13g2_decap_8 FILLER_86_746 ();
 sg13g2_decap_8 FILLER_86_753 ();
 sg13g2_decap_8 FILLER_86_760 ();
 sg13g2_decap_8 FILLER_86_767 ();
 sg13g2_decap_8 FILLER_86_774 ();
 sg13g2_decap_8 FILLER_86_781 ();
 sg13g2_decap_8 FILLER_86_788 ();
 sg13g2_decap_8 FILLER_86_795 ();
 sg13g2_decap_8 FILLER_86_802 ();
 sg13g2_decap_8 FILLER_86_809 ();
 sg13g2_decap_8 FILLER_86_816 ();
 sg13g2_decap_8 FILLER_86_823 ();
 sg13g2_decap_8 FILLER_86_830 ();
 sg13g2_decap_8 FILLER_86_837 ();
 sg13g2_decap_8 FILLER_86_844 ();
 sg13g2_decap_8 FILLER_86_851 ();
 sg13g2_decap_8 FILLER_86_858 ();
 sg13g2_decap_8 FILLER_86_865 ();
 sg13g2_decap_8 FILLER_86_872 ();
 sg13g2_decap_8 FILLER_86_879 ();
 sg13g2_decap_8 FILLER_86_886 ();
 sg13g2_decap_8 FILLER_86_893 ();
 sg13g2_decap_8 FILLER_86_900 ();
 sg13g2_decap_8 FILLER_86_907 ();
 sg13g2_decap_8 FILLER_86_914 ();
 sg13g2_decap_8 FILLER_86_921 ();
 sg13g2_decap_8 FILLER_86_928 ();
 sg13g2_decap_8 FILLER_86_935 ();
 sg13g2_decap_8 FILLER_86_942 ();
 sg13g2_decap_8 FILLER_86_949 ();
 sg13g2_decap_8 FILLER_86_956 ();
 sg13g2_decap_8 FILLER_86_963 ();
 sg13g2_decap_8 FILLER_86_970 ();
 sg13g2_decap_8 FILLER_86_977 ();
 sg13g2_decap_8 FILLER_86_984 ();
 sg13g2_decap_8 FILLER_86_991 ();
 sg13g2_decap_8 FILLER_86_998 ();
 sg13g2_decap_8 FILLER_86_1005 ();
 sg13g2_decap_8 FILLER_86_1012 ();
 sg13g2_decap_8 FILLER_86_1019 ();
 sg13g2_fill_2 FILLER_86_1026 ();
 sg13g2_fill_1 FILLER_86_1028 ();
 sg13g2_decap_8 FILLER_87_0 ();
 sg13g2_decap_8 FILLER_87_7 ();
 sg13g2_decap_8 FILLER_87_14 ();
 sg13g2_decap_8 FILLER_87_21 ();
 sg13g2_decap_8 FILLER_87_28 ();
 sg13g2_decap_8 FILLER_87_35 ();
 sg13g2_decap_8 FILLER_87_42 ();
 sg13g2_decap_8 FILLER_87_49 ();
 sg13g2_decap_8 FILLER_87_56 ();
 sg13g2_decap_8 FILLER_87_63 ();
 sg13g2_decap_8 FILLER_87_70 ();
 sg13g2_decap_8 FILLER_87_77 ();
 sg13g2_decap_8 FILLER_87_84 ();
 sg13g2_decap_8 FILLER_87_91 ();
 sg13g2_decap_8 FILLER_87_98 ();
 sg13g2_decap_8 FILLER_87_105 ();
 sg13g2_decap_8 FILLER_87_112 ();
 sg13g2_decap_8 FILLER_87_119 ();
 sg13g2_decap_8 FILLER_87_126 ();
 sg13g2_decap_8 FILLER_87_133 ();
 sg13g2_decap_8 FILLER_87_140 ();
 sg13g2_decap_8 FILLER_87_147 ();
 sg13g2_decap_8 FILLER_87_154 ();
 sg13g2_decap_8 FILLER_87_161 ();
 sg13g2_decap_8 FILLER_87_168 ();
 sg13g2_decap_8 FILLER_87_175 ();
 sg13g2_decap_8 FILLER_87_182 ();
 sg13g2_decap_8 FILLER_87_189 ();
 sg13g2_decap_8 FILLER_87_196 ();
 sg13g2_decap_8 FILLER_87_203 ();
 sg13g2_decap_8 FILLER_87_210 ();
 sg13g2_decap_8 FILLER_87_217 ();
 sg13g2_decap_8 FILLER_87_224 ();
 sg13g2_decap_8 FILLER_87_231 ();
 sg13g2_decap_8 FILLER_87_238 ();
 sg13g2_decap_8 FILLER_87_245 ();
 sg13g2_decap_8 FILLER_87_252 ();
 sg13g2_decap_8 FILLER_87_259 ();
 sg13g2_decap_8 FILLER_87_266 ();
 sg13g2_decap_8 FILLER_87_273 ();
 sg13g2_decap_8 FILLER_87_280 ();
 sg13g2_decap_8 FILLER_87_287 ();
 sg13g2_decap_8 FILLER_87_294 ();
 sg13g2_decap_8 FILLER_87_301 ();
 sg13g2_decap_8 FILLER_87_308 ();
 sg13g2_decap_8 FILLER_87_315 ();
 sg13g2_decap_8 FILLER_87_322 ();
 sg13g2_decap_8 FILLER_87_329 ();
 sg13g2_decap_8 FILLER_87_336 ();
 sg13g2_decap_8 FILLER_87_343 ();
 sg13g2_decap_8 FILLER_87_350 ();
 sg13g2_decap_8 FILLER_87_357 ();
 sg13g2_decap_8 FILLER_87_364 ();
 sg13g2_decap_8 FILLER_87_371 ();
 sg13g2_decap_8 FILLER_87_378 ();
 sg13g2_decap_8 FILLER_87_385 ();
 sg13g2_decap_8 FILLER_87_392 ();
 sg13g2_decap_8 FILLER_87_399 ();
 sg13g2_decap_8 FILLER_87_406 ();
 sg13g2_decap_8 FILLER_87_413 ();
 sg13g2_decap_8 FILLER_87_420 ();
 sg13g2_decap_8 FILLER_87_427 ();
 sg13g2_decap_8 FILLER_87_434 ();
 sg13g2_decap_8 FILLER_87_441 ();
 sg13g2_decap_8 FILLER_87_448 ();
 sg13g2_decap_8 FILLER_87_455 ();
 sg13g2_decap_8 FILLER_87_462 ();
 sg13g2_decap_8 FILLER_87_469 ();
 sg13g2_decap_8 FILLER_87_476 ();
 sg13g2_decap_8 FILLER_87_483 ();
 sg13g2_decap_8 FILLER_87_490 ();
 sg13g2_decap_8 FILLER_87_497 ();
 sg13g2_decap_8 FILLER_87_504 ();
 sg13g2_decap_8 FILLER_87_511 ();
 sg13g2_decap_8 FILLER_87_518 ();
 sg13g2_decap_8 FILLER_87_525 ();
 sg13g2_decap_8 FILLER_87_532 ();
 sg13g2_decap_8 FILLER_87_539 ();
 sg13g2_decap_8 FILLER_87_546 ();
 sg13g2_decap_8 FILLER_87_553 ();
 sg13g2_decap_8 FILLER_87_560 ();
 sg13g2_decap_8 FILLER_87_567 ();
 sg13g2_decap_8 FILLER_87_574 ();
 sg13g2_decap_8 FILLER_87_581 ();
 sg13g2_decap_8 FILLER_87_588 ();
 sg13g2_decap_8 FILLER_87_595 ();
 sg13g2_decap_8 FILLER_87_602 ();
 sg13g2_decap_8 FILLER_87_609 ();
 sg13g2_decap_8 FILLER_87_616 ();
 sg13g2_decap_8 FILLER_87_623 ();
 sg13g2_decap_8 FILLER_87_630 ();
 sg13g2_decap_8 FILLER_87_637 ();
 sg13g2_decap_8 FILLER_87_644 ();
 sg13g2_decap_8 FILLER_87_651 ();
 sg13g2_decap_8 FILLER_87_658 ();
 sg13g2_decap_8 FILLER_87_665 ();
 sg13g2_decap_8 FILLER_87_672 ();
 sg13g2_decap_8 FILLER_87_679 ();
 sg13g2_decap_8 FILLER_87_686 ();
 sg13g2_decap_8 FILLER_87_693 ();
 sg13g2_decap_8 FILLER_87_700 ();
 sg13g2_decap_8 FILLER_87_707 ();
 sg13g2_decap_8 FILLER_87_714 ();
 sg13g2_decap_8 FILLER_87_721 ();
 sg13g2_decap_8 FILLER_87_728 ();
 sg13g2_decap_8 FILLER_87_735 ();
 sg13g2_decap_8 FILLER_87_742 ();
 sg13g2_decap_8 FILLER_87_749 ();
 sg13g2_decap_8 FILLER_87_756 ();
 sg13g2_decap_8 FILLER_87_763 ();
 sg13g2_decap_8 FILLER_87_770 ();
 sg13g2_decap_8 FILLER_87_777 ();
 sg13g2_decap_8 FILLER_87_784 ();
 sg13g2_decap_8 FILLER_87_791 ();
 sg13g2_decap_8 FILLER_87_798 ();
 sg13g2_decap_8 FILLER_87_805 ();
 sg13g2_decap_8 FILLER_87_812 ();
 sg13g2_decap_8 FILLER_87_819 ();
 sg13g2_decap_8 FILLER_87_826 ();
 sg13g2_decap_8 FILLER_87_833 ();
 sg13g2_decap_8 FILLER_87_840 ();
 sg13g2_decap_8 FILLER_87_847 ();
 sg13g2_decap_8 FILLER_87_854 ();
 sg13g2_decap_8 FILLER_87_861 ();
 sg13g2_decap_8 FILLER_87_868 ();
 sg13g2_decap_8 FILLER_87_875 ();
 sg13g2_decap_8 FILLER_87_882 ();
 sg13g2_decap_8 FILLER_87_889 ();
 sg13g2_decap_8 FILLER_87_896 ();
 sg13g2_decap_8 FILLER_87_903 ();
 sg13g2_decap_8 FILLER_87_910 ();
 sg13g2_decap_8 FILLER_87_917 ();
 sg13g2_decap_8 FILLER_87_924 ();
 sg13g2_decap_8 FILLER_87_931 ();
 sg13g2_decap_8 FILLER_87_938 ();
 sg13g2_decap_8 FILLER_87_945 ();
 sg13g2_decap_8 FILLER_87_952 ();
 sg13g2_decap_8 FILLER_87_959 ();
 sg13g2_decap_8 FILLER_87_966 ();
 sg13g2_decap_8 FILLER_87_973 ();
 sg13g2_decap_8 FILLER_87_980 ();
 sg13g2_decap_8 FILLER_87_987 ();
 sg13g2_decap_8 FILLER_87_994 ();
 sg13g2_decap_8 FILLER_87_1001 ();
 sg13g2_decap_8 FILLER_87_1008 ();
 sg13g2_decap_8 FILLER_87_1015 ();
 sg13g2_decap_8 FILLER_87_1022 ();
 sg13g2_decap_8 FILLER_88_4 ();
 sg13g2_decap_8 FILLER_88_11 ();
 sg13g2_decap_8 FILLER_88_18 ();
 sg13g2_decap_8 FILLER_88_25 ();
 sg13g2_decap_8 FILLER_88_32 ();
 sg13g2_decap_8 FILLER_88_39 ();
 sg13g2_decap_8 FILLER_88_46 ();
 sg13g2_decap_8 FILLER_88_53 ();
 sg13g2_decap_8 FILLER_88_60 ();
 sg13g2_decap_8 FILLER_88_67 ();
 sg13g2_decap_8 FILLER_88_74 ();
 sg13g2_decap_8 FILLER_88_81 ();
 sg13g2_decap_8 FILLER_88_88 ();
 sg13g2_decap_8 FILLER_88_95 ();
 sg13g2_decap_8 FILLER_88_102 ();
 sg13g2_decap_8 FILLER_88_109 ();
 sg13g2_decap_8 FILLER_88_116 ();
 sg13g2_decap_8 FILLER_88_123 ();
 sg13g2_decap_8 FILLER_88_130 ();
 sg13g2_decap_8 FILLER_88_137 ();
 sg13g2_decap_8 FILLER_88_144 ();
 sg13g2_decap_8 FILLER_88_151 ();
 sg13g2_decap_8 FILLER_88_158 ();
 sg13g2_decap_8 FILLER_88_165 ();
 sg13g2_decap_8 FILLER_88_172 ();
 sg13g2_decap_8 FILLER_88_179 ();
 sg13g2_decap_8 FILLER_88_186 ();
 sg13g2_decap_8 FILLER_88_193 ();
 sg13g2_decap_8 FILLER_88_200 ();
 sg13g2_decap_8 FILLER_88_207 ();
 sg13g2_decap_8 FILLER_88_214 ();
 sg13g2_decap_8 FILLER_88_221 ();
 sg13g2_decap_8 FILLER_88_228 ();
 sg13g2_decap_8 FILLER_88_235 ();
 sg13g2_decap_8 FILLER_88_242 ();
 sg13g2_decap_8 FILLER_88_249 ();
 sg13g2_decap_8 FILLER_88_256 ();
 sg13g2_decap_8 FILLER_88_263 ();
 sg13g2_decap_8 FILLER_88_270 ();
 sg13g2_decap_8 FILLER_88_277 ();
 sg13g2_decap_8 FILLER_88_284 ();
 sg13g2_decap_8 FILLER_88_291 ();
 sg13g2_decap_8 FILLER_88_298 ();
 sg13g2_decap_8 FILLER_88_305 ();
 sg13g2_decap_8 FILLER_88_312 ();
 sg13g2_decap_8 FILLER_88_319 ();
 sg13g2_decap_8 FILLER_88_326 ();
 sg13g2_decap_8 FILLER_88_333 ();
 sg13g2_decap_8 FILLER_88_340 ();
 sg13g2_decap_8 FILLER_88_347 ();
 sg13g2_decap_8 FILLER_88_354 ();
 sg13g2_decap_8 FILLER_88_361 ();
 sg13g2_decap_8 FILLER_88_368 ();
 sg13g2_decap_8 FILLER_88_375 ();
 sg13g2_decap_8 FILLER_88_382 ();
 sg13g2_decap_8 FILLER_88_389 ();
 sg13g2_decap_8 FILLER_88_396 ();
 sg13g2_decap_8 FILLER_88_403 ();
 sg13g2_decap_8 FILLER_88_410 ();
 sg13g2_decap_8 FILLER_88_417 ();
 sg13g2_decap_8 FILLER_88_424 ();
 sg13g2_decap_8 FILLER_88_431 ();
 sg13g2_decap_8 FILLER_88_438 ();
 sg13g2_decap_8 FILLER_88_445 ();
 sg13g2_decap_8 FILLER_88_452 ();
 sg13g2_decap_8 FILLER_88_459 ();
 sg13g2_decap_8 FILLER_88_466 ();
 sg13g2_decap_8 FILLER_88_473 ();
 sg13g2_decap_8 FILLER_88_480 ();
 sg13g2_decap_8 FILLER_88_487 ();
 sg13g2_decap_8 FILLER_88_494 ();
 sg13g2_decap_8 FILLER_88_501 ();
 sg13g2_decap_8 FILLER_88_508 ();
 sg13g2_decap_8 FILLER_88_515 ();
 sg13g2_decap_8 FILLER_88_522 ();
 sg13g2_decap_8 FILLER_88_529 ();
 sg13g2_decap_8 FILLER_88_536 ();
 sg13g2_decap_8 FILLER_88_543 ();
 sg13g2_decap_8 FILLER_88_550 ();
 sg13g2_decap_8 FILLER_88_557 ();
 sg13g2_decap_8 FILLER_88_564 ();
 sg13g2_decap_8 FILLER_88_571 ();
 sg13g2_decap_8 FILLER_88_578 ();
 sg13g2_decap_8 FILLER_88_585 ();
 sg13g2_decap_8 FILLER_88_592 ();
 sg13g2_decap_8 FILLER_88_599 ();
 sg13g2_decap_8 FILLER_88_606 ();
 sg13g2_decap_8 FILLER_88_613 ();
 sg13g2_decap_8 FILLER_88_620 ();
 sg13g2_decap_8 FILLER_88_627 ();
 sg13g2_decap_8 FILLER_88_634 ();
 sg13g2_decap_8 FILLER_88_641 ();
 sg13g2_decap_8 FILLER_88_648 ();
 sg13g2_decap_8 FILLER_88_655 ();
 sg13g2_decap_8 FILLER_88_662 ();
 sg13g2_decap_8 FILLER_88_669 ();
 sg13g2_decap_8 FILLER_88_676 ();
 sg13g2_decap_8 FILLER_88_683 ();
 sg13g2_decap_8 FILLER_88_690 ();
 sg13g2_decap_8 FILLER_88_697 ();
 sg13g2_decap_8 FILLER_88_704 ();
 sg13g2_decap_8 FILLER_88_711 ();
 sg13g2_decap_8 FILLER_88_718 ();
 sg13g2_decap_8 FILLER_88_725 ();
 sg13g2_decap_8 FILLER_88_732 ();
 sg13g2_decap_8 FILLER_88_739 ();
 sg13g2_decap_8 FILLER_88_746 ();
 sg13g2_decap_8 FILLER_88_753 ();
 sg13g2_decap_8 FILLER_88_760 ();
 sg13g2_decap_8 FILLER_88_767 ();
 sg13g2_decap_8 FILLER_88_774 ();
 sg13g2_decap_8 FILLER_88_781 ();
 sg13g2_decap_8 FILLER_88_788 ();
 sg13g2_decap_8 FILLER_88_795 ();
 sg13g2_decap_8 FILLER_88_802 ();
 sg13g2_decap_8 FILLER_88_809 ();
 sg13g2_decap_8 FILLER_88_816 ();
 sg13g2_decap_8 FILLER_88_823 ();
 sg13g2_decap_8 FILLER_88_830 ();
 sg13g2_decap_8 FILLER_88_837 ();
 sg13g2_decap_8 FILLER_88_844 ();
 sg13g2_decap_8 FILLER_88_851 ();
 sg13g2_decap_8 FILLER_88_858 ();
 sg13g2_decap_8 FILLER_88_865 ();
 sg13g2_decap_8 FILLER_88_872 ();
 sg13g2_decap_8 FILLER_88_879 ();
 sg13g2_decap_8 FILLER_88_886 ();
 sg13g2_decap_8 FILLER_88_893 ();
 sg13g2_decap_8 FILLER_88_900 ();
 sg13g2_decap_8 FILLER_88_907 ();
 sg13g2_decap_8 FILLER_88_914 ();
 sg13g2_decap_8 FILLER_88_921 ();
 sg13g2_decap_8 FILLER_88_928 ();
 sg13g2_decap_8 FILLER_88_935 ();
 sg13g2_decap_8 FILLER_88_942 ();
 sg13g2_decap_8 FILLER_88_949 ();
 sg13g2_decap_8 FILLER_88_956 ();
 sg13g2_decap_8 FILLER_88_963 ();
 sg13g2_decap_8 FILLER_88_970 ();
 sg13g2_decap_8 FILLER_88_977 ();
 sg13g2_decap_8 FILLER_88_984 ();
 sg13g2_decap_8 FILLER_88_991 ();
 sg13g2_decap_8 FILLER_88_998 ();
 sg13g2_decap_8 FILLER_88_1005 ();
 sg13g2_decap_8 FILLER_88_1012 ();
 sg13g2_decap_8 FILLER_88_1019 ();
 sg13g2_fill_2 FILLER_88_1026 ();
 sg13g2_fill_1 FILLER_88_1028 ();
 sg13g2_decap_8 FILLER_89_0 ();
 sg13g2_decap_8 FILLER_89_7 ();
 sg13g2_decap_8 FILLER_89_14 ();
 sg13g2_decap_8 FILLER_89_21 ();
 sg13g2_decap_8 FILLER_89_28 ();
 sg13g2_decap_8 FILLER_89_35 ();
 sg13g2_decap_8 FILLER_89_42 ();
 sg13g2_decap_8 FILLER_89_49 ();
 sg13g2_decap_8 FILLER_89_56 ();
 sg13g2_decap_8 FILLER_89_63 ();
 sg13g2_decap_8 FILLER_89_70 ();
 sg13g2_decap_8 FILLER_89_77 ();
 sg13g2_decap_8 FILLER_89_84 ();
 sg13g2_decap_8 FILLER_89_91 ();
 sg13g2_decap_8 FILLER_89_98 ();
 sg13g2_decap_8 FILLER_89_105 ();
 sg13g2_decap_8 FILLER_89_112 ();
 sg13g2_decap_8 FILLER_89_119 ();
 sg13g2_decap_8 FILLER_89_126 ();
 sg13g2_decap_8 FILLER_89_133 ();
 sg13g2_decap_8 FILLER_89_140 ();
 sg13g2_decap_8 FILLER_89_147 ();
 sg13g2_decap_8 FILLER_89_154 ();
 sg13g2_decap_8 FILLER_89_161 ();
 sg13g2_decap_8 FILLER_89_168 ();
 sg13g2_decap_8 FILLER_89_175 ();
 sg13g2_decap_8 FILLER_89_182 ();
 sg13g2_decap_8 FILLER_89_189 ();
 sg13g2_decap_8 FILLER_89_196 ();
 sg13g2_decap_8 FILLER_89_203 ();
 sg13g2_decap_8 FILLER_89_210 ();
 sg13g2_decap_8 FILLER_89_217 ();
 sg13g2_decap_8 FILLER_89_224 ();
 sg13g2_decap_8 FILLER_89_231 ();
 sg13g2_decap_8 FILLER_89_238 ();
 sg13g2_decap_8 FILLER_89_245 ();
 sg13g2_decap_8 FILLER_89_252 ();
 sg13g2_decap_8 FILLER_89_259 ();
 sg13g2_decap_8 FILLER_89_266 ();
 sg13g2_decap_8 FILLER_89_273 ();
 sg13g2_decap_8 FILLER_89_280 ();
 sg13g2_decap_8 FILLER_89_287 ();
 sg13g2_decap_8 FILLER_89_294 ();
 sg13g2_decap_8 FILLER_89_301 ();
 sg13g2_decap_8 FILLER_89_308 ();
 sg13g2_decap_8 FILLER_89_315 ();
 sg13g2_decap_8 FILLER_89_322 ();
 sg13g2_decap_8 FILLER_89_329 ();
 sg13g2_decap_8 FILLER_89_336 ();
 sg13g2_decap_8 FILLER_89_343 ();
 sg13g2_decap_8 FILLER_89_350 ();
 sg13g2_decap_8 FILLER_89_357 ();
 sg13g2_decap_8 FILLER_89_364 ();
 sg13g2_decap_8 FILLER_89_371 ();
 sg13g2_decap_8 FILLER_89_378 ();
 sg13g2_decap_8 FILLER_89_385 ();
 sg13g2_decap_8 FILLER_89_392 ();
 sg13g2_decap_8 FILLER_89_399 ();
 sg13g2_decap_8 FILLER_89_406 ();
 sg13g2_decap_8 FILLER_89_413 ();
 sg13g2_decap_8 FILLER_89_420 ();
 sg13g2_decap_8 FILLER_89_427 ();
 sg13g2_decap_8 FILLER_89_434 ();
 sg13g2_decap_8 FILLER_89_441 ();
 sg13g2_decap_8 FILLER_89_448 ();
 sg13g2_decap_8 FILLER_89_455 ();
 sg13g2_decap_8 FILLER_89_462 ();
 sg13g2_decap_8 FILLER_89_469 ();
 sg13g2_decap_8 FILLER_89_476 ();
 sg13g2_decap_8 FILLER_89_483 ();
 sg13g2_decap_8 FILLER_89_490 ();
 sg13g2_decap_8 FILLER_89_497 ();
 sg13g2_decap_8 FILLER_89_504 ();
 sg13g2_decap_8 FILLER_89_511 ();
 sg13g2_decap_8 FILLER_89_518 ();
 sg13g2_decap_8 FILLER_89_525 ();
 sg13g2_decap_8 FILLER_89_532 ();
 sg13g2_decap_8 FILLER_89_539 ();
 sg13g2_decap_8 FILLER_89_546 ();
 sg13g2_decap_8 FILLER_89_553 ();
 sg13g2_decap_8 FILLER_89_560 ();
 sg13g2_decap_8 FILLER_89_567 ();
 sg13g2_decap_8 FILLER_89_574 ();
 sg13g2_decap_8 FILLER_89_581 ();
 sg13g2_decap_8 FILLER_89_588 ();
 sg13g2_decap_8 FILLER_89_595 ();
 sg13g2_decap_8 FILLER_89_602 ();
 sg13g2_decap_8 FILLER_89_609 ();
 sg13g2_decap_8 FILLER_89_616 ();
 sg13g2_decap_8 FILLER_89_623 ();
 sg13g2_decap_8 FILLER_89_630 ();
 sg13g2_decap_8 FILLER_89_637 ();
 sg13g2_decap_8 FILLER_89_644 ();
 sg13g2_decap_8 FILLER_89_651 ();
 sg13g2_decap_8 FILLER_89_658 ();
 sg13g2_decap_8 FILLER_89_665 ();
 sg13g2_decap_8 FILLER_89_672 ();
 sg13g2_decap_8 FILLER_89_679 ();
 sg13g2_decap_8 FILLER_89_686 ();
 sg13g2_decap_8 FILLER_89_693 ();
 sg13g2_decap_8 FILLER_89_700 ();
 sg13g2_decap_8 FILLER_89_707 ();
 sg13g2_decap_8 FILLER_89_714 ();
 sg13g2_decap_8 FILLER_89_721 ();
 sg13g2_decap_8 FILLER_89_728 ();
 sg13g2_decap_8 FILLER_89_735 ();
 sg13g2_decap_8 FILLER_89_742 ();
 sg13g2_decap_8 FILLER_89_749 ();
 sg13g2_decap_8 FILLER_89_756 ();
 sg13g2_decap_8 FILLER_89_763 ();
 sg13g2_decap_8 FILLER_89_770 ();
 sg13g2_decap_8 FILLER_89_777 ();
 sg13g2_decap_8 FILLER_89_784 ();
 sg13g2_decap_8 FILLER_89_791 ();
 sg13g2_decap_8 FILLER_89_798 ();
 sg13g2_decap_8 FILLER_89_805 ();
 sg13g2_decap_8 FILLER_89_812 ();
 sg13g2_decap_8 FILLER_89_819 ();
 sg13g2_decap_8 FILLER_89_826 ();
 sg13g2_decap_8 FILLER_89_833 ();
 sg13g2_decap_8 FILLER_89_840 ();
 sg13g2_decap_8 FILLER_89_847 ();
 sg13g2_decap_8 FILLER_89_854 ();
 sg13g2_decap_8 FILLER_89_861 ();
 sg13g2_decap_8 FILLER_89_868 ();
 sg13g2_decap_8 FILLER_89_875 ();
 sg13g2_decap_8 FILLER_89_882 ();
 sg13g2_decap_8 FILLER_89_889 ();
 sg13g2_decap_8 FILLER_89_896 ();
 sg13g2_decap_8 FILLER_89_903 ();
 sg13g2_decap_8 FILLER_89_910 ();
 sg13g2_decap_8 FILLER_89_917 ();
 sg13g2_decap_8 FILLER_89_924 ();
 sg13g2_decap_8 FILLER_89_931 ();
 sg13g2_decap_8 FILLER_89_938 ();
 sg13g2_decap_8 FILLER_89_945 ();
 sg13g2_decap_8 FILLER_89_952 ();
 sg13g2_decap_8 FILLER_89_959 ();
 sg13g2_decap_8 FILLER_89_966 ();
 sg13g2_decap_8 FILLER_89_973 ();
 sg13g2_decap_8 FILLER_89_980 ();
 sg13g2_decap_8 FILLER_89_987 ();
 sg13g2_decap_8 FILLER_89_994 ();
 sg13g2_decap_8 FILLER_89_1001 ();
 sg13g2_decap_8 FILLER_89_1008 ();
 sg13g2_decap_8 FILLER_89_1015 ();
 sg13g2_decap_8 FILLER_89_1022 ();
 sg13g2_decap_8 FILLER_90_4 ();
 sg13g2_decap_8 FILLER_90_11 ();
 sg13g2_decap_8 FILLER_90_18 ();
 sg13g2_decap_8 FILLER_90_25 ();
 sg13g2_decap_8 FILLER_90_32 ();
 sg13g2_decap_8 FILLER_90_39 ();
 sg13g2_decap_8 FILLER_90_46 ();
 sg13g2_decap_8 FILLER_90_53 ();
 sg13g2_decap_8 FILLER_90_60 ();
 sg13g2_decap_8 FILLER_90_67 ();
 sg13g2_decap_8 FILLER_90_74 ();
 sg13g2_decap_8 FILLER_90_81 ();
 sg13g2_decap_8 FILLER_90_88 ();
 sg13g2_decap_8 FILLER_90_95 ();
 sg13g2_decap_8 FILLER_90_102 ();
 sg13g2_decap_8 FILLER_90_109 ();
 sg13g2_decap_8 FILLER_90_116 ();
 sg13g2_decap_8 FILLER_90_123 ();
 sg13g2_decap_8 FILLER_90_130 ();
 sg13g2_decap_8 FILLER_90_137 ();
 sg13g2_decap_8 FILLER_90_144 ();
 sg13g2_decap_8 FILLER_90_151 ();
 sg13g2_decap_8 FILLER_90_158 ();
 sg13g2_decap_8 FILLER_90_165 ();
 sg13g2_decap_8 FILLER_90_172 ();
 sg13g2_decap_8 FILLER_90_179 ();
 sg13g2_decap_8 FILLER_90_186 ();
 sg13g2_decap_8 FILLER_90_193 ();
 sg13g2_decap_8 FILLER_90_200 ();
 sg13g2_decap_8 FILLER_90_207 ();
 sg13g2_decap_8 FILLER_90_214 ();
 sg13g2_decap_8 FILLER_90_221 ();
 sg13g2_decap_8 FILLER_90_228 ();
 sg13g2_decap_8 FILLER_90_235 ();
 sg13g2_decap_8 FILLER_90_242 ();
 sg13g2_decap_8 FILLER_90_249 ();
 sg13g2_decap_8 FILLER_90_256 ();
 sg13g2_decap_8 FILLER_90_263 ();
 sg13g2_decap_8 FILLER_90_270 ();
 sg13g2_decap_8 FILLER_90_277 ();
 sg13g2_decap_8 FILLER_90_284 ();
 sg13g2_decap_8 FILLER_90_291 ();
 sg13g2_decap_8 FILLER_90_298 ();
 sg13g2_decap_8 FILLER_90_305 ();
 sg13g2_decap_8 FILLER_90_312 ();
 sg13g2_decap_8 FILLER_90_319 ();
 sg13g2_decap_8 FILLER_90_326 ();
 sg13g2_decap_8 FILLER_90_333 ();
 sg13g2_decap_8 FILLER_90_340 ();
 sg13g2_decap_8 FILLER_90_347 ();
 sg13g2_decap_8 FILLER_90_354 ();
 sg13g2_decap_8 FILLER_90_361 ();
 sg13g2_decap_8 FILLER_90_368 ();
 sg13g2_decap_8 FILLER_90_375 ();
 sg13g2_decap_8 FILLER_90_382 ();
 sg13g2_decap_8 FILLER_90_389 ();
 sg13g2_decap_8 FILLER_90_396 ();
 sg13g2_decap_8 FILLER_90_403 ();
 sg13g2_decap_8 FILLER_90_410 ();
 sg13g2_decap_8 FILLER_90_417 ();
 sg13g2_decap_8 FILLER_90_424 ();
 sg13g2_decap_8 FILLER_90_431 ();
 sg13g2_decap_8 FILLER_90_438 ();
 sg13g2_decap_8 FILLER_90_445 ();
 sg13g2_decap_8 FILLER_90_452 ();
 sg13g2_decap_8 FILLER_90_459 ();
 sg13g2_decap_8 FILLER_90_466 ();
 sg13g2_decap_8 FILLER_90_473 ();
 sg13g2_decap_8 FILLER_90_480 ();
 sg13g2_decap_8 FILLER_90_487 ();
 sg13g2_decap_8 FILLER_90_494 ();
 sg13g2_decap_8 FILLER_90_501 ();
 sg13g2_decap_8 FILLER_90_508 ();
 sg13g2_decap_8 FILLER_90_515 ();
 sg13g2_decap_8 FILLER_90_522 ();
 sg13g2_decap_8 FILLER_90_529 ();
 sg13g2_decap_8 FILLER_90_536 ();
 sg13g2_decap_8 FILLER_90_543 ();
 sg13g2_decap_8 FILLER_90_550 ();
 sg13g2_decap_8 FILLER_90_557 ();
 sg13g2_decap_8 FILLER_90_564 ();
 sg13g2_decap_8 FILLER_90_571 ();
 sg13g2_decap_8 FILLER_90_578 ();
 sg13g2_decap_8 FILLER_90_585 ();
 sg13g2_decap_8 FILLER_90_592 ();
 sg13g2_decap_8 FILLER_90_599 ();
 sg13g2_decap_8 FILLER_90_606 ();
 sg13g2_decap_8 FILLER_90_613 ();
 sg13g2_decap_8 FILLER_90_620 ();
 sg13g2_decap_8 FILLER_90_627 ();
 sg13g2_decap_8 FILLER_90_634 ();
 sg13g2_decap_8 FILLER_90_641 ();
 sg13g2_decap_8 FILLER_90_648 ();
 sg13g2_decap_8 FILLER_90_655 ();
 sg13g2_decap_8 FILLER_90_662 ();
 sg13g2_decap_8 FILLER_90_669 ();
 sg13g2_decap_8 FILLER_90_676 ();
 sg13g2_decap_8 FILLER_90_683 ();
 sg13g2_decap_8 FILLER_90_690 ();
 sg13g2_decap_8 FILLER_90_697 ();
 sg13g2_decap_8 FILLER_90_704 ();
 sg13g2_decap_8 FILLER_90_711 ();
 sg13g2_decap_8 FILLER_90_718 ();
 sg13g2_decap_8 FILLER_90_725 ();
 sg13g2_decap_8 FILLER_90_732 ();
 sg13g2_decap_8 FILLER_90_739 ();
 sg13g2_decap_8 FILLER_90_746 ();
 sg13g2_decap_8 FILLER_90_753 ();
 sg13g2_decap_8 FILLER_90_760 ();
 sg13g2_decap_8 FILLER_90_767 ();
 sg13g2_decap_8 FILLER_90_774 ();
 sg13g2_decap_8 FILLER_90_781 ();
 sg13g2_decap_8 FILLER_90_788 ();
 sg13g2_decap_8 FILLER_90_795 ();
 sg13g2_decap_8 FILLER_90_802 ();
 sg13g2_decap_8 FILLER_90_809 ();
 sg13g2_decap_8 FILLER_90_816 ();
 sg13g2_decap_8 FILLER_90_823 ();
 sg13g2_decap_8 FILLER_90_830 ();
 sg13g2_decap_8 FILLER_90_837 ();
 sg13g2_decap_8 FILLER_90_844 ();
 sg13g2_decap_8 FILLER_90_851 ();
 sg13g2_decap_8 FILLER_90_858 ();
 sg13g2_decap_8 FILLER_90_865 ();
 sg13g2_decap_8 FILLER_90_872 ();
 sg13g2_decap_8 FILLER_90_879 ();
 sg13g2_decap_8 FILLER_90_886 ();
 sg13g2_decap_8 FILLER_90_893 ();
 sg13g2_decap_8 FILLER_90_900 ();
 sg13g2_decap_8 FILLER_90_907 ();
 sg13g2_decap_8 FILLER_90_914 ();
 sg13g2_decap_8 FILLER_90_921 ();
 sg13g2_decap_8 FILLER_90_928 ();
 sg13g2_decap_8 FILLER_90_935 ();
 sg13g2_decap_8 FILLER_90_942 ();
 sg13g2_decap_8 FILLER_90_949 ();
 sg13g2_decap_8 FILLER_90_956 ();
 sg13g2_decap_8 FILLER_90_963 ();
 sg13g2_decap_8 FILLER_90_970 ();
 sg13g2_decap_8 FILLER_90_977 ();
 sg13g2_decap_8 FILLER_90_984 ();
 sg13g2_decap_8 FILLER_90_991 ();
 sg13g2_decap_8 FILLER_90_998 ();
 sg13g2_decap_8 FILLER_90_1005 ();
 sg13g2_decap_8 FILLER_90_1012 ();
 sg13g2_decap_8 FILLER_90_1019 ();
 sg13g2_fill_2 FILLER_90_1026 ();
 sg13g2_fill_1 FILLER_90_1028 ();
 sg13g2_decap_8 FILLER_91_0 ();
 sg13g2_decap_8 FILLER_91_7 ();
 sg13g2_decap_8 FILLER_91_14 ();
 sg13g2_decap_8 FILLER_91_21 ();
 sg13g2_decap_8 FILLER_91_28 ();
 sg13g2_decap_8 FILLER_91_35 ();
 sg13g2_decap_8 FILLER_91_42 ();
 sg13g2_decap_8 FILLER_91_49 ();
 sg13g2_decap_8 FILLER_91_56 ();
 sg13g2_decap_8 FILLER_91_63 ();
 sg13g2_decap_8 FILLER_91_70 ();
 sg13g2_decap_8 FILLER_91_77 ();
 sg13g2_decap_8 FILLER_91_84 ();
 sg13g2_decap_8 FILLER_91_91 ();
 sg13g2_decap_8 FILLER_91_98 ();
 sg13g2_decap_8 FILLER_91_105 ();
 sg13g2_decap_8 FILLER_91_112 ();
 sg13g2_decap_8 FILLER_91_119 ();
 sg13g2_decap_8 FILLER_91_126 ();
 sg13g2_decap_8 FILLER_91_133 ();
 sg13g2_decap_8 FILLER_91_140 ();
 sg13g2_decap_8 FILLER_91_147 ();
 sg13g2_decap_8 FILLER_91_154 ();
 sg13g2_decap_8 FILLER_91_161 ();
 sg13g2_decap_8 FILLER_91_168 ();
 sg13g2_decap_8 FILLER_91_175 ();
 sg13g2_decap_8 FILLER_91_182 ();
 sg13g2_decap_8 FILLER_91_189 ();
 sg13g2_decap_8 FILLER_91_196 ();
 sg13g2_decap_8 FILLER_91_203 ();
 sg13g2_decap_8 FILLER_91_210 ();
 sg13g2_decap_8 FILLER_91_217 ();
 sg13g2_decap_8 FILLER_91_224 ();
 sg13g2_decap_8 FILLER_91_231 ();
 sg13g2_decap_8 FILLER_91_238 ();
 sg13g2_decap_8 FILLER_91_245 ();
 sg13g2_decap_8 FILLER_91_252 ();
 sg13g2_decap_8 FILLER_91_259 ();
 sg13g2_decap_8 FILLER_91_266 ();
 sg13g2_decap_8 FILLER_91_273 ();
 sg13g2_decap_8 FILLER_91_280 ();
 sg13g2_decap_8 FILLER_91_287 ();
 sg13g2_decap_8 FILLER_91_294 ();
 sg13g2_decap_8 FILLER_91_301 ();
 sg13g2_decap_8 FILLER_91_308 ();
 sg13g2_decap_8 FILLER_91_315 ();
 sg13g2_decap_8 FILLER_91_322 ();
 sg13g2_decap_8 FILLER_91_329 ();
 sg13g2_decap_8 FILLER_91_336 ();
 sg13g2_decap_8 FILLER_91_343 ();
 sg13g2_decap_8 FILLER_91_350 ();
 sg13g2_decap_8 FILLER_91_357 ();
 sg13g2_decap_8 FILLER_91_364 ();
 sg13g2_decap_8 FILLER_91_371 ();
 sg13g2_decap_8 FILLER_91_378 ();
 sg13g2_decap_8 FILLER_91_385 ();
 sg13g2_decap_8 FILLER_91_392 ();
 sg13g2_decap_8 FILLER_91_399 ();
 sg13g2_decap_8 FILLER_91_406 ();
 sg13g2_decap_8 FILLER_91_413 ();
 sg13g2_decap_8 FILLER_91_420 ();
 sg13g2_decap_8 FILLER_91_427 ();
 sg13g2_decap_8 FILLER_91_434 ();
 sg13g2_decap_8 FILLER_91_441 ();
 sg13g2_decap_8 FILLER_91_448 ();
 sg13g2_decap_8 FILLER_91_455 ();
 sg13g2_decap_8 FILLER_91_462 ();
 sg13g2_decap_8 FILLER_91_469 ();
 sg13g2_decap_8 FILLER_91_476 ();
 sg13g2_decap_8 FILLER_91_483 ();
 sg13g2_decap_8 FILLER_91_490 ();
 sg13g2_decap_8 FILLER_91_497 ();
 sg13g2_decap_8 FILLER_91_504 ();
 sg13g2_decap_8 FILLER_91_511 ();
 sg13g2_decap_8 FILLER_91_518 ();
 sg13g2_decap_8 FILLER_91_525 ();
 sg13g2_decap_8 FILLER_91_532 ();
 sg13g2_decap_8 FILLER_91_539 ();
 sg13g2_decap_8 FILLER_91_546 ();
 sg13g2_decap_8 FILLER_91_553 ();
 sg13g2_decap_8 FILLER_91_560 ();
 sg13g2_decap_8 FILLER_91_567 ();
 sg13g2_decap_8 FILLER_91_574 ();
 sg13g2_decap_8 FILLER_91_581 ();
 sg13g2_decap_8 FILLER_91_588 ();
 sg13g2_decap_8 FILLER_91_595 ();
 sg13g2_decap_8 FILLER_91_602 ();
 sg13g2_decap_8 FILLER_91_609 ();
 sg13g2_decap_8 FILLER_91_616 ();
 sg13g2_decap_8 FILLER_91_623 ();
 sg13g2_decap_8 FILLER_91_630 ();
 sg13g2_decap_8 FILLER_91_637 ();
 sg13g2_decap_8 FILLER_91_644 ();
 sg13g2_decap_8 FILLER_91_651 ();
 sg13g2_decap_8 FILLER_91_658 ();
 sg13g2_decap_8 FILLER_91_665 ();
 sg13g2_decap_8 FILLER_91_672 ();
 sg13g2_decap_8 FILLER_91_679 ();
 sg13g2_decap_8 FILLER_91_686 ();
 sg13g2_decap_8 FILLER_91_693 ();
 sg13g2_decap_8 FILLER_91_700 ();
 sg13g2_decap_8 FILLER_91_707 ();
 sg13g2_decap_8 FILLER_91_714 ();
 sg13g2_decap_8 FILLER_91_721 ();
 sg13g2_decap_8 FILLER_91_728 ();
 sg13g2_decap_8 FILLER_91_735 ();
 sg13g2_decap_8 FILLER_91_742 ();
 sg13g2_decap_8 FILLER_91_749 ();
 sg13g2_decap_8 FILLER_91_756 ();
 sg13g2_decap_8 FILLER_91_763 ();
 sg13g2_decap_8 FILLER_91_770 ();
 sg13g2_decap_8 FILLER_91_777 ();
 sg13g2_decap_8 FILLER_91_784 ();
 sg13g2_decap_8 FILLER_91_791 ();
 sg13g2_decap_8 FILLER_91_798 ();
 sg13g2_decap_8 FILLER_91_805 ();
 sg13g2_decap_8 FILLER_91_812 ();
 sg13g2_decap_8 FILLER_91_819 ();
 sg13g2_decap_8 FILLER_91_826 ();
 sg13g2_decap_8 FILLER_91_833 ();
 sg13g2_decap_8 FILLER_91_840 ();
 sg13g2_decap_8 FILLER_91_847 ();
 sg13g2_decap_8 FILLER_91_854 ();
 sg13g2_decap_8 FILLER_91_861 ();
 sg13g2_decap_8 FILLER_91_868 ();
 sg13g2_decap_8 FILLER_91_875 ();
 sg13g2_decap_8 FILLER_91_882 ();
 sg13g2_decap_8 FILLER_91_889 ();
 sg13g2_decap_8 FILLER_91_896 ();
 sg13g2_decap_8 FILLER_91_903 ();
 sg13g2_decap_8 FILLER_91_910 ();
 sg13g2_decap_8 FILLER_91_917 ();
 sg13g2_decap_8 FILLER_91_924 ();
 sg13g2_decap_8 FILLER_91_931 ();
 sg13g2_decap_8 FILLER_91_938 ();
 sg13g2_decap_8 FILLER_91_945 ();
 sg13g2_decap_8 FILLER_91_952 ();
 sg13g2_decap_8 FILLER_91_959 ();
 sg13g2_decap_8 FILLER_91_966 ();
 sg13g2_decap_8 FILLER_91_973 ();
 sg13g2_decap_8 FILLER_91_980 ();
 sg13g2_decap_8 FILLER_91_987 ();
 sg13g2_decap_8 FILLER_91_994 ();
 sg13g2_decap_8 FILLER_91_1001 ();
 sg13g2_decap_8 FILLER_91_1008 ();
 sg13g2_decap_8 FILLER_91_1015 ();
 sg13g2_decap_8 FILLER_91_1022 ();
 sg13g2_decap_8 FILLER_92_0 ();
 sg13g2_decap_8 FILLER_92_7 ();
 sg13g2_decap_8 FILLER_92_14 ();
 sg13g2_decap_8 FILLER_92_21 ();
 sg13g2_decap_8 FILLER_92_28 ();
 sg13g2_decap_8 FILLER_92_35 ();
 sg13g2_decap_8 FILLER_92_42 ();
 sg13g2_decap_8 FILLER_92_49 ();
 sg13g2_decap_8 FILLER_92_56 ();
 sg13g2_decap_8 FILLER_92_63 ();
 sg13g2_decap_8 FILLER_92_70 ();
 sg13g2_decap_8 FILLER_92_77 ();
 sg13g2_decap_8 FILLER_92_84 ();
 sg13g2_decap_8 FILLER_92_91 ();
 sg13g2_decap_8 FILLER_92_98 ();
 sg13g2_decap_8 FILLER_92_105 ();
 sg13g2_decap_8 FILLER_92_112 ();
 sg13g2_decap_8 FILLER_92_119 ();
 sg13g2_decap_8 FILLER_92_126 ();
 sg13g2_decap_8 FILLER_92_133 ();
 sg13g2_decap_8 FILLER_92_140 ();
 sg13g2_decap_8 FILLER_92_147 ();
 sg13g2_decap_8 FILLER_92_154 ();
 sg13g2_decap_8 FILLER_92_161 ();
 sg13g2_decap_8 FILLER_92_168 ();
 sg13g2_decap_8 FILLER_92_175 ();
 sg13g2_decap_8 FILLER_92_182 ();
 sg13g2_decap_8 FILLER_92_189 ();
 sg13g2_decap_8 FILLER_92_196 ();
 sg13g2_decap_8 FILLER_92_203 ();
 sg13g2_decap_8 FILLER_92_210 ();
 sg13g2_decap_8 FILLER_92_217 ();
 sg13g2_decap_8 FILLER_92_224 ();
 sg13g2_decap_8 FILLER_92_231 ();
 sg13g2_decap_8 FILLER_92_238 ();
 sg13g2_decap_8 FILLER_92_245 ();
 sg13g2_decap_8 FILLER_92_252 ();
 sg13g2_decap_8 FILLER_92_259 ();
 sg13g2_decap_8 FILLER_92_266 ();
 sg13g2_decap_8 FILLER_92_273 ();
 sg13g2_decap_8 FILLER_92_280 ();
 sg13g2_decap_8 FILLER_92_287 ();
 sg13g2_decap_8 FILLER_92_294 ();
 sg13g2_decap_8 FILLER_92_301 ();
 sg13g2_decap_8 FILLER_92_308 ();
 sg13g2_decap_8 FILLER_92_315 ();
 sg13g2_decap_8 FILLER_92_322 ();
 sg13g2_decap_8 FILLER_92_329 ();
 sg13g2_decap_8 FILLER_92_336 ();
 sg13g2_decap_8 FILLER_92_343 ();
 sg13g2_decap_8 FILLER_92_350 ();
 sg13g2_decap_8 FILLER_92_357 ();
 sg13g2_decap_8 FILLER_92_364 ();
 sg13g2_decap_8 FILLER_92_371 ();
 sg13g2_decap_8 FILLER_92_378 ();
 sg13g2_decap_8 FILLER_92_385 ();
 sg13g2_decap_8 FILLER_92_392 ();
 sg13g2_decap_8 FILLER_92_399 ();
 sg13g2_decap_8 FILLER_92_406 ();
 sg13g2_decap_8 FILLER_92_413 ();
 sg13g2_decap_8 FILLER_92_420 ();
 sg13g2_decap_8 FILLER_92_427 ();
 sg13g2_decap_8 FILLER_92_434 ();
 sg13g2_decap_8 FILLER_92_441 ();
 sg13g2_decap_8 FILLER_92_448 ();
 sg13g2_decap_8 FILLER_92_455 ();
 sg13g2_decap_8 FILLER_92_462 ();
 sg13g2_decap_8 FILLER_92_469 ();
 sg13g2_decap_8 FILLER_92_476 ();
 sg13g2_decap_8 FILLER_92_483 ();
 sg13g2_decap_8 FILLER_92_490 ();
 sg13g2_decap_8 FILLER_92_497 ();
 sg13g2_decap_8 FILLER_92_504 ();
 sg13g2_decap_8 FILLER_92_511 ();
 sg13g2_decap_8 FILLER_92_518 ();
 sg13g2_decap_8 FILLER_92_525 ();
 sg13g2_decap_8 FILLER_92_532 ();
 sg13g2_decap_8 FILLER_92_539 ();
 sg13g2_decap_8 FILLER_92_546 ();
 sg13g2_decap_8 FILLER_92_553 ();
 sg13g2_decap_8 FILLER_92_560 ();
 sg13g2_decap_8 FILLER_92_567 ();
 sg13g2_decap_8 FILLER_92_574 ();
 sg13g2_decap_8 FILLER_92_581 ();
 sg13g2_decap_8 FILLER_92_588 ();
 sg13g2_decap_8 FILLER_92_595 ();
 sg13g2_decap_8 FILLER_92_602 ();
 sg13g2_decap_8 FILLER_92_609 ();
 sg13g2_decap_8 FILLER_92_616 ();
 sg13g2_decap_8 FILLER_92_623 ();
 sg13g2_decap_8 FILLER_92_630 ();
 sg13g2_decap_8 FILLER_92_637 ();
 sg13g2_decap_8 FILLER_92_644 ();
 sg13g2_decap_8 FILLER_92_651 ();
 sg13g2_decap_8 FILLER_92_658 ();
 sg13g2_decap_8 FILLER_92_665 ();
 sg13g2_decap_8 FILLER_92_672 ();
 sg13g2_decap_8 FILLER_92_679 ();
 sg13g2_decap_8 FILLER_92_686 ();
 sg13g2_decap_8 FILLER_92_693 ();
 sg13g2_decap_8 FILLER_92_700 ();
 sg13g2_decap_8 FILLER_92_707 ();
 sg13g2_decap_8 FILLER_92_714 ();
 sg13g2_decap_8 FILLER_92_721 ();
 sg13g2_decap_8 FILLER_92_728 ();
 sg13g2_decap_8 FILLER_92_735 ();
 sg13g2_decap_8 FILLER_92_742 ();
 sg13g2_decap_8 FILLER_92_749 ();
 sg13g2_decap_8 FILLER_92_756 ();
 sg13g2_decap_8 FILLER_92_763 ();
 sg13g2_decap_8 FILLER_92_770 ();
 sg13g2_decap_8 FILLER_92_777 ();
 sg13g2_decap_8 FILLER_92_784 ();
 sg13g2_decap_8 FILLER_92_791 ();
 sg13g2_decap_8 FILLER_92_798 ();
 sg13g2_decap_8 FILLER_92_805 ();
 sg13g2_decap_8 FILLER_92_812 ();
 sg13g2_decap_8 FILLER_92_819 ();
 sg13g2_decap_8 FILLER_92_826 ();
 sg13g2_decap_8 FILLER_92_833 ();
 sg13g2_decap_8 FILLER_92_840 ();
 sg13g2_decap_8 FILLER_92_847 ();
 sg13g2_decap_8 FILLER_92_854 ();
 sg13g2_decap_8 FILLER_92_861 ();
 sg13g2_decap_8 FILLER_92_868 ();
 sg13g2_decap_8 FILLER_92_875 ();
 sg13g2_decap_8 FILLER_92_882 ();
 sg13g2_decap_8 FILLER_92_889 ();
 sg13g2_decap_8 FILLER_92_896 ();
 sg13g2_decap_8 FILLER_92_903 ();
 sg13g2_decap_8 FILLER_92_910 ();
 sg13g2_decap_8 FILLER_92_917 ();
 sg13g2_decap_8 FILLER_92_924 ();
 sg13g2_decap_8 FILLER_92_931 ();
 sg13g2_decap_8 FILLER_92_938 ();
 sg13g2_decap_8 FILLER_92_945 ();
 sg13g2_decap_8 FILLER_92_952 ();
 sg13g2_decap_8 FILLER_92_959 ();
 sg13g2_decap_8 FILLER_92_966 ();
 sg13g2_decap_8 FILLER_92_973 ();
 sg13g2_decap_8 FILLER_92_980 ();
 sg13g2_decap_8 FILLER_92_987 ();
 sg13g2_decap_8 FILLER_92_994 ();
 sg13g2_decap_8 FILLER_92_1001 ();
 sg13g2_decap_8 FILLER_92_1008 ();
 sg13g2_decap_8 FILLER_92_1015 ();
 sg13g2_decap_8 FILLER_92_1022 ();
 sg13g2_decap_8 FILLER_93_5 ();
 sg13g2_decap_8 FILLER_93_12 ();
 sg13g2_decap_8 FILLER_93_19 ();
 sg13g2_decap_8 FILLER_93_26 ();
 sg13g2_decap_8 FILLER_93_33 ();
 sg13g2_decap_8 FILLER_93_40 ();
 sg13g2_decap_8 FILLER_93_47 ();
 sg13g2_decap_8 FILLER_93_54 ();
 sg13g2_decap_8 FILLER_93_61 ();
 sg13g2_decap_8 FILLER_93_68 ();
 sg13g2_decap_8 FILLER_93_75 ();
 sg13g2_decap_8 FILLER_93_82 ();
 sg13g2_decap_8 FILLER_93_89 ();
 sg13g2_decap_8 FILLER_93_96 ();
 sg13g2_decap_8 FILLER_93_103 ();
 sg13g2_decap_8 FILLER_93_110 ();
 sg13g2_decap_8 FILLER_93_117 ();
 sg13g2_decap_8 FILLER_93_124 ();
 sg13g2_decap_8 FILLER_93_131 ();
 sg13g2_decap_8 FILLER_93_138 ();
 sg13g2_decap_8 FILLER_93_145 ();
 sg13g2_decap_8 FILLER_93_152 ();
 sg13g2_decap_8 FILLER_93_159 ();
 sg13g2_decap_8 FILLER_93_166 ();
 sg13g2_decap_8 FILLER_93_173 ();
 sg13g2_decap_8 FILLER_93_180 ();
 sg13g2_decap_8 FILLER_93_187 ();
 sg13g2_decap_8 FILLER_93_194 ();
 sg13g2_decap_8 FILLER_93_201 ();
 sg13g2_decap_8 FILLER_93_208 ();
 sg13g2_decap_8 FILLER_93_215 ();
 sg13g2_decap_8 FILLER_93_222 ();
 sg13g2_decap_8 FILLER_93_229 ();
 sg13g2_decap_8 FILLER_93_236 ();
 sg13g2_decap_8 FILLER_93_243 ();
 sg13g2_decap_8 FILLER_93_250 ();
 sg13g2_decap_8 FILLER_93_257 ();
 sg13g2_decap_8 FILLER_93_264 ();
 sg13g2_decap_8 FILLER_93_271 ();
 sg13g2_decap_8 FILLER_93_278 ();
 sg13g2_decap_8 FILLER_93_285 ();
 sg13g2_decap_8 FILLER_93_292 ();
 sg13g2_decap_8 FILLER_93_299 ();
 sg13g2_decap_8 FILLER_93_306 ();
 sg13g2_decap_8 FILLER_93_313 ();
 sg13g2_decap_8 FILLER_93_320 ();
 sg13g2_decap_8 FILLER_93_327 ();
 sg13g2_decap_8 FILLER_93_334 ();
 sg13g2_decap_8 FILLER_93_341 ();
 sg13g2_decap_8 FILLER_93_348 ();
 sg13g2_decap_8 FILLER_93_355 ();
 sg13g2_decap_8 FILLER_93_362 ();
 sg13g2_decap_8 FILLER_93_369 ();
 sg13g2_decap_8 FILLER_93_376 ();
 sg13g2_decap_8 FILLER_93_383 ();
 sg13g2_decap_8 FILLER_93_390 ();
 sg13g2_decap_8 FILLER_93_397 ();
 sg13g2_decap_8 FILLER_93_404 ();
 sg13g2_decap_8 FILLER_93_411 ();
 sg13g2_decap_8 FILLER_93_418 ();
 sg13g2_decap_8 FILLER_93_425 ();
 sg13g2_decap_8 FILLER_93_432 ();
 sg13g2_decap_8 FILLER_93_439 ();
 sg13g2_decap_8 FILLER_93_446 ();
 sg13g2_decap_8 FILLER_93_453 ();
 sg13g2_decap_8 FILLER_93_460 ();
 sg13g2_decap_8 FILLER_93_467 ();
 sg13g2_decap_8 FILLER_93_474 ();
 sg13g2_decap_8 FILLER_93_481 ();
 sg13g2_decap_8 FILLER_93_488 ();
 sg13g2_decap_8 FILLER_93_495 ();
 sg13g2_decap_8 FILLER_93_502 ();
 sg13g2_decap_8 FILLER_93_509 ();
 sg13g2_decap_8 FILLER_93_516 ();
 sg13g2_decap_8 FILLER_93_523 ();
 sg13g2_decap_8 FILLER_93_530 ();
 sg13g2_decap_8 FILLER_93_537 ();
 sg13g2_decap_8 FILLER_93_544 ();
 sg13g2_decap_8 FILLER_93_551 ();
 sg13g2_decap_8 FILLER_93_558 ();
 sg13g2_decap_8 FILLER_93_565 ();
 sg13g2_decap_8 FILLER_93_572 ();
 sg13g2_decap_8 FILLER_93_579 ();
 sg13g2_decap_8 FILLER_93_586 ();
 sg13g2_decap_8 FILLER_93_593 ();
 sg13g2_decap_8 FILLER_93_600 ();
 sg13g2_decap_8 FILLER_93_607 ();
 sg13g2_decap_8 FILLER_93_614 ();
 sg13g2_decap_8 FILLER_93_621 ();
 sg13g2_decap_8 FILLER_93_628 ();
 sg13g2_decap_8 FILLER_93_635 ();
 sg13g2_decap_8 FILLER_93_642 ();
 sg13g2_decap_8 FILLER_93_649 ();
 sg13g2_decap_8 FILLER_93_656 ();
 sg13g2_decap_8 FILLER_93_663 ();
 sg13g2_decap_8 FILLER_93_670 ();
 sg13g2_decap_8 FILLER_93_677 ();
 sg13g2_decap_8 FILLER_93_684 ();
 sg13g2_decap_8 FILLER_93_691 ();
 sg13g2_decap_8 FILLER_93_698 ();
 sg13g2_decap_8 FILLER_93_705 ();
 sg13g2_decap_8 FILLER_93_712 ();
 sg13g2_decap_8 FILLER_93_719 ();
 sg13g2_decap_8 FILLER_93_726 ();
 sg13g2_decap_8 FILLER_93_733 ();
 sg13g2_decap_8 FILLER_93_740 ();
 sg13g2_decap_8 FILLER_93_747 ();
 sg13g2_decap_8 FILLER_93_754 ();
 sg13g2_decap_8 FILLER_93_761 ();
 sg13g2_decap_8 FILLER_93_768 ();
 sg13g2_decap_8 FILLER_93_775 ();
 sg13g2_decap_8 FILLER_93_782 ();
 sg13g2_decap_8 FILLER_93_789 ();
 sg13g2_decap_8 FILLER_93_796 ();
 sg13g2_decap_8 FILLER_93_803 ();
 sg13g2_decap_8 FILLER_93_810 ();
 sg13g2_decap_8 FILLER_93_817 ();
 sg13g2_decap_8 FILLER_93_824 ();
 sg13g2_decap_8 FILLER_93_831 ();
 sg13g2_decap_8 FILLER_93_838 ();
 sg13g2_decap_8 FILLER_93_845 ();
 sg13g2_decap_8 FILLER_93_852 ();
 sg13g2_decap_8 FILLER_93_859 ();
 sg13g2_decap_8 FILLER_93_866 ();
 sg13g2_decap_8 FILLER_93_873 ();
 sg13g2_decap_8 FILLER_93_880 ();
 sg13g2_decap_8 FILLER_93_887 ();
 sg13g2_decap_8 FILLER_93_894 ();
 sg13g2_decap_8 FILLER_93_901 ();
 sg13g2_decap_8 FILLER_93_908 ();
 sg13g2_decap_8 FILLER_93_915 ();
 sg13g2_decap_8 FILLER_93_922 ();
 sg13g2_decap_8 FILLER_93_929 ();
 sg13g2_decap_8 FILLER_93_936 ();
 sg13g2_decap_8 FILLER_93_943 ();
 sg13g2_decap_8 FILLER_93_950 ();
 sg13g2_decap_8 FILLER_93_957 ();
 sg13g2_decap_8 FILLER_93_964 ();
 sg13g2_decap_8 FILLER_93_971 ();
 sg13g2_decap_8 FILLER_93_978 ();
 sg13g2_decap_8 FILLER_93_985 ();
 sg13g2_decap_8 FILLER_93_992 ();
 sg13g2_decap_8 FILLER_93_999 ();
 sg13g2_decap_8 FILLER_93_1006 ();
 sg13g2_decap_8 FILLER_93_1013 ();
 sg13g2_decap_8 FILLER_93_1020 ();
 sg13g2_fill_2 FILLER_93_1027 ();
 sg13g2_decap_8 FILLER_94_0 ();
 sg13g2_decap_8 FILLER_94_7 ();
 sg13g2_decap_8 FILLER_94_14 ();
 sg13g2_decap_8 FILLER_94_21 ();
 sg13g2_decap_8 FILLER_94_28 ();
 sg13g2_decap_8 FILLER_94_35 ();
 sg13g2_decap_8 FILLER_94_42 ();
 sg13g2_decap_8 FILLER_94_49 ();
 sg13g2_decap_8 FILLER_94_56 ();
 sg13g2_decap_8 FILLER_94_63 ();
 sg13g2_decap_8 FILLER_94_70 ();
 sg13g2_decap_8 FILLER_94_77 ();
 sg13g2_decap_8 FILLER_94_84 ();
 sg13g2_decap_8 FILLER_94_91 ();
 sg13g2_decap_8 FILLER_94_98 ();
 sg13g2_decap_8 FILLER_94_105 ();
 sg13g2_decap_8 FILLER_94_112 ();
 sg13g2_decap_8 FILLER_94_119 ();
 sg13g2_decap_8 FILLER_94_126 ();
 sg13g2_decap_8 FILLER_94_133 ();
 sg13g2_decap_8 FILLER_94_140 ();
 sg13g2_decap_8 FILLER_94_147 ();
 sg13g2_decap_8 FILLER_94_154 ();
 sg13g2_decap_8 FILLER_94_161 ();
 sg13g2_decap_8 FILLER_94_168 ();
 sg13g2_decap_8 FILLER_94_175 ();
 sg13g2_decap_8 FILLER_94_182 ();
 sg13g2_decap_8 FILLER_94_189 ();
 sg13g2_decap_8 FILLER_94_196 ();
 sg13g2_decap_8 FILLER_94_203 ();
 sg13g2_decap_8 FILLER_94_210 ();
 sg13g2_decap_8 FILLER_94_217 ();
 sg13g2_decap_8 FILLER_94_224 ();
 sg13g2_decap_8 FILLER_94_231 ();
 sg13g2_decap_8 FILLER_94_238 ();
 sg13g2_decap_8 FILLER_94_245 ();
 sg13g2_decap_8 FILLER_94_252 ();
 sg13g2_decap_8 FILLER_94_259 ();
 sg13g2_decap_8 FILLER_94_266 ();
 sg13g2_decap_8 FILLER_94_273 ();
 sg13g2_decap_8 FILLER_94_280 ();
 sg13g2_decap_8 FILLER_94_287 ();
 sg13g2_decap_8 FILLER_94_294 ();
 sg13g2_decap_8 FILLER_94_301 ();
 sg13g2_decap_8 FILLER_94_308 ();
 sg13g2_decap_8 FILLER_94_315 ();
 sg13g2_decap_8 FILLER_94_322 ();
 sg13g2_decap_8 FILLER_94_329 ();
 sg13g2_decap_8 FILLER_94_336 ();
 sg13g2_decap_8 FILLER_94_343 ();
 sg13g2_decap_8 FILLER_94_350 ();
 sg13g2_decap_8 FILLER_94_357 ();
 sg13g2_decap_8 FILLER_94_364 ();
 sg13g2_decap_8 FILLER_94_371 ();
 sg13g2_decap_8 FILLER_94_378 ();
 sg13g2_decap_8 FILLER_94_385 ();
 sg13g2_decap_8 FILLER_94_392 ();
 sg13g2_decap_8 FILLER_94_399 ();
 sg13g2_decap_8 FILLER_94_406 ();
 sg13g2_decap_8 FILLER_94_413 ();
 sg13g2_decap_8 FILLER_94_420 ();
 sg13g2_decap_8 FILLER_94_427 ();
 sg13g2_decap_8 FILLER_94_434 ();
 sg13g2_decap_8 FILLER_94_441 ();
 sg13g2_decap_8 FILLER_94_448 ();
 sg13g2_decap_8 FILLER_94_455 ();
 sg13g2_decap_8 FILLER_94_462 ();
 sg13g2_decap_8 FILLER_94_469 ();
 sg13g2_decap_8 FILLER_94_476 ();
 sg13g2_decap_8 FILLER_94_483 ();
 sg13g2_decap_8 FILLER_94_490 ();
 sg13g2_decap_8 FILLER_94_497 ();
 sg13g2_decap_8 FILLER_94_504 ();
 sg13g2_decap_8 FILLER_94_511 ();
 sg13g2_decap_8 FILLER_94_518 ();
 sg13g2_decap_8 FILLER_94_525 ();
 sg13g2_decap_8 FILLER_94_532 ();
 sg13g2_decap_8 FILLER_94_539 ();
 sg13g2_decap_8 FILLER_94_546 ();
 sg13g2_decap_8 FILLER_94_553 ();
 sg13g2_decap_8 FILLER_94_560 ();
 sg13g2_decap_8 FILLER_94_567 ();
 sg13g2_decap_8 FILLER_94_574 ();
 sg13g2_decap_8 FILLER_94_581 ();
 sg13g2_decap_8 FILLER_94_588 ();
 sg13g2_decap_8 FILLER_94_595 ();
 sg13g2_decap_8 FILLER_94_602 ();
 sg13g2_decap_8 FILLER_94_609 ();
 sg13g2_decap_8 FILLER_94_616 ();
 sg13g2_decap_8 FILLER_94_623 ();
 sg13g2_decap_8 FILLER_94_630 ();
 sg13g2_decap_8 FILLER_94_637 ();
 sg13g2_decap_8 FILLER_94_644 ();
 sg13g2_decap_8 FILLER_94_651 ();
 sg13g2_decap_8 FILLER_94_658 ();
 sg13g2_decap_8 FILLER_94_665 ();
 sg13g2_decap_8 FILLER_94_672 ();
 sg13g2_decap_8 FILLER_94_679 ();
 sg13g2_decap_8 FILLER_94_686 ();
 sg13g2_decap_8 FILLER_94_693 ();
 sg13g2_decap_8 FILLER_94_700 ();
 sg13g2_decap_8 FILLER_94_707 ();
 sg13g2_decap_8 FILLER_94_714 ();
 sg13g2_decap_8 FILLER_94_721 ();
 sg13g2_decap_8 FILLER_94_728 ();
 sg13g2_decap_8 FILLER_94_735 ();
 sg13g2_decap_8 FILLER_94_742 ();
 sg13g2_decap_8 FILLER_94_749 ();
 sg13g2_decap_8 FILLER_94_756 ();
 sg13g2_decap_8 FILLER_94_763 ();
 sg13g2_decap_8 FILLER_94_770 ();
 sg13g2_decap_8 FILLER_94_777 ();
 sg13g2_decap_8 FILLER_94_784 ();
 sg13g2_decap_8 FILLER_94_791 ();
 sg13g2_decap_8 FILLER_94_798 ();
 sg13g2_decap_8 FILLER_94_805 ();
 sg13g2_decap_8 FILLER_94_812 ();
 sg13g2_decap_8 FILLER_94_819 ();
 sg13g2_decap_8 FILLER_94_826 ();
 sg13g2_decap_8 FILLER_94_833 ();
 sg13g2_decap_8 FILLER_94_840 ();
 sg13g2_decap_8 FILLER_94_847 ();
 sg13g2_decap_8 FILLER_94_854 ();
 sg13g2_decap_8 FILLER_94_861 ();
 sg13g2_decap_8 FILLER_94_868 ();
 sg13g2_decap_8 FILLER_94_875 ();
 sg13g2_decap_8 FILLER_94_882 ();
 sg13g2_decap_8 FILLER_94_889 ();
 sg13g2_decap_8 FILLER_94_896 ();
 sg13g2_decap_8 FILLER_94_903 ();
 sg13g2_decap_8 FILLER_94_910 ();
 sg13g2_decap_8 FILLER_94_917 ();
 sg13g2_decap_8 FILLER_94_924 ();
 sg13g2_decap_8 FILLER_94_931 ();
 sg13g2_decap_8 FILLER_94_938 ();
 sg13g2_decap_8 FILLER_94_945 ();
 sg13g2_decap_8 FILLER_94_952 ();
 sg13g2_decap_8 FILLER_94_959 ();
 sg13g2_decap_8 FILLER_94_966 ();
 sg13g2_decap_8 FILLER_94_973 ();
 sg13g2_decap_8 FILLER_94_980 ();
 sg13g2_decap_8 FILLER_94_987 ();
 sg13g2_decap_8 FILLER_94_994 ();
 sg13g2_decap_8 FILLER_94_1001 ();
 sg13g2_decap_8 FILLER_94_1008 ();
 sg13g2_decap_8 FILLER_94_1015 ();
 sg13g2_decap_8 FILLER_94_1022 ();
 sg13g2_decap_8 FILLER_95_4 ();
 sg13g2_decap_8 FILLER_95_11 ();
 sg13g2_decap_8 FILLER_95_18 ();
 sg13g2_decap_8 FILLER_95_25 ();
 sg13g2_decap_8 FILLER_95_32 ();
 sg13g2_decap_8 FILLER_95_39 ();
 sg13g2_decap_8 FILLER_95_46 ();
 sg13g2_decap_8 FILLER_95_53 ();
 sg13g2_decap_8 FILLER_95_60 ();
 sg13g2_decap_8 FILLER_95_67 ();
 sg13g2_decap_8 FILLER_95_74 ();
 sg13g2_decap_8 FILLER_95_81 ();
 sg13g2_decap_8 FILLER_95_88 ();
 sg13g2_decap_8 FILLER_95_95 ();
 sg13g2_decap_8 FILLER_95_102 ();
 sg13g2_decap_8 FILLER_95_109 ();
 sg13g2_decap_8 FILLER_95_116 ();
 sg13g2_decap_8 FILLER_95_123 ();
 sg13g2_decap_8 FILLER_95_130 ();
 sg13g2_decap_8 FILLER_95_137 ();
 sg13g2_decap_8 FILLER_95_144 ();
 sg13g2_decap_8 FILLER_95_151 ();
 sg13g2_decap_8 FILLER_95_158 ();
 sg13g2_decap_8 FILLER_95_165 ();
 sg13g2_decap_8 FILLER_95_172 ();
 sg13g2_decap_8 FILLER_95_179 ();
 sg13g2_decap_8 FILLER_95_186 ();
 sg13g2_decap_8 FILLER_95_193 ();
 sg13g2_decap_8 FILLER_95_200 ();
 sg13g2_decap_8 FILLER_95_207 ();
 sg13g2_decap_8 FILLER_95_214 ();
 sg13g2_decap_8 FILLER_95_221 ();
 sg13g2_decap_8 FILLER_95_228 ();
 sg13g2_decap_8 FILLER_95_235 ();
 sg13g2_decap_8 FILLER_95_242 ();
 sg13g2_decap_8 FILLER_95_249 ();
 sg13g2_decap_8 FILLER_95_256 ();
 sg13g2_decap_8 FILLER_95_263 ();
 sg13g2_decap_8 FILLER_95_270 ();
 sg13g2_decap_8 FILLER_95_277 ();
 sg13g2_decap_8 FILLER_95_284 ();
 sg13g2_decap_8 FILLER_95_291 ();
 sg13g2_decap_8 FILLER_95_298 ();
 sg13g2_decap_8 FILLER_95_305 ();
 sg13g2_decap_8 FILLER_95_312 ();
 sg13g2_decap_8 FILLER_95_319 ();
 sg13g2_decap_8 FILLER_95_326 ();
 sg13g2_decap_8 FILLER_95_333 ();
 sg13g2_decap_8 FILLER_95_340 ();
 sg13g2_decap_8 FILLER_95_347 ();
 sg13g2_decap_8 FILLER_95_354 ();
 sg13g2_decap_8 FILLER_95_361 ();
 sg13g2_decap_8 FILLER_95_368 ();
 sg13g2_decap_8 FILLER_95_375 ();
 sg13g2_decap_8 FILLER_95_382 ();
 sg13g2_decap_8 FILLER_95_389 ();
 sg13g2_decap_8 FILLER_95_396 ();
 sg13g2_decap_8 FILLER_95_403 ();
 sg13g2_decap_8 FILLER_95_410 ();
 sg13g2_decap_8 FILLER_95_417 ();
 sg13g2_decap_8 FILLER_95_424 ();
 sg13g2_decap_8 FILLER_95_431 ();
 sg13g2_decap_8 FILLER_95_438 ();
 sg13g2_decap_8 FILLER_95_445 ();
 sg13g2_decap_8 FILLER_95_452 ();
 sg13g2_decap_8 FILLER_95_459 ();
 sg13g2_decap_8 FILLER_95_466 ();
 sg13g2_decap_8 FILLER_95_473 ();
 sg13g2_decap_8 FILLER_95_480 ();
 sg13g2_decap_8 FILLER_95_487 ();
 sg13g2_decap_8 FILLER_95_494 ();
 sg13g2_decap_8 FILLER_95_501 ();
 sg13g2_decap_8 FILLER_95_508 ();
 sg13g2_decap_8 FILLER_95_515 ();
 sg13g2_decap_8 FILLER_95_522 ();
 sg13g2_decap_8 FILLER_95_529 ();
 sg13g2_decap_8 FILLER_95_536 ();
 sg13g2_decap_8 FILLER_95_543 ();
 sg13g2_decap_8 FILLER_95_550 ();
 sg13g2_decap_8 FILLER_95_557 ();
 sg13g2_decap_8 FILLER_95_564 ();
 sg13g2_decap_8 FILLER_95_571 ();
 sg13g2_decap_8 FILLER_95_578 ();
 sg13g2_decap_8 FILLER_95_585 ();
 sg13g2_decap_8 FILLER_95_592 ();
 sg13g2_decap_8 FILLER_95_599 ();
 sg13g2_decap_8 FILLER_95_606 ();
 sg13g2_decap_8 FILLER_95_613 ();
 sg13g2_decap_8 FILLER_95_620 ();
 sg13g2_decap_8 FILLER_95_627 ();
 sg13g2_decap_8 FILLER_95_634 ();
 sg13g2_decap_8 FILLER_95_641 ();
 sg13g2_decap_8 FILLER_95_648 ();
 sg13g2_decap_8 FILLER_95_655 ();
 sg13g2_decap_8 FILLER_95_662 ();
 sg13g2_decap_8 FILLER_95_669 ();
 sg13g2_decap_8 FILLER_95_676 ();
 sg13g2_decap_8 FILLER_95_683 ();
 sg13g2_decap_8 FILLER_95_690 ();
 sg13g2_decap_8 FILLER_95_697 ();
 sg13g2_decap_8 FILLER_95_704 ();
 sg13g2_decap_8 FILLER_95_711 ();
 sg13g2_decap_8 FILLER_95_718 ();
 sg13g2_decap_8 FILLER_95_725 ();
 sg13g2_decap_8 FILLER_95_732 ();
 sg13g2_decap_8 FILLER_95_739 ();
 sg13g2_decap_8 FILLER_95_746 ();
 sg13g2_decap_8 FILLER_95_753 ();
 sg13g2_decap_8 FILLER_95_760 ();
 sg13g2_decap_8 FILLER_95_767 ();
 sg13g2_decap_8 FILLER_95_774 ();
 sg13g2_decap_8 FILLER_95_781 ();
 sg13g2_decap_8 FILLER_95_788 ();
 sg13g2_decap_8 FILLER_95_795 ();
 sg13g2_decap_8 FILLER_95_802 ();
 sg13g2_decap_8 FILLER_95_809 ();
 sg13g2_decap_8 FILLER_95_816 ();
 sg13g2_decap_8 FILLER_95_823 ();
 sg13g2_decap_8 FILLER_95_830 ();
 sg13g2_decap_8 FILLER_95_837 ();
 sg13g2_decap_8 FILLER_95_844 ();
 sg13g2_decap_8 FILLER_95_851 ();
 sg13g2_decap_8 FILLER_95_858 ();
 sg13g2_decap_8 FILLER_95_865 ();
 sg13g2_decap_8 FILLER_95_872 ();
 sg13g2_decap_8 FILLER_95_879 ();
 sg13g2_decap_8 FILLER_95_886 ();
 sg13g2_decap_8 FILLER_95_893 ();
 sg13g2_decap_8 FILLER_95_900 ();
 sg13g2_decap_8 FILLER_95_907 ();
 sg13g2_decap_8 FILLER_95_914 ();
 sg13g2_decap_8 FILLER_95_921 ();
 sg13g2_decap_8 FILLER_95_928 ();
 sg13g2_decap_8 FILLER_95_935 ();
 sg13g2_decap_8 FILLER_95_942 ();
 sg13g2_decap_8 FILLER_95_949 ();
 sg13g2_decap_8 FILLER_95_956 ();
 sg13g2_decap_8 FILLER_95_963 ();
 sg13g2_decap_8 FILLER_95_970 ();
 sg13g2_decap_8 FILLER_95_977 ();
 sg13g2_decap_8 FILLER_95_984 ();
 sg13g2_decap_8 FILLER_95_991 ();
 sg13g2_decap_8 FILLER_95_998 ();
 sg13g2_decap_8 FILLER_95_1005 ();
 sg13g2_decap_8 FILLER_95_1012 ();
 sg13g2_decap_8 FILLER_95_1019 ();
 sg13g2_fill_2 FILLER_95_1026 ();
 sg13g2_fill_1 FILLER_95_1028 ();
 sg13g2_decap_8 FILLER_96_0 ();
 sg13g2_decap_8 FILLER_96_7 ();
 sg13g2_decap_8 FILLER_96_14 ();
 sg13g2_decap_8 FILLER_96_21 ();
 sg13g2_decap_8 FILLER_96_28 ();
 sg13g2_decap_8 FILLER_96_35 ();
 sg13g2_decap_8 FILLER_96_42 ();
 sg13g2_decap_8 FILLER_96_49 ();
 sg13g2_decap_8 FILLER_96_56 ();
 sg13g2_decap_8 FILLER_96_63 ();
 sg13g2_decap_8 FILLER_96_70 ();
 sg13g2_decap_8 FILLER_96_77 ();
 sg13g2_decap_8 FILLER_96_84 ();
 sg13g2_decap_8 FILLER_96_91 ();
 sg13g2_decap_8 FILLER_96_98 ();
 sg13g2_decap_8 FILLER_96_105 ();
 sg13g2_decap_8 FILLER_96_112 ();
 sg13g2_decap_8 FILLER_96_119 ();
 sg13g2_decap_8 FILLER_96_126 ();
 sg13g2_decap_8 FILLER_96_133 ();
 sg13g2_decap_8 FILLER_96_140 ();
 sg13g2_decap_8 FILLER_96_147 ();
 sg13g2_decap_8 FILLER_96_154 ();
 sg13g2_decap_8 FILLER_96_161 ();
 sg13g2_decap_8 FILLER_96_168 ();
 sg13g2_decap_8 FILLER_96_175 ();
 sg13g2_decap_8 FILLER_96_182 ();
 sg13g2_decap_8 FILLER_96_189 ();
 sg13g2_decap_8 FILLER_96_196 ();
 sg13g2_decap_8 FILLER_96_203 ();
 sg13g2_decap_8 FILLER_96_210 ();
 sg13g2_decap_8 FILLER_96_217 ();
 sg13g2_decap_8 FILLER_96_224 ();
 sg13g2_decap_8 FILLER_96_231 ();
 sg13g2_decap_8 FILLER_96_238 ();
 sg13g2_decap_8 FILLER_96_245 ();
 sg13g2_decap_8 FILLER_96_252 ();
 sg13g2_decap_8 FILLER_96_259 ();
 sg13g2_decap_8 FILLER_96_266 ();
 sg13g2_decap_8 FILLER_96_273 ();
 sg13g2_decap_8 FILLER_96_280 ();
 sg13g2_decap_8 FILLER_96_287 ();
 sg13g2_decap_8 FILLER_96_294 ();
 sg13g2_decap_8 FILLER_96_301 ();
 sg13g2_decap_8 FILLER_96_308 ();
 sg13g2_decap_8 FILLER_96_315 ();
 sg13g2_decap_8 FILLER_96_322 ();
 sg13g2_decap_8 FILLER_96_329 ();
 sg13g2_decap_8 FILLER_96_336 ();
 sg13g2_decap_8 FILLER_96_343 ();
 sg13g2_decap_8 FILLER_96_350 ();
 sg13g2_decap_8 FILLER_96_357 ();
 sg13g2_decap_8 FILLER_96_364 ();
 sg13g2_decap_8 FILLER_96_371 ();
 sg13g2_decap_8 FILLER_96_378 ();
 sg13g2_decap_8 FILLER_96_385 ();
 sg13g2_decap_8 FILLER_96_392 ();
 sg13g2_decap_8 FILLER_96_399 ();
 sg13g2_decap_8 FILLER_96_406 ();
 sg13g2_decap_8 FILLER_96_413 ();
 sg13g2_decap_8 FILLER_96_420 ();
 sg13g2_decap_8 FILLER_96_427 ();
 sg13g2_decap_8 FILLER_96_434 ();
 sg13g2_decap_8 FILLER_96_441 ();
 sg13g2_decap_8 FILLER_96_448 ();
 sg13g2_decap_8 FILLER_96_455 ();
 sg13g2_decap_8 FILLER_96_462 ();
 sg13g2_decap_8 FILLER_96_469 ();
 sg13g2_decap_8 FILLER_96_476 ();
 sg13g2_decap_8 FILLER_96_483 ();
 sg13g2_decap_8 FILLER_96_490 ();
 sg13g2_decap_8 FILLER_96_497 ();
 sg13g2_decap_8 FILLER_96_504 ();
 sg13g2_decap_8 FILLER_96_511 ();
 sg13g2_decap_8 FILLER_96_518 ();
 sg13g2_decap_8 FILLER_96_525 ();
 sg13g2_decap_8 FILLER_96_532 ();
 sg13g2_decap_8 FILLER_96_539 ();
 sg13g2_decap_8 FILLER_96_546 ();
 sg13g2_decap_8 FILLER_96_553 ();
 sg13g2_decap_8 FILLER_96_560 ();
 sg13g2_decap_8 FILLER_96_567 ();
 sg13g2_decap_8 FILLER_96_574 ();
 sg13g2_decap_8 FILLER_96_581 ();
 sg13g2_decap_8 FILLER_96_588 ();
 sg13g2_decap_8 FILLER_96_595 ();
 sg13g2_decap_8 FILLER_96_602 ();
 sg13g2_decap_8 FILLER_96_609 ();
 sg13g2_decap_8 FILLER_96_616 ();
 sg13g2_decap_8 FILLER_96_623 ();
 sg13g2_decap_8 FILLER_96_630 ();
 sg13g2_decap_8 FILLER_96_637 ();
 sg13g2_decap_8 FILLER_96_644 ();
 sg13g2_decap_8 FILLER_96_651 ();
 sg13g2_decap_8 FILLER_96_658 ();
 sg13g2_decap_8 FILLER_96_665 ();
 sg13g2_decap_8 FILLER_96_672 ();
 sg13g2_decap_8 FILLER_96_679 ();
 sg13g2_decap_8 FILLER_96_686 ();
 sg13g2_decap_8 FILLER_96_693 ();
 sg13g2_decap_8 FILLER_96_700 ();
 sg13g2_decap_8 FILLER_96_707 ();
 sg13g2_decap_8 FILLER_96_714 ();
 sg13g2_decap_8 FILLER_96_721 ();
 sg13g2_decap_8 FILLER_96_728 ();
 sg13g2_decap_8 FILLER_96_735 ();
 sg13g2_decap_8 FILLER_96_742 ();
 sg13g2_decap_8 FILLER_96_749 ();
 sg13g2_decap_8 FILLER_96_756 ();
 sg13g2_decap_8 FILLER_96_763 ();
 sg13g2_decap_8 FILLER_96_770 ();
 sg13g2_decap_8 FILLER_96_777 ();
 sg13g2_decap_8 FILLER_96_784 ();
 sg13g2_decap_8 FILLER_96_791 ();
 sg13g2_decap_8 FILLER_96_798 ();
 sg13g2_decap_8 FILLER_96_805 ();
 sg13g2_decap_8 FILLER_96_812 ();
 sg13g2_decap_8 FILLER_96_819 ();
 sg13g2_decap_8 FILLER_96_826 ();
 sg13g2_decap_8 FILLER_96_833 ();
 sg13g2_decap_8 FILLER_96_840 ();
 sg13g2_decap_8 FILLER_96_847 ();
 sg13g2_decap_8 FILLER_96_854 ();
 sg13g2_decap_8 FILLER_96_861 ();
 sg13g2_decap_8 FILLER_96_868 ();
 sg13g2_decap_8 FILLER_96_875 ();
 sg13g2_decap_8 FILLER_96_882 ();
 sg13g2_decap_8 FILLER_96_889 ();
 sg13g2_decap_8 FILLER_96_896 ();
 sg13g2_decap_8 FILLER_96_903 ();
 sg13g2_decap_8 FILLER_96_910 ();
 sg13g2_decap_8 FILLER_96_917 ();
 sg13g2_decap_8 FILLER_96_924 ();
 sg13g2_decap_8 FILLER_96_931 ();
 sg13g2_decap_8 FILLER_96_938 ();
 sg13g2_decap_8 FILLER_96_945 ();
 sg13g2_decap_8 FILLER_96_952 ();
 sg13g2_decap_8 FILLER_96_959 ();
 sg13g2_decap_8 FILLER_96_966 ();
 sg13g2_decap_8 FILLER_96_973 ();
 sg13g2_decap_8 FILLER_96_980 ();
 sg13g2_decap_8 FILLER_96_987 ();
 sg13g2_decap_8 FILLER_96_994 ();
 sg13g2_decap_8 FILLER_96_1001 ();
 sg13g2_decap_8 FILLER_96_1008 ();
 sg13g2_decap_8 FILLER_96_1015 ();
 sg13g2_decap_8 FILLER_96_1022 ();
 sg13g2_decap_8 FILLER_97_0 ();
 sg13g2_decap_8 FILLER_97_7 ();
 sg13g2_decap_8 FILLER_97_14 ();
 sg13g2_decap_8 FILLER_97_21 ();
 sg13g2_decap_8 FILLER_97_28 ();
 sg13g2_decap_8 FILLER_97_35 ();
 sg13g2_decap_8 FILLER_97_42 ();
 sg13g2_decap_8 FILLER_97_49 ();
 sg13g2_decap_8 FILLER_97_56 ();
 sg13g2_decap_8 FILLER_97_63 ();
 sg13g2_decap_8 FILLER_97_70 ();
 sg13g2_decap_8 FILLER_97_77 ();
 sg13g2_decap_8 FILLER_97_84 ();
 sg13g2_decap_8 FILLER_97_91 ();
 sg13g2_decap_8 FILLER_97_98 ();
 sg13g2_decap_8 FILLER_97_105 ();
 sg13g2_decap_8 FILLER_97_112 ();
 sg13g2_decap_8 FILLER_97_119 ();
 sg13g2_decap_8 FILLER_97_126 ();
 sg13g2_decap_8 FILLER_97_133 ();
 sg13g2_decap_8 FILLER_97_140 ();
 sg13g2_decap_8 FILLER_97_147 ();
 sg13g2_decap_8 FILLER_97_154 ();
 sg13g2_decap_8 FILLER_97_161 ();
 sg13g2_decap_8 FILLER_97_168 ();
 sg13g2_decap_8 FILLER_97_175 ();
 sg13g2_decap_8 FILLER_97_182 ();
 sg13g2_decap_8 FILLER_97_189 ();
 sg13g2_decap_8 FILLER_97_196 ();
 sg13g2_decap_8 FILLER_97_203 ();
 sg13g2_decap_8 FILLER_97_210 ();
 sg13g2_decap_8 FILLER_97_217 ();
 sg13g2_decap_8 FILLER_97_224 ();
 sg13g2_decap_8 FILLER_97_231 ();
 sg13g2_decap_8 FILLER_97_238 ();
 sg13g2_decap_8 FILLER_97_245 ();
 sg13g2_decap_8 FILLER_97_252 ();
 sg13g2_decap_8 FILLER_97_259 ();
 sg13g2_decap_8 FILLER_97_266 ();
 sg13g2_decap_8 FILLER_97_273 ();
 sg13g2_decap_8 FILLER_97_280 ();
 sg13g2_decap_8 FILLER_97_287 ();
 sg13g2_decap_8 FILLER_97_294 ();
 sg13g2_decap_8 FILLER_97_301 ();
 sg13g2_decap_8 FILLER_97_308 ();
 sg13g2_decap_8 FILLER_97_315 ();
 sg13g2_decap_8 FILLER_97_322 ();
 sg13g2_decap_8 FILLER_97_329 ();
 sg13g2_decap_8 FILLER_97_336 ();
 sg13g2_decap_8 FILLER_97_343 ();
 sg13g2_decap_8 FILLER_97_350 ();
 sg13g2_decap_8 FILLER_97_357 ();
 sg13g2_decap_8 FILLER_97_364 ();
 sg13g2_decap_8 FILLER_97_371 ();
 sg13g2_decap_8 FILLER_97_378 ();
 sg13g2_decap_8 FILLER_97_385 ();
 sg13g2_decap_8 FILLER_97_392 ();
 sg13g2_decap_8 FILLER_97_399 ();
 sg13g2_decap_8 FILLER_97_406 ();
 sg13g2_decap_8 FILLER_97_413 ();
 sg13g2_decap_8 FILLER_97_420 ();
 sg13g2_decap_8 FILLER_97_427 ();
 sg13g2_decap_8 FILLER_97_434 ();
 sg13g2_decap_8 FILLER_97_441 ();
 sg13g2_decap_8 FILLER_97_448 ();
 sg13g2_decap_8 FILLER_97_455 ();
 sg13g2_decap_8 FILLER_97_462 ();
 sg13g2_decap_8 FILLER_97_469 ();
 sg13g2_decap_8 FILLER_97_476 ();
 sg13g2_decap_8 FILLER_97_483 ();
 sg13g2_decap_8 FILLER_97_490 ();
 sg13g2_decap_8 FILLER_97_497 ();
 sg13g2_decap_8 FILLER_97_504 ();
 sg13g2_decap_8 FILLER_97_511 ();
 sg13g2_decap_8 FILLER_97_518 ();
 sg13g2_decap_8 FILLER_97_525 ();
 sg13g2_decap_8 FILLER_97_532 ();
 sg13g2_decap_8 FILLER_97_539 ();
 sg13g2_decap_8 FILLER_97_546 ();
 sg13g2_decap_8 FILLER_97_553 ();
 sg13g2_decap_8 FILLER_97_560 ();
 sg13g2_decap_8 FILLER_97_567 ();
 sg13g2_decap_8 FILLER_97_574 ();
 sg13g2_decap_8 FILLER_97_581 ();
 sg13g2_decap_8 FILLER_97_588 ();
 sg13g2_decap_8 FILLER_97_595 ();
 sg13g2_decap_8 FILLER_97_602 ();
 sg13g2_decap_8 FILLER_97_609 ();
 sg13g2_decap_8 FILLER_97_616 ();
 sg13g2_decap_8 FILLER_97_623 ();
 sg13g2_decap_8 FILLER_97_630 ();
 sg13g2_decap_8 FILLER_97_637 ();
 sg13g2_decap_8 FILLER_97_644 ();
 sg13g2_decap_8 FILLER_97_651 ();
 sg13g2_decap_8 FILLER_97_658 ();
 sg13g2_decap_8 FILLER_97_665 ();
 sg13g2_decap_8 FILLER_97_672 ();
 sg13g2_decap_8 FILLER_97_679 ();
 sg13g2_decap_8 FILLER_97_686 ();
 sg13g2_decap_8 FILLER_97_693 ();
 sg13g2_decap_8 FILLER_97_700 ();
 sg13g2_decap_8 FILLER_97_707 ();
 sg13g2_decap_8 FILLER_97_714 ();
 sg13g2_decap_8 FILLER_97_721 ();
 sg13g2_decap_8 FILLER_97_728 ();
 sg13g2_decap_8 FILLER_97_735 ();
 sg13g2_decap_8 FILLER_97_742 ();
 sg13g2_decap_8 FILLER_97_749 ();
 sg13g2_decap_8 FILLER_97_756 ();
 sg13g2_decap_8 FILLER_97_763 ();
 sg13g2_decap_8 FILLER_97_770 ();
 sg13g2_decap_8 FILLER_97_777 ();
 sg13g2_decap_8 FILLER_97_784 ();
 sg13g2_decap_8 FILLER_97_791 ();
 sg13g2_decap_8 FILLER_97_798 ();
 sg13g2_decap_8 FILLER_97_805 ();
 sg13g2_decap_8 FILLER_97_812 ();
 sg13g2_decap_8 FILLER_97_819 ();
 sg13g2_decap_8 FILLER_97_826 ();
 sg13g2_decap_8 FILLER_97_833 ();
 sg13g2_decap_8 FILLER_97_840 ();
 sg13g2_decap_8 FILLER_97_847 ();
 sg13g2_decap_8 FILLER_97_854 ();
 sg13g2_decap_8 FILLER_97_861 ();
 sg13g2_decap_8 FILLER_97_868 ();
 sg13g2_decap_8 FILLER_97_875 ();
 sg13g2_decap_8 FILLER_97_882 ();
 sg13g2_decap_8 FILLER_97_889 ();
 sg13g2_decap_8 FILLER_97_896 ();
 sg13g2_decap_8 FILLER_97_903 ();
 sg13g2_decap_8 FILLER_97_910 ();
 sg13g2_decap_8 FILLER_97_917 ();
 sg13g2_decap_8 FILLER_97_924 ();
 sg13g2_decap_8 FILLER_97_931 ();
 sg13g2_decap_8 FILLER_97_938 ();
 sg13g2_decap_8 FILLER_97_945 ();
 sg13g2_decap_8 FILLER_97_952 ();
 sg13g2_decap_8 FILLER_97_959 ();
 sg13g2_decap_8 FILLER_97_966 ();
 sg13g2_decap_8 FILLER_97_973 ();
 sg13g2_decap_8 FILLER_97_980 ();
 sg13g2_decap_8 FILLER_97_987 ();
 sg13g2_decap_8 FILLER_97_994 ();
 sg13g2_decap_8 FILLER_97_1001 ();
 sg13g2_decap_8 FILLER_97_1008 ();
 sg13g2_decap_8 FILLER_97_1015 ();
 sg13g2_decap_8 FILLER_97_1022 ();
 sg13g2_decap_8 FILLER_98_4 ();
 sg13g2_decap_8 FILLER_98_11 ();
 sg13g2_decap_8 FILLER_98_18 ();
 sg13g2_decap_8 FILLER_98_25 ();
 sg13g2_decap_8 FILLER_98_32 ();
 sg13g2_decap_8 FILLER_98_39 ();
 sg13g2_decap_8 FILLER_98_46 ();
 sg13g2_decap_8 FILLER_98_53 ();
 sg13g2_decap_8 FILLER_98_60 ();
 sg13g2_decap_8 FILLER_98_67 ();
 sg13g2_decap_8 FILLER_98_74 ();
 sg13g2_decap_8 FILLER_98_81 ();
 sg13g2_decap_8 FILLER_98_88 ();
 sg13g2_decap_8 FILLER_98_95 ();
 sg13g2_decap_8 FILLER_98_102 ();
 sg13g2_decap_8 FILLER_98_109 ();
 sg13g2_decap_8 FILLER_98_116 ();
 sg13g2_decap_8 FILLER_98_123 ();
 sg13g2_decap_8 FILLER_98_130 ();
 sg13g2_decap_8 FILLER_98_137 ();
 sg13g2_decap_8 FILLER_98_144 ();
 sg13g2_decap_8 FILLER_98_151 ();
 sg13g2_decap_8 FILLER_98_158 ();
 sg13g2_decap_8 FILLER_98_165 ();
 sg13g2_decap_8 FILLER_98_172 ();
 sg13g2_decap_8 FILLER_98_179 ();
 sg13g2_decap_8 FILLER_98_186 ();
 sg13g2_decap_8 FILLER_98_193 ();
 sg13g2_decap_8 FILLER_98_200 ();
 sg13g2_decap_8 FILLER_98_207 ();
 sg13g2_decap_8 FILLER_98_214 ();
 sg13g2_decap_8 FILLER_98_221 ();
 sg13g2_decap_8 FILLER_98_228 ();
 sg13g2_decap_8 FILLER_98_235 ();
 sg13g2_decap_8 FILLER_98_242 ();
 sg13g2_decap_8 FILLER_98_249 ();
 sg13g2_decap_8 FILLER_98_256 ();
 sg13g2_decap_8 FILLER_98_263 ();
 sg13g2_decap_8 FILLER_98_270 ();
 sg13g2_decap_8 FILLER_98_277 ();
 sg13g2_decap_8 FILLER_98_284 ();
 sg13g2_decap_8 FILLER_98_291 ();
 sg13g2_decap_8 FILLER_98_298 ();
 sg13g2_decap_8 FILLER_98_305 ();
 sg13g2_decap_8 FILLER_98_312 ();
 sg13g2_decap_8 FILLER_98_319 ();
 sg13g2_decap_8 FILLER_98_326 ();
 sg13g2_decap_8 FILLER_98_333 ();
 sg13g2_decap_8 FILLER_98_340 ();
 sg13g2_decap_8 FILLER_98_347 ();
 sg13g2_decap_8 FILLER_98_354 ();
 sg13g2_decap_8 FILLER_98_361 ();
 sg13g2_decap_8 FILLER_98_368 ();
 sg13g2_decap_8 FILLER_98_375 ();
 sg13g2_decap_8 FILLER_98_382 ();
 sg13g2_decap_8 FILLER_98_389 ();
 sg13g2_decap_8 FILLER_98_396 ();
 sg13g2_decap_8 FILLER_98_403 ();
 sg13g2_decap_8 FILLER_98_410 ();
 sg13g2_decap_8 FILLER_98_417 ();
 sg13g2_decap_8 FILLER_98_424 ();
 sg13g2_decap_8 FILLER_98_431 ();
 sg13g2_decap_8 FILLER_98_438 ();
 sg13g2_decap_8 FILLER_98_445 ();
 sg13g2_decap_8 FILLER_98_452 ();
 sg13g2_decap_8 FILLER_98_459 ();
 sg13g2_decap_8 FILLER_98_466 ();
 sg13g2_decap_8 FILLER_98_473 ();
 sg13g2_decap_8 FILLER_98_480 ();
 sg13g2_decap_8 FILLER_98_487 ();
 sg13g2_decap_8 FILLER_98_494 ();
 sg13g2_decap_8 FILLER_98_501 ();
 sg13g2_decap_8 FILLER_98_508 ();
 sg13g2_decap_8 FILLER_98_515 ();
 sg13g2_decap_8 FILLER_98_522 ();
 sg13g2_decap_8 FILLER_98_529 ();
 sg13g2_decap_8 FILLER_98_536 ();
 sg13g2_decap_8 FILLER_98_543 ();
 sg13g2_decap_8 FILLER_98_550 ();
 sg13g2_decap_8 FILLER_98_557 ();
 sg13g2_decap_8 FILLER_98_564 ();
 sg13g2_decap_8 FILLER_98_571 ();
 sg13g2_decap_8 FILLER_98_578 ();
 sg13g2_decap_8 FILLER_98_585 ();
 sg13g2_decap_8 FILLER_98_592 ();
 sg13g2_decap_8 FILLER_98_599 ();
 sg13g2_decap_8 FILLER_98_606 ();
 sg13g2_decap_8 FILLER_98_613 ();
 sg13g2_decap_8 FILLER_98_620 ();
 sg13g2_decap_8 FILLER_98_627 ();
 sg13g2_decap_8 FILLER_98_634 ();
 sg13g2_decap_8 FILLER_98_641 ();
 sg13g2_decap_8 FILLER_98_648 ();
 sg13g2_decap_8 FILLER_98_655 ();
 sg13g2_decap_8 FILLER_98_662 ();
 sg13g2_decap_8 FILLER_98_669 ();
 sg13g2_decap_8 FILLER_98_676 ();
 sg13g2_decap_8 FILLER_98_683 ();
 sg13g2_decap_8 FILLER_98_690 ();
 sg13g2_decap_8 FILLER_98_697 ();
 sg13g2_decap_8 FILLER_98_704 ();
 sg13g2_decap_8 FILLER_98_711 ();
 sg13g2_decap_8 FILLER_98_718 ();
 sg13g2_decap_8 FILLER_98_725 ();
 sg13g2_decap_8 FILLER_98_732 ();
 sg13g2_decap_8 FILLER_98_739 ();
 sg13g2_decap_8 FILLER_98_746 ();
 sg13g2_decap_8 FILLER_98_753 ();
 sg13g2_decap_8 FILLER_98_760 ();
 sg13g2_decap_8 FILLER_98_767 ();
 sg13g2_decap_8 FILLER_98_774 ();
 sg13g2_decap_8 FILLER_98_781 ();
 sg13g2_decap_8 FILLER_98_788 ();
 sg13g2_decap_8 FILLER_98_795 ();
 sg13g2_decap_8 FILLER_98_802 ();
 sg13g2_decap_8 FILLER_98_809 ();
 sg13g2_decap_8 FILLER_98_816 ();
 sg13g2_decap_8 FILLER_98_823 ();
 sg13g2_decap_8 FILLER_98_830 ();
 sg13g2_decap_8 FILLER_98_837 ();
 sg13g2_decap_8 FILLER_98_844 ();
 sg13g2_decap_8 FILLER_98_851 ();
 sg13g2_decap_8 FILLER_98_858 ();
 sg13g2_decap_8 FILLER_98_865 ();
 sg13g2_decap_8 FILLER_98_872 ();
 sg13g2_decap_8 FILLER_98_879 ();
 sg13g2_decap_8 FILLER_98_886 ();
 sg13g2_decap_8 FILLER_98_893 ();
 sg13g2_decap_8 FILLER_98_900 ();
 sg13g2_decap_8 FILLER_98_907 ();
 sg13g2_decap_8 FILLER_98_914 ();
 sg13g2_decap_8 FILLER_98_921 ();
 sg13g2_decap_8 FILLER_98_928 ();
 sg13g2_decap_8 FILLER_98_935 ();
 sg13g2_decap_8 FILLER_98_942 ();
 sg13g2_decap_8 FILLER_98_949 ();
 sg13g2_decap_8 FILLER_98_956 ();
 sg13g2_decap_8 FILLER_98_963 ();
 sg13g2_decap_8 FILLER_98_970 ();
 sg13g2_decap_8 FILLER_98_977 ();
 sg13g2_decap_8 FILLER_98_984 ();
 sg13g2_decap_8 FILLER_98_991 ();
 sg13g2_decap_8 FILLER_98_998 ();
 sg13g2_decap_8 FILLER_98_1005 ();
 sg13g2_decap_8 FILLER_98_1012 ();
 sg13g2_decap_8 FILLER_98_1019 ();
 sg13g2_fill_2 FILLER_98_1026 ();
 sg13g2_fill_1 FILLER_98_1028 ();
 sg13g2_decap_8 FILLER_99_0 ();
 sg13g2_decap_8 FILLER_99_7 ();
 sg13g2_decap_8 FILLER_99_14 ();
 sg13g2_decap_8 FILLER_99_21 ();
 sg13g2_decap_8 FILLER_99_28 ();
 sg13g2_decap_8 FILLER_99_35 ();
 sg13g2_decap_8 FILLER_99_42 ();
 sg13g2_decap_8 FILLER_99_49 ();
 sg13g2_decap_8 FILLER_99_56 ();
 sg13g2_decap_8 FILLER_99_63 ();
 sg13g2_decap_8 FILLER_99_70 ();
 sg13g2_decap_8 FILLER_99_77 ();
 sg13g2_decap_8 FILLER_99_84 ();
 sg13g2_decap_8 FILLER_99_91 ();
 sg13g2_decap_8 FILLER_99_98 ();
 sg13g2_decap_8 FILLER_99_105 ();
 sg13g2_decap_8 FILLER_99_112 ();
 sg13g2_decap_8 FILLER_99_119 ();
 sg13g2_decap_8 FILLER_99_126 ();
 sg13g2_decap_8 FILLER_99_133 ();
 sg13g2_decap_8 FILLER_99_140 ();
 sg13g2_decap_8 FILLER_99_147 ();
 sg13g2_decap_8 FILLER_99_154 ();
 sg13g2_decap_8 FILLER_99_161 ();
 sg13g2_decap_8 FILLER_99_168 ();
 sg13g2_decap_8 FILLER_99_175 ();
 sg13g2_decap_8 FILLER_99_182 ();
 sg13g2_decap_8 FILLER_99_189 ();
 sg13g2_decap_8 FILLER_99_196 ();
 sg13g2_decap_8 FILLER_99_203 ();
 sg13g2_decap_8 FILLER_99_210 ();
 sg13g2_decap_8 FILLER_99_217 ();
 sg13g2_decap_8 FILLER_99_224 ();
 sg13g2_decap_8 FILLER_99_231 ();
 sg13g2_decap_8 FILLER_99_238 ();
 sg13g2_decap_8 FILLER_99_245 ();
 sg13g2_decap_8 FILLER_99_252 ();
 sg13g2_decap_8 FILLER_99_259 ();
 sg13g2_decap_8 FILLER_99_266 ();
 sg13g2_decap_8 FILLER_99_273 ();
 sg13g2_decap_8 FILLER_99_280 ();
 sg13g2_decap_8 FILLER_99_287 ();
 sg13g2_decap_8 FILLER_99_294 ();
 sg13g2_decap_8 FILLER_99_301 ();
 sg13g2_decap_8 FILLER_99_308 ();
 sg13g2_decap_8 FILLER_99_315 ();
 sg13g2_decap_8 FILLER_99_322 ();
 sg13g2_decap_8 FILLER_99_329 ();
 sg13g2_decap_8 FILLER_99_336 ();
 sg13g2_decap_8 FILLER_99_343 ();
 sg13g2_decap_8 FILLER_99_350 ();
 sg13g2_decap_8 FILLER_99_357 ();
 sg13g2_decap_8 FILLER_99_364 ();
 sg13g2_decap_8 FILLER_99_371 ();
 sg13g2_decap_8 FILLER_99_378 ();
 sg13g2_decap_8 FILLER_99_385 ();
 sg13g2_decap_8 FILLER_99_392 ();
 sg13g2_decap_8 FILLER_99_399 ();
 sg13g2_decap_8 FILLER_99_406 ();
 sg13g2_decap_8 FILLER_99_413 ();
 sg13g2_decap_8 FILLER_99_420 ();
 sg13g2_decap_8 FILLER_99_427 ();
 sg13g2_decap_8 FILLER_99_434 ();
 sg13g2_decap_8 FILLER_99_441 ();
 sg13g2_decap_8 FILLER_99_448 ();
 sg13g2_decap_8 FILLER_99_455 ();
 sg13g2_decap_8 FILLER_99_462 ();
 sg13g2_decap_8 FILLER_99_469 ();
 sg13g2_decap_8 FILLER_99_476 ();
 sg13g2_decap_8 FILLER_99_483 ();
 sg13g2_decap_8 FILLER_99_490 ();
 sg13g2_decap_8 FILLER_99_497 ();
 sg13g2_decap_8 FILLER_99_504 ();
 sg13g2_decap_8 FILLER_99_511 ();
 sg13g2_decap_8 FILLER_99_518 ();
 sg13g2_decap_8 FILLER_99_525 ();
 sg13g2_decap_8 FILLER_99_532 ();
 sg13g2_decap_8 FILLER_99_539 ();
 sg13g2_decap_8 FILLER_99_546 ();
 sg13g2_decap_8 FILLER_99_553 ();
 sg13g2_decap_8 FILLER_99_560 ();
 sg13g2_decap_8 FILLER_99_567 ();
 sg13g2_decap_8 FILLER_99_574 ();
 sg13g2_decap_8 FILLER_99_581 ();
 sg13g2_decap_8 FILLER_99_588 ();
 sg13g2_decap_8 FILLER_99_595 ();
 sg13g2_decap_8 FILLER_99_602 ();
 sg13g2_decap_8 FILLER_99_609 ();
 sg13g2_decap_8 FILLER_99_616 ();
 sg13g2_decap_8 FILLER_99_623 ();
 sg13g2_decap_8 FILLER_99_630 ();
 sg13g2_decap_8 FILLER_99_637 ();
 sg13g2_decap_8 FILLER_99_644 ();
 sg13g2_decap_8 FILLER_99_651 ();
 sg13g2_decap_8 FILLER_99_658 ();
 sg13g2_decap_8 FILLER_99_665 ();
 sg13g2_decap_8 FILLER_99_672 ();
 sg13g2_decap_8 FILLER_99_679 ();
 sg13g2_decap_8 FILLER_99_686 ();
 sg13g2_decap_8 FILLER_99_693 ();
 sg13g2_decap_8 FILLER_99_700 ();
 sg13g2_decap_8 FILLER_99_707 ();
 sg13g2_decap_8 FILLER_99_714 ();
 sg13g2_decap_8 FILLER_99_721 ();
 sg13g2_decap_8 FILLER_99_728 ();
 sg13g2_decap_8 FILLER_99_735 ();
 sg13g2_decap_8 FILLER_99_742 ();
 sg13g2_decap_8 FILLER_99_749 ();
 sg13g2_decap_8 FILLER_99_756 ();
 sg13g2_decap_8 FILLER_99_763 ();
 sg13g2_decap_8 FILLER_99_770 ();
 sg13g2_decap_8 FILLER_99_777 ();
 sg13g2_decap_8 FILLER_99_784 ();
 sg13g2_decap_8 FILLER_99_791 ();
 sg13g2_decap_8 FILLER_99_798 ();
 sg13g2_decap_8 FILLER_99_805 ();
 sg13g2_decap_8 FILLER_99_812 ();
 sg13g2_decap_8 FILLER_99_819 ();
 sg13g2_decap_8 FILLER_99_826 ();
 sg13g2_decap_8 FILLER_99_833 ();
 sg13g2_decap_8 FILLER_99_840 ();
 sg13g2_decap_8 FILLER_99_847 ();
 sg13g2_decap_8 FILLER_99_854 ();
 sg13g2_decap_8 FILLER_99_861 ();
 sg13g2_decap_8 FILLER_99_868 ();
 sg13g2_decap_8 FILLER_99_875 ();
 sg13g2_decap_8 FILLER_99_882 ();
 sg13g2_decap_8 FILLER_99_889 ();
 sg13g2_decap_8 FILLER_99_896 ();
 sg13g2_decap_8 FILLER_99_903 ();
 sg13g2_decap_8 FILLER_99_910 ();
 sg13g2_decap_8 FILLER_99_917 ();
 sg13g2_decap_8 FILLER_99_924 ();
 sg13g2_decap_8 FILLER_99_931 ();
 sg13g2_decap_8 FILLER_99_938 ();
 sg13g2_decap_8 FILLER_99_945 ();
 sg13g2_decap_8 FILLER_99_952 ();
 sg13g2_decap_8 FILLER_99_959 ();
 sg13g2_decap_8 FILLER_99_966 ();
 sg13g2_decap_8 FILLER_99_973 ();
 sg13g2_decap_8 FILLER_99_980 ();
 sg13g2_decap_8 FILLER_99_987 ();
 sg13g2_decap_8 FILLER_99_994 ();
 sg13g2_decap_8 FILLER_99_1001 ();
 sg13g2_decap_8 FILLER_99_1008 ();
 sg13g2_decap_8 FILLER_99_1015 ();
 sg13g2_decap_8 FILLER_99_1022 ();
 sg13g2_decap_8 FILLER_100_0 ();
 sg13g2_decap_8 FILLER_100_7 ();
 sg13g2_decap_8 FILLER_100_14 ();
 sg13g2_decap_8 FILLER_100_21 ();
 sg13g2_decap_8 FILLER_100_28 ();
 sg13g2_decap_8 FILLER_100_35 ();
 sg13g2_decap_8 FILLER_100_42 ();
 sg13g2_decap_8 FILLER_100_49 ();
 sg13g2_decap_8 FILLER_100_56 ();
 sg13g2_decap_8 FILLER_100_63 ();
 sg13g2_decap_8 FILLER_100_70 ();
 sg13g2_decap_8 FILLER_100_77 ();
 sg13g2_decap_8 FILLER_100_84 ();
 sg13g2_decap_8 FILLER_100_91 ();
 sg13g2_decap_8 FILLER_100_98 ();
 sg13g2_decap_8 FILLER_100_105 ();
 sg13g2_decap_8 FILLER_100_112 ();
 sg13g2_decap_8 FILLER_100_119 ();
 sg13g2_decap_8 FILLER_100_126 ();
 sg13g2_decap_8 FILLER_100_133 ();
 sg13g2_decap_8 FILLER_100_140 ();
 sg13g2_decap_8 FILLER_100_147 ();
 sg13g2_decap_8 FILLER_100_154 ();
 sg13g2_decap_8 FILLER_100_161 ();
 sg13g2_decap_8 FILLER_100_168 ();
 sg13g2_decap_8 FILLER_100_175 ();
 sg13g2_decap_8 FILLER_100_182 ();
 sg13g2_decap_8 FILLER_100_189 ();
 sg13g2_decap_8 FILLER_100_196 ();
 sg13g2_decap_8 FILLER_100_203 ();
 sg13g2_decap_8 FILLER_100_210 ();
 sg13g2_decap_8 FILLER_100_217 ();
 sg13g2_decap_8 FILLER_100_224 ();
 sg13g2_decap_8 FILLER_100_231 ();
 sg13g2_decap_8 FILLER_100_238 ();
 sg13g2_decap_8 FILLER_100_245 ();
 sg13g2_decap_8 FILLER_100_252 ();
 sg13g2_decap_8 FILLER_100_259 ();
 sg13g2_decap_8 FILLER_100_266 ();
 sg13g2_decap_8 FILLER_100_273 ();
 sg13g2_decap_8 FILLER_100_280 ();
 sg13g2_decap_8 FILLER_100_287 ();
 sg13g2_decap_8 FILLER_100_294 ();
 sg13g2_decap_8 FILLER_100_301 ();
 sg13g2_decap_8 FILLER_100_308 ();
 sg13g2_decap_8 FILLER_100_315 ();
 sg13g2_decap_8 FILLER_100_322 ();
 sg13g2_decap_8 FILLER_100_329 ();
 sg13g2_decap_8 FILLER_100_336 ();
 sg13g2_decap_8 FILLER_100_343 ();
 sg13g2_decap_8 FILLER_100_350 ();
 sg13g2_decap_8 FILLER_100_357 ();
 sg13g2_decap_8 FILLER_100_364 ();
 sg13g2_decap_8 FILLER_100_371 ();
 sg13g2_decap_8 FILLER_100_378 ();
 sg13g2_decap_8 FILLER_100_385 ();
 sg13g2_decap_8 FILLER_100_392 ();
 sg13g2_decap_8 FILLER_100_399 ();
 sg13g2_decap_8 FILLER_100_406 ();
 sg13g2_decap_8 FILLER_100_413 ();
 sg13g2_decap_8 FILLER_100_420 ();
 sg13g2_decap_8 FILLER_100_427 ();
 sg13g2_decap_8 FILLER_100_434 ();
 sg13g2_decap_8 FILLER_100_441 ();
 sg13g2_decap_8 FILLER_100_448 ();
 sg13g2_decap_8 FILLER_100_455 ();
 sg13g2_decap_8 FILLER_100_462 ();
 sg13g2_decap_8 FILLER_100_469 ();
 sg13g2_decap_8 FILLER_100_476 ();
 sg13g2_decap_8 FILLER_100_483 ();
 sg13g2_decap_8 FILLER_100_490 ();
 sg13g2_decap_8 FILLER_100_497 ();
 sg13g2_decap_8 FILLER_100_504 ();
 sg13g2_decap_8 FILLER_100_511 ();
 sg13g2_decap_8 FILLER_100_518 ();
 sg13g2_decap_8 FILLER_100_525 ();
 sg13g2_decap_8 FILLER_100_532 ();
 sg13g2_decap_8 FILLER_100_539 ();
 sg13g2_decap_8 FILLER_100_546 ();
 sg13g2_decap_8 FILLER_100_553 ();
 sg13g2_decap_8 FILLER_100_560 ();
 sg13g2_decap_8 FILLER_100_567 ();
 sg13g2_decap_8 FILLER_100_574 ();
 sg13g2_decap_8 FILLER_100_581 ();
 sg13g2_decap_8 FILLER_100_588 ();
 sg13g2_decap_8 FILLER_100_595 ();
 sg13g2_decap_8 FILLER_100_602 ();
 sg13g2_decap_8 FILLER_100_609 ();
 sg13g2_decap_8 FILLER_100_616 ();
 sg13g2_decap_8 FILLER_100_623 ();
 sg13g2_decap_8 FILLER_100_630 ();
 sg13g2_decap_8 FILLER_100_637 ();
 sg13g2_decap_8 FILLER_100_644 ();
 sg13g2_decap_8 FILLER_100_651 ();
 sg13g2_decap_8 FILLER_100_658 ();
 sg13g2_decap_8 FILLER_100_665 ();
 sg13g2_decap_8 FILLER_100_672 ();
 sg13g2_decap_8 FILLER_100_679 ();
 sg13g2_decap_8 FILLER_100_686 ();
 sg13g2_decap_8 FILLER_100_693 ();
 sg13g2_decap_8 FILLER_100_700 ();
 sg13g2_decap_8 FILLER_100_707 ();
 sg13g2_decap_8 FILLER_100_714 ();
 sg13g2_decap_8 FILLER_100_721 ();
 sg13g2_decap_8 FILLER_100_728 ();
 sg13g2_decap_8 FILLER_100_735 ();
 sg13g2_decap_8 FILLER_100_742 ();
 sg13g2_decap_8 FILLER_100_749 ();
 sg13g2_decap_8 FILLER_100_756 ();
 sg13g2_decap_8 FILLER_100_763 ();
 sg13g2_decap_8 FILLER_100_770 ();
 sg13g2_decap_8 FILLER_100_777 ();
 sg13g2_decap_8 FILLER_100_784 ();
 sg13g2_decap_8 FILLER_100_791 ();
 sg13g2_decap_8 FILLER_100_798 ();
 sg13g2_decap_8 FILLER_100_805 ();
 sg13g2_decap_8 FILLER_100_812 ();
 sg13g2_decap_8 FILLER_100_819 ();
 sg13g2_decap_8 FILLER_100_826 ();
 sg13g2_decap_8 FILLER_100_833 ();
 sg13g2_decap_8 FILLER_100_840 ();
 sg13g2_decap_8 FILLER_100_847 ();
 sg13g2_decap_8 FILLER_100_854 ();
 sg13g2_decap_8 FILLER_100_861 ();
 sg13g2_decap_8 FILLER_100_868 ();
 sg13g2_decap_8 FILLER_100_875 ();
 sg13g2_decap_8 FILLER_100_882 ();
 sg13g2_decap_8 FILLER_100_889 ();
 sg13g2_decap_8 FILLER_100_896 ();
 sg13g2_decap_8 FILLER_100_903 ();
 sg13g2_decap_8 FILLER_100_910 ();
 sg13g2_decap_8 FILLER_100_917 ();
 sg13g2_decap_8 FILLER_100_924 ();
 sg13g2_decap_8 FILLER_100_931 ();
 sg13g2_decap_8 FILLER_100_938 ();
 sg13g2_decap_8 FILLER_100_945 ();
 sg13g2_decap_8 FILLER_100_952 ();
 sg13g2_decap_8 FILLER_100_959 ();
 sg13g2_decap_8 FILLER_100_966 ();
 sg13g2_decap_8 FILLER_100_973 ();
 sg13g2_decap_8 FILLER_100_980 ();
 sg13g2_decap_8 FILLER_100_987 ();
 sg13g2_decap_8 FILLER_100_994 ();
 sg13g2_decap_8 FILLER_100_1001 ();
 sg13g2_decap_8 FILLER_100_1008 ();
 sg13g2_decap_8 FILLER_100_1015 ();
 sg13g2_decap_8 FILLER_100_1022 ();
 sg13g2_decap_8 FILLER_101_0 ();
 sg13g2_decap_8 FILLER_101_7 ();
 sg13g2_decap_8 FILLER_101_14 ();
 sg13g2_decap_8 FILLER_101_21 ();
 sg13g2_decap_8 FILLER_101_28 ();
 sg13g2_decap_8 FILLER_101_35 ();
 sg13g2_decap_8 FILLER_101_42 ();
 sg13g2_decap_8 FILLER_101_49 ();
 sg13g2_decap_8 FILLER_101_56 ();
 sg13g2_decap_8 FILLER_101_63 ();
 sg13g2_decap_8 FILLER_101_70 ();
 sg13g2_decap_8 FILLER_101_77 ();
 sg13g2_decap_8 FILLER_101_84 ();
 sg13g2_decap_8 FILLER_101_91 ();
 sg13g2_decap_8 FILLER_101_98 ();
 sg13g2_decap_8 FILLER_101_105 ();
 sg13g2_decap_8 FILLER_101_112 ();
 sg13g2_decap_8 FILLER_101_119 ();
 sg13g2_decap_8 FILLER_101_126 ();
 sg13g2_decap_8 FILLER_101_133 ();
 sg13g2_decap_8 FILLER_101_140 ();
 sg13g2_decap_8 FILLER_101_147 ();
 sg13g2_decap_8 FILLER_101_154 ();
 sg13g2_decap_8 FILLER_101_161 ();
 sg13g2_decap_8 FILLER_101_168 ();
 sg13g2_decap_8 FILLER_101_175 ();
 sg13g2_decap_8 FILLER_101_182 ();
 sg13g2_decap_8 FILLER_101_189 ();
 sg13g2_decap_8 FILLER_101_196 ();
 sg13g2_decap_8 FILLER_101_203 ();
 sg13g2_decap_8 FILLER_101_210 ();
 sg13g2_decap_8 FILLER_101_217 ();
 sg13g2_decap_8 FILLER_101_224 ();
 sg13g2_decap_8 FILLER_101_231 ();
 sg13g2_decap_8 FILLER_101_238 ();
 sg13g2_decap_8 FILLER_101_245 ();
 sg13g2_decap_8 FILLER_101_252 ();
 sg13g2_decap_8 FILLER_101_259 ();
 sg13g2_decap_8 FILLER_101_266 ();
 sg13g2_decap_8 FILLER_101_273 ();
 sg13g2_decap_8 FILLER_101_280 ();
 sg13g2_decap_8 FILLER_101_287 ();
 sg13g2_decap_8 FILLER_101_294 ();
 sg13g2_decap_8 FILLER_101_301 ();
 sg13g2_decap_8 FILLER_101_308 ();
 sg13g2_decap_8 FILLER_101_315 ();
 sg13g2_decap_8 FILLER_101_322 ();
 sg13g2_decap_8 FILLER_101_329 ();
 sg13g2_decap_8 FILLER_101_336 ();
 sg13g2_decap_8 FILLER_101_343 ();
 sg13g2_decap_8 FILLER_101_350 ();
 sg13g2_decap_8 FILLER_101_357 ();
 sg13g2_decap_8 FILLER_101_364 ();
 sg13g2_decap_8 FILLER_101_371 ();
 sg13g2_decap_8 FILLER_101_378 ();
 sg13g2_decap_8 FILLER_101_385 ();
 sg13g2_decap_8 FILLER_101_392 ();
 sg13g2_decap_8 FILLER_101_399 ();
 sg13g2_decap_8 FILLER_101_406 ();
 sg13g2_decap_8 FILLER_101_413 ();
 sg13g2_decap_8 FILLER_101_420 ();
 sg13g2_decap_8 FILLER_101_427 ();
 sg13g2_decap_8 FILLER_101_434 ();
 sg13g2_decap_8 FILLER_101_441 ();
 sg13g2_decap_8 FILLER_101_448 ();
 sg13g2_decap_8 FILLER_101_455 ();
 sg13g2_decap_8 FILLER_101_462 ();
 sg13g2_decap_8 FILLER_101_469 ();
 sg13g2_decap_8 FILLER_101_476 ();
 sg13g2_decap_8 FILLER_101_483 ();
 sg13g2_decap_8 FILLER_101_490 ();
 sg13g2_decap_8 FILLER_101_497 ();
 sg13g2_decap_8 FILLER_101_504 ();
 sg13g2_decap_8 FILLER_101_511 ();
 sg13g2_decap_8 FILLER_101_518 ();
 sg13g2_decap_8 FILLER_101_525 ();
 sg13g2_decap_8 FILLER_101_532 ();
 sg13g2_decap_8 FILLER_101_539 ();
 sg13g2_decap_8 FILLER_101_546 ();
 sg13g2_decap_8 FILLER_101_553 ();
 sg13g2_decap_8 FILLER_101_560 ();
 sg13g2_decap_8 FILLER_101_567 ();
 sg13g2_decap_8 FILLER_101_574 ();
 sg13g2_decap_8 FILLER_101_581 ();
 sg13g2_decap_8 FILLER_101_588 ();
 sg13g2_decap_8 FILLER_101_595 ();
 sg13g2_decap_8 FILLER_101_602 ();
 sg13g2_decap_8 FILLER_101_609 ();
 sg13g2_decap_8 FILLER_101_616 ();
 sg13g2_decap_8 FILLER_101_623 ();
 sg13g2_decap_8 FILLER_101_630 ();
 sg13g2_decap_8 FILLER_101_637 ();
 sg13g2_decap_8 FILLER_101_644 ();
 sg13g2_decap_8 FILLER_101_651 ();
 sg13g2_decap_8 FILLER_101_658 ();
 sg13g2_decap_8 FILLER_101_665 ();
 sg13g2_decap_8 FILLER_101_672 ();
 sg13g2_decap_8 FILLER_101_679 ();
 sg13g2_decap_8 FILLER_101_686 ();
 sg13g2_decap_8 FILLER_101_693 ();
 sg13g2_decap_8 FILLER_101_700 ();
 sg13g2_decap_8 FILLER_101_707 ();
 sg13g2_decap_8 FILLER_101_714 ();
 sg13g2_decap_8 FILLER_101_721 ();
 sg13g2_decap_8 FILLER_101_728 ();
 sg13g2_decap_8 FILLER_101_735 ();
 sg13g2_decap_8 FILLER_101_742 ();
 sg13g2_decap_8 FILLER_101_749 ();
 sg13g2_decap_8 FILLER_101_756 ();
 sg13g2_decap_8 FILLER_101_763 ();
 sg13g2_decap_8 FILLER_101_770 ();
 sg13g2_decap_8 FILLER_101_777 ();
 sg13g2_decap_8 FILLER_101_784 ();
 sg13g2_decap_8 FILLER_101_791 ();
 sg13g2_decap_8 FILLER_101_798 ();
 sg13g2_decap_8 FILLER_101_805 ();
 sg13g2_decap_8 FILLER_101_812 ();
 sg13g2_decap_8 FILLER_101_819 ();
 sg13g2_decap_8 FILLER_101_826 ();
 sg13g2_decap_8 FILLER_101_833 ();
 sg13g2_decap_8 FILLER_101_840 ();
 sg13g2_decap_8 FILLER_101_847 ();
 sg13g2_decap_8 FILLER_101_854 ();
 sg13g2_decap_8 FILLER_101_861 ();
 sg13g2_decap_8 FILLER_101_868 ();
 sg13g2_decap_8 FILLER_101_875 ();
 sg13g2_decap_8 FILLER_101_882 ();
 sg13g2_decap_8 FILLER_101_889 ();
 sg13g2_decap_8 FILLER_101_896 ();
 sg13g2_decap_8 FILLER_101_903 ();
 sg13g2_decap_8 FILLER_101_910 ();
 sg13g2_decap_8 FILLER_101_917 ();
 sg13g2_decap_8 FILLER_101_924 ();
 sg13g2_decap_8 FILLER_101_931 ();
 sg13g2_decap_8 FILLER_101_938 ();
 sg13g2_decap_8 FILLER_101_945 ();
 sg13g2_decap_8 FILLER_101_952 ();
 sg13g2_decap_8 FILLER_101_959 ();
 sg13g2_decap_8 FILLER_101_966 ();
 sg13g2_decap_8 FILLER_101_973 ();
 sg13g2_decap_8 FILLER_101_980 ();
 sg13g2_decap_8 FILLER_101_987 ();
 sg13g2_decap_8 FILLER_101_994 ();
 sg13g2_decap_8 FILLER_101_1001 ();
 sg13g2_decap_8 FILLER_101_1008 ();
 sg13g2_decap_8 FILLER_101_1015 ();
 sg13g2_decap_8 FILLER_101_1022 ();
 sg13g2_decap_8 FILLER_102_0 ();
 sg13g2_decap_8 FILLER_102_7 ();
 sg13g2_decap_8 FILLER_102_14 ();
 sg13g2_decap_8 FILLER_102_21 ();
 sg13g2_decap_8 FILLER_102_28 ();
 sg13g2_decap_8 FILLER_102_35 ();
 sg13g2_decap_8 FILLER_102_42 ();
 sg13g2_decap_8 FILLER_102_49 ();
 sg13g2_decap_8 FILLER_102_56 ();
 sg13g2_decap_8 FILLER_102_63 ();
 sg13g2_decap_8 FILLER_102_70 ();
 sg13g2_decap_8 FILLER_102_77 ();
 sg13g2_decap_8 FILLER_102_84 ();
 sg13g2_decap_8 FILLER_102_91 ();
 sg13g2_decap_8 FILLER_102_98 ();
 sg13g2_decap_8 FILLER_102_105 ();
 sg13g2_decap_8 FILLER_102_112 ();
 sg13g2_decap_8 FILLER_102_119 ();
 sg13g2_decap_8 FILLER_102_126 ();
 sg13g2_decap_8 FILLER_102_133 ();
 sg13g2_decap_8 FILLER_102_140 ();
 sg13g2_decap_8 FILLER_102_147 ();
 sg13g2_decap_8 FILLER_102_154 ();
 sg13g2_decap_8 FILLER_102_161 ();
 sg13g2_decap_8 FILLER_102_168 ();
 sg13g2_decap_8 FILLER_102_175 ();
 sg13g2_decap_8 FILLER_102_182 ();
 sg13g2_decap_8 FILLER_102_189 ();
 sg13g2_decap_8 FILLER_102_196 ();
 sg13g2_decap_8 FILLER_102_203 ();
 sg13g2_decap_8 FILLER_102_210 ();
 sg13g2_decap_8 FILLER_102_217 ();
 sg13g2_decap_8 FILLER_102_224 ();
 sg13g2_decap_8 FILLER_102_231 ();
 sg13g2_decap_8 FILLER_102_238 ();
 sg13g2_decap_8 FILLER_102_245 ();
 sg13g2_decap_8 FILLER_102_252 ();
 sg13g2_decap_8 FILLER_102_259 ();
 sg13g2_decap_8 FILLER_102_266 ();
 sg13g2_decap_8 FILLER_102_273 ();
 sg13g2_decap_8 FILLER_102_280 ();
 sg13g2_decap_8 FILLER_102_287 ();
 sg13g2_decap_8 FILLER_102_294 ();
 sg13g2_decap_8 FILLER_102_301 ();
 sg13g2_decap_8 FILLER_102_308 ();
 sg13g2_decap_8 FILLER_102_315 ();
 sg13g2_decap_8 FILLER_102_322 ();
 sg13g2_decap_8 FILLER_102_329 ();
 sg13g2_decap_8 FILLER_102_336 ();
 sg13g2_decap_8 FILLER_102_343 ();
 sg13g2_decap_8 FILLER_102_350 ();
 sg13g2_decap_8 FILLER_102_357 ();
 sg13g2_decap_8 FILLER_102_364 ();
 sg13g2_decap_8 FILLER_102_371 ();
 sg13g2_decap_8 FILLER_102_378 ();
 sg13g2_decap_8 FILLER_102_385 ();
 sg13g2_decap_8 FILLER_102_392 ();
 sg13g2_decap_8 FILLER_102_399 ();
 sg13g2_decap_8 FILLER_102_406 ();
 sg13g2_decap_8 FILLER_102_413 ();
 sg13g2_decap_8 FILLER_102_420 ();
 sg13g2_decap_8 FILLER_102_427 ();
 sg13g2_decap_8 FILLER_102_434 ();
 sg13g2_decap_8 FILLER_102_441 ();
 sg13g2_decap_8 FILLER_102_448 ();
 sg13g2_decap_8 FILLER_102_455 ();
 sg13g2_decap_8 FILLER_102_462 ();
 sg13g2_decap_8 FILLER_102_469 ();
 sg13g2_decap_8 FILLER_102_476 ();
 sg13g2_decap_8 FILLER_102_483 ();
 sg13g2_decap_8 FILLER_102_490 ();
 sg13g2_decap_8 FILLER_102_497 ();
 sg13g2_decap_8 FILLER_102_504 ();
 sg13g2_decap_8 FILLER_102_511 ();
 sg13g2_decap_8 FILLER_102_518 ();
 sg13g2_decap_8 FILLER_102_525 ();
 sg13g2_decap_8 FILLER_102_532 ();
 sg13g2_decap_8 FILLER_102_539 ();
 sg13g2_decap_8 FILLER_102_546 ();
 sg13g2_decap_8 FILLER_102_553 ();
 sg13g2_decap_8 FILLER_102_560 ();
 sg13g2_decap_8 FILLER_102_567 ();
 sg13g2_decap_8 FILLER_102_574 ();
 sg13g2_decap_8 FILLER_102_581 ();
 sg13g2_decap_8 FILLER_102_588 ();
 sg13g2_decap_8 FILLER_102_595 ();
 sg13g2_decap_8 FILLER_102_602 ();
 sg13g2_decap_8 FILLER_102_609 ();
 sg13g2_decap_8 FILLER_102_616 ();
 sg13g2_decap_8 FILLER_102_623 ();
 sg13g2_decap_8 FILLER_102_630 ();
 sg13g2_decap_8 FILLER_102_637 ();
 sg13g2_decap_8 FILLER_102_644 ();
 sg13g2_decap_8 FILLER_102_651 ();
 sg13g2_decap_8 FILLER_102_658 ();
 sg13g2_decap_8 FILLER_102_665 ();
 sg13g2_decap_8 FILLER_102_672 ();
 sg13g2_decap_8 FILLER_102_679 ();
 sg13g2_decap_8 FILLER_102_686 ();
 sg13g2_decap_8 FILLER_102_693 ();
 sg13g2_decap_8 FILLER_102_700 ();
 sg13g2_decap_8 FILLER_102_707 ();
 sg13g2_decap_8 FILLER_102_714 ();
 sg13g2_decap_8 FILLER_102_721 ();
 sg13g2_decap_8 FILLER_102_728 ();
 sg13g2_decap_8 FILLER_102_735 ();
 sg13g2_decap_8 FILLER_102_742 ();
 sg13g2_decap_8 FILLER_102_749 ();
 sg13g2_decap_8 FILLER_102_756 ();
 sg13g2_decap_8 FILLER_102_763 ();
 sg13g2_decap_8 FILLER_102_770 ();
 sg13g2_decap_8 FILLER_102_777 ();
 sg13g2_decap_8 FILLER_102_784 ();
 sg13g2_decap_8 FILLER_102_791 ();
 sg13g2_decap_8 FILLER_102_798 ();
 sg13g2_decap_8 FILLER_102_805 ();
 sg13g2_decap_8 FILLER_102_812 ();
 sg13g2_decap_8 FILLER_102_819 ();
 sg13g2_decap_8 FILLER_102_826 ();
 sg13g2_decap_8 FILLER_102_833 ();
 sg13g2_decap_8 FILLER_102_840 ();
 sg13g2_decap_8 FILLER_102_847 ();
 sg13g2_decap_8 FILLER_102_854 ();
 sg13g2_decap_8 FILLER_102_861 ();
 sg13g2_decap_8 FILLER_102_868 ();
 sg13g2_decap_8 FILLER_102_875 ();
 sg13g2_decap_8 FILLER_102_882 ();
 sg13g2_decap_8 FILLER_102_889 ();
 sg13g2_decap_8 FILLER_102_896 ();
 sg13g2_decap_8 FILLER_102_903 ();
 sg13g2_decap_8 FILLER_102_910 ();
 sg13g2_decap_8 FILLER_102_917 ();
 sg13g2_decap_8 FILLER_102_924 ();
 sg13g2_decap_8 FILLER_102_931 ();
 sg13g2_decap_8 FILLER_102_938 ();
 sg13g2_decap_8 FILLER_102_945 ();
 sg13g2_decap_8 FILLER_102_952 ();
 sg13g2_decap_8 FILLER_102_959 ();
 sg13g2_decap_8 FILLER_102_966 ();
 sg13g2_decap_8 FILLER_102_973 ();
 sg13g2_decap_8 FILLER_102_980 ();
 sg13g2_decap_8 FILLER_102_987 ();
 sg13g2_decap_8 FILLER_102_994 ();
 sg13g2_decap_8 FILLER_102_1001 ();
 sg13g2_decap_8 FILLER_102_1008 ();
 sg13g2_decap_8 FILLER_102_1015 ();
 sg13g2_decap_8 FILLER_102_1022 ();
 sg13g2_decap_8 FILLER_103_0 ();
 sg13g2_decap_8 FILLER_103_7 ();
 sg13g2_decap_8 FILLER_103_14 ();
 sg13g2_decap_8 FILLER_103_21 ();
 sg13g2_decap_8 FILLER_103_28 ();
 sg13g2_decap_8 FILLER_103_35 ();
 sg13g2_decap_8 FILLER_103_42 ();
 sg13g2_decap_8 FILLER_103_49 ();
 sg13g2_decap_8 FILLER_103_56 ();
 sg13g2_decap_8 FILLER_103_63 ();
 sg13g2_decap_8 FILLER_103_70 ();
 sg13g2_decap_8 FILLER_103_77 ();
 sg13g2_decap_8 FILLER_103_84 ();
 sg13g2_decap_8 FILLER_103_91 ();
 sg13g2_decap_8 FILLER_103_98 ();
 sg13g2_decap_8 FILLER_103_105 ();
 sg13g2_decap_8 FILLER_103_112 ();
 sg13g2_decap_8 FILLER_103_119 ();
 sg13g2_decap_8 FILLER_103_126 ();
 sg13g2_decap_8 FILLER_103_133 ();
 sg13g2_decap_8 FILLER_103_140 ();
 sg13g2_decap_8 FILLER_103_147 ();
 sg13g2_decap_8 FILLER_103_154 ();
 sg13g2_decap_8 FILLER_103_161 ();
 sg13g2_decap_8 FILLER_103_168 ();
 sg13g2_decap_8 FILLER_103_175 ();
 sg13g2_decap_8 FILLER_103_182 ();
 sg13g2_decap_8 FILLER_103_189 ();
 sg13g2_decap_8 FILLER_103_196 ();
 sg13g2_decap_8 FILLER_103_203 ();
 sg13g2_decap_8 FILLER_103_210 ();
 sg13g2_decap_8 FILLER_103_217 ();
 sg13g2_decap_8 FILLER_103_224 ();
 sg13g2_decap_8 FILLER_103_231 ();
 sg13g2_decap_8 FILLER_103_238 ();
 sg13g2_decap_8 FILLER_103_245 ();
 sg13g2_decap_8 FILLER_103_252 ();
 sg13g2_decap_8 FILLER_103_259 ();
 sg13g2_decap_8 FILLER_103_266 ();
 sg13g2_decap_8 FILLER_103_273 ();
 sg13g2_decap_8 FILLER_103_280 ();
 sg13g2_decap_8 FILLER_103_287 ();
 sg13g2_decap_8 FILLER_103_294 ();
 sg13g2_decap_8 FILLER_103_301 ();
 sg13g2_decap_8 FILLER_103_308 ();
 sg13g2_decap_8 FILLER_103_315 ();
 sg13g2_decap_8 FILLER_103_322 ();
 sg13g2_decap_8 FILLER_103_329 ();
 sg13g2_decap_8 FILLER_103_336 ();
 sg13g2_decap_8 FILLER_103_343 ();
 sg13g2_decap_8 FILLER_103_350 ();
 sg13g2_decap_8 FILLER_103_357 ();
 sg13g2_decap_8 FILLER_103_364 ();
 sg13g2_decap_8 FILLER_103_371 ();
 sg13g2_decap_8 FILLER_103_378 ();
 sg13g2_decap_8 FILLER_103_385 ();
 sg13g2_decap_8 FILLER_103_392 ();
 sg13g2_decap_8 FILLER_103_399 ();
 sg13g2_decap_8 FILLER_103_406 ();
 sg13g2_decap_8 FILLER_103_413 ();
 sg13g2_decap_8 FILLER_103_420 ();
 sg13g2_decap_8 FILLER_103_427 ();
 sg13g2_decap_8 FILLER_103_434 ();
 sg13g2_decap_8 FILLER_103_441 ();
 sg13g2_decap_8 FILLER_103_448 ();
 sg13g2_decap_8 FILLER_103_455 ();
 sg13g2_decap_8 FILLER_103_462 ();
 sg13g2_decap_8 FILLER_103_469 ();
 sg13g2_decap_8 FILLER_103_476 ();
 sg13g2_decap_8 FILLER_103_483 ();
 sg13g2_decap_8 FILLER_103_490 ();
 sg13g2_decap_8 FILLER_103_497 ();
 sg13g2_decap_8 FILLER_103_504 ();
 sg13g2_decap_8 FILLER_103_511 ();
 sg13g2_decap_8 FILLER_103_518 ();
 sg13g2_decap_8 FILLER_103_525 ();
 sg13g2_decap_8 FILLER_103_532 ();
 sg13g2_decap_8 FILLER_103_539 ();
 sg13g2_decap_8 FILLER_103_546 ();
 sg13g2_decap_8 FILLER_103_553 ();
 sg13g2_decap_8 FILLER_103_560 ();
 sg13g2_decap_8 FILLER_103_567 ();
 sg13g2_decap_8 FILLER_103_574 ();
 sg13g2_decap_8 FILLER_103_581 ();
 sg13g2_decap_8 FILLER_103_588 ();
 sg13g2_decap_8 FILLER_103_595 ();
 sg13g2_decap_8 FILLER_103_602 ();
 sg13g2_decap_8 FILLER_103_609 ();
 sg13g2_decap_8 FILLER_103_616 ();
 sg13g2_decap_8 FILLER_103_623 ();
 sg13g2_decap_8 FILLER_103_630 ();
 sg13g2_decap_8 FILLER_103_637 ();
 sg13g2_decap_8 FILLER_103_644 ();
 sg13g2_decap_8 FILLER_103_651 ();
 sg13g2_decap_8 FILLER_103_658 ();
 sg13g2_decap_8 FILLER_103_665 ();
 sg13g2_decap_8 FILLER_103_672 ();
 sg13g2_decap_8 FILLER_103_679 ();
 sg13g2_decap_8 FILLER_103_686 ();
 sg13g2_decap_8 FILLER_103_693 ();
 sg13g2_decap_8 FILLER_103_700 ();
 sg13g2_decap_8 FILLER_103_707 ();
 sg13g2_decap_8 FILLER_103_714 ();
 sg13g2_decap_8 FILLER_103_721 ();
 sg13g2_decap_8 FILLER_103_728 ();
 sg13g2_decap_8 FILLER_103_735 ();
 sg13g2_decap_8 FILLER_103_742 ();
 sg13g2_decap_8 FILLER_103_749 ();
 sg13g2_decap_8 FILLER_103_756 ();
 sg13g2_decap_8 FILLER_103_763 ();
 sg13g2_decap_8 FILLER_103_770 ();
 sg13g2_decap_8 FILLER_103_777 ();
 sg13g2_decap_8 FILLER_103_784 ();
 sg13g2_decap_8 FILLER_103_791 ();
 sg13g2_decap_8 FILLER_103_798 ();
 sg13g2_decap_8 FILLER_103_805 ();
 sg13g2_decap_8 FILLER_103_812 ();
 sg13g2_decap_8 FILLER_103_819 ();
 sg13g2_decap_8 FILLER_103_826 ();
 sg13g2_decap_8 FILLER_103_833 ();
 sg13g2_decap_8 FILLER_103_840 ();
 sg13g2_decap_8 FILLER_103_847 ();
 sg13g2_decap_8 FILLER_103_854 ();
 sg13g2_decap_8 FILLER_103_861 ();
 sg13g2_decap_8 FILLER_103_868 ();
 sg13g2_decap_8 FILLER_103_875 ();
 sg13g2_decap_8 FILLER_103_882 ();
 sg13g2_decap_8 FILLER_103_889 ();
 sg13g2_decap_8 FILLER_103_896 ();
 sg13g2_decap_8 FILLER_103_903 ();
 sg13g2_decap_8 FILLER_103_910 ();
 sg13g2_decap_8 FILLER_103_917 ();
 sg13g2_decap_8 FILLER_103_924 ();
 sg13g2_decap_8 FILLER_103_931 ();
 sg13g2_decap_8 FILLER_103_938 ();
 sg13g2_decap_8 FILLER_103_945 ();
 sg13g2_decap_8 FILLER_103_952 ();
 sg13g2_decap_8 FILLER_103_959 ();
 sg13g2_decap_8 FILLER_103_966 ();
 sg13g2_decap_8 FILLER_103_973 ();
 sg13g2_decap_8 FILLER_103_980 ();
 sg13g2_decap_8 FILLER_103_987 ();
 sg13g2_decap_8 FILLER_103_994 ();
 sg13g2_decap_8 FILLER_103_1001 ();
 sg13g2_decap_8 FILLER_103_1008 ();
 sg13g2_decap_8 FILLER_103_1015 ();
 sg13g2_decap_8 FILLER_103_1022 ();
 sg13g2_decap_8 FILLER_104_0 ();
 sg13g2_decap_8 FILLER_104_7 ();
 sg13g2_decap_8 FILLER_104_14 ();
 sg13g2_decap_8 FILLER_104_21 ();
 sg13g2_decap_8 FILLER_104_28 ();
 sg13g2_decap_8 FILLER_104_35 ();
 sg13g2_decap_8 FILLER_104_42 ();
 sg13g2_decap_8 FILLER_104_49 ();
 sg13g2_decap_8 FILLER_104_56 ();
 sg13g2_decap_8 FILLER_104_63 ();
 sg13g2_decap_8 FILLER_104_70 ();
 sg13g2_decap_8 FILLER_104_77 ();
 sg13g2_decap_8 FILLER_104_84 ();
 sg13g2_decap_8 FILLER_104_91 ();
 sg13g2_decap_8 FILLER_104_98 ();
 sg13g2_decap_8 FILLER_104_105 ();
 sg13g2_decap_8 FILLER_104_112 ();
 sg13g2_decap_8 FILLER_104_119 ();
 sg13g2_decap_8 FILLER_104_126 ();
 sg13g2_decap_8 FILLER_104_133 ();
 sg13g2_decap_8 FILLER_104_140 ();
 sg13g2_decap_8 FILLER_104_147 ();
 sg13g2_decap_8 FILLER_104_154 ();
 sg13g2_decap_8 FILLER_104_161 ();
 sg13g2_decap_8 FILLER_104_168 ();
 sg13g2_decap_8 FILLER_104_175 ();
 sg13g2_decap_8 FILLER_104_182 ();
 sg13g2_decap_8 FILLER_104_189 ();
 sg13g2_decap_8 FILLER_104_196 ();
 sg13g2_decap_8 FILLER_104_203 ();
 sg13g2_decap_8 FILLER_104_210 ();
 sg13g2_decap_8 FILLER_104_217 ();
 sg13g2_decap_8 FILLER_104_224 ();
 sg13g2_decap_8 FILLER_104_231 ();
 sg13g2_decap_8 FILLER_104_238 ();
 sg13g2_decap_8 FILLER_104_245 ();
 sg13g2_decap_8 FILLER_104_252 ();
 sg13g2_decap_8 FILLER_104_259 ();
 sg13g2_decap_8 FILLER_104_266 ();
 sg13g2_decap_8 FILLER_104_273 ();
 sg13g2_decap_8 FILLER_104_280 ();
 sg13g2_decap_8 FILLER_104_287 ();
 sg13g2_decap_8 FILLER_104_294 ();
 sg13g2_decap_8 FILLER_104_301 ();
 sg13g2_decap_8 FILLER_104_308 ();
 sg13g2_decap_8 FILLER_104_315 ();
 sg13g2_decap_8 FILLER_104_322 ();
 sg13g2_decap_8 FILLER_104_329 ();
 sg13g2_decap_8 FILLER_104_336 ();
 sg13g2_decap_8 FILLER_104_343 ();
 sg13g2_decap_8 FILLER_104_350 ();
 sg13g2_decap_8 FILLER_104_357 ();
 sg13g2_decap_8 FILLER_104_364 ();
 sg13g2_decap_8 FILLER_104_371 ();
 sg13g2_decap_8 FILLER_104_378 ();
 sg13g2_decap_8 FILLER_104_385 ();
 sg13g2_decap_8 FILLER_104_392 ();
 sg13g2_decap_8 FILLER_104_399 ();
 sg13g2_decap_8 FILLER_104_406 ();
 sg13g2_decap_8 FILLER_104_413 ();
 sg13g2_decap_8 FILLER_104_420 ();
 sg13g2_decap_8 FILLER_104_427 ();
 sg13g2_decap_8 FILLER_104_434 ();
 sg13g2_decap_8 FILLER_104_441 ();
 sg13g2_decap_8 FILLER_104_448 ();
 sg13g2_decap_8 FILLER_104_455 ();
 sg13g2_decap_8 FILLER_104_462 ();
 sg13g2_decap_8 FILLER_104_469 ();
 sg13g2_decap_8 FILLER_104_476 ();
 sg13g2_decap_8 FILLER_104_483 ();
 sg13g2_decap_8 FILLER_104_490 ();
 sg13g2_decap_8 FILLER_104_497 ();
 sg13g2_decap_8 FILLER_104_504 ();
 sg13g2_decap_8 FILLER_104_511 ();
 sg13g2_decap_8 FILLER_104_518 ();
 sg13g2_decap_8 FILLER_104_525 ();
 sg13g2_decap_8 FILLER_104_532 ();
 sg13g2_decap_8 FILLER_104_539 ();
 sg13g2_decap_8 FILLER_104_546 ();
 sg13g2_decap_8 FILLER_104_553 ();
 sg13g2_decap_8 FILLER_104_560 ();
 sg13g2_decap_8 FILLER_104_567 ();
 sg13g2_decap_8 FILLER_104_574 ();
 sg13g2_decap_8 FILLER_104_581 ();
 sg13g2_decap_8 FILLER_104_588 ();
 sg13g2_decap_8 FILLER_104_595 ();
 sg13g2_decap_8 FILLER_104_602 ();
 sg13g2_decap_8 FILLER_104_609 ();
 sg13g2_decap_8 FILLER_104_616 ();
 sg13g2_decap_8 FILLER_104_623 ();
 sg13g2_decap_8 FILLER_104_630 ();
 sg13g2_decap_8 FILLER_104_637 ();
 sg13g2_decap_8 FILLER_104_644 ();
 sg13g2_decap_8 FILLER_104_651 ();
 sg13g2_decap_8 FILLER_104_658 ();
 sg13g2_decap_8 FILLER_104_665 ();
 sg13g2_decap_8 FILLER_104_672 ();
 sg13g2_decap_8 FILLER_104_679 ();
 sg13g2_decap_8 FILLER_104_686 ();
 sg13g2_decap_8 FILLER_104_693 ();
 sg13g2_decap_8 FILLER_104_700 ();
 sg13g2_decap_8 FILLER_104_707 ();
 sg13g2_decap_8 FILLER_104_714 ();
 sg13g2_decap_8 FILLER_104_721 ();
 sg13g2_decap_8 FILLER_104_728 ();
 sg13g2_decap_8 FILLER_104_735 ();
 sg13g2_decap_8 FILLER_104_742 ();
 sg13g2_decap_8 FILLER_104_749 ();
 sg13g2_decap_8 FILLER_104_756 ();
 sg13g2_decap_8 FILLER_104_763 ();
 sg13g2_decap_8 FILLER_104_770 ();
 sg13g2_decap_8 FILLER_104_777 ();
 sg13g2_decap_8 FILLER_104_784 ();
 sg13g2_decap_8 FILLER_104_791 ();
 sg13g2_decap_8 FILLER_104_798 ();
 sg13g2_decap_8 FILLER_104_805 ();
 sg13g2_decap_8 FILLER_104_812 ();
 sg13g2_decap_8 FILLER_104_819 ();
 sg13g2_decap_8 FILLER_104_826 ();
 sg13g2_decap_8 FILLER_104_833 ();
 sg13g2_decap_8 FILLER_104_840 ();
 sg13g2_decap_8 FILLER_104_847 ();
 sg13g2_decap_8 FILLER_104_854 ();
 sg13g2_decap_8 FILLER_104_861 ();
 sg13g2_decap_8 FILLER_104_868 ();
 sg13g2_decap_8 FILLER_104_875 ();
 sg13g2_decap_8 FILLER_104_882 ();
 sg13g2_decap_8 FILLER_104_889 ();
 sg13g2_decap_8 FILLER_104_896 ();
 sg13g2_decap_8 FILLER_104_903 ();
 sg13g2_decap_8 FILLER_104_910 ();
 sg13g2_decap_8 FILLER_104_917 ();
 sg13g2_decap_8 FILLER_104_924 ();
 sg13g2_decap_8 FILLER_104_931 ();
 sg13g2_decap_8 FILLER_104_938 ();
 sg13g2_decap_8 FILLER_104_945 ();
 sg13g2_decap_8 FILLER_104_952 ();
 sg13g2_decap_8 FILLER_104_959 ();
 sg13g2_decap_8 FILLER_104_966 ();
 sg13g2_decap_8 FILLER_104_973 ();
 sg13g2_decap_8 FILLER_104_980 ();
 sg13g2_decap_8 FILLER_104_987 ();
 sg13g2_decap_8 FILLER_104_994 ();
 sg13g2_decap_8 FILLER_104_1001 ();
 sg13g2_decap_8 FILLER_104_1008 ();
 sg13g2_decap_8 FILLER_104_1015 ();
 sg13g2_decap_8 FILLER_104_1022 ();
 sg13g2_decap_8 FILLER_105_0 ();
 sg13g2_decap_8 FILLER_105_7 ();
 sg13g2_decap_8 FILLER_105_14 ();
 sg13g2_decap_8 FILLER_105_21 ();
 sg13g2_decap_8 FILLER_105_28 ();
 sg13g2_decap_8 FILLER_105_35 ();
 sg13g2_decap_8 FILLER_105_42 ();
 sg13g2_decap_8 FILLER_105_49 ();
 sg13g2_decap_8 FILLER_105_56 ();
 sg13g2_decap_8 FILLER_105_63 ();
 sg13g2_decap_8 FILLER_105_70 ();
 sg13g2_decap_8 FILLER_105_77 ();
 sg13g2_decap_8 FILLER_105_84 ();
 sg13g2_decap_8 FILLER_105_91 ();
 sg13g2_decap_8 FILLER_105_98 ();
 sg13g2_decap_8 FILLER_105_105 ();
 sg13g2_decap_8 FILLER_105_112 ();
 sg13g2_decap_8 FILLER_105_119 ();
 sg13g2_decap_8 FILLER_105_126 ();
 sg13g2_decap_8 FILLER_105_133 ();
 sg13g2_decap_8 FILLER_105_140 ();
 sg13g2_decap_8 FILLER_105_147 ();
 sg13g2_decap_8 FILLER_105_154 ();
 sg13g2_decap_8 FILLER_105_161 ();
 sg13g2_decap_8 FILLER_105_168 ();
 sg13g2_decap_8 FILLER_105_175 ();
 sg13g2_decap_8 FILLER_105_182 ();
 sg13g2_decap_8 FILLER_105_189 ();
 sg13g2_decap_8 FILLER_105_196 ();
 sg13g2_decap_8 FILLER_105_203 ();
 sg13g2_decap_8 FILLER_105_210 ();
 sg13g2_decap_8 FILLER_105_217 ();
 sg13g2_decap_8 FILLER_105_224 ();
 sg13g2_decap_8 FILLER_105_231 ();
 sg13g2_decap_8 FILLER_105_238 ();
 sg13g2_decap_8 FILLER_105_245 ();
 sg13g2_decap_8 FILLER_105_252 ();
 sg13g2_decap_8 FILLER_105_259 ();
 sg13g2_decap_8 FILLER_105_266 ();
 sg13g2_decap_8 FILLER_105_273 ();
 sg13g2_decap_8 FILLER_105_280 ();
 sg13g2_decap_8 FILLER_105_287 ();
 sg13g2_decap_8 FILLER_105_294 ();
 sg13g2_decap_8 FILLER_105_301 ();
 sg13g2_decap_8 FILLER_105_308 ();
 sg13g2_decap_8 FILLER_105_315 ();
 sg13g2_decap_8 FILLER_105_322 ();
 sg13g2_decap_8 FILLER_105_329 ();
 sg13g2_decap_8 FILLER_105_336 ();
 sg13g2_decap_8 FILLER_105_343 ();
 sg13g2_decap_8 FILLER_105_350 ();
 sg13g2_decap_8 FILLER_105_357 ();
 sg13g2_decap_8 FILLER_105_364 ();
 sg13g2_decap_8 FILLER_105_371 ();
 sg13g2_decap_8 FILLER_105_378 ();
 sg13g2_decap_8 FILLER_105_385 ();
 sg13g2_decap_8 FILLER_105_392 ();
 sg13g2_decap_8 FILLER_105_399 ();
 sg13g2_decap_8 FILLER_105_406 ();
 sg13g2_decap_8 FILLER_105_413 ();
 sg13g2_decap_8 FILLER_105_420 ();
 sg13g2_decap_8 FILLER_105_427 ();
 sg13g2_decap_8 FILLER_105_434 ();
 sg13g2_decap_8 FILLER_105_441 ();
 sg13g2_decap_8 FILLER_105_448 ();
 sg13g2_decap_8 FILLER_105_455 ();
 sg13g2_decap_8 FILLER_105_462 ();
 sg13g2_decap_8 FILLER_105_469 ();
 sg13g2_decap_8 FILLER_105_476 ();
 sg13g2_decap_8 FILLER_105_483 ();
 sg13g2_decap_8 FILLER_105_490 ();
 sg13g2_decap_8 FILLER_105_497 ();
 sg13g2_decap_8 FILLER_105_504 ();
 sg13g2_decap_8 FILLER_105_511 ();
 sg13g2_decap_8 FILLER_105_518 ();
 sg13g2_decap_8 FILLER_105_525 ();
 sg13g2_decap_8 FILLER_105_532 ();
 sg13g2_decap_8 FILLER_105_539 ();
 sg13g2_decap_8 FILLER_105_546 ();
 sg13g2_decap_8 FILLER_105_553 ();
 sg13g2_decap_8 FILLER_105_560 ();
 sg13g2_decap_8 FILLER_105_567 ();
 sg13g2_decap_8 FILLER_105_574 ();
 sg13g2_decap_8 FILLER_105_581 ();
 sg13g2_decap_8 FILLER_105_588 ();
 sg13g2_decap_8 FILLER_105_595 ();
 sg13g2_decap_8 FILLER_105_602 ();
 sg13g2_decap_8 FILLER_105_609 ();
 sg13g2_decap_8 FILLER_105_616 ();
 sg13g2_decap_8 FILLER_105_623 ();
 sg13g2_decap_8 FILLER_105_630 ();
 sg13g2_decap_8 FILLER_105_637 ();
 sg13g2_decap_8 FILLER_105_644 ();
 sg13g2_decap_8 FILLER_105_651 ();
 sg13g2_decap_8 FILLER_105_658 ();
 sg13g2_decap_8 FILLER_105_665 ();
 sg13g2_decap_8 FILLER_105_672 ();
 sg13g2_decap_8 FILLER_105_679 ();
 sg13g2_decap_8 FILLER_105_686 ();
 sg13g2_decap_8 FILLER_105_693 ();
 sg13g2_decap_8 FILLER_105_700 ();
 sg13g2_decap_8 FILLER_105_707 ();
 sg13g2_decap_8 FILLER_105_714 ();
 sg13g2_decap_8 FILLER_105_721 ();
 sg13g2_decap_8 FILLER_105_728 ();
 sg13g2_decap_8 FILLER_105_735 ();
 sg13g2_decap_8 FILLER_105_742 ();
 sg13g2_decap_8 FILLER_105_749 ();
 sg13g2_decap_8 FILLER_105_756 ();
 sg13g2_decap_8 FILLER_105_763 ();
 sg13g2_decap_8 FILLER_105_770 ();
 sg13g2_decap_8 FILLER_105_777 ();
 sg13g2_decap_8 FILLER_105_784 ();
 sg13g2_decap_8 FILLER_105_791 ();
 sg13g2_decap_8 FILLER_105_798 ();
 sg13g2_decap_8 FILLER_105_805 ();
 sg13g2_decap_8 FILLER_105_812 ();
 sg13g2_decap_8 FILLER_105_819 ();
 sg13g2_decap_8 FILLER_105_826 ();
 sg13g2_decap_8 FILLER_105_833 ();
 sg13g2_decap_8 FILLER_105_840 ();
 sg13g2_decap_8 FILLER_105_847 ();
 sg13g2_decap_8 FILLER_105_854 ();
 sg13g2_decap_8 FILLER_105_861 ();
 sg13g2_decap_8 FILLER_105_868 ();
 sg13g2_decap_8 FILLER_105_875 ();
 sg13g2_decap_8 FILLER_105_882 ();
 sg13g2_decap_8 FILLER_105_889 ();
 sg13g2_decap_8 FILLER_105_896 ();
 sg13g2_decap_8 FILLER_105_903 ();
 sg13g2_decap_8 FILLER_105_910 ();
 sg13g2_decap_8 FILLER_105_917 ();
 sg13g2_decap_8 FILLER_105_924 ();
 sg13g2_decap_8 FILLER_105_931 ();
 sg13g2_decap_8 FILLER_105_938 ();
 sg13g2_decap_8 FILLER_105_945 ();
 sg13g2_decap_8 FILLER_105_952 ();
 sg13g2_decap_8 FILLER_105_959 ();
 sg13g2_decap_8 FILLER_105_966 ();
 sg13g2_decap_8 FILLER_105_973 ();
 sg13g2_decap_8 FILLER_105_980 ();
 sg13g2_decap_8 FILLER_105_987 ();
 sg13g2_decap_8 FILLER_105_994 ();
 sg13g2_decap_8 FILLER_105_1001 ();
 sg13g2_decap_8 FILLER_105_1008 ();
 sg13g2_decap_8 FILLER_105_1015 ();
 sg13g2_decap_8 FILLER_105_1022 ();
 sg13g2_decap_8 FILLER_106_0 ();
 sg13g2_decap_8 FILLER_106_7 ();
 sg13g2_decap_8 FILLER_106_14 ();
 sg13g2_decap_8 FILLER_106_21 ();
 sg13g2_decap_8 FILLER_106_28 ();
 sg13g2_decap_8 FILLER_106_35 ();
 sg13g2_decap_8 FILLER_106_42 ();
 sg13g2_decap_8 FILLER_106_49 ();
 sg13g2_decap_8 FILLER_106_56 ();
 sg13g2_decap_8 FILLER_106_63 ();
 sg13g2_decap_8 FILLER_106_70 ();
 sg13g2_decap_8 FILLER_106_77 ();
 sg13g2_decap_8 FILLER_106_84 ();
 sg13g2_decap_8 FILLER_106_91 ();
 sg13g2_decap_8 FILLER_106_98 ();
 sg13g2_decap_8 FILLER_106_105 ();
 sg13g2_decap_8 FILLER_106_112 ();
 sg13g2_decap_8 FILLER_106_119 ();
 sg13g2_decap_8 FILLER_106_126 ();
 sg13g2_decap_8 FILLER_106_133 ();
 sg13g2_decap_8 FILLER_106_140 ();
 sg13g2_decap_8 FILLER_106_147 ();
 sg13g2_decap_8 FILLER_106_154 ();
 sg13g2_decap_8 FILLER_106_161 ();
 sg13g2_decap_8 FILLER_106_168 ();
 sg13g2_decap_8 FILLER_106_175 ();
 sg13g2_decap_8 FILLER_106_182 ();
 sg13g2_decap_8 FILLER_106_189 ();
 sg13g2_decap_8 FILLER_106_196 ();
 sg13g2_decap_8 FILLER_106_203 ();
 sg13g2_decap_8 FILLER_106_210 ();
 sg13g2_decap_8 FILLER_106_217 ();
 sg13g2_decap_8 FILLER_106_224 ();
 sg13g2_decap_8 FILLER_106_231 ();
 sg13g2_decap_8 FILLER_106_238 ();
 sg13g2_decap_8 FILLER_106_245 ();
 sg13g2_decap_8 FILLER_106_252 ();
 sg13g2_decap_8 FILLER_106_259 ();
 sg13g2_decap_8 FILLER_106_266 ();
 sg13g2_decap_8 FILLER_106_273 ();
 sg13g2_decap_8 FILLER_106_280 ();
 sg13g2_decap_8 FILLER_106_287 ();
 sg13g2_decap_8 FILLER_106_294 ();
 sg13g2_decap_8 FILLER_106_301 ();
 sg13g2_decap_8 FILLER_106_308 ();
 sg13g2_decap_8 FILLER_106_315 ();
 sg13g2_decap_8 FILLER_106_322 ();
 sg13g2_decap_8 FILLER_106_329 ();
 sg13g2_decap_8 FILLER_106_336 ();
 sg13g2_decap_8 FILLER_106_343 ();
 sg13g2_decap_8 FILLER_106_350 ();
 sg13g2_decap_8 FILLER_106_357 ();
 sg13g2_decap_8 FILLER_106_364 ();
 sg13g2_decap_8 FILLER_106_371 ();
 sg13g2_decap_8 FILLER_106_378 ();
 sg13g2_decap_8 FILLER_106_385 ();
 sg13g2_decap_8 FILLER_106_392 ();
 sg13g2_decap_8 FILLER_106_399 ();
 sg13g2_decap_8 FILLER_106_406 ();
 sg13g2_decap_8 FILLER_106_413 ();
 sg13g2_decap_8 FILLER_106_420 ();
 sg13g2_decap_8 FILLER_106_427 ();
 sg13g2_decap_8 FILLER_106_434 ();
 sg13g2_decap_8 FILLER_106_441 ();
 sg13g2_decap_8 FILLER_106_448 ();
 sg13g2_decap_8 FILLER_106_455 ();
 sg13g2_decap_8 FILLER_106_462 ();
 sg13g2_decap_8 FILLER_106_469 ();
 sg13g2_decap_8 FILLER_106_476 ();
 sg13g2_decap_8 FILLER_106_483 ();
 sg13g2_decap_8 FILLER_106_490 ();
 sg13g2_decap_8 FILLER_106_497 ();
 sg13g2_decap_8 FILLER_106_504 ();
 sg13g2_decap_8 FILLER_106_511 ();
 sg13g2_decap_8 FILLER_106_518 ();
 sg13g2_decap_8 FILLER_106_525 ();
 sg13g2_decap_8 FILLER_106_532 ();
 sg13g2_decap_8 FILLER_106_539 ();
 sg13g2_decap_8 FILLER_106_546 ();
 sg13g2_decap_8 FILLER_106_553 ();
 sg13g2_decap_8 FILLER_106_560 ();
 sg13g2_decap_8 FILLER_106_567 ();
 sg13g2_decap_8 FILLER_106_574 ();
 sg13g2_decap_8 FILLER_106_581 ();
 sg13g2_decap_8 FILLER_106_588 ();
 sg13g2_decap_8 FILLER_106_595 ();
 sg13g2_decap_8 FILLER_106_602 ();
 sg13g2_decap_8 FILLER_106_609 ();
 sg13g2_decap_8 FILLER_106_616 ();
 sg13g2_decap_8 FILLER_106_623 ();
 sg13g2_decap_8 FILLER_106_630 ();
 sg13g2_decap_8 FILLER_106_637 ();
 sg13g2_decap_8 FILLER_106_644 ();
 sg13g2_decap_8 FILLER_106_651 ();
 sg13g2_decap_8 FILLER_106_658 ();
 sg13g2_decap_8 FILLER_106_665 ();
 sg13g2_decap_8 FILLER_106_672 ();
 sg13g2_decap_8 FILLER_106_679 ();
 sg13g2_decap_8 FILLER_106_686 ();
 sg13g2_decap_8 FILLER_106_693 ();
 sg13g2_decap_8 FILLER_106_700 ();
 sg13g2_decap_8 FILLER_106_707 ();
 sg13g2_decap_8 FILLER_106_714 ();
 sg13g2_decap_8 FILLER_106_721 ();
 sg13g2_decap_8 FILLER_106_728 ();
 sg13g2_decap_8 FILLER_106_735 ();
 sg13g2_decap_8 FILLER_106_742 ();
 sg13g2_decap_8 FILLER_106_749 ();
 sg13g2_decap_8 FILLER_106_756 ();
 sg13g2_decap_8 FILLER_106_763 ();
 sg13g2_decap_8 FILLER_106_770 ();
 sg13g2_decap_8 FILLER_106_777 ();
 sg13g2_decap_8 FILLER_106_784 ();
 sg13g2_decap_8 FILLER_106_791 ();
 sg13g2_decap_8 FILLER_106_798 ();
 sg13g2_decap_8 FILLER_106_805 ();
 sg13g2_decap_8 FILLER_106_812 ();
 sg13g2_decap_8 FILLER_106_819 ();
 sg13g2_decap_8 FILLER_106_826 ();
 sg13g2_decap_8 FILLER_106_833 ();
 sg13g2_decap_8 FILLER_106_840 ();
 sg13g2_decap_8 FILLER_106_847 ();
 sg13g2_decap_8 FILLER_106_854 ();
 sg13g2_decap_8 FILLER_106_861 ();
 sg13g2_decap_8 FILLER_106_868 ();
 sg13g2_decap_8 FILLER_106_875 ();
 sg13g2_decap_8 FILLER_106_882 ();
 sg13g2_decap_8 FILLER_106_889 ();
 sg13g2_decap_8 FILLER_106_896 ();
 sg13g2_decap_8 FILLER_106_903 ();
 sg13g2_decap_8 FILLER_106_910 ();
 sg13g2_decap_8 FILLER_106_917 ();
 sg13g2_decap_8 FILLER_106_924 ();
 sg13g2_decap_8 FILLER_106_931 ();
 sg13g2_decap_8 FILLER_106_938 ();
 sg13g2_decap_8 FILLER_106_945 ();
 sg13g2_decap_8 FILLER_106_952 ();
 sg13g2_decap_8 FILLER_106_959 ();
 sg13g2_decap_8 FILLER_106_966 ();
 sg13g2_decap_8 FILLER_106_973 ();
 sg13g2_decap_8 FILLER_106_980 ();
 sg13g2_decap_8 FILLER_106_987 ();
 sg13g2_decap_8 FILLER_106_994 ();
 sg13g2_decap_8 FILLER_106_1001 ();
 sg13g2_decap_8 FILLER_106_1008 ();
 sg13g2_decap_8 FILLER_106_1015 ();
 sg13g2_decap_8 FILLER_106_1022 ();
 assign uio_oe[0] = net25;
 assign uio_oe[1] = net26;
 assign uio_oe[2] = net27;
 assign uio_oe[3] = net28;
 assign uio_oe[4] = net29;
 assign uio_oe[5] = net30;
 assign uio_oe[6] = net31;
 assign uio_oe[7] = net32;
 assign uio_out[0] = net33;
 assign uio_out[1] = net34;
 assign uio_out[2] = net35;
 assign uio_out[3] = net36;
 assign uio_out[4] = net37;
 assign uio_out[5] = net38;
 assign uio_out[6] = net39;
 assign uio_out[7] = net40;
endmodule
