magic
tech ihp-sg13g2
magscale 1 2
timestamp 1754573650
<< metal1 >>
rect 1152 41600 20452 41624
rect 1152 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20452 41600
rect 1152 41536 20452 41560
rect 19467 41432 19509 41441
rect 19467 41392 19468 41432
rect 19508 41392 19509 41432
rect 19467 41383 19509 41392
rect 19851 41432 19893 41441
rect 19851 41392 19852 41432
rect 19892 41392 19893 41432
rect 19851 41383 19893 41392
rect 1603 41264 1661 41265
rect 1603 41224 1612 41264
rect 1652 41224 1661 41264
rect 1603 41223 1661 41224
rect 2851 41264 2909 41265
rect 2851 41224 2860 41264
rect 2900 41224 2909 41264
rect 2851 41223 2909 41224
rect 3235 41264 3293 41265
rect 3235 41224 3244 41264
rect 3284 41224 3293 41264
rect 3235 41223 3293 41224
rect 4483 41264 4541 41265
rect 4483 41224 4492 41264
rect 4532 41224 4541 41264
rect 4483 41223 4541 41224
rect 4963 41264 5021 41265
rect 4963 41224 4972 41264
rect 5012 41224 5021 41264
rect 4963 41223 5021 41224
rect 5067 41264 5109 41273
rect 5067 41224 5068 41264
rect 5108 41224 5109 41264
rect 5067 41215 5109 41224
rect 5259 41264 5301 41273
rect 5259 41224 5260 41264
rect 5300 41224 5301 41264
rect 5259 41215 5301 41224
rect 5635 41264 5693 41265
rect 5635 41224 5644 41264
rect 5684 41224 5693 41264
rect 5635 41223 5693 41224
rect 6883 41264 6941 41265
rect 6883 41224 6892 41264
rect 6932 41224 6941 41264
rect 6883 41223 6941 41224
rect 7075 41264 7133 41265
rect 7075 41224 7084 41264
rect 7124 41224 7133 41264
rect 7075 41223 7133 41224
rect 8323 41264 8381 41265
rect 8323 41224 8332 41264
rect 8372 41224 8381 41264
rect 8323 41223 8381 41224
rect 8899 41264 8957 41265
rect 8899 41224 8908 41264
rect 8948 41224 8957 41264
rect 8899 41223 8957 41224
rect 10147 41264 10205 41265
rect 10147 41224 10156 41264
rect 10196 41224 10205 41264
rect 10147 41223 10205 41224
rect 10723 41264 10781 41265
rect 10723 41224 10732 41264
rect 10772 41224 10781 41264
rect 10723 41223 10781 41224
rect 11971 41264 12029 41265
rect 11971 41224 11980 41264
rect 12020 41224 12029 41264
rect 11971 41223 12029 41224
rect 12355 41264 12413 41265
rect 12355 41224 12364 41264
rect 12404 41224 12413 41264
rect 12355 41223 12413 41224
rect 13603 41264 13661 41265
rect 13603 41224 13612 41264
rect 13652 41224 13661 41264
rect 13603 41223 13661 41224
rect 13987 41264 14045 41265
rect 13987 41224 13996 41264
rect 14036 41224 14045 41264
rect 13987 41223 14045 41224
rect 15235 41264 15293 41265
rect 15235 41224 15244 41264
rect 15284 41224 15293 41264
rect 15235 41223 15293 41224
rect 15619 41264 15677 41265
rect 15619 41224 15628 41264
rect 15668 41224 15677 41264
rect 15619 41223 15677 41224
rect 16867 41264 16925 41265
rect 16867 41224 16876 41264
rect 16916 41224 16925 41264
rect 16867 41223 16925 41224
rect 17067 41264 17109 41273
rect 17067 41224 17068 41264
rect 17108 41224 17109 41264
rect 17067 41215 17109 41224
rect 17259 41264 17301 41273
rect 17259 41224 17260 41264
rect 17300 41224 17301 41264
rect 17259 41215 17301 41224
rect 17347 41264 17405 41265
rect 17347 41224 17356 41264
rect 17396 41224 17405 41264
rect 17347 41223 17405 41224
rect 1219 41180 1277 41181
rect 1219 41140 1228 41180
rect 1268 41140 1277 41180
rect 1219 41139 1277 41140
rect 17731 41180 17789 41181
rect 17731 41140 17740 41180
rect 17780 41140 17789 41180
rect 17731 41139 17789 41140
rect 18115 41180 18173 41181
rect 18115 41140 18124 41180
rect 18164 41140 18173 41180
rect 18115 41139 18173 41140
rect 18499 41180 18557 41181
rect 18499 41140 18508 41180
rect 18548 41140 18557 41180
rect 18499 41139 18557 41140
rect 18883 41180 18941 41181
rect 18883 41140 18892 41180
rect 18932 41140 18941 41180
rect 18883 41139 18941 41140
rect 19267 41180 19325 41181
rect 19267 41140 19276 41180
rect 19316 41140 19325 41180
rect 19267 41139 19325 41140
rect 19651 41180 19709 41181
rect 19651 41140 19660 41180
rect 19700 41140 19709 41180
rect 19651 41139 19709 41140
rect 20035 41180 20093 41181
rect 20035 41140 20044 41180
rect 20084 41140 20093 41180
rect 20035 41139 20093 41140
rect 3051 41096 3093 41105
rect 3051 41056 3052 41096
rect 3092 41056 3093 41096
rect 3051 41047 3093 41056
rect 17931 41096 17973 41105
rect 17931 41056 17932 41096
rect 17972 41056 17973 41096
rect 17931 41047 17973 41056
rect 1419 41012 1461 41021
rect 1419 40972 1420 41012
rect 1460 40972 1461 41012
rect 1419 40963 1461 40972
rect 4683 41012 4725 41021
rect 4683 40972 4684 41012
rect 4724 40972 4725 41012
rect 4683 40963 4725 40972
rect 5259 41012 5301 41021
rect 5259 40972 5260 41012
rect 5300 40972 5301 41012
rect 5259 40963 5301 40972
rect 5451 41012 5493 41021
rect 5451 40972 5452 41012
rect 5492 40972 5493 41012
rect 5451 40963 5493 40972
rect 8523 41012 8565 41021
rect 8523 40972 8524 41012
rect 8564 40972 8565 41012
rect 8523 40963 8565 40972
rect 10347 41012 10389 41021
rect 10347 40972 10348 41012
rect 10388 40972 10389 41012
rect 10347 40963 10389 40972
rect 10539 41012 10581 41021
rect 10539 40972 10540 41012
rect 10580 40972 10581 41012
rect 10539 40963 10581 40972
rect 12171 41012 12213 41021
rect 12171 40972 12172 41012
rect 12212 40972 12213 41012
rect 12171 40963 12213 40972
rect 13803 41012 13845 41021
rect 13803 40972 13804 41012
rect 13844 40972 13845 41012
rect 13803 40963 13845 40972
rect 15435 41012 15477 41021
rect 15435 40972 15436 41012
rect 15476 40972 15477 41012
rect 15435 40963 15477 40972
rect 17067 41012 17109 41021
rect 17067 40972 17068 41012
rect 17108 40972 17109 41012
rect 17067 40963 17109 40972
rect 17547 41012 17589 41021
rect 17547 40972 17548 41012
rect 17588 40972 17589 41012
rect 17547 40963 17589 40972
rect 18315 41012 18357 41021
rect 18315 40972 18316 41012
rect 18356 40972 18357 41012
rect 18315 40963 18357 40972
rect 18699 41012 18741 41021
rect 18699 40972 18700 41012
rect 18740 40972 18741 41012
rect 18699 40963 18741 40972
rect 19083 41012 19125 41021
rect 19083 40972 19084 41012
rect 19124 40972 19125 41012
rect 19083 40963 19125 40972
rect 1152 40844 20352 40868
rect 1152 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 20352 40844
rect 1152 40780 20352 40804
rect 6699 40676 6741 40685
rect 6699 40636 6700 40676
rect 6740 40636 6741 40676
rect 6699 40627 6741 40636
rect 10347 40676 10389 40685
rect 10347 40636 10348 40676
rect 10388 40636 10389 40676
rect 10347 40627 10389 40636
rect 12171 40676 12213 40685
rect 12171 40636 12172 40676
rect 12212 40636 12213 40676
rect 12171 40627 12213 40636
rect 18507 40676 18549 40685
rect 18507 40636 18508 40676
rect 18548 40636 18549 40676
rect 18507 40627 18549 40636
rect 19371 40676 19413 40685
rect 19371 40636 19372 40676
rect 19412 40636 19413 40676
rect 19371 40627 19413 40636
rect 19755 40676 19797 40685
rect 19755 40636 19756 40676
rect 19796 40636 19797 40676
rect 19755 40627 19797 40636
rect 13123 40592 13181 40593
rect 13123 40552 13132 40592
rect 13172 40552 13181 40592
rect 13123 40551 13181 40552
rect 18123 40592 18165 40601
rect 18123 40552 18124 40592
rect 18164 40552 18165 40592
rect 18123 40543 18165 40552
rect 18987 40592 19029 40601
rect 18987 40552 18988 40592
rect 19028 40552 19029 40592
rect 18987 40543 19029 40552
rect 6499 40508 6557 40509
rect 6499 40468 6508 40508
rect 6548 40468 6557 40508
rect 6499 40467 6557 40468
rect 10531 40508 10589 40509
rect 10531 40468 10540 40508
rect 10580 40468 10589 40508
rect 10531 40467 10589 40468
rect 13315 40508 13373 40509
rect 13315 40468 13324 40508
rect 13364 40468 13373 40508
rect 13315 40467 13373 40468
rect 17923 40508 17981 40509
rect 17923 40468 17932 40508
rect 17972 40468 17981 40508
rect 17923 40467 17981 40468
rect 18307 40508 18365 40509
rect 18307 40468 18316 40508
rect 18356 40468 18365 40508
rect 18307 40467 18365 40468
rect 18691 40508 18749 40509
rect 18691 40468 18700 40508
rect 18740 40468 18749 40508
rect 18691 40467 18749 40468
rect 19171 40508 19229 40509
rect 19171 40468 19180 40508
rect 19220 40468 19229 40508
rect 19171 40467 19229 40468
rect 19555 40508 19613 40509
rect 19555 40468 19564 40508
rect 19604 40468 19613 40508
rect 19555 40467 19613 40468
rect 19939 40508 19997 40509
rect 19939 40468 19948 40508
rect 19988 40468 19997 40508
rect 19939 40467 19997 40468
rect 1315 40424 1373 40425
rect 1315 40384 1324 40424
rect 1364 40384 1373 40424
rect 1315 40383 1373 40384
rect 2563 40424 2621 40425
rect 2563 40384 2572 40424
rect 2612 40384 2621 40424
rect 2563 40383 2621 40384
rect 2947 40424 3005 40425
rect 2947 40384 2956 40424
rect 2996 40384 3005 40424
rect 2947 40383 3005 40384
rect 4195 40424 4253 40425
rect 4195 40384 4204 40424
rect 4244 40384 4253 40424
rect 4195 40383 4253 40384
rect 4867 40424 4925 40425
rect 4867 40384 4876 40424
rect 4916 40384 4925 40424
rect 4867 40383 4925 40384
rect 6115 40424 6173 40425
rect 6115 40384 6124 40424
rect 6164 40384 6173 40424
rect 6115 40383 6173 40384
rect 6883 40424 6941 40425
rect 6883 40384 6892 40424
rect 6932 40384 6941 40424
rect 6883 40383 6941 40384
rect 8131 40424 8189 40425
rect 8131 40384 8140 40424
rect 8180 40384 8189 40424
rect 8131 40383 8189 40384
rect 8707 40424 8765 40425
rect 8707 40384 8716 40424
rect 8756 40384 8765 40424
rect 8707 40383 8765 40384
rect 9955 40424 10013 40425
rect 9955 40384 9964 40424
rect 10004 40384 10013 40424
rect 9955 40383 10013 40384
rect 10723 40424 10781 40425
rect 10723 40384 10732 40424
rect 10772 40384 10781 40424
rect 10723 40383 10781 40384
rect 11971 40424 12029 40425
rect 11971 40384 11980 40424
rect 12020 40384 12029 40424
rect 11971 40383 12029 40384
rect 12451 40424 12509 40425
rect 12451 40384 12460 40424
rect 12500 40384 12509 40424
rect 12451 40383 12509 40384
rect 12747 40424 12789 40433
rect 12747 40384 12748 40424
rect 12788 40384 12789 40424
rect 12747 40375 12789 40384
rect 13699 40424 13757 40425
rect 13699 40384 13708 40424
rect 13748 40384 13757 40424
rect 13699 40383 13757 40384
rect 14947 40424 15005 40425
rect 14947 40384 14956 40424
rect 14996 40384 15005 40424
rect 14947 40383 15005 40384
rect 15339 40424 15381 40433
rect 15339 40384 15340 40424
rect 15380 40384 15381 40424
rect 15339 40375 15381 40384
rect 15435 40424 15477 40433
rect 15435 40384 15436 40424
rect 15476 40384 15477 40424
rect 15435 40375 15477 40384
rect 15531 40424 15573 40433
rect 15531 40384 15532 40424
rect 15572 40384 15573 40424
rect 15531 40375 15573 40384
rect 15627 40424 15669 40433
rect 15627 40384 15628 40424
rect 15668 40384 15669 40424
rect 15627 40375 15669 40384
rect 15915 40424 15957 40433
rect 15915 40384 15916 40424
rect 15956 40384 15957 40424
rect 15915 40375 15957 40384
rect 16011 40424 16053 40433
rect 16011 40384 16012 40424
rect 16052 40384 16053 40424
rect 16395 40424 16437 40433
rect 16011 40375 16053 40384
rect 16107 40403 16149 40412
rect 16107 40363 16108 40403
rect 16148 40363 16149 40403
rect 16395 40384 16396 40424
rect 16436 40384 16437 40424
rect 16395 40375 16437 40384
rect 16491 40424 16533 40433
rect 16491 40384 16492 40424
rect 16532 40384 16533 40424
rect 16491 40375 16533 40384
rect 16587 40424 16629 40433
rect 16587 40384 16588 40424
rect 16628 40384 16629 40424
rect 16587 40375 16629 40384
rect 16875 40424 16917 40433
rect 16875 40384 16876 40424
rect 16916 40384 16917 40424
rect 16875 40375 16917 40384
rect 16971 40424 17013 40433
rect 16971 40384 16972 40424
rect 17012 40384 17013 40424
rect 16971 40375 17013 40384
rect 17067 40424 17109 40433
rect 17067 40384 17068 40424
rect 17108 40384 17109 40424
rect 17067 40375 17109 40384
rect 17259 40424 17301 40433
rect 17259 40384 17260 40424
rect 17300 40384 17301 40424
rect 17259 40375 17301 40384
rect 17451 40424 17493 40433
rect 17451 40384 17452 40424
rect 17492 40384 17493 40424
rect 17451 40375 17493 40384
rect 17539 40424 17597 40425
rect 17539 40384 17548 40424
rect 17588 40384 17597 40424
rect 17539 40383 17597 40384
rect 20227 40424 20285 40425
rect 20227 40384 20236 40424
rect 20276 40384 20285 40424
rect 20227 40383 20285 40384
rect 16107 40354 16149 40363
rect 12843 40340 12885 40349
rect 12843 40300 12844 40340
rect 12884 40300 12885 40340
rect 12843 40291 12885 40300
rect 20139 40340 20181 40349
rect 20139 40300 20140 40340
rect 20180 40300 20181 40340
rect 20139 40291 20181 40300
rect 2763 40256 2805 40265
rect 2763 40216 2764 40256
rect 2804 40216 2805 40256
rect 2763 40207 2805 40216
rect 4395 40256 4437 40265
rect 4395 40216 4396 40256
rect 4436 40216 4437 40256
rect 4395 40207 4437 40216
rect 4675 40256 4733 40257
rect 4675 40216 4684 40256
rect 4724 40216 4733 40256
rect 4675 40215 4733 40216
rect 6315 40256 6357 40265
rect 6315 40216 6316 40256
rect 6356 40216 6357 40256
rect 6315 40207 6357 40216
rect 8331 40256 8373 40265
rect 8331 40216 8332 40256
rect 8372 40216 8373 40256
rect 8331 40207 8373 40216
rect 10155 40256 10197 40265
rect 10155 40216 10156 40256
rect 10196 40216 10197 40256
rect 10155 40207 10197 40216
rect 13515 40256 13557 40265
rect 13515 40216 13516 40256
rect 13556 40216 13557 40256
rect 13515 40207 13557 40216
rect 15147 40256 15189 40265
rect 15147 40216 15148 40256
rect 15188 40216 15189 40256
rect 15147 40207 15189 40216
rect 15811 40256 15869 40257
rect 15811 40216 15820 40256
rect 15860 40216 15869 40256
rect 15811 40215 15869 40216
rect 16291 40256 16349 40257
rect 16291 40216 16300 40256
rect 16340 40216 16349 40256
rect 16291 40215 16349 40216
rect 16771 40256 16829 40257
rect 16771 40216 16780 40256
rect 16820 40216 16829 40256
rect 16771 40215 16829 40216
rect 17347 40256 17405 40257
rect 17347 40216 17356 40256
rect 17396 40216 17405 40256
rect 17347 40215 17405 40216
rect 17739 40256 17781 40265
rect 17739 40216 17740 40256
rect 17780 40216 17781 40256
rect 17739 40207 17781 40216
rect 1152 40088 20452 40112
rect 1152 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20452 40088
rect 1152 40024 20452 40048
rect 7467 39920 7509 39929
rect 7467 39880 7468 39920
rect 7508 39880 7509 39920
rect 7467 39871 7509 39880
rect 8235 39920 8277 39929
rect 8235 39880 8236 39920
rect 8276 39880 8277 39920
rect 8235 39871 8277 39880
rect 18699 39920 18741 39929
rect 18699 39880 18700 39920
rect 18740 39880 18741 39920
rect 18699 39871 18741 39880
rect 19179 39920 19221 39929
rect 19179 39880 19180 39920
rect 19220 39880 19221 39920
rect 19179 39871 19221 39880
rect 19467 39920 19509 39929
rect 19467 39880 19468 39920
rect 19508 39880 19509 39920
rect 19467 39871 19509 39880
rect 19851 39920 19893 39929
rect 19851 39880 19852 39920
rect 19892 39880 19893 39920
rect 19851 39871 19893 39880
rect 6603 39836 6645 39845
rect 6603 39796 6604 39836
rect 6644 39796 6645 39836
rect 6603 39787 6645 39796
rect 10443 39836 10485 39845
rect 10443 39796 10444 39836
rect 10484 39796 10485 39836
rect 10443 39787 10485 39796
rect 12075 39836 12117 39845
rect 12075 39796 12076 39836
rect 12116 39796 12117 39836
rect 12075 39787 12117 39796
rect 17739 39836 17781 39845
rect 17739 39796 17740 39836
rect 17780 39796 17781 39836
rect 17739 39787 17781 39796
rect 1219 39752 1277 39753
rect 1219 39712 1228 39752
rect 1268 39712 1277 39752
rect 1219 39711 1277 39712
rect 2467 39752 2525 39753
rect 2467 39712 2476 39752
rect 2516 39712 2525 39752
rect 2467 39711 2525 39712
rect 3139 39752 3197 39753
rect 3139 39712 3148 39752
rect 3188 39712 3197 39752
rect 3139 39711 3197 39712
rect 4387 39752 4445 39753
rect 4387 39712 4396 39752
rect 4436 39712 4445 39752
rect 4387 39711 4445 39712
rect 4875 39752 4917 39761
rect 4875 39712 4876 39752
rect 4916 39712 4917 39752
rect 4875 39703 4917 39712
rect 4971 39752 5013 39761
rect 4971 39712 4972 39752
rect 5012 39712 5013 39752
rect 4971 39703 5013 39712
rect 5923 39752 5981 39753
rect 5923 39712 5932 39752
rect 5972 39712 5981 39752
rect 5923 39711 5981 39712
rect 6411 39747 6453 39756
rect 6411 39707 6412 39747
rect 6452 39707 6453 39747
rect 6411 39698 6453 39707
rect 8715 39752 8757 39761
rect 8715 39712 8716 39752
rect 8756 39712 8757 39752
rect 8715 39703 8757 39712
rect 8811 39752 8853 39761
rect 8811 39712 8812 39752
rect 8852 39712 8853 39752
rect 8811 39703 8853 39712
rect 9291 39752 9333 39761
rect 9291 39712 9292 39752
rect 9332 39712 9333 39752
rect 9291 39703 9333 39712
rect 9763 39752 9821 39753
rect 9763 39712 9772 39752
rect 9812 39712 9821 39752
rect 9763 39711 9821 39712
rect 10251 39747 10293 39756
rect 10251 39707 10252 39747
rect 10292 39707 10293 39747
rect 10627 39752 10685 39753
rect 10627 39712 10636 39752
rect 10676 39712 10685 39752
rect 10627 39711 10685 39712
rect 11875 39752 11933 39753
rect 11875 39712 11884 39752
rect 11924 39712 11933 39752
rect 11875 39711 11933 39712
rect 12355 39752 12413 39753
rect 12355 39712 12364 39752
rect 12404 39712 12413 39752
rect 12355 39711 12413 39712
rect 12651 39752 12693 39761
rect 12651 39712 12652 39752
rect 12692 39712 12693 39752
rect 10251 39698 10293 39707
rect 12651 39703 12693 39712
rect 12747 39752 12789 39761
rect 12747 39712 12748 39752
rect 12788 39712 12789 39752
rect 12747 39703 12789 39712
rect 13315 39752 13373 39753
rect 13315 39712 13324 39752
rect 13364 39712 13373 39752
rect 13315 39711 13373 39712
rect 14563 39752 14621 39753
rect 14563 39712 14572 39752
rect 14612 39712 14621 39752
rect 14563 39711 14621 39712
rect 14947 39752 15005 39753
rect 14947 39712 14956 39752
rect 14996 39712 15005 39752
rect 14947 39711 15005 39712
rect 15051 39752 15093 39761
rect 15051 39712 15052 39752
rect 15092 39712 15093 39752
rect 15051 39703 15093 39712
rect 15243 39752 15285 39761
rect 15243 39712 15244 39752
rect 15284 39712 15285 39752
rect 15243 39703 15285 39712
rect 15523 39752 15581 39753
rect 15523 39712 15532 39752
rect 15572 39712 15581 39752
rect 15523 39711 15581 39712
rect 15627 39752 15669 39761
rect 15627 39712 15628 39752
rect 15668 39712 15669 39752
rect 15627 39703 15669 39712
rect 15819 39752 15861 39761
rect 15819 39712 15820 39752
rect 15860 39712 15861 39752
rect 15819 39703 15861 39712
rect 16291 39752 16349 39753
rect 16291 39712 16300 39752
rect 16340 39712 16349 39752
rect 16291 39711 16349 39712
rect 17539 39752 17597 39753
rect 17539 39712 17548 39752
rect 17588 39712 17597 39752
rect 17539 39711 17597 39712
rect 19083 39752 19125 39761
rect 19083 39712 19084 39752
rect 19124 39712 19125 39752
rect 19083 39703 19125 39712
rect 19275 39752 19317 39761
rect 19275 39712 19276 39752
rect 19316 39712 19317 39752
rect 19275 39703 19317 39712
rect 5355 39668 5397 39677
rect 5355 39628 5356 39668
rect 5396 39628 5397 39668
rect 5355 39619 5397 39628
rect 5451 39668 5493 39677
rect 5451 39628 5452 39668
rect 5492 39628 5493 39668
rect 5451 39619 5493 39628
rect 6891 39668 6933 39677
rect 6891 39628 6892 39668
rect 6932 39628 6933 39668
rect 6891 39619 6933 39628
rect 7075 39668 7133 39669
rect 7075 39628 7084 39668
rect 7124 39628 7133 39668
rect 7075 39627 7133 39628
rect 7651 39668 7709 39669
rect 7651 39628 7660 39668
rect 7700 39628 7709 39668
rect 7651 39627 7709 39628
rect 7843 39668 7901 39669
rect 7843 39628 7852 39668
rect 7892 39628 7901 39668
rect 7843 39627 7901 39628
rect 8419 39668 8477 39669
rect 8419 39628 8428 39668
rect 8468 39628 8477 39668
rect 8419 39627 8477 39628
rect 9195 39668 9237 39677
rect 9195 39628 9196 39668
rect 9236 39628 9237 39668
rect 9195 39619 9237 39628
rect 16011 39668 16053 39677
rect 16011 39628 16012 39668
rect 16052 39628 16053 39668
rect 16011 39619 16053 39628
rect 17923 39668 17981 39669
rect 17923 39628 17932 39668
rect 17972 39628 17981 39668
rect 17923 39627 17981 39628
rect 18499 39668 18557 39669
rect 18499 39628 18508 39668
rect 18548 39628 18557 39668
rect 18499 39627 18557 39628
rect 18883 39668 18941 39669
rect 18883 39628 18892 39668
rect 18932 39628 18941 39668
rect 18883 39627 18941 39628
rect 19651 39668 19709 39669
rect 19651 39628 19660 39668
rect 19700 39628 19709 39668
rect 19651 39627 19709 39628
rect 20035 39668 20093 39669
rect 20035 39628 20044 39668
rect 20084 39628 20093 39668
rect 20035 39627 20093 39628
rect 2859 39584 2901 39593
rect 2859 39544 2860 39584
rect 2900 39544 2901 39584
rect 2859 39535 2901 39544
rect 7275 39584 7317 39593
rect 7275 39544 7276 39584
rect 7316 39544 7317 39584
rect 7275 39535 7317 39544
rect 13027 39584 13085 39585
rect 13027 39544 13036 39584
rect 13076 39544 13085 39584
rect 13027 39543 13085 39544
rect 18123 39584 18165 39593
rect 18123 39544 18124 39584
rect 18164 39544 18165 39584
rect 18123 39535 18165 39544
rect 2667 39500 2709 39509
rect 2667 39460 2668 39500
rect 2708 39460 2709 39500
rect 2667 39451 2709 39460
rect 4587 39500 4629 39509
rect 4587 39460 4588 39500
rect 4628 39460 4629 39500
rect 4587 39451 4629 39460
rect 8043 39500 8085 39509
rect 8043 39460 8044 39500
rect 8084 39460 8085 39500
rect 8043 39451 8085 39460
rect 14763 39500 14805 39509
rect 14763 39460 14764 39500
rect 14804 39460 14805 39500
rect 14763 39451 14805 39460
rect 15243 39500 15285 39509
rect 15243 39460 15244 39500
rect 15284 39460 15285 39500
rect 15243 39451 15285 39460
rect 15819 39500 15861 39509
rect 15819 39460 15820 39500
rect 15860 39460 15861 39500
rect 15819 39451 15861 39460
rect 18315 39500 18357 39509
rect 18315 39460 18316 39500
rect 18356 39460 18357 39500
rect 18315 39451 18357 39460
rect 1152 39332 20352 39356
rect 1152 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 20352 39332
rect 1152 39268 20352 39292
rect 4971 39080 5013 39089
rect 4971 39040 4972 39080
rect 5012 39040 5013 39080
rect 4971 39031 5013 39040
rect 6699 39080 6741 39089
rect 6699 39040 6700 39080
rect 6740 39040 6741 39080
rect 15339 39080 15381 39089
rect 6699 39031 6741 39040
rect 13899 39054 13941 39063
rect 13899 39014 13900 39054
rect 13940 39014 13941 39054
rect 15339 39040 15340 39080
rect 15380 39040 15381 39080
rect 15339 39031 15381 39040
rect 15531 39080 15573 39089
rect 15531 39040 15532 39080
rect 15572 39040 15573 39080
rect 15531 39031 15573 39040
rect 15723 39080 15765 39089
rect 15723 39040 15724 39080
rect 15764 39040 15765 39080
rect 15723 39031 15765 39040
rect 18411 39080 18453 39089
rect 18411 39040 18412 39080
rect 18452 39040 18453 39080
rect 18411 39031 18453 39040
rect 18891 39080 18933 39089
rect 18891 39040 18892 39080
rect 18932 39040 18933 39080
rect 18891 39031 18933 39040
rect 19851 39080 19893 39089
rect 19851 39040 19852 39080
rect 19892 39040 19893 39080
rect 19851 39031 19893 39040
rect 13899 39005 13941 39014
rect 1315 38996 1373 38997
rect 1315 38956 1324 38996
rect 1364 38956 1373 38996
rect 1315 38955 1373 38956
rect 3331 38996 3389 38997
rect 3331 38956 3340 38996
rect 3380 38956 3389 38996
rect 3331 38955 3389 38956
rect 4387 38996 4445 38997
rect 4387 38956 4396 38996
rect 4436 38956 4445 38996
rect 4387 38955 4445 38956
rect 4771 38996 4829 38997
rect 4771 38956 4780 38996
rect 4820 38956 4829 38996
rect 4771 38955 4829 38956
rect 9195 38996 9237 39005
rect 9195 38956 9196 38996
rect 9236 38956 9237 38996
rect 1699 38954 1757 38955
rect 1699 38914 1708 38954
rect 1748 38914 1757 38954
rect 9195 38947 9237 38956
rect 16299 38996 16341 39005
rect 16299 38956 16300 38996
rect 16340 38956 16341 38996
rect 16299 38947 16341 38956
rect 18315 38996 18357 39005
rect 18315 38956 18316 38996
rect 18356 38956 18357 38996
rect 18315 38947 18357 38956
rect 18507 38996 18549 39005
rect 18507 38956 18508 38996
rect 18548 38956 18549 38996
rect 18507 38947 18549 38956
rect 19075 38996 19133 38997
rect 19075 38956 19084 38996
rect 19124 38956 19133 38996
rect 19075 38955 19133 38956
rect 19459 38996 19517 38997
rect 19459 38956 19468 38996
rect 19508 38956 19517 38996
rect 19459 38955 19517 38956
rect 20035 38996 20093 38997
rect 20035 38956 20044 38996
rect 20084 38956 20093 38996
rect 20035 38955 20093 38956
rect 10155 38926 10197 38935
rect 1699 38913 1757 38914
rect 2947 38912 3005 38913
rect 2947 38872 2956 38912
rect 2996 38872 3005 38912
rect 2947 38871 3005 38872
rect 5251 38912 5309 38913
rect 5251 38872 5260 38912
rect 5300 38872 5309 38912
rect 5251 38871 5309 38872
rect 6499 38912 6557 38913
rect 6499 38872 6508 38912
rect 6548 38872 6557 38912
rect 6499 38871 6557 38872
rect 6883 38912 6941 38913
rect 6883 38872 6892 38912
rect 6932 38872 6941 38912
rect 6883 38871 6941 38872
rect 8131 38912 8189 38913
rect 8131 38872 8140 38912
rect 8180 38872 8189 38912
rect 8131 38871 8189 38872
rect 8619 38912 8661 38921
rect 8619 38872 8620 38912
rect 8660 38872 8661 38912
rect 8619 38863 8661 38872
rect 8715 38912 8757 38921
rect 8715 38872 8716 38912
rect 8756 38872 8757 38912
rect 8715 38863 8757 38872
rect 9099 38912 9141 38921
rect 9099 38872 9100 38912
rect 9140 38872 9141 38912
rect 9099 38863 9141 38872
rect 9667 38912 9725 38913
rect 9667 38872 9676 38912
rect 9716 38872 9725 38912
rect 10155 38886 10156 38926
rect 10196 38886 10197 38926
rect 10155 38877 10197 38886
rect 10531 38912 10589 38913
rect 9667 38871 9725 38872
rect 10531 38872 10540 38912
rect 10580 38872 10589 38912
rect 10531 38871 10589 38872
rect 11779 38912 11837 38913
rect 11779 38872 11788 38912
rect 11828 38872 11837 38912
rect 11779 38871 11837 38872
rect 12355 38912 12413 38913
rect 12355 38872 12364 38912
rect 12404 38872 12413 38912
rect 12355 38871 12413 38872
rect 13603 38912 13661 38913
rect 13603 38872 13612 38912
rect 13652 38872 13661 38912
rect 13603 38871 13661 38872
rect 13899 38904 13941 38913
rect 13899 38864 13900 38904
rect 13940 38864 13941 38904
rect 13899 38855 13941 38864
rect 14283 38912 14325 38921
rect 14283 38872 14284 38912
rect 14324 38872 14325 38912
rect 14283 38863 14325 38872
rect 14379 38912 14421 38921
rect 14379 38872 14380 38912
rect 14420 38872 14421 38912
rect 14379 38863 14421 38872
rect 14475 38912 14517 38921
rect 14475 38872 14476 38912
rect 14516 38872 14517 38912
rect 14475 38863 14517 38872
rect 14571 38912 14613 38921
rect 14571 38872 14572 38912
rect 14612 38872 14613 38912
rect 14571 38863 14613 38872
rect 14755 38912 14813 38913
rect 14755 38872 14764 38912
rect 14804 38872 14813 38912
rect 14755 38871 14813 38872
rect 14859 38912 14901 38921
rect 14859 38872 14860 38912
rect 14900 38872 14901 38912
rect 14859 38863 14901 38872
rect 15051 38912 15093 38921
rect 15051 38872 15052 38912
rect 15092 38872 15093 38912
rect 15051 38863 15093 38872
rect 15339 38912 15381 38921
rect 15339 38872 15340 38912
rect 15380 38872 15381 38912
rect 15339 38863 15381 38872
rect 15723 38912 15765 38921
rect 15723 38872 15724 38912
rect 15764 38872 15765 38912
rect 15723 38863 15765 38872
rect 15915 38912 15957 38921
rect 15915 38872 15916 38912
rect 15956 38872 15957 38912
rect 15915 38863 15957 38872
rect 16003 38912 16061 38913
rect 16003 38872 16012 38912
rect 16052 38872 16061 38912
rect 16003 38871 16061 38872
rect 16203 38912 16245 38921
rect 16203 38872 16204 38912
rect 16244 38872 16245 38912
rect 16203 38863 16245 38872
rect 16395 38912 16437 38921
rect 16395 38872 16396 38912
rect 16436 38872 16437 38912
rect 16395 38863 16437 38872
rect 16579 38912 16637 38913
rect 16579 38872 16588 38912
rect 16628 38872 16637 38912
rect 16579 38871 16637 38872
rect 17827 38912 17885 38913
rect 17827 38872 17836 38912
rect 17876 38872 17885 38912
rect 17827 38871 17885 38872
rect 18219 38912 18261 38921
rect 18219 38872 18220 38912
rect 18260 38872 18261 38912
rect 18219 38863 18261 38872
rect 18595 38912 18653 38913
rect 18595 38872 18604 38912
rect 18644 38872 18653 38912
rect 18595 38871 18653 38872
rect 18787 38912 18845 38913
rect 18787 38872 18796 38912
rect 18836 38872 18845 38912
rect 18787 38871 18845 38872
rect 10347 38828 10389 38837
rect 10347 38788 10348 38828
rect 10388 38788 10389 38828
rect 10347 38779 10389 38788
rect 11979 38828 12021 38837
rect 11979 38788 11980 38828
rect 12020 38788 12021 38828
rect 11979 38779 12021 38788
rect 14955 38828 14997 38837
rect 14955 38788 14956 38828
rect 14996 38788 14997 38828
rect 14955 38779 14997 38788
rect 1515 38744 1557 38753
rect 1515 38704 1516 38744
rect 1556 38704 1557 38744
rect 1515 38695 1557 38704
rect 3147 38744 3189 38753
rect 3147 38704 3148 38744
rect 3188 38704 3189 38744
rect 3147 38695 3189 38704
rect 3531 38744 3573 38753
rect 3531 38704 3532 38744
rect 3572 38704 3573 38744
rect 3531 38695 3573 38704
rect 3811 38744 3869 38745
rect 3811 38704 3820 38744
rect 3860 38704 3869 38744
rect 3811 38703 3869 38704
rect 4011 38744 4053 38753
rect 4011 38704 4012 38744
rect 4052 38704 4053 38744
rect 4011 38695 4053 38704
rect 4587 38744 4629 38753
rect 4587 38704 4588 38744
rect 4628 38704 4629 38744
rect 4587 38695 4629 38704
rect 8331 38744 8373 38753
rect 8331 38704 8332 38744
rect 8372 38704 8373 38744
rect 8331 38695 8373 38704
rect 12171 38744 12213 38753
rect 12171 38704 12172 38744
rect 12212 38704 12213 38744
rect 12171 38695 12213 38704
rect 14091 38744 14133 38753
rect 14091 38704 14092 38744
rect 14132 38704 14133 38744
rect 14091 38695 14133 38704
rect 18027 38744 18069 38753
rect 18027 38704 18028 38744
rect 18068 38704 18069 38744
rect 18027 38695 18069 38704
rect 19275 38744 19317 38753
rect 19275 38704 19276 38744
rect 19316 38704 19317 38744
rect 19275 38695 19317 38704
rect 19659 38744 19701 38753
rect 19659 38704 19660 38744
rect 19700 38704 19701 38744
rect 19659 38695 19701 38704
rect 1152 38576 20452 38600
rect 1152 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20452 38576
rect 1152 38512 20452 38536
rect 1515 38408 1557 38417
rect 1515 38368 1516 38408
rect 1556 38368 1557 38408
rect 1515 38359 1557 38368
rect 1899 38408 1941 38417
rect 1899 38368 1900 38408
rect 1940 38368 1941 38408
rect 1899 38359 1941 38368
rect 4203 38408 4245 38417
rect 4203 38368 4204 38408
rect 4244 38368 4245 38408
rect 4203 38359 4245 38368
rect 4395 38408 4437 38417
rect 4395 38368 4396 38408
rect 4436 38368 4437 38408
rect 4395 38359 4437 38368
rect 14851 38408 14909 38409
rect 14851 38368 14860 38408
rect 14900 38368 14909 38408
rect 14851 38367 14909 38368
rect 17835 38408 17877 38417
rect 17835 38368 17836 38408
rect 17876 38368 17877 38408
rect 17835 38359 17877 38368
rect 5067 38324 5109 38333
rect 5067 38284 5068 38324
rect 5108 38284 5109 38324
rect 5067 38275 5109 38284
rect 14379 38324 14421 38333
rect 14379 38284 14380 38324
rect 14420 38284 14421 38324
rect 14379 38275 14421 38284
rect 2563 38240 2621 38241
rect 2563 38200 2572 38240
rect 2612 38200 2621 38240
rect 2563 38199 2621 38200
rect 3811 38240 3869 38241
rect 3811 38200 3820 38240
rect 3860 38200 3869 38240
rect 3811 38199 3869 38200
rect 4779 38240 4821 38249
rect 4779 38200 4780 38240
rect 4820 38200 4821 38240
rect 4779 38191 4821 38200
rect 5259 38235 5301 38244
rect 5259 38195 5260 38235
rect 5300 38195 5301 38235
rect 5731 38240 5789 38241
rect 5731 38200 5740 38240
rect 5780 38200 5789 38240
rect 5731 38199 5789 38200
rect 6699 38240 6741 38249
rect 6699 38200 6700 38240
rect 6740 38200 6741 38240
rect 5259 38186 5301 38195
rect 6699 38191 6741 38200
rect 6795 38240 6837 38249
rect 6795 38200 6796 38240
rect 6836 38200 6837 38240
rect 6795 38191 6837 38200
rect 7651 38240 7709 38241
rect 7651 38200 7660 38240
rect 7700 38200 7709 38240
rect 7651 38199 7709 38200
rect 8899 38240 8957 38241
rect 8899 38200 8908 38240
rect 8948 38200 8957 38240
rect 8899 38199 8957 38200
rect 9283 38240 9341 38241
rect 9283 38200 9292 38240
rect 9332 38200 9341 38240
rect 9283 38199 9341 38200
rect 10531 38240 10589 38241
rect 10531 38200 10540 38240
rect 10580 38200 10589 38240
rect 10531 38199 10589 38200
rect 11107 38240 11165 38241
rect 11107 38200 11116 38240
rect 11156 38200 11165 38240
rect 11107 38199 11165 38200
rect 12355 38240 12413 38241
rect 12355 38200 12364 38240
rect 12404 38200 12413 38240
rect 12355 38199 12413 38200
rect 12555 38240 12597 38249
rect 12555 38200 12556 38240
rect 12596 38200 12597 38240
rect 12555 38191 12597 38200
rect 12747 38240 12789 38249
rect 12747 38200 12748 38240
rect 12788 38200 12789 38240
rect 12747 38191 12789 38200
rect 12931 38240 12989 38241
rect 12931 38200 12940 38240
rect 12980 38200 12989 38240
rect 12931 38199 12989 38200
rect 14179 38240 14237 38241
rect 14179 38200 14188 38240
rect 14228 38200 14237 38240
rect 14179 38199 14237 38200
rect 14571 38240 14613 38249
rect 14571 38200 14572 38240
rect 14612 38200 14613 38240
rect 14571 38191 14613 38200
rect 14667 38240 14709 38249
rect 14667 38200 14668 38240
rect 14708 38200 14709 38240
rect 14667 38191 14709 38200
rect 14763 38240 14805 38249
rect 14763 38200 14764 38240
rect 14804 38200 14805 38240
rect 14763 38191 14805 38200
rect 15139 38240 15197 38241
rect 15139 38200 15148 38240
rect 15188 38200 15197 38240
rect 15139 38199 15197 38200
rect 15435 38240 15477 38249
rect 15435 38200 15436 38240
rect 15476 38200 15477 38240
rect 15435 38191 15477 38200
rect 15531 38240 15573 38249
rect 15531 38200 15532 38240
rect 15572 38200 15573 38240
rect 15531 38191 15573 38200
rect 16387 38240 16445 38241
rect 16387 38200 16396 38240
rect 16436 38200 16445 38240
rect 16387 38199 16445 38200
rect 17635 38240 17693 38241
rect 17635 38200 17644 38240
rect 17684 38200 17693 38240
rect 17635 38199 17693 38200
rect 18211 38240 18269 38241
rect 18211 38200 18220 38240
rect 18260 38200 18269 38240
rect 18507 38240 18549 38249
rect 18211 38199 18269 38200
rect 18355 38230 18413 38231
rect 18355 38190 18364 38230
rect 18404 38190 18413 38230
rect 18507 38200 18508 38240
rect 18548 38200 18549 38240
rect 18507 38191 18549 38200
rect 18603 38240 18645 38249
rect 18603 38200 18604 38240
rect 18644 38200 18645 38240
rect 18603 38191 18645 38200
rect 18696 38240 18754 38241
rect 18696 38200 18705 38240
rect 18745 38200 18754 38240
rect 18696 38199 18754 38200
rect 18979 38240 19037 38241
rect 18979 38200 18988 38240
rect 19028 38200 19037 38240
rect 18979 38199 19037 38200
rect 19371 38240 19413 38249
rect 19371 38200 19372 38240
rect 19412 38200 19413 38240
rect 19371 38191 19413 38200
rect 18355 38189 18413 38190
rect 1315 38156 1373 38157
rect 1315 38116 1324 38156
rect 1364 38116 1373 38156
rect 1315 38115 1373 38116
rect 1699 38156 1757 38157
rect 1699 38116 1708 38156
rect 1748 38116 1757 38156
rect 1699 38115 1757 38116
rect 2187 38156 2229 38165
rect 2187 38116 2188 38156
rect 2228 38116 2229 38156
rect 2187 38107 2229 38116
rect 4003 38156 4061 38157
rect 4003 38116 4012 38156
rect 4052 38116 4061 38156
rect 4003 38115 4061 38116
rect 4579 38156 4637 38157
rect 4579 38116 4588 38156
rect 4628 38116 4637 38156
rect 4579 38115 4637 38116
rect 6219 38156 6261 38165
rect 6219 38116 6220 38156
rect 6260 38116 6261 38156
rect 6219 38107 6261 38116
rect 6315 38156 6357 38165
rect 6315 38116 6316 38156
rect 6356 38116 6357 38156
rect 6315 38107 6357 38116
rect 7267 38156 7325 38157
rect 7267 38116 7276 38156
rect 7316 38116 7325 38156
rect 7267 38115 7325 38116
rect 16003 38156 16061 38157
rect 16003 38116 16012 38156
rect 16052 38116 16061 38156
rect 16003 38115 16061 38116
rect 19083 38156 19125 38165
rect 19083 38116 19084 38156
rect 19124 38116 19125 38156
rect 19083 38107 19125 38116
rect 19275 38156 19317 38165
rect 19275 38116 19276 38156
rect 19316 38116 19317 38156
rect 19275 38107 19317 38116
rect 19555 38156 19613 38157
rect 19555 38116 19564 38156
rect 19604 38116 19613 38156
rect 19555 38115 19613 38116
rect 19939 38156 19997 38157
rect 19939 38116 19948 38156
rect 19988 38116 19997 38156
rect 19939 38115 19997 38116
rect 12747 38072 12789 38081
rect 12747 38032 12748 38072
rect 12788 38032 12789 38072
rect 12747 38023 12789 38032
rect 15811 38072 15869 38073
rect 15811 38032 15820 38072
rect 15860 38032 15869 38072
rect 15811 38031 15869 38032
rect 16203 38072 16245 38081
rect 16203 38032 16204 38072
rect 16244 38032 16245 38072
rect 16203 38023 16245 38032
rect 19179 38072 19221 38081
rect 19179 38032 19180 38072
rect 19220 38032 19221 38072
rect 19179 38023 19221 38032
rect 2379 37988 2421 37997
rect 2379 37948 2380 37988
rect 2420 37948 2421 37988
rect 2379 37939 2421 37948
rect 7467 37988 7509 37997
rect 7467 37948 7468 37988
rect 7508 37948 7509 37988
rect 7467 37939 7509 37948
rect 9099 37988 9141 37997
rect 9099 37948 9100 37988
rect 9140 37948 9141 37988
rect 9099 37939 9141 37948
rect 10731 37988 10773 37997
rect 10731 37948 10732 37988
rect 10772 37948 10773 37988
rect 10731 37939 10773 37948
rect 10923 37988 10965 37997
rect 10923 37948 10924 37988
rect 10964 37948 10965 37988
rect 10923 37939 10965 37948
rect 18219 37988 18261 37997
rect 18219 37948 18220 37988
rect 18260 37948 18261 37988
rect 18219 37939 18261 37948
rect 19755 37988 19797 37997
rect 19755 37948 19756 37988
rect 19796 37948 19797 37988
rect 19755 37939 19797 37948
rect 20139 37988 20181 37997
rect 20139 37948 20140 37988
rect 20180 37948 20181 37988
rect 20139 37939 20181 37948
rect 1152 37820 20352 37844
rect 1152 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 20352 37820
rect 1152 37756 20352 37780
rect 1419 37652 1461 37661
rect 1419 37612 1420 37652
rect 1460 37612 1461 37652
rect 1419 37603 1461 37612
rect 7179 37652 7221 37661
rect 7179 37612 7180 37652
rect 7220 37612 7221 37652
rect 7179 37603 7221 37612
rect 9579 37652 9621 37661
rect 9579 37612 9580 37652
rect 9620 37612 9621 37652
rect 9579 37603 9621 37612
rect 9963 37652 10005 37661
rect 9963 37612 9964 37652
rect 10004 37612 10005 37652
rect 9963 37603 10005 37612
rect 13707 37652 13749 37661
rect 13707 37612 13708 37652
rect 13748 37612 13749 37652
rect 13707 37603 13749 37612
rect 14379 37652 14421 37661
rect 14379 37612 14380 37652
rect 14420 37612 14421 37652
rect 14379 37603 14421 37612
rect 14667 37652 14709 37661
rect 14667 37612 14668 37652
rect 14708 37612 14709 37652
rect 14667 37603 14709 37612
rect 16107 37652 16149 37661
rect 16107 37612 16108 37652
rect 16148 37612 16149 37652
rect 16107 37603 16149 37612
rect 17163 37652 17205 37661
rect 17163 37612 17164 37652
rect 17204 37612 17205 37652
rect 17163 37603 17205 37612
rect 18307 37652 18365 37653
rect 18307 37612 18316 37652
rect 18356 37612 18365 37652
rect 18307 37611 18365 37612
rect 18499 37652 18557 37653
rect 18499 37612 18508 37652
rect 18548 37612 18557 37652
rect 18499 37611 18557 37612
rect 20235 37652 20277 37661
rect 20235 37612 20236 37652
rect 20276 37612 20277 37652
rect 20235 37603 20277 37612
rect 4779 37568 4821 37577
rect 4779 37528 4780 37568
rect 4820 37528 4821 37568
rect 4779 37519 4821 37528
rect 15723 37568 15765 37577
rect 15723 37528 15724 37568
rect 15764 37528 15765 37568
rect 15723 37519 15765 37528
rect 1219 37484 1277 37485
rect 1219 37444 1228 37484
rect 1268 37444 1277 37484
rect 1219 37443 1277 37444
rect 3619 37484 3677 37485
rect 3619 37444 3628 37484
rect 3668 37444 3677 37484
rect 3619 37443 3677 37444
rect 4291 37484 4349 37485
rect 4291 37444 4300 37484
rect 4340 37444 4349 37484
rect 4291 37443 4349 37444
rect 4963 37484 5021 37485
rect 4963 37444 4972 37484
rect 5012 37444 5021 37484
rect 4963 37443 5021 37444
rect 6979 37484 7037 37485
rect 6979 37444 6988 37484
rect 7028 37444 7037 37484
rect 6979 37443 7037 37444
rect 9379 37484 9437 37485
rect 9379 37444 9388 37484
rect 9428 37444 9437 37484
rect 9379 37443 9437 37444
rect 9763 37484 9821 37485
rect 9763 37444 9772 37484
rect 9812 37444 9821 37484
rect 9763 37443 9821 37444
rect 15627 37484 15669 37493
rect 15627 37444 15628 37484
rect 15668 37444 15669 37484
rect 15627 37435 15669 37444
rect 15819 37484 15861 37493
rect 15819 37444 15820 37484
rect 15860 37444 15861 37484
rect 15819 37435 15861 37444
rect 17347 37484 17405 37485
rect 17347 37444 17356 37484
rect 17396 37444 17405 37484
rect 19747 37484 19805 37485
rect 17347 37443 17405 37444
rect 16675 37442 16733 37443
rect 1803 37414 1845 37423
rect 1803 37374 1804 37414
rect 1844 37374 1845 37414
rect 9003 37414 9045 37423
rect 1803 37365 1845 37374
rect 2275 37400 2333 37401
rect 2275 37360 2284 37400
rect 2324 37360 2333 37400
rect 2275 37359 2333 37360
rect 2763 37400 2805 37409
rect 2763 37360 2764 37400
rect 2804 37360 2805 37400
rect 2763 37351 2805 37360
rect 2859 37400 2901 37409
rect 2859 37360 2860 37400
rect 2900 37360 2901 37400
rect 3339 37400 3381 37409
rect 2859 37351 2901 37360
rect 3243 37380 3285 37389
rect 3243 37340 3244 37380
rect 3284 37340 3285 37380
rect 3339 37360 3340 37400
rect 3380 37360 3381 37400
rect 3339 37351 3381 37360
rect 5347 37400 5405 37401
rect 5347 37360 5356 37400
rect 5396 37360 5405 37400
rect 5347 37359 5405 37360
rect 6595 37400 6653 37401
rect 6595 37360 6604 37400
rect 6644 37360 6653 37400
rect 6595 37359 6653 37360
rect 7467 37400 7509 37409
rect 7467 37360 7468 37400
rect 7508 37360 7509 37400
rect 7467 37351 7509 37360
rect 7563 37400 7605 37409
rect 7563 37360 7564 37400
rect 7604 37360 7605 37400
rect 7563 37351 7605 37360
rect 7947 37400 7989 37409
rect 7947 37360 7948 37400
rect 7988 37360 7989 37400
rect 7947 37351 7989 37360
rect 8043 37400 8085 37409
rect 8043 37360 8044 37400
rect 8084 37360 8085 37400
rect 8043 37351 8085 37360
rect 8515 37400 8573 37401
rect 8515 37360 8524 37400
rect 8564 37360 8573 37400
rect 9003 37374 9004 37414
rect 9044 37374 9045 37414
rect 9003 37365 9045 37374
rect 10243 37400 10301 37401
rect 8515 37359 8573 37360
rect 10243 37360 10252 37400
rect 10292 37360 10301 37400
rect 10243 37359 10301 37360
rect 10435 37400 10493 37401
rect 10435 37360 10444 37400
rect 10484 37360 10493 37400
rect 10435 37359 10493 37360
rect 11683 37400 11741 37401
rect 11683 37360 11692 37400
rect 11732 37360 11741 37400
rect 11683 37359 11741 37360
rect 12259 37400 12317 37401
rect 12259 37360 12268 37400
rect 12308 37360 12317 37400
rect 12259 37359 12317 37360
rect 13507 37400 13565 37401
rect 13507 37360 13516 37400
rect 13556 37360 13565 37400
rect 13507 37359 13565 37360
rect 13707 37400 13749 37409
rect 13707 37360 13708 37400
rect 13748 37360 13749 37400
rect 13707 37351 13749 37360
rect 13899 37400 13941 37409
rect 13899 37360 13900 37400
rect 13940 37360 13941 37400
rect 13899 37351 13941 37360
rect 14083 37400 14141 37401
rect 14083 37360 14092 37400
rect 14132 37360 14141 37400
rect 14083 37359 14141 37360
rect 14187 37400 14229 37409
rect 14187 37360 14188 37400
rect 14228 37360 14229 37400
rect 14187 37351 14229 37360
rect 14379 37400 14421 37409
rect 14379 37360 14380 37400
rect 14420 37360 14421 37400
rect 14379 37351 14421 37360
rect 14563 37400 14621 37401
rect 14563 37360 14572 37400
rect 14612 37360 14621 37400
rect 14563 37359 14621 37360
rect 14859 37400 14901 37409
rect 14859 37360 14860 37400
rect 14900 37360 14901 37400
rect 14859 37351 14901 37360
rect 14955 37400 14997 37409
rect 14955 37360 14956 37400
rect 14996 37360 14997 37400
rect 14955 37351 14997 37360
rect 15051 37400 15093 37409
rect 15051 37360 15052 37400
rect 15092 37360 15093 37400
rect 15051 37351 15093 37360
rect 15523 37400 15581 37401
rect 15523 37360 15532 37400
rect 15572 37360 15581 37400
rect 15523 37359 15581 37360
rect 15915 37400 15957 37409
rect 15915 37360 15916 37400
rect 15956 37360 15957 37400
rect 15915 37351 15957 37360
rect 16099 37400 16157 37401
rect 16099 37360 16108 37400
rect 16148 37360 16157 37400
rect 16099 37359 16157 37360
rect 16299 37400 16341 37409
rect 16675 37402 16684 37442
rect 16724 37402 16733 37442
rect 17931 37442 17973 37451
rect 19747 37444 19756 37484
rect 19796 37444 19805 37484
rect 19747 37443 19805 37444
rect 16675 37401 16733 37402
rect 16299 37360 16300 37400
rect 16340 37360 16341 37400
rect 16299 37351 16341 37360
rect 16387 37400 16445 37401
rect 16387 37360 16396 37400
rect 16436 37360 16445 37400
rect 16387 37359 16445 37360
rect 16779 37400 16821 37409
rect 16779 37360 16780 37400
rect 16820 37360 16821 37400
rect 16779 37351 16821 37360
rect 16875 37400 16917 37409
rect 16875 37360 16876 37400
rect 16916 37360 16917 37400
rect 17931 37402 17932 37442
rect 17972 37402 17973 37442
rect 17931 37393 17973 37402
rect 18891 37400 18933 37409
rect 16875 37351 16917 37360
rect 17617 37385 17675 37386
rect 17617 37345 17626 37385
rect 17666 37345 17675 37385
rect 18891 37360 18892 37400
rect 18932 37360 18933 37400
rect 18891 37351 18933 37360
rect 19171 37400 19229 37401
rect 19171 37360 19180 37400
rect 19220 37360 19229 37400
rect 19171 37359 19229 37360
rect 19459 37400 19517 37401
rect 19459 37360 19468 37400
rect 19508 37360 19517 37400
rect 19459 37359 19517 37360
rect 20126 37389 20168 37398
rect 17617 37344 17675 37345
rect 20126 37349 20127 37389
rect 20167 37349 20168 37389
rect 20126 37340 20168 37349
rect 3243 37331 3285 37340
rect 18027 37316 18069 37325
rect 18027 37276 18028 37316
rect 18068 37276 18069 37316
rect 18027 37267 18069 37276
rect 18795 37316 18837 37325
rect 18795 37276 18796 37316
rect 18836 37276 18837 37316
rect 18795 37267 18837 37276
rect 1611 37232 1653 37241
rect 1611 37192 1612 37232
rect 1652 37192 1653 37232
rect 1611 37183 1653 37192
rect 3819 37232 3861 37241
rect 3819 37192 3820 37232
rect 3860 37192 3861 37232
rect 3819 37183 3861 37192
rect 4099 37232 4157 37233
rect 4099 37192 4108 37232
rect 4148 37192 4157 37232
rect 4099 37191 4157 37192
rect 4491 37232 4533 37241
rect 4491 37192 4492 37232
rect 4532 37192 4533 37232
rect 4491 37183 4533 37192
rect 5163 37232 5205 37241
rect 5163 37192 5164 37232
rect 5204 37192 5205 37232
rect 5163 37183 5205 37192
rect 6795 37232 6837 37241
rect 6795 37192 6796 37232
rect 6836 37192 6837 37232
rect 6795 37183 6837 37192
rect 9195 37232 9237 37241
rect 9195 37192 9196 37232
rect 9236 37192 9237 37232
rect 9195 37183 9237 37192
rect 10155 37232 10197 37241
rect 10155 37192 10156 37232
rect 10196 37192 10197 37232
rect 10155 37183 10197 37192
rect 11883 37232 11925 37241
rect 11883 37192 11884 37232
rect 11924 37192 11925 37232
rect 11883 37183 11925 37192
rect 12075 37232 12117 37241
rect 12075 37192 12076 37232
rect 12116 37192 12117 37232
rect 12075 37183 12117 37192
rect 15139 37232 15197 37233
rect 15139 37192 15148 37232
rect 15188 37192 15197 37232
rect 15139 37191 15197 37192
rect 16579 37232 16637 37233
rect 16579 37192 16588 37232
rect 16628 37192 16637 37232
rect 16579 37191 16637 37192
rect 19563 37232 19605 37241
rect 19563 37192 19564 37232
rect 19604 37192 19605 37232
rect 19563 37183 19605 37192
rect 19947 37232 19989 37241
rect 19947 37192 19948 37232
rect 19988 37192 19989 37232
rect 19947 37183 19989 37192
rect 1152 37064 20452 37088
rect 1152 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20452 37064
rect 1152 37000 20452 37024
rect 1515 36896 1557 36905
rect 1515 36856 1516 36896
rect 1556 36856 1557 36896
rect 1515 36847 1557 36856
rect 5739 36896 5781 36905
rect 5739 36856 5740 36896
rect 5780 36856 5781 36896
rect 5739 36847 5781 36856
rect 9387 36896 9429 36905
rect 9387 36856 9388 36896
rect 9428 36856 9429 36896
rect 9387 36847 9429 36856
rect 15531 36896 15573 36905
rect 15531 36856 15532 36896
rect 15572 36856 15573 36896
rect 15531 36847 15573 36856
rect 18123 36896 18165 36905
rect 18123 36856 18124 36896
rect 18164 36856 18165 36896
rect 18123 36847 18165 36856
rect 19275 36896 19317 36905
rect 19275 36856 19276 36896
rect 19316 36856 19317 36896
rect 19275 36847 19317 36856
rect 5163 36812 5205 36821
rect 5163 36772 5164 36812
rect 5204 36772 5205 36812
rect 5163 36763 5205 36772
rect 11787 36812 11829 36821
rect 11787 36772 11788 36812
rect 11828 36772 11829 36812
rect 11787 36763 11829 36772
rect 13803 36812 13845 36821
rect 13803 36772 13804 36812
rect 13844 36772 13845 36812
rect 13803 36763 13845 36772
rect 15907 36812 15965 36813
rect 15907 36772 15916 36812
rect 15956 36772 15965 36812
rect 15907 36771 15965 36772
rect 3531 36748 3573 36757
rect 1699 36728 1757 36729
rect 1699 36688 1708 36728
rect 1748 36688 1757 36728
rect 3435 36728 3477 36737
rect 1699 36687 1757 36688
rect 2947 36707 3005 36708
rect 2947 36667 2956 36707
rect 2996 36667 3005 36707
rect 3435 36688 3436 36728
rect 3476 36688 3477 36728
rect 3531 36708 3532 36748
rect 3572 36708 3573 36748
rect 3531 36699 3573 36708
rect 3915 36728 3957 36737
rect 3435 36679 3477 36688
rect 3915 36688 3916 36728
rect 3956 36688 3957 36728
rect 3915 36679 3957 36688
rect 4483 36728 4541 36729
rect 4483 36688 4492 36728
rect 4532 36688 4541 36728
rect 4483 36687 4541 36688
rect 4971 36723 5013 36732
rect 4971 36683 4972 36723
rect 5012 36683 5013 36723
rect 5923 36728 5981 36729
rect 5923 36688 5932 36728
rect 5972 36688 5981 36728
rect 5923 36687 5981 36688
rect 7171 36728 7229 36729
rect 7171 36688 7180 36728
rect 7220 36688 7229 36728
rect 7171 36687 7229 36688
rect 7659 36728 7701 36737
rect 7659 36688 7660 36728
rect 7700 36688 7701 36728
rect 4971 36674 5013 36683
rect 7659 36679 7701 36688
rect 7755 36728 7797 36737
rect 7755 36688 7756 36728
rect 7796 36688 7797 36728
rect 7755 36679 7797 36688
rect 8139 36728 8181 36737
rect 8139 36688 8140 36728
rect 8180 36688 8181 36728
rect 8139 36679 8181 36688
rect 8707 36728 8765 36729
rect 8707 36688 8716 36728
rect 8756 36688 8765 36728
rect 8707 36687 8765 36688
rect 9195 36723 9237 36732
rect 9195 36683 9196 36723
rect 9236 36683 9237 36723
rect 9195 36674 9237 36683
rect 10059 36728 10101 36737
rect 10059 36688 10060 36728
rect 10100 36688 10101 36728
rect 10059 36679 10101 36688
rect 10155 36728 10197 36737
rect 10155 36688 10156 36728
rect 10196 36688 10197 36728
rect 10155 36679 10197 36688
rect 10539 36728 10581 36737
rect 10539 36688 10540 36728
rect 10580 36688 10581 36728
rect 10539 36679 10581 36688
rect 10635 36728 10677 36737
rect 10635 36688 10636 36728
rect 10676 36688 10677 36728
rect 10635 36679 10677 36688
rect 11107 36728 11165 36729
rect 11107 36688 11116 36728
rect 11156 36688 11165 36728
rect 12075 36728 12117 36737
rect 11107 36687 11165 36688
rect 11595 36714 11637 36723
rect 11595 36674 11596 36714
rect 11636 36674 11637 36714
rect 12075 36688 12076 36728
rect 12116 36688 12117 36728
rect 12075 36679 12117 36688
rect 12171 36728 12213 36737
rect 12171 36688 12172 36728
rect 12212 36688 12213 36728
rect 12171 36679 12213 36688
rect 12555 36728 12597 36737
rect 12555 36688 12556 36728
rect 12596 36688 12597 36728
rect 12555 36679 12597 36688
rect 13123 36728 13181 36729
rect 13123 36688 13132 36728
rect 13172 36688 13181 36728
rect 14083 36728 14141 36729
rect 13123 36687 13181 36688
rect 13659 36686 13701 36695
rect 14083 36688 14092 36728
rect 14132 36688 14141 36728
rect 14083 36687 14141 36688
rect 15331 36728 15389 36729
rect 15331 36688 15340 36728
rect 15380 36688 15389 36728
rect 16003 36728 16061 36729
rect 15331 36687 15389 36688
rect 15915 36705 15957 36714
rect 2947 36666 3005 36667
rect 11595 36665 11637 36674
rect 1315 36644 1373 36645
rect 1315 36604 1324 36644
rect 1364 36604 1373 36644
rect 1315 36603 1373 36604
rect 4011 36644 4053 36653
rect 4011 36604 4012 36644
rect 4052 36604 4053 36644
rect 4011 36595 4053 36604
rect 5539 36644 5597 36645
rect 5539 36604 5548 36644
rect 5588 36604 5597 36644
rect 5539 36603 5597 36604
rect 8235 36644 8277 36653
rect 8235 36604 8236 36644
rect 8276 36604 8277 36644
rect 8235 36595 8277 36604
rect 9571 36644 9629 36645
rect 9571 36604 9580 36644
rect 9620 36604 9629 36644
rect 9571 36603 9629 36604
rect 12651 36644 12693 36653
rect 12651 36604 12652 36644
rect 12692 36604 12693 36644
rect 13659 36646 13660 36686
rect 13700 36646 13701 36686
rect 15915 36665 15916 36705
rect 15956 36665 15957 36705
rect 16003 36688 16012 36728
rect 16052 36688 16061 36728
rect 16299 36728 16341 36737
rect 16003 36687 16061 36688
rect 16203 36713 16245 36722
rect 15915 36656 15957 36665
rect 16203 36673 16204 36713
rect 16244 36673 16245 36713
rect 16299 36688 16300 36728
rect 16340 36688 16341 36728
rect 16675 36728 16733 36729
rect 16299 36679 16341 36688
rect 16456 36713 16498 36722
rect 16203 36664 16245 36673
rect 16456 36673 16457 36713
rect 16497 36673 16498 36713
rect 16675 36688 16684 36728
rect 16724 36688 16733 36728
rect 16675 36687 16733 36688
rect 17067 36728 17109 36737
rect 17067 36688 17068 36728
rect 17108 36688 17109 36728
rect 17067 36679 17109 36688
rect 17259 36728 17301 36737
rect 17259 36688 17260 36728
rect 17300 36688 17301 36728
rect 17259 36679 17301 36688
rect 17451 36728 17493 36737
rect 17451 36688 17452 36728
rect 17492 36688 17493 36728
rect 17451 36679 17493 36688
rect 17827 36728 17885 36729
rect 17827 36688 17836 36728
rect 17876 36688 17885 36728
rect 17827 36687 17885 36688
rect 17931 36728 17973 36737
rect 17931 36688 17932 36728
rect 17972 36688 17973 36728
rect 17931 36679 17973 36688
rect 18115 36728 18173 36729
rect 18115 36688 18124 36728
rect 18164 36688 18173 36728
rect 18115 36687 18173 36688
rect 18315 36728 18357 36737
rect 18315 36688 18316 36728
rect 18356 36688 18357 36728
rect 18315 36679 18357 36688
rect 18507 36728 18549 36737
rect 18507 36688 18508 36728
rect 18548 36688 18549 36728
rect 18507 36679 18549 36688
rect 16456 36664 16498 36673
rect 13659 36637 13701 36646
rect 16779 36644 16821 36653
rect 12651 36595 12693 36604
rect 16779 36604 16780 36644
rect 16820 36604 16821 36644
rect 16779 36595 16821 36604
rect 16971 36644 17013 36653
rect 16971 36604 16972 36644
rect 17012 36604 17013 36644
rect 16971 36595 17013 36604
rect 17355 36644 17397 36653
rect 17355 36604 17356 36644
rect 17396 36604 17397 36644
rect 17355 36595 17397 36604
rect 18411 36644 18453 36653
rect 18411 36604 18412 36644
rect 18452 36604 18453 36644
rect 18411 36595 18453 36604
rect 18691 36644 18749 36645
rect 18691 36604 18700 36644
rect 18740 36604 18749 36644
rect 18691 36603 18749 36604
rect 19075 36644 19133 36645
rect 19075 36604 19084 36644
rect 19124 36604 19133 36644
rect 19075 36603 19133 36604
rect 19459 36644 19517 36645
rect 19459 36604 19468 36644
rect 19508 36604 19517 36644
rect 19459 36603 19517 36604
rect 19843 36644 19901 36645
rect 19843 36604 19852 36644
rect 19892 36604 19901 36644
rect 19843 36603 19901 36604
rect 9771 36560 9813 36569
rect 9771 36520 9772 36560
rect 9812 36520 9813 36560
rect 9771 36511 9813 36520
rect 16875 36560 16917 36569
rect 16875 36520 16876 36560
rect 16916 36520 16917 36560
rect 16875 36511 16917 36520
rect 18891 36560 18933 36569
rect 18891 36520 18892 36560
rect 18932 36520 18933 36560
rect 18891 36511 18933 36520
rect 20043 36560 20085 36569
rect 20043 36520 20044 36560
rect 20084 36520 20085 36560
rect 20043 36511 20085 36520
rect 3147 36476 3189 36485
rect 3147 36436 3148 36476
rect 3188 36436 3189 36476
rect 3147 36427 3189 36436
rect 7371 36476 7413 36485
rect 7371 36436 7372 36476
rect 7412 36436 7413 36476
rect 7371 36427 7413 36436
rect 19659 36476 19701 36485
rect 19659 36436 19660 36476
rect 19700 36436 19701 36476
rect 19659 36427 19701 36436
rect 1152 36308 20352 36332
rect 1152 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 20352 36308
rect 1152 36244 20352 36268
rect 16579 36182 16637 36183
rect 1611 36140 1653 36149
rect 1611 36100 1612 36140
rect 1652 36100 1653 36140
rect 1611 36091 1653 36100
rect 2571 36140 2613 36149
rect 2571 36100 2572 36140
rect 2612 36100 2613 36140
rect 2571 36091 2613 36100
rect 11979 36140 12021 36149
rect 11979 36100 11980 36140
rect 12020 36100 12021 36140
rect 11979 36091 12021 36100
rect 13803 36140 13845 36149
rect 13803 36100 13804 36140
rect 13844 36100 13845 36140
rect 13803 36091 13845 36100
rect 15435 36140 15477 36149
rect 16579 36142 16588 36182
rect 16628 36142 16637 36182
rect 16579 36141 16637 36142
rect 15435 36100 15436 36140
rect 15476 36100 15477 36140
rect 15435 36091 15477 36100
rect 16387 36056 16445 36057
rect 16387 36016 16396 36056
rect 16436 36016 16445 36056
rect 16387 36015 16445 36016
rect 1411 35972 1469 35973
rect 1411 35932 1420 35972
rect 1460 35932 1469 35972
rect 1411 35931 1469 35932
rect 1795 35972 1853 35973
rect 1795 35932 1804 35972
rect 1844 35932 1853 35972
rect 1795 35931 1853 35932
rect 2371 35972 2429 35973
rect 2371 35932 2380 35972
rect 2420 35932 2429 35972
rect 2371 35931 2429 35932
rect 3915 35972 3957 35981
rect 3915 35932 3916 35972
rect 3956 35932 3957 35972
rect 3915 35923 3957 35932
rect 9187 35972 9245 35973
rect 9187 35932 9196 35972
rect 9236 35932 9245 35972
rect 9187 35931 9245 35932
rect 19363 35972 19421 35973
rect 19363 35932 19372 35972
rect 19412 35932 19421 35972
rect 19363 35931 19421 35932
rect 19747 35972 19805 35973
rect 19747 35932 19756 35972
rect 19796 35932 19805 35972
rect 19747 35931 19805 35932
rect 2955 35902 2997 35911
rect 2955 35862 2956 35902
rect 2996 35862 2997 35902
rect 2955 35853 2997 35862
rect 3427 35888 3485 35889
rect 3427 35848 3436 35888
rect 3476 35848 3485 35888
rect 3427 35847 3485 35848
rect 4011 35888 4053 35897
rect 4011 35848 4012 35888
rect 4052 35848 4053 35888
rect 4011 35839 4053 35848
rect 4395 35888 4437 35897
rect 4395 35848 4396 35888
rect 4436 35848 4437 35888
rect 4395 35839 4437 35848
rect 4491 35888 4533 35897
rect 4491 35848 4492 35888
rect 4532 35848 4533 35888
rect 4491 35839 4533 35848
rect 5067 35888 5109 35897
rect 5067 35848 5068 35888
rect 5108 35848 5109 35888
rect 5067 35839 5109 35848
rect 5259 35888 5301 35897
rect 5259 35848 5260 35888
rect 5300 35848 5301 35888
rect 5259 35839 5301 35848
rect 5347 35888 5405 35889
rect 5347 35848 5356 35888
rect 5396 35848 5405 35888
rect 5347 35847 5405 35848
rect 5539 35888 5597 35889
rect 5539 35848 5548 35888
rect 5588 35848 5597 35888
rect 5539 35847 5597 35848
rect 6787 35888 6845 35889
rect 6787 35848 6796 35888
rect 6836 35848 6845 35888
rect 6787 35847 6845 35848
rect 7275 35888 7317 35897
rect 7275 35848 7276 35888
rect 7316 35848 7317 35888
rect 7275 35839 7317 35848
rect 7371 35888 7413 35897
rect 7371 35848 7372 35888
rect 7412 35848 7413 35888
rect 7371 35839 7413 35848
rect 7755 35888 7797 35897
rect 7755 35848 7756 35888
rect 7796 35848 7797 35888
rect 7755 35839 7797 35848
rect 7851 35888 7893 35897
rect 8811 35893 8853 35902
rect 7851 35848 7852 35888
rect 7892 35848 7893 35888
rect 7851 35839 7893 35848
rect 8323 35888 8381 35889
rect 8323 35848 8332 35888
rect 8372 35848 8381 35888
rect 8323 35847 8381 35848
rect 8811 35853 8812 35893
rect 8852 35853 8853 35893
rect 8811 35844 8853 35853
rect 9675 35888 9717 35897
rect 9675 35848 9676 35888
rect 9716 35848 9717 35888
rect 9675 35839 9717 35848
rect 9771 35888 9813 35897
rect 9771 35848 9772 35888
rect 9812 35848 9813 35888
rect 9771 35839 9813 35848
rect 9867 35888 9909 35897
rect 9867 35848 9868 35888
rect 9908 35848 9909 35888
rect 9867 35839 9909 35848
rect 10059 35888 10101 35897
rect 10059 35848 10060 35888
rect 10100 35848 10101 35888
rect 10059 35839 10101 35848
rect 10155 35888 10197 35897
rect 10155 35848 10156 35888
rect 10196 35848 10197 35888
rect 10155 35839 10197 35848
rect 10251 35888 10293 35897
rect 10251 35848 10252 35888
rect 10292 35848 10293 35888
rect 10251 35839 10293 35848
rect 10347 35888 10389 35897
rect 10347 35848 10348 35888
rect 10388 35848 10389 35888
rect 10347 35839 10389 35848
rect 10531 35888 10589 35889
rect 10531 35848 10540 35888
rect 10580 35848 10589 35888
rect 10531 35847 10589 35848
rect 11779 35888 11837 35889
rect 11779 35848 11788 35888
rect 11828 35848 11837 35888
rect 11779 35847 11837 35848
rect 12355 35888 12413 35889
rect 12355 35848 12364 35888
rect 12404 35848 12413 35888
rect 12355 35847 12413 35848
rect 13603 35888 13661 35889
rect 13603 35848 13612 35888
rect 13652 35848 13661 35888
rect 13603 35847 13661 35848
rect 13987 35888 14045 35889
rect 13987 35848 13996 35888
rect 14036 35848 14045 35888
rect 13987 35847 14045 35848
rect 15235 35888 15293 35889
rect 15235 35848 15244 35888
rect 15284 35848 15293 35888
rect 15235 35847 15293 35848
rect 15715 35888 15773 35889
rect 15715 35848 15724 35888
rect 15764 35848 15773 35888
rect 15715 35847 15773 35848
rect 16011 35888 16053 35897
rect 16011 35848 16012 35888
rect 16052 35848 16053 35888
rect 16011 35839 16053 35848
rect 16971 35888 17013 35897
rect 16971 35848 16972 35888
rect 17012 35848 17013 35888
rect 16971 35839 17013 35848
rect 17251 35888 17309 35889
rect 17251 35848 17260 35888
rect 17300 35848 17309 35888
rect 17251 35847 17309 35848
rect 17731 35888 17789 35889
rect 17731 35848 17740 35888
rect 17780 35848 17789 35888
rect 17731 35847 17789 35848
rect 18979 35888 19037 35889
rect 18979 35848 18988 35888
rect 19028 35848 19037 35888
rect 18979 35847 19037 35848
rect 20126 35888 20168 35897
rect 20126 35848 20127 35888
rect 20167 35848 20168 35888
rect 20126 35839 20168 35848
rect 2763 35804 2805 35813
rect 2763 35764 2764 35804
rect 2804 35764 2805 35804
rect 2763 35755 2805 35764
rect 5163 35804 5205 35813
rect 5163 35764 5164 35804
rect 5204 35764 5205 35804
rect 5163 35755 5205 35764
rect 6987 35804 7029 35813
rect 6987 35764 6988 35804
rect 7028 35764 7029 35804
rect 6987 35755 7029 35764
rect 16107 35804 16149 35813
rect 16107 35764 16108 35804
rect 16148 35764 16149 35804
rect 16107 35755 16149 35764
rect 16875 35804 16917 35813
rect 16875 35764 16876 35804
rect 16916 35764 16917 35804
rect 16875 35755 16917 35764
rect 20235 35804 20277 35813
rect 20235 35764 20236 35804
rect 20276 35764 20277 35804
rect 20235 35755 20277 35764
rect 1995 35720 2037 35729
rect 1995 35680 1996 35720
rect 2036 35680 2037 35720
rect 1995 35671 2037 35680
rect 4779 35720 4821 35729
rect 4779 35680 4780 35720
rect 4820 35680 4821 35720
rect 4779 35671 4821 35680
rect 9003 35720 9045 35729
rect 9003 35680 9004 35720
rect 9044 35680 9045 35720
rect 9003 35671 9045 35680
rect 9387 35720 9429 35729
rect 9387 35680 9388 35720
rect 9428 35680 9429 35720
rect 9387 35671 9429 35680
rect 9571 35720 9629 35721
rect 9571 35680 9580 35720
rect 9620 35680 9629 35720
rect 9571 35679 9629 35680
rect 19179 35720 19221 35729
rect 19179 35680 19180 35720
rect 19220 35680 19221 35720
rect 19179 35671 19221 35680
rect 19563 35720 19605 35729
rect 19563 35680 19564 35720
rect 19604 35680 19605 35720
rect 19563 35671 19605 35680
rect 19947 35720 19989 35729
rect 19947 35680 19948 35720
rect 19988 35680 19989 35720
rect 19947 35671 19989 35680
rect 1152 35552 20452 35576
rect 1152 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20452 35552
rect 1152 35488 20452 35512
rect 9867 35384 9909 35393
rect 9867 35344 9868 35384
rect 9908 35344 9909 35384
rect 9867 35335 9909 35344
rect 7659 35300 7701 35309
rect 7659 35260 7660 35300
rect 7700 35260 7701 35300
rect 7659 35251 7701 35260
rect 12451 35300 12509 35301
rect 12451 35260 12460 35300
rect 12500 35260 12509 35300
rect 12451 35259 12509 35260
rect 17163 35300 17205 35309
rect 17163 35260 17164 35300
rect 17204 35260 17205 35300
rect 17163 35251 17205 35260
rect 19179 35300 19221 35309
rect 19179 35260 19180 35300
rect 19220 35260 19221 35300
rect 19179 35251 19221 35260
rect 1891 35216 1949 35217
rect 1891 35176 1900 35216
rect 1940 35176 1949 35216
rect 1891 35175 1949 35176
rect 3139 35216 3197 35217
rect 3139 35176 3148 35216
rect 3188 35176 3197 35216
rect 3139 35175 3197 35176
rect 4195 35216 4253 35217
rect 4195 35176 4204 35216
rect 4244 35176 4253 35216
rect 4195 35175 4253 35176
rect 5443 35216 5501 35217
rect 5443 35176 5452 35216
rect 5492 35176 5501 35216
rect 5443 35175 5501 35176
rect 5931 35216 5973 35225
rect 5931 35176 5932 35216
rect 5972 35176 5973 35216
rect 5931 35167 5973 35176
rect 6027 35216 6069 35225
rect 6027 35176 6028 35216
rect 6068 35176 6069 35216
rect 6027 35167 6069 35176
rect 6979 35216 7037 35217
rect 6979 35176 6988 35216
rect 7028 35176 7037 35216
rect 7851 35216 7893 35225
rect 6979 35175 7037 35176
rect 7467 35202 7509 35211
rect 7467 35162 7468 35202
rect 7508 35162 7509 35202
rect 7851 35176 7852 35216
rect 7892 35176 7893 35216
rect 7851 35167 7893 35176
rect 8035 35216 8093 35217
rect 8035 35176 8044 35216
rect 8084 35176 8093 35216
rect 8035 35175 8093 35176
rect 8227 35216 8285 35217
rect 8227 35176 8236 35216
rect 8276 35176 8285 35216
rect 8227 35175 8285 35176
rect 9475 35216 9533 35217
rect 9475 35176 9484 35216
rect 9524 35176 9533 35216
rect 11299 35216 11357 35217
rect 9475 35175 9533 35176
rect 10051 35195 10109 35196
rect 7467 35153 7509 35162
rect 10051 35155 10060 35195
rect 10100 35155 10109 35195
rect 11299 35176 11308 35216
rect 11348 35176 11357 35216
rect 11299 35175 11357 35176
rect 11587 35216 11645 35217
rect 11587 35176 11596 35216
rect 11636 35176 11645 35216
rect 11587 35175 11645 35176
rect 12835 35216 12893 35217
rect 12835 35176 12844 35216
rect 12884 35176 12893 35216
rect 12835 35175 12893 35176
rect 13131 35216 13173 35225
rect 13131 35176 13132 35216
rect 13172 35176 13173 35216
rect 13131 35167 13173 35176
rect 13227 35216 13269 35225
rect 13227 35176 13228 35216
rect 13268 35176 13269 35216
rect 13227 35167 13269 35176
rect 13699 35216 13757 35217
rect 13699 35176 13708 35216
rect 13748 35176 13757 35216
rect 13699 35175 13757 35176
rect 14947 35216 15005 35217
rect 14947 35176 14956 35216
rect 14996 35176 15005 35216
rect 14947 35175 15005 35176
rect 15339 35216 15381 35225
rect 15339 35176 15340 35216
rect 15380 35176 15381 35216
rect 15339 35167 15381 35176
rect 15531 35216 15573 35225
rect 15531 35176 15532 35216
rect 15572 35176 15573 35216
rect 15531 35167 15573 35176
rect 15715 35216 15773 35217
rect 15715 35176 15724 35216
rect 15764 35176 15773 35216
rect 15715 35175 15773 35176
rect 16963 35216 17021 35217
rect 16963 35176 16972 35216
rect 17012 35176 17021 35216
rect 16963 35175 17021 35176
rect 17451 35216 17493 35225
rect 17451 35176 17452 35216
rect 17492 35176 17493 35216
rect 17451 35167 17493 35176
rect 17547 35216 17589 35225
rect 17547 35176 17548 35216
rect 17588 35176 17589 35216
rect 17547 35167 17589 35176
rect 18499 35216 18557 35217
rect 18499 35176 18508 35216
rect 18548 35176 18557 35216
rect 18499 35175 18557 35176
rect 19035 35206 19077 35215
rect 19035 35166 19036 35206
rect 19076 35166 19077 35206
rect 19035 35157 19077 35166
rect 10051 35154 10109 35155
rect 1507 35132 1565 35133
rect 1507 35092 1516 35132
rect 1556 35092 1565 35132
rect 1507 35091 1565 35092
rect 3811 35132 3869 35133
rect 3811 35092 3820 35132
rect 3860 35092 3869 35132
rect 3811 35091 3869 35092
rect 6411 35132 6453 35141
rect 6411 35092 6412 35132
rect 6452 35092 6453 35132
rect 6411 35083 6453 35092
rect 6507 35132 6549 35141
rect 6507 35092 6508 35132
rect 6548 35092 6549 35132
rect 6507 35083 6549 35092
rect 17931 35132 17973 35141
rect 17931 35092 17932 35132
rect 17972 35092 17973 35132
rect 17931 35083 17973 35092
rect 18027 35132 18069 35141
rect 18027 35092 18028 35132
rect 18068 35092 18069 35132
rect 18027 35083 18069 35092
rect 19651 35132 19709 35133
rect 19651 35092 19660 35132
rect 19700 35092 19709 35132
rect 19651 35091 19709 35092
rect 19843 35132 19901 35133
rect 19843 35092 19852 35132
rect 19892 35092 19901 35132
rect 19843 35091 19901 35092
rect 1323 35048 1365 35057
rect 1323 35008 1324 35048
rect 1364 35008 1365 35048
rect 1323 34999 1365 35008
rect 1707 35048 1749 35057
rect 1707 35008 1708 35048
rect 1748 35008 1749 35048
rect 1707 34999 1749 35008
rect 3531 35048 3573 35057
rect 3531 35008 3532 35048
rect 3572 35008 3573 35048
rect 3531 34999 3573 35008
rect 4011 35048 4053 35057
rect 4011 35008 4012 35048
rect 4052 35008 4053 35048
rect 4011 34999 4053 35008
rect 5643 35048 5685 35057
rect 5643 35008 5644 35048
rect 5684 35008 5685 35048
rect 5643 34999 5685 35008
rect 19467 35048 19509 35057
rect 19467 35008 19468 35048
rect 19508 35008 19509 35048
rect 19467 34999 19509 35008
rect 3339 34964 3381 34973
rect 3339 34924 3340 34964
rect 3380 34924 3381 34964
rect 3339 34915 3381 34924
rect 7947 34964 7989 34973
rect 7947 34924 7948 34964
rect 7988 34924 7989 34964
rect 7947 34915 7989 34924
rect 9675 34964 9717 34973
rect 9675 34924 9676 34964
rect 9716 34924 9717 34964
rect 9675 34915 9717 34924
rect 13507 34964 13565 34965
rect 13507 34924 13516 34964
rect 13556 34924 13565 34964
rect 13507 34923 13565 34924
rect 15147 34964 15189 34973
rect 15147 34924 15148 34964
rect 15188 34924 15189 34964
rect 15147 34915 15189 34924
rect 15339 34964 15381 34973
rect 15339 34924 15340 34964
rect 15380 34924 15381 34964
rect 15339 34915 15381 34924
rect 20043 34964 20085 34973
rect 20043 34924 20044 34964
rect 20084 34924 20085 34964
rect 20043 34915 20085 34924
rect 1152 34796 20352 34820
rect 1152 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 20352 34796
rect 1152 34732 20352 34756
rect 3339 34628 3381 34637
rect 3339 34588 3340 34628
rect 3380 34588 3381 34628
rect 3339 34579 3381 34588
rect 7179 34628 7221 34637
rect 7179 34588 7180 34628
rect 7220 34588 7221 34628
rect 7179 34579 7221 34588
rect 14475 34628 14517 34637
rect 14475 34588 14476 34628
rect 14516 34588 14517 34628
rect 14475 34579 14517 34588
rect 14667 34628 14709 34637
rect 14667 34588 14668 34628
rect 14708 34588 14709 34628
rect 14667 34579 14709 34588
rect 4683 34460 4725 34469
rect 3139 34447 3197 34448
rect 3139 34407 3148 34447
rect 3188 34407 3197 34447
rect 3139 34406 3197 34407
rect 3675 34418 3717 34427
rect 3675 34378 3676 34418
rect 3716 34378 3717 34418
rect 4683 34420 4684 34460
rect 4724 34420 4725 34460
rect 4683 34411 4725 34420
rect 8427 34460 8469 34469
rect 8427 34420 8428 34460
rect 8468 34420 8469 34460
rect 8427 34411 8469 34420
rect 8523 34460 8565 34469
rect 8523 34420 8524 34460
rect 8564 34420 8565 34460
rect 11499 34460 11541 34469
rect 8523 34411 8565 34420
rect 9531 34418 9573 34427
rect 1315 34376 1373 34377
rect 1315 34336 1324 34376
rect 1364 34336 1373 34376
rect 1315 34335 1373 34336
rect 1507 34376 1565 34377
rect 1507 34336 1516 34376
rect 1556 34336 1565 34376
rect 1507 34335 1565 34336
rect 2755 34376 2813 34377
rect 2755 34336 2764 34376
rect 2804 34336 2813 34376
rect 3675 34369 3717 34378
rect 4195 34376 4253 34377
rect 2755 34335 2813 34336
rect 4195 34336 4204 34376
rect 4244 34336 4253 34376
rect 4195 34335 4253 34336
rect 4779 34376 4821 34385
rect 4779 34336 4780 34376
rect 4820 34336 4821 34376
rect 4779 34327 4821 34336
rect 5163 34376 5205 34385
rect 5163 34336 5164 34376
rect 5204 34336 5205 34376
rect 5163 34327 5205 34336
rect 5259 34376 5301 34385
rect 5259 34336 5260 34376
rect 5300 34336 5301 34376
rect 5259 34327 5301 34336
rect 5731 34376 5789 34377
rect 5731 34336 5740 34376
rect 5780 34336 5789 34376
rect 5731 34335 5789 34336
rect 6979 34376 7037 34377
rect 6979 34336 6988 34376
rect 7028 34336 7037 34376
rect 7659 34376 7701 34385
rect 6979 34335 7037 34336
rect 7467 34355 7509 34364
rect 7467 34315 7468 34355
rect 7508 34315 7509 34355
rect 7467 34306 7509 34315
rect 7563 34355 7605 34364
rect 7563 34315 7564 34355
rect 7604 34315 7605 34355
rect 7659 34336 7660 34376
rect 7700 34336 7701 34376
rect 7659 34327 7701 34336
rect 7947 34376 7989 34385
rect 7947 34336 7948 34376
rect 7988 34336 7989 34376
rect 7947 34327 7989 34336
rect 8043 34376 8085 34385
rect 9531 34378 9532 34418
rect 9572 34378 9573 34418
rect 11499 34420 11500 34460
rect 11540 34420 11541 34460
rect 11499 34411 11541 34420
rect 19939 34397 19997 34398
rect 8043 34336 8044 34376
rect 8084 34336 8085 34376
rect 8043 34327 8085 34336
rect 8995 34376 9053 34377
rect 8995 34336 9004 34376
rect 9044 34336 9053 34376
rect 9531 34369 9573 34378
rect 9963 34376 10005 34385
rect 8995 34335 9053 34336
rect 9963 34336 9964 34376
rect 10004 34336 10005 34376
rect 9963 34327 10005 34336
rect 10059 34376 10101 34385
rect 10059 34336 10060 34376
rect 10100 34336 10101 34376
rect 10059 34327 10101 34336
rect 10155 34376 10197 34385
rect 10155 34336 10156 34376
rect 10196 34336 10197 34376
rect 10155 34327 10197 34336
rect 10347 34376 10389 34385
rect 10347 34336 10348 34376
rect 10388 34336 10389 34376
rect 10347 34327 10389 34336
rect 10443 34376 10485 34385
rect 10443 34336 10444 34376
rect 10484 34336 10485 34376
rect 10443 34327 10485 34336
rect 10539 34376 10581 34385
rect 10539 34336 10540 34376
rect 10580 34336 10581 34376
rect 10539 34327 10581 34336
rect 10923 34376 10965 34385
rect 10923 34336 10924 34376
rect 10964 34336 10965 34376
rect 10923 34327 10965 34336
rect 11019 34376 11061 34385
rect 11019 34336 11020 34376
rect 11060 34336 11061 34376
rect 11019 34327 11061 34336
rect 11403 34376 11445 34385
rect 12459 34381 12501 34390
rect 11403 34336 11404 34376
rect 11444 34336 11445 34376
rect 11403 34327 11445 34336
rect 11971 34376 12029 34377
rect 11971 34336 11980 34376
rect 12020 34336 12029 34376
rect 11971 34335 12029 34336
rect 12459 34341 12460 34381
rect 12500 34341 12501 34381
rect 12459 34332 12501 34341
rect 13027 34376 13085 34377
rect 13027 34336 13036 34376
rect 13076 34336 13085 34376
rect 13027 34335 13085 34336
rect 14275 34376 14333 34377
rect 14275 34336 14284 34376
rect 14324 34336 14333 34376
rect 14275 34335 14333 34336
rect 14667 34376 14709 34385
rect 14667 34336 14668 34376
rect 14708 34336 14709 34376
rect 14667 34327 14709 34336
rect 14859 34376 14901 34385
rect 14859 34336 14860 34376
rect 14900 34336 14901 34376
rect 14859 34327 14901 34336
rect 14947 34376 15005 34377
rect 14947 34336 14956 34376
rect 14996 34336 15005 34376
rect 14947 34335 15005 34336
rect 16675 34376 16733 34377
rect 16675 34336 16684 34376
rect 16724 34336 16733 34376
rect 16675 34335 16733 34336
rect 17059 34376 17117 34377
rect 17059 34336 17068 34376
rect 17108 34336 17117 34376
rect 17059 34335 17117 34336
rect 18307 34376 18365 34377
rect 18307 34336 18316 34376
rect 18356 34336 18365 34376
rect 18307 34335 18365 34336
rect 18691 34376 18749 34377
rect 18691 34336 18700 34376
rect 18740 34336 18749 34376
rect 19939 34357 19948 34397
rect 19988 34357 19997 34397
rect 19939 34356 19997 34357
rect 18691 34335 18749 34336
rect 15427 34334 15485 34335
rect 7563 34306 7605 34315
rect 3531 34292 3573 34301
rect 3531 34252 3532 34292
rect 3572 34252 3573 34292
rect 3531 34243 3573 34252
rect 12651 34292 12693 34301
rect 15427 34294 15436 34334
rect 15476 34294 15485 34334
rect 15427 34293 15485 34294
rect 12651 34252 12652 34292
rect 12692 34252 12693 34292
rect 12651 34243 12693 34252
rect 1227 34208 1269 34217
rect 1227 34168 1228 34208
rect 1268 34168 1269 34208
rect 1227 34159 1269 34168
rect 2955 34208 2997 34217
rect 2955 34168 2956 34208
rect 2996 34168 2997 34208
rect 2955 34159 2997 34168
rect 7363 34208 7421 34209
rect 7363 34168 7372 34208
rect 7412 34168 7421 34208
rect 7363 34167 7421 34168
rect 9675 34208 9717 34217
rect 9675 34168 9676 34208
rect 9716 34168 9717 34208
rect 9675 34159 9717 34168
rect 9859 34208 9917 34209
rect 9859 34168 9868 34208
rect 9908 34168 9917 34208
rect 9859 34167 9917 34168
rect 10627 34208 10685 34209
rect 10627 34168 10636 34208
rect 10676 34168 10685 34208
rect 10627 34167 10685 34168
rect 15139 34208 15197 34209
rect 15139 34168 15148 34208
rect 15188 34168 15197 34208
rect 15139 34167 15197 34168
rect 16875 34208 16917 34217
rect 16875 34168 16876 34208
rect 16916 34168 16917 34208
rect 16875 34159 16917 34168
rect 18507 34208 18549 34217
rect 18507 34168 18508 34208
rect 18548 34168 18549 34208
rect 18507 34159 18549 34168
rect 20139 34208 20181 34217
rect 20139 34168 20140 34208
rect 20180 34168 20181 34208
rect 20139 34159 20181 34168
rect 1152 34040 20452 34064
rect 1152 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20452 34040
rect 1152 33976 20452 34000
rect 3523 33872 3581 33873
rect 3523 33832 3532 33872
rect 3572 33832 3581 33872
rect 3523 33831 3581 33832
rect 3811 33872 3869 33873
rect 3811 33832 3820 33872
rect 3860 33832 3869 33872
rect 3811 33831 3869 33832
rect 4395 33872 4437 33881
rect 4395 33832 4396 33872
rect 4436 33832 4437 33872
rect 4395 33823 4437 33832
rect 4675 33872 4733 33873
rect 4675 33832 4684 33872
rect 4724 33832 4733 33872
rect 4675 33831 4733 33832
rect 11979 33872 12021 33881
rect 11979 33832 11980 33872
rect 12020 33832 12021 33872
rect 11979 33823 12021 33832
rect 15435 33872 15477 33881
rect 15435 33832 15436 33872
rect 15476 33832 15477 33872
rect 15435 33823 15477 33832
rect 19275 33872 19317 33881
rect 19275 33832 19276 33872
rect 19316 33832 19317 33872
rect 19275 33823 19317 33832
rect 1323 33704 1365 33713
rect 1323 33664 1324 33704
rect 1364 33664 1365 33704
rect 1323 33655 1365 33664
rect 1419 33704 1461 33713
rect 1419 33664 1420 33704
rect 1460 33664 1461 33704
rect 1419 33655 1461 33664
rect 1611 33704 1653 33713
rect 1611 33664 1612 33704
rect 1652 33664 1653 33704
rect 1611 33655 1653 33664
rect 1891 33704 1949 33705
rect 1891 33664 1900 33704
rect 1940 33664 1949 33704
rect 1891 33663 1949 33664
rect 3139 33704 3197 33705
rect 3139 33664 3148 33704
rect 3188 33664 3197 33704
rect 3139 33663 3197 33664
rect 4011 33704 4053 33713
rect 4011 33664 4012 33704
rect 4052 33664 4053 33704
rect 4011 33655 4053 33664
rect 4107 33704 4149 33713
rect 4107 33664 4108 33704
rect 4148 33664 4149 33704
rect 4107 33655 4149 33664
rect 4867 33704 4925 33705
rect 4867 33664 4876 33704
rect 4916 33664 4925 33704
rect 4867 33663 4925 33664
rect 6115 33704 6173 33705
rect 6115 33664 6124 33704
rect 6164 33664 6173 33704
rect 6115 33663 6173 33664
rect 6499 33704 6557 33705
rect 6499 33664 6508 33704
rect 6548 33664 6557 33704
rect 6499 33663 6557 33664
rect 6603 33704 6645 33713
rect 6603 33664 6604 33704
rect 6644 33664 6645 33704
rect 6603 33655 6645 33664
rect 6795 33704 6837 33713
rect 6795 33664 6796 33704
rect 6836 33664 6837 33704
rect 6795 33655 6837 33664
rect 7267 33704 7325 33705
rect 7267 33664 7276 33704
rect 7316 33664 7325 33704
rect 7267 33663 7325 33664
rect 8515 33704 8573 33705
rect 8515 33664 8524 33704
rect 8564 33664 8573 33704
rect 8515 33663 8573 33664
rect 8899 33704 8957 33705
rect 8899 33664 8908 33704
rect 8948 33664 8957 33704
rect 8899 33663 8957 33664
rect 10147 33704 10205 33705
rect 10147 33664 10156 33704
rect 10196 33664 10205 33704
rect 10147 33663 10205 33664
rect 10531 33704 10589 33705
rect 10531 33664 10540 33704
rect 10580 33664 10589 33704
rect 12355 33704 12413 33705
rect 10531 33663 10589 33664
rect 11779 33683 11837 33684
rect 11779 33643 11788 33683
rect 11828 33643 11837 33683
rect 12355 33664 12364 33704
rect 12404 33664 12413 33704
rect 12355 33663 12413 33664
rect 13603 33704 13661 33705
rect 13603 33664 13612 33704
rect 13652 33664 13661 33704
rect 13603 33663 13661 33664
rect 13987 33704 14045 33705
rect 13987 33664 13996 33704
rect 14036 33664 14045 33704
rect 13987 33663 14045 33664
rect 15235 33704 15293 33705
rect 15235 33664 15244 33704
rect 15284 33664 15293 33704
rect 15235 33663 15293 33664
rect 15619 33704 15677 33705
rect 15619 33664 15628 33704
rect 15668 33664 15677 33704
rect 15619 33663 15677 33664
rect 16867 33704 16925 33705
rect 16867 33664 16876 33704
rect 16916 33664 16925 33704
rect 16867 33663 16925 33664
rect 17547 33704 17589 33713
rect 17547 33664 17548 33704
rect 17588 33664 17589 33704
rect 17547 33655 17589 33664
rect 17643 33704 17685 33713
rect 17643 33664 17644 33704
rect 17684 33664 17685 33704
rect 17643 33655 17685 33664
rect 18595 33704 18653 33705
rect 18595 33664 18604 33704
rect 18644 33664 18653 33704
rect 18595 33663 18653 33664
rect 19083 33699 19125 33708
rect 19083 33659 19084 33699
rect 19124 33659 19125 33699
rect 19083 33650 19125 33659
rect 11779 33642 11837 33643
rect 18027 33620 18069 33629
rect 18027 33580 18028 33620
rect 18068 33580 18069 33620
rect 18027 33571 18069 33580
rect 18123 33620 18165 33629
rect 18123 33580 18124 33620
rect 18164 33580 18165 33620
rect 18123 33571 18165 33580
rect 19467 33620 19509 33629
rect 19467 33580 19468 33620
rect 19508 33580 19509 33620
rect 19467 33571 19509 33580
rect 19747 33620 19805 33621
rect 19747 33580 19756 33620
rect 19796 33580 19805 33620
rect 19747 33579 19805 33580
rect 1411 33536 1469 33537
rect 1411 33496 1420 33536
rect 1460 33496 1469 33536
rect 1411 33495 1469 33496
rect 20139 33536 20181 33545
rect 20139 33496 20140 33536
rect 20180 33496 20181 33536
rect 20139 33487 20181 33496
rect 3339 33452 3381 33461
rect 3339 33412 3340 33452
rect 3380 33412 3381 33452
rect 3339 33403 3381 33412
rect 6315 33452 6357 33461
rect 6315 33412 6316 33452
rect 6356 33412 6357 33452
rect 6315 33403 6357 33412
rect 6795 33452 6837 33461
rect 6795 33412 6796 33452
rect 6836 33412 6837 33452
rect 6795 33403 6837 33412
rect 7083 33452 7125 33461
rect 7083 33412 7084 33452
rect 7124 33412 7125 33452
rect 7083 33403 7125 33412
rect 10347 33452 10389 33461
rect 10347 33412 10348 33452
rect 10388 33412 10389 33452
rect 10347 33403 10389 33412
rect 13803 33452 13845 33461
rect 13803 33412 13804 33452
rect 13844 33412 13845 33452
rect 13803 33403 13845 33412
rect 17067 33452 17109 33461
rect 17067 33412 17068 33452
rect 17108 33412 17109 33452
rect 17067 33403 17109 33412
rect 19947 33452 19989 33461
rect 19947 33412 19948 33452
rect 19988 33412 19989 33452
rect 19947 33403 19989 33412
rect 1152 33284 20352 33308
rect 1152 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 20352 33284
rect 1152 33220 20352 33244
rect 2379 33116 2421 33125
rect 2379 33076 2380 33116
rect 2420 33076 2421 33116
rect 2379 33067 2421 33076
rect 10443 33116 10485 33125
rect 10443 33076 10444 33116
rect 10484 33076 10485 33116
rect 10443 33067 10485 33076
rect 11307 33116 11349 33125
rect 11307 33076 11308 33116
rect 11348 33076 11349 33116
rect 11307 33067 11349 33076
rect 16107 33116 16149 33125
rect 16107 33076 16108 33116
rect 16148 33076 16149 33116
rect 16107 33067 16149 33076
rect 19083 33116 19125 33125
rect 19083 33076 19084 33116
rect 19124 33076 19125 33116
rect 19083 33067 19125 33076
rect 4683 33032 4725 33041
rect 4683 32992 4684 33032
rect 4724 32992 4725 33032
rect 4683 32983 4725 32992
rect 12363 33032 12405 33041
rect 12363 32992 12364 33032
rect 12404 32992 12405 33032
rect 12363 32983 12405 32992
rect 20139 33032 20181 33041
rect 20139 32992 20140 33032
rect 20180 32992 20181 33032
rect 20139 32983 20181 32992
rect 2179 32948 2237 32949
rect 2179 32908 2188 32948
rect 2228 32908 2237 32948
rect 2179 32907 2237 32908
rect 3147 32948 3189 32957
rect 3147 32908 3148 32948
rect 3188 32908 3189 32948
rect 14283 32948 14325 32957
rect 3147 32899 3189 32908
rect 6651 32906 6693 32915
rect 1960 32879 2002 32888
rect 1411 32864 1469 32865
rect 1411 32824 1420 32864
rect 1460 32824 1469 32864
rect 1411 32823 1469 32824
rect 1507 32864 1565 32865
rect 1507 32824 1516 32864
rect 1556 32824 1565 32864
rect 1507 32823 1565 32824
rect 1707 32864 1749 32873
rect 1707 32824 1708 32864
rect 1748 32824 1749 32864
rect 1707 32815 1749 32824
rect 1803 32864 1845 32873
rect 1803 32824 1804 32864
rect 1844 32824 1845 32864
rect 1960 32839 1961 32879
rect 2001 32839 2002 32879
rect 4203 32878 4245 32887
rect 1960 32830 2002 32839
rect 2667 32864 2709 32873
rect 1803 32815 1845 32824
rect 2667 32824 2668 32864
rect 2708 32824 2709 32864
rect 2667 32815 2709 32824
rect 2763 32864 2805 32873
rect 2763 32824 2764 32864
rect 2804 32824 2805 32864
rect 2763 32815 2805 32824
rect 3243 32864 3285 32873
rect 3243 32824 3244 32864
rect 3284 32824 3285 32864
rect 3243 32815 3285 32824
rect 3715 32864 3773 32865
rect 3715 32824 3724 32864
rect 3764 32824 3773 32864
rect 4203 32838 4204 32878
rect 4244 32838 4245 32878
rect 6651 32866 6652 32906
rect 6692 32866 6693 32906
rect 14283 32908 14284 32948
rect 14324 32908 14325 32948
rect 14283 32899 14325 32908
rect 19363 32948 19421 32949
rect 19363 32908 19372 32948
rect 19412 32908 19421 32948
rect 19363 32907 19421 32908
rect 19747 32948 19805 32949
rect 19747 32908 19756 32948
rect 19796 32908 19805 32948
rect 19747 32907 19805 32908
rect 15243 32878 15285 32887
rect 4203 32829 4245 32838
rect 4867 32864 4925 32865
rect 3715 32823 3773 32824
rect 4867 32824 4876 32864
rect 4916 32824 4925 32864
rect 4867 32823 4925 32824
rect 6115 32864 6173 32865
rect 6115 32824 6124 32864
rect 6164 32824 6173 32864
rect 6651 32857 6693 32866
rect 7171 32864 7229 32865
rect 6115 32823 6173 32824
rect 7171 32824 7180 32864
rect 7220 32824 7229 32864
rect 7171 32823 7229 32824
rect 7659 32864 7701 32873
rect 7659 32824 7660 32864
rect 7700 32824 7701 32864
rect 7659 32815 7701 32824
rect 7755 32864 7797 32873
rect 7755 32824 7756 32864
rect 7796 32824 7797 32864
rect 7755 32815 7797 32824
rect 8139 32864 8181 32873
rect 8139 32824 8140 32864
rect 8180 32824 8181 32864
rect 8139 32815 8181 32824
rect 8235 32864 8277 32873
rect 8235 32824 8236 32864
rect 8276 32824 8277 32864
rect 8235 32815 8277 32824
rect 8715 32864 8757 32873
rect 8715 32824 8716 32864
rect 8756 32824 8757 32864
rect 8715 32815 8757 32824
rect 8811 32864 8853 32873
rect 8811 32824 8812 32864
rect 8852 32824 8853 32864
rect 8811 32815 8853 32824
rect 8995 32864 9053 32865
rect 8995 32824 9004 32864
rect 9044 32824 9053 32864
rect 8995 32823 9053 32824
rect 10243 32864 10301 32865
rect 10243 32824 10252 32864
rect 10292 32824 10301 32864
rect 10243 32823 10301 32824
rect 10627 32864 10685 32865
rect 10627 32824 10636 32864
rect 10676 32824 10685 32864
rect 10627 32823 10685 32824
rect 11587 32864 11645 32865
rect 11587 32824 11596 32864
rect 11636 32824 11645 32864
rect 11587 32823 11645 32824
rect 11971 32864 12029 32865
rect 11971 32824 11980 32864
rect 12020 32824 12029 32864
rect 11971 32823 12029 32824
rect 12075 32864 12117 32873
rect 12075 32824 12076 32864
rect 12116 32824 12117 32864
rect 12075 32815 12117 32824
rect 12747 32864 12789 32873
rect 12747 32824 12748 32864
rect 12788 32824 12789 32864
rect 12747 32815 12789 32824
rect 12843 32864 12885 32873
rect 12843 32824 12844 32864
rect 12884 32824 12885 32864
rect 12843 32815 12885 32824
rect 13035 32864 13077 32873
rect 13035 32824 13036 32864
rect 13076 32824 13077 32864
rect 13035 32815 13077 32824
rect 13323 32864 13365 32873
rect 13323 32824 13324 32864
rect 13364 32824 13365 32864
rect 13323 32815 13365 32824
rect 13707 32864 13749 32873
rect 13707 32824 13708 32864
rect 13748 32824 13749 32864
rect 13707 32815 13749 32824
rect 13803 32864 13845 32873
rect 13803 32824 13804 32864
rect 13844 32824 13845 32864
rect 13803 32815 13845 32824
rect 14187 32864 14229 32873
rect 14187 32824 14188 32864
rect 14228 32824 14229 32864
rect 14187 32815 14229 32824
rect 14755 32864 14813 32865
rect 14755 32824 14764 32864
rect 14804 32824 14813 32864
rect 15243 32838 15244 32878
rect 15284 32838 15285 32878
rect 18507 32878 18549 32887
rect 15243 32829 15285 32838
rect 15627 32864 15669 32873
rect 14755 32823 14813 32824
rect 15627 32824 15628 32864
rect 15668 32824 15669 32864
rect 15627 32815 15669 32824
rect 15723 32864 15765 32873
rect 15723 32824 15724 32864
rect 15764 32824 15765 32864
rect 15915 32864 15957 32873
rect 15723 32815 15765 32824
rect 15819 32843 15861 32852
rect 15819 32803 15820 32843
rect 15860 32803 15861 32843
rect 15915 32824 15916 32864
rect 15956 32824 15957 32864
rect 15915 32815 15957 32824
rect 16107 32864 16149 32873
rect 16107 32824 16108 32864
rect 16148 32824 16149 32864
rect 16387 32864 16445 32865
rect 16107 32815 16149 32824
rect 16299 32822 16341 32831
rect 16387 32824 16396 32864
rect 16436 32824 16445 32864
rect 16387 32823 16445 32824
rect 16971 32864 17013 32873
rect 16971 32824 16972 32864
rect 17012 32824 17013 32864
rect 15819 32794 15861 32803
rect 4395 32780 4437 32789
rect 4395 32740 4396 32780
rect 4436 32740 4437 32780
rect 4395 32731 4437 32740
rect 6315 32780 6357 32789
rect 6315 32740 6316 32780
rect 6356 32740 6357 32780
rect 6315 32731 6357 32740
rect 13131 32780 13173 32789
rect 13131 32740 13132 32780
rect 13172 32740 13173 32780
rect 13131 32731 13173 32740
rect 15435 32780 15477 32789
rect 15435 32740 15436 32780
rect 15476 32740 15477 32780
rect 16299 32782 16300 32822
rect 16340 32782 16341 32822
rect 16971 32815 17013 32824
rect 17067 32864 17109 32873
rect 17067 32824 17068 32864
rect 17108 32824 17109 32864
rect 17067 32815 17109 32824
rect 17451 32864 17493 32873
rect 17451 32824 17452 32864
rect 17492 32824 17493 32864
rect 17451 32815 17493 32824
rect 17547 32864 17589 32873
rect 17547 32824 17548 32864
rect 17588 32824 17589 32864
rect 17547 32815 17589 32824
rect 18019 32864 18077 32865
rect 18019 32824 18028 32864
rect 18068 32824 18077 32864
rect 18507 32838 18508 32878
rect 18548 32838 18549 32878
rect 18507 32829 18549 32838
rect 18891 32864 18933 32873
rect 18019 32823 18077 32824
rect 18891 32824 18892 32864
rect 18932 32824 18933 32864
rect 18891 32815 18933 32824
rect 19083 32864 19125 32873
rect 19083 32824 19084 32864
rect 19124 32824 19125 32864
rect 19083 32815 19125 32824
rect 16299 32773 16341 32782
rect 18699 32780 18741 32789
rect 15435 32731 15477 32740
rect 18699 32740 18700 32780
rect 18740 32740 18741 32780
rect 18699 32731 18741 32740
rect 1891 32696 1949 32697
rect 1891 32656 1900 32696
rect 1940 32656 1949 32696
rect 8515 32696 8573 32697
rect 1891 32655 1949 32656
rect 6507 32654 6549 32663
rect 8515 32656 8524 32696
rect 8564 32656 8573 32696
rect 8515 32655 8573 32656
rect 10443 32696 10485 32705
rect 10443 32656 10444 32696
rect 10484 32656 10485 32696
rect 6507 32614 6508 32654
rect 6548 32614 6549 32654
rect 10443 32647 10485 32656
rect 12547 32696 12605 32697
rect 12547 32656 12556 32696
rect 12596 32656 12605 32696
rect 12547 32655 12605 32656
rect 19563 32696 19605 32705
rect 19563 32656 19564 32696
rect 19604 32656 19605 32696
rect 19563 32647 19605 32656
rect 19947 32696 19989 32705
rect 19947 32656 19948 32696
rect 19988 32656 19989 32696
rect 19947 32647 19989 32656
rect 6507 32605 6549 32614
rect 11883 32638 11925 32647
rect 11883 32598 11884 32638
rect 11924 32598 11925 32638
rect 11883 32589 11925 32598
rect 1152 32528 20452 32552
rect 1152 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20452 32528
rect 1152 32464 20452 32488
rect 2859 32360 2901 32369
rect 2859 32320 2860 32360
rect 2900 32320 2901 32360
rect 2859 32311 2901 32320
rect 3243 32360 3285 32369
rect 3243 32320 3244 32360
rect 3284 32320 3285 32360
rect 3243 32311 3285 32320
rect 10539 32360 10581 32369
rect 10539 32320 10540 32360
rect 10580 32320 10581 32360
rect 10539 32311 10581 32320
rect 12259 32360 12317 32361
rect 12259 32320 12268 32360
rect 12308 32320 12317 32360
rect 12259 32319 12317 32320
rect 13131 32360 13173 32369
rect 13131 32320 13132 32360
rect 13172 32320 13173 32360
rect 13131 32311 13173 32320
rect 14467 32360 14525 32361
rect 14467 32320 14476 32360
rect 14516 32320 14525 32360
rect 14467 32319 14525 32320
rect 19179 32360 19221 32369
rect 19179 32320 19180 32360
rect 19220 32320 19221 32360
rect 19179 32311 19221 32320
rect 6699 32276 6741 32285
rect 6699 32236 6700 32276
rect 6740 32236 6741 32276
rect 6699 32227 6741 32236
rect 6891 32276 6933 32285
rect 6891 32236 6892 32276
rect 6932 32236 6933 32276
rect 6891 32227 6933 32236
rect 1219 32192 1277 32193
rect 1219 32152 1228 32192
rect 1268 32152 1277 32192
rect 1219 32151 1277 32152
rect 2467 32192 2525 32193
rect 2467 32152 2476 32192
rect 2516 32152 2525 32192
rect 2467 32151 2525 32152
rect 3435 32187 3477 32196
rect 3435 32147 3436 32187
rect 3476 32147 3477 32187
rect 3907 32192 3965 32193
rect 3907 32152 3916 32192
rect 3956 32152 3965 32192
rect 3907 32151 3965 32152
rect 4875 32192 4917 32201
rect 4875 32152 4876 32192
rect 4916 32152 4917 32192
rect 3435 32138 3477 32147
rect 4875 32143 4917 32152
rect 4971 32192 5013 32201
rect 4971 32152 4972 32192
rect 5012 32152 5013 32192
rect 4971 32143 5013 32152
rect 5251 32192 5309 32193
rect 5251 32152 5260 32192
rect 5300 32152 5309 32192
rect 5251 32151 5309 32152
rect 6499 32192 6557 32193
rect 6499 32152 6508 32192
rect 6548 32152 6557 32192
rect 6499 32151 6557 32152
rect 7083 32187 7125 32196
rect 7083 32147 7084 32187
rect 7124 32147 7125 32187
rect 7555 32192 7613 32193
rect 7555 32152 7564 32192
rect 7604 32152 7613 32192
rect 7555 32151 7613 32152
rect 8043 32192 8085 32201
rect 8043 32152 8044 32192
rect 8084 32152 8085 32192
rect 7083 32138 7125 32147
rect 8043 32143 8085 32152
rect 8523 32192 8565 32201
rect 8523 32152 8524 32192
rect 8564 32152 8565 32192
rect 8523 32143 8565 32152
rect 8619 32192 8661 32201
rect 8619 32152 8620 32192
rect 8660 32152 8661 32192
rect 8619 32143 8661 32152
rect 9091 32192 9149 32193
rect 9091 32152 9100 32192
rect 9140 32152 9149 32192
rect 9091 32151 9149 32152
rect 10339 32192 10397 32193
rect 10339 32152 10348 32192
rect 10388 32152 10397 32192
rect 10339 32151 10397 32152
rect 10819 32192 10877 32193
rect 10819 32152 10828 32192
rect 10868 32152 10877 32192
rect 10819 32151 10877 32152
rect 11115 32192 11157 32201
rect 11115 32152 11116 32192
rect 11156 32152 11157 32192
rect 11115 32143 11157 32152
rect 11211 32192 11253 32201
rect 11211 32152 11212 32192
rect 11252 32152 11253 32192
rect 11211 32143 11253 32152
rect 11691 32192 11733 32201
rect 11691 32152 11692 32192
rect 11732 32152 11733 32192
rect 11691 32143 11733 32152
rect 11883 32192 11925 32201
rect 11883 32152 11884 32192
rect 11924 32152 11925 32192
rect 11883 32143 11925 32152
rect 11971 32192 12029 32193
rect 11971 32152 11980 32192
rect 12020 32152 12029 32192
rect 11971 32151 12029 32152
rect 12171 32192 12213 32201
rect 12171 32152 12172 32192
rect 12212 32152 12213 32192
rect 12171 32143 12213 32152
rect 12363 32192 12405 32201
rect 12363 32152 12364 32192
rect 12404 32152 12405 32192
rect 12363 32143 12405 32152
rect 12451 32192 12509 32193
rect 12451 32152 12460 32192
rect 12500 32152 12509 32192
rect 12451 32151 12509 32152
rect 12643 32192 12701 32193
rect 12643 32152 12652 32192
rect 12692 32152 12701 32192
rect 12643 32151 12701 32152
rect 12747 32192 12789 32201
rect 12747 32152 12748 32192
rect 12788 32152 12789 32192
rect 12747 32143 12789 32152
rect 12939 32192 12981 32201
rect 12939 32152 12940 32192
rect 12980 32152 12981 32192
rect 12939 32143 12981 32152
rect 13323 32192 13365 32201
rect 13323 32152 13324 32192
rect 13364 32152 13365 32192
rect 13323 32143 13365 32152
rect 13707 32192 13749 32201
rect 13707 32152 13708 32192
rect 13748 32152 13749 32192
rect 13707 32143 13749 32152
rect 13995 32192 14037 32201
rect 13995 32152 13996 32192
rect 14036 32152 14037 32192
rect 13995 32143 14037 32152
rect 14379 32192 14421 32201
rect 14379 32152 14380 32192
rect 14420 32152 14421 32192
rect 14379 32143 14421 32152
rect 14571 32192 14613 32201
rect 14571 32152 14572 32192
rect 14612 32152 14613 32192
rect 14571 32143 14613 32152
rect 14659 32192 14717 32193
rect 14659 32152 14668 32192
rect 14708 32152 14717 32192
rect 14659 32151 14717 32152
rect 15051 32192 15093 32201
rect 15051 32152 15052 32192
rect 15092 32152 15093 32192
rect 15051 32143 15093 32152
rect 15147 32192 15189 32201
rect 15147 32152 15148 32192
rect 15188 32152 15189 32192
rect 15147 32143 15189 32152
rect 15243 32192 15285 32201
rect 15243 32152 15244 32192
rect 15284 32152 15285 32192
rect 15243 32143 15285 32152
rect 15339 32192 15381 32201
rect 15339 32152 15340 32192
rect 15380 32152 15381 32192
rect 15339 32143 15381 32152
rect 15531 32192 15573 32201
rect 15531 32152 15532 32192
rect 15572 32152 15573 32192
rect 15531 32143 15573 32152
rect 15723 32192 15765 32201
rect 15723 32152 15724 32192
rect 15764 32152 15765 32192
rect 15723 32143 15765 32152
rect 15811 32192 15869 32193
rect 15811 32152 15820 32192
rect 15860 32152 15869 32192
rect 15811 32151 15869 32152
rect 16195 32192 16253 32193
rect 16195 32152 16204 32192
rect 16244 32152 16253 32192
rect 17835 32192 17877 32201
rect 16195 32151 16253 32152
rect 17443 32171 17501 32172
rect 17443 32131 17452 32171
rect 17492 32131 17501 32171
rect 17835 32152 17836 32192
rect 17876 32152 17877 32192
rect 17835 32143 17877 32152
rect 18027 32192 18069 32201
rect 18027 32152 18028 32192
rect 18068 32152 18069 32192
rect 18027 32143 18069 32152
rect 18219 32192 18261 32201
rect 18219 32152 18220 32192
rect 18260 32152 18261 32192
rect 18219 32143 18261 32152
rect 18411 32192 18453 32201
rect 18411 32152 18412 32192
rect 18452 32152 18453 32192
rect 18411 32143 18453 32152
rect 17443 32130 17501 32131
rect 3043 32108 3101 32109
rect 3043 32068 3052 32108
rect 3092 32068 3101 32108
rect 3043 32067 3101 32068
rect 4395 32108 4437 32117
rect 4395 32068 4396 32108
rect 4436 32068 4437 32108
rect 4395 32059 4437 32068
rect 4491 32108 4533 32117
rect 4491 32068 4492 32108
rect 4532 32068 4533 32108
rect 4491 32059 4533 32068
rect 8139 32108 8181 32117
rect 8139 32068 8140 32108
rect 8180 32068 8181 32108
rect 8139 32059 8181 32068
rect 18595 32108 18653 32109
rect 18595 32068 18604 32108
rect 18644 32068 18653 32108
rect 18595 32067 18653 32068
rect 18979 32108 19037 32109
rect 18979 32068 18988 32108
rect 19028 32068 19037 32108
rect 18979 32067 19037 32068
rect 19363 32108 19421 32109
rect 19363 32068 19372 32108
rect 19412 32068 19421 32108
rect 19363 32067 19421 32068
rect 19747 32108 19805 32109
rect 19747 32068 19756 32108
rect 19796 32068 19805 32108
rect 19747 32067 19805 32068
rect 11491 32024 11549 32025
rect 11491 31984 11500 32024
rect 11540 31984 11549 32024
rect 11491 31983 11549 31984
rect 13323 32024 13365 32033
rect 13323 31984 13324 32024
rect 13364 31984 13365 32024
rect 13323 31975 13365 31984
rect 13995 32024 14037 32033
rect 13995 31984 13996 32024
rect 14036 31984 14037 32024
rect 13995 31975 14037 31984
rect 18027 32024 18069 32033
rect 18027 31984 18028 32024
rect 18068 31984 18069 32024
rect 18027 31975 18069 31984
rect 18219 32024 18261 32033
rect 18219 31984 18220 32024
rect 18260 31984 18261 32024
rect 18219 31975 18261 31984
rect 2667 31940 2709 31949
rect 2667 31900 2668 31940
rect 2708 31900 2709 31940
rect 2667 31891 2709 31900
rect 11691 31940 11733 31949
rect 11691 31900 11692 31940
rect 11732 31900 11733 31940
rect 11691 31891 11733 31900
rect 12939 31940 12981 31949
rect 12939 31900 12940 31940
rect 12980 31900 12981 31940
rect 12939 31891 12981 31900
rect 15531 31940 15573 31949
rect 15531 31900 15532 31940
rect 15572 31900 15573 31940
rect 15531 31891 15573 31900
rect 17643 31940 17685 31949
rect 17643 31900 17644 31940
rect 17684 31900 17685 31940
rect 17643 31891 17685 31900
rect 18795 31940 18837 31949
rect 18795 31900 18796 31940
rect 18836 31900 18837 31940
rect 18795 31891 18837 31900
rect 19563 31940 19605 31949
rect 19563 31900 19564 31940
rect 19604 31900 19605 31940
rect 19563 31891 19605 31900
rect 19947 31940 19989 31949
rect 19947 31900 19948 31940
rect 19988 31900 19989 31940
rect 19947 31891 19989 31900
rect 1152 31772 20352 31796
rect 1152 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 20352 31772
rect 1152 31708 20352 31732
rect 4587 31604 4629 31613
rect 4587 31564 4588 31604
rect 4628 31564 4629 31604
rect 4587 31555 4629 31564
rect 4779 31604 4821 31613
rect 4779 31564 4780 31604
rect 4820 31564 4821 31604
rect 4779 31555 4821 31564
rect 17067 31604 17109 31613
rect 17067 31564 17068 31604
rect 17108 31564 17109 31604
rect 17067 31555 17109 31564
rect 8043 31520 8085 31529
rect 8043 31480 8044 31520
rect 8084 31480 8085 31520
rect 8043 31471 8085 31480
rect 8427 31520 8469 31529
rect 8427 31480 8428 31520
rect 8468 31480 8469 31520
rect 8427 31471 8469 31480
rect 8811 31520 8853 31529
rect 8811 31480 8812 31520
rect 8852 31480 8853 31520
rect 8811 31471 8853 31480
rect 10539 31520 10581 31529
rect 10539 31480 10540 31520
rect 10580 31480 10581 31520
rect 10539 31471 10581 31480
rect 16299 31520 16341 31529
rect 16299 31480 16300 31520
rect 16340 31480 16341 31520
rect 16299 31471 16341 31480
rect 8331 31436 8373 31445
rect 8331 31396 8332 31436
rect 8372 31396 8373 31436
rect 8331 31387 8373 31396
rect 8523 31436 8565 31445
rect 8523 31396 8524 31436
rect 8564 31396 8565 31436
rect 8523 31387 8565 31396
rect 13131 31436 13173 31445
rect 13131 31396 13132 31436
rect 13172 31396 13173 31436
rect 13131 31387 13173 31396
rect 18027 31436 18069 31445
rect 18027 31396 18028 31436
rect 18068 31396 18069 31436
rect 16675 31394 16733 31395
rect 1219 31352 1277 31353
rect 1219 31312 1228 31352
rect 1268 31312 1277 31352
rect 1219 31311 1277 31312
rect 2467 31352 2525 31353
rect 2467 31312 2476 31352
rect 2516 31312 2525 31352
rect 2467 31311 2525 31312
rect 3139 31352 3197 31353
rect 3139 31312 3148 31352
rect 3188 31312 3197 31352
rect 3139 31311 3197 31312
rect 4387 31352 4445 31353
rect 4387 31312 4396 31352
rect 4436 31312 4445 31352
rect 4387 31311 4445 31312
rect 4963 31352 5021 31353
rect 4963 31312 4972 31352
rect 5012 31312 5021 31352
rect 4963 31311 5021 31312
rect 6211 31352 6269 31353
rect 6211 31312 6220 31352
rect 6260 31312 6269 31352
rect 6211 31311 6269 31312
rect 6595 31352 6653 31353
rect 6595 31312 6604 31352
rect 6644 31312 6653 31352
rect 6595 31311 6653 31312
rect 7843 31352 7901 31353
rect 7843 31312 7852 31352
rect 7892 31312 7901 31352
rect 7843 31311 7901 31312
rect 8235 31352 8277 31361
rect 8235 31312 8236 31352
rect 8276 31312 8277 31352
rect 8235 31303 8277 31312
rect 8611 31352 8669 31353
rect 8611 31312 8620 31352
rect 8660 31312 8669 31352
rect 8611 31311 8669 31312
rect 9091 31352 9149 31353
rect 9091 31312 9100 31352
rect 9140 31312 9149 31352
rect 9091 31311 9149 31312
rect 10339 31352 10397 31353
rect 10339 31312 10348 31352
rect 10388 31312 10397 31352
rect 10339 31311 10397 31312
rect 10915 31352 10973 31353
rect 10915 31312 10924 31352
rect 10964 31312 10973 31352
rect 10915 31311 10973 31312
rect 12163 31352 12221 31353
rect 12163 31312 12172 31352
rect 12212 31312 12221 31352
rect 12163 31311 12221 31312
rect 12651 31352 12693 31361
rect 12651 31312 12652 31352
rect 12692 31312 12693 31352
rect 12651 31303 12693 31312
rect 12747 31352 12789 31361
rect 12747 31312 12748 31352
rect 12788 31312 12789 31352
rect 12747 31303 12789 31312
rect 13227 31352 13269 31361
rect 14187 31357 14229 31366
rect 13227 31312 13228 31352
rect 13268 31312 13269 31352
rect 13227 31303 13269 31312
rect 13699 31352 13757 31353
rect 13699 31312 13708 31352
rect 13748 31312 13757 31352
rect 13699 31311 13757 31312
rect 14187 31317 14188 31357
rect 14228 31317 14229 31357
rect 14187 31308 14229 31317
rect 14851 31352 14909 31353
rect 14851 31312 14860 31352
rect 14900 31312 14909 31352
rect 14851 31311 14909 31312
rect 16099 31352 16157 31353
rect 16099 31312 16108 31352
rect 16148 31312 16157 31352
rect 16099 31311 16157 31312
rect 16491 31352 16533 31361
rect 16491 31312 16492 31352
rect 16532 31312 16533 31352
rect 16491 31303 16533 31312
rect 16587 31352 16629 31361
rect 16675 31354 16684 31394
rect 16724 31354 16733 31394
rect 18027 31387 18069 31396
rect 18123 31436 18165 31445
rect 18123 31396 18124 31436
rect 18164 31396 18165 31436
rect 18123 31387 18165 31396
rect 19459 31436 19517 31437
rect 19459 31396 19468 31436
rect 19508 31396 19517 31436
rect 19459 31395 19517 31396
rect 19843 31436 19901 31437
rect 19843 31396 19852 31436
rect 19892 31396 19901 31436
rect 19843 31395 19901 31396
rect 19131 31361 19173 31370
rect 16675 31353 16733 31354
rect 16587 31312 16588 31352
rect 16628 31312 16629 31352
rect 16587 31303 16629 31312
rect 16963 31352 17021 31353
rect 16963 31312 16972 31352
rect 17012 31312 17021 31352
rect 17547 31352 17589 31361
rect 16963 31311 17021 31312
rect 17163 31339 17205 31348
rect 17163 31299 17164 31339
rect 17204 31299 17205 31339
rect 17547 31312 17548 31352
rect 17588 31312 17589 31352
rect 17547 31303 17589 31312
rect 17643 31352 17685 31361
rect 17643 31312 17644 31352
rect 17684 31312 17685 31352
rect 17643 31303 17685 31312
rect 18595 31352 18653 31353
rect 18595 31312 18604 31352
rect 18644 31312 18653 31352
rect 19131 31321 19132 31361
rect 19172 31321 19173 31361
rect 19131 31312 19173 31321
rect 18595 31311 18653 31312
rect 17163 31290 17205 31299
rect 12363 31268 12405 31277
rect 12363 31228 12364 31268
rect 12404 31228 12405 31268
rect 12363 31219 12405 31228
rect 14379 31268 14421 31277
rect 14379 31228 14380 31268
rect 14420 31228 14421 31268
rect 14379 31219 14421 31228
rect 19275 31268 19317 31277
rect 19275 31228 19276 31268
rect 19316 31228 19317 31268
rect 19275 31219 19317 31228
rect 2667 31184 2709 31193
rect 2667 31144 2668 31184
rect 2708 31144 2709 31184
rect 2667 31135 2709 31144
rect 2947 31184 3005 31185
rect 2947 31144 2956 31184
rect 2996 31144 3005 31184
rect 2947 31143 3005 31144
rect 4587 31184 4629 31193
rect 4587 31144 4588 31184
rect 4628 31144 4629 31184
rect 4587 31135 4629 31144
rect 16771 31184 16829 31185
rect 16771 31144 16780 31184
rect 16820 31144 16829 31184
rect 16771 31143 16829 31144
rect 19659 31184 19701 31193
rect 19659 31144 19660 31184
rect 19700 31144 19701 31184
rect 19659 31135 19701 31144
rect 20043 31184 20085 31193
rect 20043 31144 20044 31184
rect 20084 31144 20085 31184
rect 20043 31135 20085 31144
rect 1152 31016 20452 31040
rect 1152 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20452 31016
rect 1152 30952 20452 30976
rect 1419 30848 1461 30857
rect 1419 30808 1420 30848
rect 1460 30808 1461 30848
rect 1419 30799 1461 30808
rect 4875 30848 4917 30857
rect 4875 30808 4876 30848
rect 4916 30808 4917 30848
rect 4875 30799 4917 30808
rect 7947 30848 7989 30857
rect 7947 30808 7948 30848
rect 7988 30808 7989 30848
rect 7947 30799 7989 30808
rect 12363 30848 12405 30857
rect 12363 30808 12364 30848
rect 12404 30808 12405 30848
rect 12363 30799 12405 30808
rect 13995 30848 14037 30857
rect 13995 30808 13996 30848
rect 14036 30808 14037 30848
rect 13995 30799 14037 30808
rect 16107 30848 16149 30857
rect 16107 30808 16108 30848
rect 16148 30808 16149 30848
rect 16107 30799 16149 30808
rect 19659 30848 19701 30857
rect 19659 30808 19660 30848
rect 19700 30808 19701 30848
rect 19659 30799 19701 30808
rect 1603 30680 1661 30681
rect 1603 30640 1612 30680
rect 1652 30640 1661 30680
rect 1603 30639 1661 30640
rect 2851 30680 2909 30681
rect 2851 30640 2860 30680
rect 2900 30640 2909 30680
rect 2851 30639 2909 30640
rect 3427 30680 3485 30681
rect 3427 30640 3436 30680
rect 3476 30640 3485 30680
rect 3427 30639 3485 30640
rect 4675 30680 4733 30681
rect 4675 30640 4684 30680
rect 4724 30640 4733 30680
rect 4675 30639 4733 30640
rect 5347 30680 5405 30681
rect 5347 30640 5356 30680
rect 5396 30640 5405 30680
rect 5347 30639 5405 30640
rect 5643 30680 5685 30689
rect 5643 30640 5644 30680
rect 5684 30640 5685 30680
rect 5643 30631 5685 30640
rect 5739 30680 5781 30689
rect 5739 30640 5740 30680
rect 5780 30640 5781 30680
rect 5739 30631 5781 30640
rect 6211 30680 6269 30681
rect 6211 30640 6220 30680
rect 6260 30640 6269 30680
rect 6211 30639 6269 30640
rect 6499 30680 6557 30681
rect 6499 30640 6508 30680
rect 6548 30640 6557 30680
rect 6499 30639 6557 30640
rect 7747 30680 7805 30681
rect 7747 30640 7756 30680
rect 7796 30640 7805 30680
rect 7747 30639 7805 30640
rect 9091 30680 9149 30681
rect 9091 30640 9100 30680
rect 9140 30640 9149 30680
rect 9091 30639 9149 30640
rect 9387 30680 9429 30689
rect 9387 30640 9388 30680
rect 9428 30640 9429 30680
rect 9387 30631 9429 30640
rect 9763 30680 9821 30681
rect 9763 30640 9772 30680
rect 9812 30640 9821 30680
rect 9763 30639 9821 30640
rect 9955 30680 10013 30681
rect 9955 30640 9964 30680
rect 10004 30640 10013 30680
rect 9955 30639 10013 30640
rect 11203 30680 11261 30681
rect 11203 30640 11212 30680
rect 11252 30640 11261 30680
rect 11203 30639 11261 30640
rect 11587 30680 11645 30681
rect 11587 30640 11596 30680
rect 11636 30640 11645 30680
rect 11587 30639 11645 30640
rect 11979 30680 12021 30689
rect 11979 30640 11980 30680
rect 12020 30640 12021 30680
rect 11979 30631 12021 30640
rect 12547 30680 12605 30681
rect 12547 30640 12556 30680
rect 12596 30640 12605 30680
rect 12547 30639 12605 30640
rect 13795 30680 13853 30681
rect 13795 30640 13804 30680
rect 13844 30640 13853 30680
rect 13795 30639 13853 30640
rect 14379 30680 14421 30689
rect 14379 30640 14380 30680
rect 14420 30640 14421 30680
rect 14379 30631 14421 30640
rect 14475 30680 14517 30689
rect 14475 30640 14476 30680
rect 14516 30640 14517 30680
rect 14475 30631 14517 30640
rect 14859 30680 14901 30689
rect 14859 30640 14860 30680
rect 14900 30640 14901 30680
rect 14859 30631 14901 30640
rect 15427 30680 15485 30681
rect 15427 30640 15436 30680
rect 15476 30640 15485 30680
rect 15427 30639 15485 30640
rect 15915 30675 15957 30684
rect 15915 30635 15916 30675
rect 15956 30635 15957 30675
rect 16291 30680 16349 30681
rect 16291 30640 16300 30680
rect 16340 30640 16349 30680
rect 16291 30639 16349 30640
rect 17539 30680 17597 30681
rect 17539 30640 17548 30680
rect 17588 30640 17597 30680
rect 17539 30639 17597 30640
rect 18211 30680 18269 30681
rect 18211 30640 18220 30680
rect 18260 30640 18269 30680
rect 18211 30639 18269 30640
rect 19459 30680 19517 30681
rect 19459 30640 19468 30680
rect 19508 30640 19517 30680
rect 19459 30639 19517 30640
rect 15915 30626 15957 30635
rect 1219 30596 1277 30597
rect 1219 30556 1228 30596
rect 1268 30556 1277 30596
rect 1219 30555 1277 30556
rect 5059 30596 5117 30597
rect 5059 30556 5068 30596
rect 5108 30556 5117 30596
rect 5059 30555 5117 30556
rect 9483 30596 9525 30605
rect 9483 30556 9484 30596
rect 9524 30556 9525 30596
rect 9483 30547 9525 30556
rect 9675 30596 9717 30605
rect 9675 30556 9676 30596
rect 9716 30556 9717 30596
rect 9675 30547 9717 30556
rect 11691 30596 11733 30605
rect 11691 30556 11692 30596
rect 11732 30556 11733 30596
rect 11691 30547 11733 30556
rect 11883 30596 11925 30605
rect 11883 30556 11884 30596
rect 11924 30556 11925 30596
rect 11883 30547 11925 30556
rect 12163 30596 12221 30597
rect 12163 30556 12172 30596
rect 12212 30556 12221 30596
rect 12163 30555 12221 30556
rect 14955 30596 14997 30605
rect 14955 30556 14956 30596
rect 14996 30556 14997 30596
rect 14955 30547 14997 30556
rect 19843 30596 19901 30597
rect 19843 30556 19852 30596
rect 19892 30556 19901 30596
rect 19843 30555 19901 30556
rect 9579 30512 9621 30521
rect 9579 30472 9580 30512
rect 9620 30472 9621 30512
rect 9579 30463 9621 30472
rect 11787 30512 11829 30521
rect 11787 30472 11788 30512
rect 11828 30472 11829 30512
rect 11787 30463 11829 30472
rect 3051 30428 3093 30437
rect 3051 30388 3052 30428
rect 3092 30388 3093 30428
rect 3051 30379 3093 30388
rect 3243 30428 3285 30437
rect 3243 30388 3244 30428
rect 3284 30388 3285 30428
rect 3243 30379 3285 30388
rect 6019 30428 6077 30429
rect 6019 30388 6028 30428
rect 6068 30388 6077 30428
rect 6019 30387 6077 30388
rect 6315 30428 6357 30437
rect 6315 30388 6316 30428
rect 6356 30388 6357 30428
rect 6315 30379 6357 30388
rect 8619 30428 8661 30437
rect 8619 30388 8620 30428
rect 8660 30388 8661 30428
rect 8619 30379 8661 30388
rect 11403 30428 11445 30437
rect 11403 30388 11404 30428
rect 11444 30388 11445 30428
rect 11403 30379 11445 30388
rect 17739 30428 17781 30437
rect 17739 30388 17740 30428
rect 17780 30388 17781 30428
rect 17739 30379 17781 30388
rect 20043 30428 20085 30437
rect 20043 30388 20044 30428
rect 20084 30388 20085 30428
rect 20043 30379 20085 30388
rect 1152 30260 20352 30284
rect 1152 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 20352 30260
rect 1152 30196 20352 30220
rect 9867 30092 9909 30101
rect 9867 30052 9868 30092
rect 9908 30052 9909 30092
rect 9867 30043 9909 30052
rect 12939 30092 12981 30101
rect 12939 30052 12940 30092
rect 12980 30052 12981 30092
rect 12939 30043 12981 30052
rect 16203 30092 16245 30101
rect 16203 30052 16204 30092
rect 16244 30052 16245 30092
rect 16203 30043 16245 30052
rect 16395 30092 16437 30101
rect 16395 30052 16396 30092
rect 16436 30052 16437 30092
rect 16395 30043 16437 30052
rect 17067 30092 17109 30101
rect 17067 30052 17068 30092
rect 17108 30052 17109 30092
rect 17067 30043 17109 30052
rect 8139 30008 8181 30017
rect 8139 29968 8140 30008
rect 8180 29968 8181 30008
rect 8139 29959 8181 29968
rect 9187 30008 9245 30009
rect 9187 29968 9196 30008
rect 9236 29968 9245 30008
rect 9187 29967 9245 29968
rect 11779 30008 11837 30009
rect 11779 29968 11788 30008
rect 11828 29968 11837 30008
rect 11779 29967 11837 29968
rect 12739 29924 12797 29925
rect 12739 29884 12748 29924
rect 12788 29884 12797 29924
rect 12739 29883 12797 29884
rect 17835 29924 17877 29933
rect 17835 29884 17836 29924
rect 17876 29884 17877 29924
rect 17835 29875 17877 29884
rect 19363 29924 19421 29925
rect 19363 29884 19372 29924
rect 19412 29884 19421 29924
rect 19363 29883 19421 29884
rect 19747 29924 19805 29925
rect 19747 29884 19756 29924
rect 19796 29884 19805 29924
rect 19747 29883 19805 29884
rect 18939 29849 18981 29858
rect 1315 29840 1373 29841
rect 1315 29800 1324 29840
rect 1364 29800 1373 29840
rect 1315 29799 1373 29800
rect 1507 29840 1565 29841
rect 1507 29800 1516 29840
rect 1556 29800 1565 29840
rect 1507 29799 1565 29800
rect 2755 29840 2813 29841
rect 2755 29800 2764 29840
rect 2804 29800 2813 29840
rect 2755 29799 2813 29800
rect 3331 29840 3389 29841
rect 3331 29800 3340 29840
rect 3380 29800 3389 29840
rect 3331 29799 3389 29800
rect 4579 29840 4637 29841
rect 4579 29800 4588 29840
rect 4628 29800 4637 29840
rect 4579 29799 4637 29800
rect 5059 29840 5117 29841
rect 5059 29800 5068 29840
rect 5108 29800 5117 29840
rect 5059 29799 5117 29800
rect 6307 29840 6365 29841
rect 6307 29800 6316 29840
rect 6356 29800 6365 29840
rect 6307 29799 6365 29800
rect 6691 29840 6749 29841
rect 6691 29800 6700 29840
rect 6740 29800 6749 29840
rect 6691 29799 6749 29800
rect 7939 29840 7997 29841
rect 7939 29800 7948 29840
rect 7988 29800 7997 29840
rect 7939 29799 7997 29800
rect 8515 29840 8573 29841
rect 8515 29800 8524 29840
rect 8564 29800 8573 29840
rect 8515 29799 8573 29800
rect 8811 29840 8853 29849
rect 8811 29800 8812 29840
rect 8852 29800 8853 29840
rect 8811 29791 8853 29800
rect 9475 29840 9533 29841
rect 9475 29800 9484 29840
rect 9524 29800 9533 29840
rect 9475 29799 9533 29800
rect 9579 29840 9621 29849
rect 9579 29800 9580 29840
rect 9620 29800 9621 29840
rect 9579 29791 9621 29800
rect 10147 29840 10205 29841
rect 10147 29800 10156 29840
rect 10196 29800 10205 29840
rect 10147 29799 10205 29800
rect 11395 29840 11453 29841
rect 11395 29800 11404 29840
rect 11444 29800 11453 29840
rect 11395 29799 11453 29800
rect 12171 29840 12213 29849
rect 12171 29800 12172 29840
rect 12212 29800 12213 29840
rect 12171 29791 12213 29800
rect 12451 29840 12509 29841
rect 12451 29800 12460 29840
rect 12500 29800 12509 29840
rect 12451 29799 12509 29800
rect 13123 29840 13181 29841
rect 13123 29800 13132 29840
rect 13172 29800 13181 29840
rect 13123 29799 13181 29800
rect 14371 29840 14429 29841
rect 14371 29800 14380 29840
rect 14420 29800 14429 29840
rect 14371 29799 14429 29800
rect 14755 29840 14813 29841
rect 14755 29800 14764 29840
rect 14804 29800 14813 29840
rect 14755 29799 14813 29800
rect 16003 29840 16061 29841
rect 16003 29800 16012 29840
rect 16052 29800 16061 29840
rect 16003 29799 16061 29800
rect 16395 29840 16437 29849
rect 16395 29800 16396 29840
rect 16436 29800 16437 29840
rect 16395 29791 16437 29800
rect 16587 29840 16629 29849
rect 16587 29800 16588 29840
rect 16628 29800 16629 29840
rect 16587 29791 16629 29800
rect 16675 29840 16733 29841
rect 16675 29800 16684 29840
rect 16724 29800 16733 29840
rect 16675 29799 16733 29800
rect 16875 29840 16917 29849
rect 16875 29800 16876 29840
rect 16916 29800 16917 29840
rect 16875 29791 16917 29800
rect 17067 29840 17109 29849
rect 17067 29800 17068 29840
rect 17108 29800 17109 29840
rect 17067 29791 17109 29800
rect 17355 29840 17397 29849
rect 17355 29800 17356 29840
rect 17396 29800 17397 29840
rect 17355 29791 17397 29800
rect 17451 29840 17493 29849
rect 17451 29800 17452 29840
rect 17492 29800 17493 29840
rect 17451 29791 17493 29800
rect 17931 29840 17973 29849
rect 17931 29800 17932 29840
rect 17972 29800 17973 29840
rect 17931 29791 17973 29800
rect 18403 29840 18461 29841
rect 18403 29800 18412 29840
rect 18452 29800 18461 29840
rect 18939 29809 18940 29849
rect 18980 29809 18981 29849
rect 18939 29800 18981 29809
rect 18403 29799 18461 29800
rect 8907 29756 8949 29765
rect 8907 29716 8908 29756
rect 8948 29716 8949 29756
rect 8907 29707 8949 29716
rect 12075 29756 12117 29765
rect 12075 29716 12076 29756
rect 12116 29716 12117 29756
rect 12075 29707 12117 29716
rect 14571 29756 14613 29765
rect 14571 29716 14572 29756
rect 14612 29716 14613 29756
rect 14571 29707 14613 29716
rect 19083 29756 19125 29765
rect 19083 29716 19084 29756
rect 19124 29716 19125 29756
rect 19083 29707 19125 29716
rect 1227 29672 1269 29681
rect 1227 29632 1228 29672
rect 1268 29632 1269 29672
rect 1227 29623 1269 29632
rect 2955 29672 2997 29681
rect 2955 29632 2956 29672
rect 2996 29632 2997 29672
rect 2955 29623 2997 29632
rect 3147 29672 3189 29681
rect 3147 29632 3148 29672
rect 3188 29632 3189 29672
rect 3147 29623 3189 29632
rect 4875 29672 4917 29681
rect 4875 29632 4876 29672
rect 4916 29632 4917 29672
rect 4875 29623 4917 29632
rect 9387 29668 9429 29677
rect 9387 29628 9388 29668
rect 9428 29628 9429 29668
rect 9387 29619 9429 29628
rect 11595 29672 11637 29681
rect 11595 29632 11596 29672
rect 11636 29632 11637 29672
rect 11595 29623 11637 29632
rect 19563 29672 19605 29681
rect 19563 29632 19564 29672
rect 19604 29632 19605 29672
rect 19563 29623 19605 29632
rect 19947 29672 19989 29681
rect 19947 29632 19948 29672
rect 19988 29632 19989 29672
rect 19947 29623 19989 29632
rect 1152 29504 20452 29528
rect 1152 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20452 29504
rect 1152 29440 20452 29464
rect 15531 29336 15573 29345
rect 15531 29296 15532 29336
rect 15572 29296 15573 29336
rect 15531 29287 15573 29296
rect 18987 29336 19029 29345
rect 18987 29296 18988 29336
rect 19028 29296 19029 29336
rect 18987 29287 19029 29296
rect 12459 29252 12501 29261
rect 12459 29212 12460 29252
rect 12500 29212 12501 29252
rect 12459 29203 12501 29212
rect 1219 29168 1277 29169
rect 1219 29128 1228 29168
rect 1268 29128 1277 29168
rect 1219 29127 1277 29128
rect 2467 29168 2525 29169
rect 2467 29128 2476 29168
rect 2516 29128 2525 29168
rect 2467 29127 2525 29128
rect 3235 29168 3293 29169
rect 3235 29128 3244 29168
rect 3284 29128 3293 29168
rect 3235 29127 3293 29128
rect 4483 29168 4541 29169
rect 4483 29128 4492 29168
rect 4532 29128 4541 29168
rect 4483 29127 4541 29128
rect 4867 29168 4925 29169
rect 4867 29128 4876 29168
rect 4916 29128 4925 29168
rect 4867 29127 4925 29128
rect 6115 29168 6173 29169
rect 6115 29128 6124 29168
rect 6164 29128 6173 29168
rect 6115 29127 6173 29128
rect 6499 29168 6557 29169
rect 6499 29128 6508 29168
rect 6548 29128 6557 29168
rect 6499 29127 6557 29128
rect 7747 29168 7805 29169
rect 7747 29128 7756 29168
rect 7796 29128 7805 29168
rect 7747 29127 7805 29128
rect 8131 29168 8189 29169
rect 8131 29128 8140 29168
rect 8180 29128 8189 29168
rect 8131 29127 8189 29128
rect 8235 29168 8277 29177
rect 8235 29128 8236 29168
rect 8276 29128 8277 29168
rect 8235 29119 8277 29128
rect 8427 29168 8469 29177
rect 8427 29128 8428 29168
rect 8468 29128 8469 29168
rect 8427 29119 8469 29128
rect 8611 29168 8669 29169
rect 8611 29128 8620 29168
rect 8660 29128 8669 29168
rect 8611 29127 8669 29128
rect 9859 29168 9917 29169
rect 9859 29128 9868 29168
rect 9908 29128 9917 29168
rect 9859 29127 9917 29128
rect 10339 29168 10397 29169
rect 10339 29128 10348 29168
rect 10388 29128 10397 29168
rect 10339 29127 10397 29128
rect 11587 29168 11645 29169
rect 11587 29128 11596 29168
rect 11636 29128 11645 29168
rect 11587 29127 11645 29128
rect 12067 29168 12125 29169
rect 12067 29128 12076 29168
rect 12116 29128 12125 29168
rect 12067 29127 12125 29128
rect 12363 29168 12405 29177
rect 12363 29128 12364 29168
rect 12404 29128 12405 29168
rect 12363 29119 12405 29128
rect 12939 29168 12981 29177
rect 12939 29128 12940 29168
rect 12980 29128 12981 29168
rect 12939 29119 12981 29128
rect 13315 29168 13373 29169
rect 13315 29128 13324 29168
rect 13364 29128 13373 29168
rect 13315 29127 13373 29128
rect 13699 29168 13757 29169
rect 13699 29128 13708 29168
rect 13748 29128 13757 29168
rect 13699 29127 13757 29128
rect 14947 29168 15005 29169
rect 14947 29128 14956 29168
rect 14996 29128 15005 29168
rect 14947 29127 15005 29128
rect 15339 29168 15381 29177
rect 15339 29128 15340 29168
rect 15380 29128 15381 29168
rect 15339 29119 15381 29128
rect 15627 29168 15669 29177
rect 15627 29128 15628 29168
rect 15668 29128 15669 29168
rect 15627 29119 15669 29128
rect 15811 29168 15869 29169
rect 15811 29128 15820 29168
rect 15860 29128 15869 29168
rect 15811 29127 15869 29128
rect 17059 29168 17117 29169
rect 17059 29128 17068 29168
rect 17108 29128 17117 29168
rect 17059 29127 17117 29128
rect 17539 29168 17597 29169
rect 17539 29128 17548 29168
rect 17588 29128 17597 29168
rect 17539 29127 17597 29128
rect 18787 29168 18845 29169
rect 18787 29128 18796 29168
rect 18836 29128 18845 29168
rect 18787 29127 18845 29128
rect 2851 29084 2909 29085
rect 2851 29044 2860 29084
rect 2900 29044 2909 29084
rect 2851 29043 2909 29044
rect 13035 29084 13077 29093
rect 13035 29044 13036 29084
rect 13076 29044 13077 29084
rect 13035 29035 13077 29044
rect 13227 29084 13269 29093
rect 13227 29044 13228 29084
rect 13268 29044 13269 29084
rect 13227 29035 13269 29044
rect 19363 29084 19421 29085
rect 19363 29044 19372 29084
rect 19412 29044 19421 29084
rect 19363 29043 19421 29044
rect 19747 29084 19805 29085
rect 19747 29044 19756 29084
rect 19796 29044 19805 29084
rect 19747 29043 19805 29044
rect 3051 29000 3093 29009
rect 3051 28960 3052 29000
rect 3092 28960 3093 29000
rect 3051 28951 3093 28960
rect 11787 29000 11829 29009
rect 11787 28960 11788 29000
rect 11828 28960 11829 29000
rect 11787 28951 11829 28960
rect 13131 29000 13173 29009
rect 13131 28960 13132 29000
rect 13172 28960 13173 29000
rect 13131 28951 13173 28960
rect 19947 29000 19989 29009
rect 19947 28960 19948 29000
rect 19988 28960 19989 29000
rect 19947 28951 19989 28960
rect 2667 28916 2709 28925
rect 2667 28876 2668 28916
rect 2708 28876 2709 28916
rect 2667 28867 2709 28876
rect 4683 28916 4725 28925
rect 4683 28876 4684 28916
rect 4724 28876 4725 28916
rect 4683 28867 4725 28876
rect 6315 28916 6357 28925
rect 6315 28876 6316 28916
rect 6356 28876 6357 28916
rect 6315 28867 6357 28876
rect 7947 28916 7989 28925
rect 7947 28876 7948 28916
rect 7988 28876 7989 28916
rect 7947 28867 7989 28876
rect 8427 28916 8469 28925
rect 8427 28876 8428 28916
rect 8468 28876 8469 28916
rect 8427 28867 8469 28876
rect 10059 28916 10101 28925
rect 10059 28876 10060 28916
rect 10100 28876 10101 28916
rect 10059 28867 10101 28876
rect 12739 28916 12797 28917
rect 12739 28876 12748 28916
rect 12788 28876 12797 28916
rect 12739 28875 12797 28876
rect 15147 28916 15189 28925
rect 15147 28876 15148 28916
rect 15188 28876 15189 28916
rect 15147 28867 15189 28876
rect 17259 28916 17301 28925
rect 17259 28876 17260 28916
rect 17300 28876 17301 28916
rect 17259 28867 17301 28876
rect 19563 28916 19605 28925
rect 19563 28876 19564 28916
rect 19604 28876 19605 28916
rect 19563 28867 19605 28876
rect 1152 28748 20352 28772
rect 1152 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 20352 28748
rect 1152 28684 20352 28708
rect 4203 28580 4245 28589
rect 4203 28540 4204 28580
rect 4244 28540 4245 28580
rect 4203 28531 4245 28540
rect 7083 28580 7125 28589
rect 7083 28540 7084 28580
rect 7124 28540 7125 28580
rect 7083 28531 7125 28540
rect 11307 28580 11349 28589
rect 11307 28540 11308 28580
rect 11348 28540 11349 28580
rect 11307 28531 11349 28540
rect 12939 28580 12981 28589
rect 12939 28540 12940 28580
rect 12980 28540 12981 28580
rect 12939 28531 12981 28540
rect 3819 28496 3861 28505
rect 3819 28456 3820 28496
rect 3860 28456 3861 28496
rect 3819 28447 3861 28456
rect 12739 28496 12797 28497
rect 12739 28456 12748 28496
rect 12788 28456 12797 28496
rect 12739 28455 12797 28456
rect 3619 28412 3677 28413
rect 3619 28372 3628 28412
rect 3668 28372 3677 28412
rect 3619 28371 3677 28372
rect 4003 28412 4061 28413
rect 4003 28372 4012 28412
rect 4052 28372 4061 28412
rect 4003 28371 4061 28372
rect 4587 28412 4629 28421
rect 4587 28372 4588 28412
rect 4628 28372 4629 28412
rect 4587 28363 4629 28372
rect 6883 28412 6941 28413
rect 6883 28372 6892 28412
rect 6932 28372 6941 28412
rect 6883 28371 6941 28372
rect 19363 28412 19421 28413
rect 19363 28372 19372 28412
rect 19412 28372 19421 28412
rect 19363 28371 19421 28372
rect 19747 28412 19805 28413
rect 19747 28372 19756 28412
rect 19796 28372 19805 28412
rect 19747 28371 19805 28372
rect 1219 28328 1277 28329
rect 1219 28288 1228 28328
rect 1268 28288 1277 28328
rect 1219 28287 1277 28288
rect 2467 28328 2525 28329
rect 2467 28288 2476 28328
rect 2516 28288 2525 28328
rect 2947 28328 3005 28329
rect 2467 28287 2525 28288
rect 2848 28324 2906 28325
rect 2848 28284 2857 28324
rect 2897 28284 2906 28324
rect 2947 28288 2956 28328
rect 2996 28288 3005 28328
rect 2947 28287 3005 28288
rect 3147 28328 3189 28337
rect 3147 28288 3148 28328
rect 3188 28288 3189 28328
rect 2848 28283 2906 28284
rect 3147 28279 3189 28288
rect 3243 28328 3285 28337
rect 3243 28288 3244 28328
rect 3284 28288 3285 28328
rect 3243 28279 3285 28288
rect 3336 28328 3394 28329
rect 3336 28288 3345 28328
rect 3385 28288 3394 28328
rect 3336 28287 3394 28288
rect 5251 28328 5309 28329
rect 5251 28288 5260 28328
rect 5300 28288 5309 28328
rect 5251 28287 5309 28288
rect 6499 28328 6557 28329
rect 6499 28288 6508 28328
rect 6548 28288 6557 28328
rect 6499 28287 6557 28288
rect 7267 28328 7325 28329
rect 7267 28288 7276 28328
rect 7316 28288 7325 28328
rect 7267 28287 7325 28288
rect 8515 28328 8573 28329
rect 8515 28288 8524 28328
rect 8564 28288 8573 28328
rect 8515 28287 8573 28288
rect 8995 28328 9053 28329
rect 8995 28288 9004 28328
rect 9044 28288 9053 28328
rect 8995 28287 9053 28288
rect 9187 28328 9245 28329
rect 9187 28288 9196 28328
rect 9236 28288 9245 28328
rect 9187 28287 9245 28288
rect 10435 28328 10493 28329
rect 10435 28288 10444 28328
rect 10484 28288 10493 28328
rect 10435 28287 10493 28288
rect 11011 28328 11069 28329
rect 11011 28288 11020 28328
rect 11060 28288 11069 28328
rect 11011 28287 11069 28288
rect 11115 28328 11157 28337
rect 11115 28288 11116 28328
rect 11156 28288 11157 28328
rect 11115 28279 11157 28288
rect 11307 28328 11349 28337
rect 11307 28288 11308 28328
rect 11348 28288 11349 28328
rect 11307 28279 11349 28288
rect 11499 28328 11541 28337
rect 11499 28288 11500 28328
rect 11540 28288 11541 28328
rect 11499 28279 11541 28288
rect 11595 28328 11637 28337
rect 11595 28288 11596 28328
rect 11636 28288 11637 28328
rect 11595 28279 11637 28288
rect 11691 28328 11733 28337
rect 11691 28288 11692 28328
rect 11732 28288 11733 28328
rect 11691 28279 11733 28288
rect 12067 28328 12125 28329
rect 12067 28288 12076 28328
rect 12116 28288 12125 28328
rect 12067 28287 12125 28288
rect 12363 28328 12405 28337
rect 12363 28288 12364 28328
rect 12404 28288 12405 28328
rect 12363 28279 12405 28288
rect 12939 28328 12981 28337
rect 12939 28288 12940 28328
rect 12980 28288 12981 28328
rect 12939 28279 12981 28288
rect 13131 28328 13173 28337
rect 13131 28288 13132 28328
rect 13172 28288 13173 28328
rect 13131 28279 13173 28288
rect 13219 28328 13277 28329
rect 13219 28288 13228 28328
rect 13268 28288 13277 28328
rect 13219 28287 13277 28288
rect 13507 28328 13565 28329
rect 13507 28288 13516 28328
rect 13556 28288 13565 28328
rect 13507 28287 13565 28288
rect 14755 28328 14813 28329
rect 14755 28288 14764 28328
rect 14804 28288 14813 28328
rect 14755 28287 14813 28288
rect 15243 28328 15285 28337
rect 15243 28288 15244 28328
rect 15284 28288 15285 28328
rect 15243 28279 15285 28288
rect 15339 28328 15381 28337
rect 15339 28288 15340 28328
rect 15380 28288 15381 28328
rect 15339 28279 15381 28288
rect 15723 28328 15765 28337
rect 15723 28288 15724 28328
rect 15764 28288 15765 28328
rect 15723 28279 15765 28288
rect 15819 28328 15861 28337
rect 16779 28333 16821 28342
rect 15819 28288 15820 28328
rect 15860 28288 15861 28328
rect 15819 28279 15861 28288
rect 16291 28328 16349 28329
rect 16291 28288 16300 28328
rect 16340 28288 16349 28328
rect 16291 28287 16349 28288
rect 16779 28293 16780 28333
rect 16820 28293 16821 28333
rect 16779 28284 16821 28293
rect 17259 28328 17301 28337
rect 17259 28288 17260 28328
rect 17300 28288 17301 28328
rect 17259 28279 17301 28288
rect 17355 28328 17397 28337
rect 17355 28288 17356 28328
rect 17396 28288 17397 28328
rect 17355 28279 17397 28288
rect 17739 28328 17781 28337
rect 17739 28288 17740 28328
rect 17780 28288 17781 28328
rect 17739 28279 17781 28288
rect 17835 28328 17877 28337
rect 18795 28333 18837 28342
rect 17835 28288 17836 28328
rect 17876 28288 17877 28328
rect 17835 28279 17877 28288
rect 18307 28328 18365 28329
rect 18307 28288 18316 28328
rect 18356 28288 18365 28328
rect 18307 28287 18365 28288
rect 18795 28293 18796 28333
rect 18836 28293 18837 28333
rect 18795 28284 18837 28293
rect 12459 28244 12501 28253
rect 12459 28204 12460 28244
rect 12500 28204 12501 28244
rect 12459 28195 12501 28204
rect 16971 28244 17013 28253
rect 16971 28204 16972 28244
rect 17012 28204 17013 28244
rect 16971 28195 17013 28204
rect 18987 28244 19029 28253
rect 18987 28204 18988 28244
rect 19028 28204 19029 28244
rect 18987 28195 19029 28204
rect 2667 28160 2709 28169
rect 2667 28120 2668 28160
rect 2708 28120 2709 28160
rect 2667 28111 2709 28120
rect 3235 28160 3293 28161
rect 3235 28120 3244 28160
rect 3284 28120 3293 28160
rect 3235 28119 3293 28120
rect 4867 28160 4925 28161
rect 4867 28120 4876 28160
rect 4916 28120 4925 28160
rect 4867 28119 4925 28120
rect 6699 28160 6741 28169
rect 6699 28120 6700 28160
rect 6740 28120 6741 28160
rect 6699 28111 6741 28120
rect 8715 28160 8757 28169
rect 8715 28120 8716 28160
rect 8756 28120 8757 28160
rect 8715 28111 8757 28120
rect 8907 28160 8949 28169
rect 8907 28120 8908 28160
rect 8948 28120 8949 28160
rect 8907 28111 8949 28120
rect 10635 28160 10677 28169
rect 10635 28120 10636 28160
rect 10676 28120 10677 28160
rect 10635 28111 10677 28120
rect 11779 28160 11837 28161
rect 11779 28120 11788 28160
rect 11828 28120 11837 28160
rect 11779 28119 11837 28120
rect 14955 28160 14997 28169
rect 14955 28120 14956 28160
rect 14996 28120 14997 28160
rect 14955 28111 14997 28120
rect 19563 28160 19605 28169
rect 19563 28120 19564 28160
rect 19604 28120 19605 28160
rect 19563 28111 19605 28120
rect 19947 28160 19989 28169
rect 19947 28120 19948 28160
rect 19988 28120 19989 28160
rect 19947 28111 19989 28120
rect 1152 27992 20452 28016
rect 1152 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20452 27992
rect 1152 27928 20452 27952
rect 11875 27824 11933 27825
rect 11875 27784 11884 27824
rect 11924 27784 11933 27824
rect 11875 27783 11933 27784
rect 12739 27824 12797 27825
rect 12739 27784 12748 27824
rect 12788 27784 12797 27824
rect 12739 27783 12797 27784
rect 16779 27824 16821 27833
rect 16779 27784 16780 27824
rect 16820 27784 16821 27824
rect 16779 27775 16821 27784
rect 5547 27740 5589 27749
rect 5547 27700 5548 27740
rect 5588 27700 5589 27740
rect 5547 27691 5589 27700
rect 6795 27740 6837 27749
rect 6795 27700 6796 27740
rect 6836 27700 6837 27740
rect 6795 27691 6837 27700
rect 8811 27740 8853 27749
rect 8811 27700 8812 27740
rect 8852 27700 8853 27740
rect 8811 27691 8853 27700
rect 9099 27740 9141 27749
rect 9099 27700 9100 27740
rect 9140 27700 9141 27740
rect 9099 27691 9141 27700
rect 9771 27740 9813 27749
rect 9771 27700 9772 27740
rect 9812 27700 9813 27740
rect 9771 27691 9813 27700
rect 15147 27740 15189 27749
rect 15147 27700 15148 27740
rect 15188 27700 15189 27740
rect 15147 27691 15189 27700
rect 19275 27740 19317 27749
rect 19275 27700 19276 27740
rect 19316 27700 19317 27740
rect 19275 27691 19317 27700
rect 1315 27656 1373 27657
rect 1315 27616 1324 27656
rect 1364 27616 1373 27656
rect 1315 27615 1373 27616
rect 1419 27656 1461 27665
rect 1419 27616 1420 27656
rect 1460 27616 1461 27656
rect 1419 27607 1461 27616
rect 1611 27656 1653 27665
rect 1611 27616 1612 27656
rect 1652 27616 1653 27656
rect 1611 27607 1653 27616
rect 1795 27656 1853 27657
rect 1795 27616 1804 27656
rect 1844 27616 1853 27656
rect 1795 27615 1853 27616
rect 3043 27656 3101 27657
rect 3043 27616 3052 27656
rect 3092 27616 3101 27656
rect 3043 27615 3101 27616
rect 3819 27656 3861 27665
rect 3819 27616 3820 27656
rect 3860 27616 3861 27656
rect 3819 27607 3861 27616
rect 3915 27656 3957 27665
rect 3915 27616 3916 27656
rect 3956 27616 3957 27656
rect 3915 27607 3957 27616
rect 4867 27656 4925 27657
rect 4867 27616 4876 27656
rect 4916 27616 4925 27656
rect 4867 27615 4925 27616
rect 5355 27651 5397 27660
rect 5355 27611 5356 27651
rect 5396 27611 5397 27651
rect 5355 27602 5397 27611
rect 6027 27656 6069 27665
rect 6027 27616 6028 27656
rect 6068 27616 6069 27656
rect 6027 27607 6069 27616
rect 6123 27656 6165 27665
rect 6123 27616 6124 27656
rect 6164 27616 6165 27656
rect 6123 27607 6165 27616
rect 6403 27656 6461 27657
rect 6403 27616 6412 27656
rect 6452 27616 6461 27656
rect 6403 27615 6461 27616
rect 6691 27656 6749 27657
rect 6691 27616 6700 27656
rect 6740 27616 6749 27656
rect 6691 27615 6749 27616
rect 7083 27656 7125 27665
rect 7083 27616 7084 27656
rect 7124 27616 7125 27656
rect 7083 27607 7125 27616
rect 7179 27656 7221 27665
rect 7179 27616 7180 27656
rect 7220 27616 7221 27656
rect 7179 27607 7221 27616
rect 8131 27656 8189 27657
rect 8131 27616 8140 27656
rect 8180 27616 8189 27656
rect 9003 27656 9045 27665
rect 8131 27615 8189 27616
rect 8667 27646 8709 27655
rect 8667 27606 8668 27646
rect 8708 27606 8709 27646
rect 9003 27616 9004 27656
rect 9044 27616 9045 27656
rect 9003 27607 9045 27616
rect 9195 27656 9237 27665
rect 9195 27616 9196 27656
rect 9236 27616 9237 27656
rect 9195 27607 9237 27616
rect 9283 27656 9341 27657
rect 9283 27616 9292 27656
rect 9332 27616 9341 27656
rect 9283 27615 9341 27616
rect 9483 27656 9525 27665
rect 9483 27616 9484 27656
rect 9524 27616 9525 27656
rect 9483 27607 9525 27616
rect 9579 27656 9621 27665
rect 9579 27616 9580 27656
rect 9620 27616 9621 27656
rect 9579 27607 9621 27616
rect 9675 27656 9717 27665
rect 9675 27616 9676 27656
rect 9716 27616 9717 27656
rect 9675 27607 9717 27616
rect 10147 27656 10205 27657
rect 10147 27616 10156 27656
rect 10196 27616 10205 27656
rect 10147 27615 10205 27616
rect 11395 27656 11453 27657
rect 11395 27616 11404 27656
rect 11444 27616 11453 27656
rect 11395 27615 11453 27616
rect 11787 27656 11829 27665
rect 11787 27616 11788 27656
rect 11828 27616 11829 27656
rect 11787 27607 11829 27616
rect 11979 27656 12021 27665
rect 11979 27616 11980 27656
rect 12020 27616 12021 27656
rect 11979 27607 12021 27616
rect 12067 27656 12125 27657
rect 12067 27616 12076 27656
rect 12116 27616 12125 27656
rect 12067 27615 12125 27616
rect 12459 27656 12501 27665
rect 12459 27616 12460 27656
rect 12500 27616 12501 27656
rect 12459 27607 12501 27616
rect 12555 27656 12597 27665
rect 12555 27616 12556 27656
rect 12596 27616 12597 27656
rect 13515 27656 13557 27665
rect 12555 27607 12597 27616
rect 13419 27637 13461 27646
rect 8667 27597 8709 27606
rect 13419 27597 13420 27637
rect 13460 27597 13461 27637
rect 13515 27616 13516 27656
rect 13556 27616 13557 27656
rect 13515 27607 13557 27616
rect 14467 27656 14525 27657
rect 14467 27616 14476 27656
rect 14516 27616 14525 27656
rect 14467 27615 14525 27616
rect 14955 27651 14997 27660
rect 14955 27611 14956 27651
rect 14996 27611 14997 27651
rect 15331 27656 15389 27657
rect 15331 27616 15340 27656
rect 15380 27616 15389 27656
rect 15331 27615 15389 27616
rect 16579 27656 16637 27657
rect 16579 27616 16588 27656
rect 16628 27616 16637 27656
rect 16579 27615 16637 27616
rect 17827 27656 17885 27657
rect 17827 27616 17836 27656
rect 17876 27616 17885 27656
rect 17827 27615 17885 27616
rect 19075 27656 19133 27657
rect 19075 27616 19084 27656
rect 19124 27616 19133 27656
rect 19075 27615 19133 27616
rect 14955 27602 14997 27611
rect 13419 27588 13461 27597
rect 4299 27572 4341 27581
rect 4299 27532 4300 27572
rect 4340 27532 4341 27572
rect 4299 27523 4341 27532
rect 4395 27572 4437 27581
rect 4395 27532 4396 27572
rect 4436 27532 4437 27572
rect 4395 27523 4437 27532
rect 7563 27572 7605 27581
rect 7563 27532 7564 27572
rect 7604 27532 7605 27572
rect 7563 27523 7605 27532
rect 7659 27572 7701 27581
rect 7659 27532 7660 27572
rect 7700 27532 7701 27572
rect 7659 27523 7701 27532
rect 12931 27572 12989 27573
rect 12931 27532 12940 27572
rect 12980 27532 12989 27572
rect 12931 27531 12989 27532
rect 13899 27572 13941 27581
rect 13899 27532 13900 27572
rect 13940 27532 13941 27572
rect 13899 27523 13941 27532
rect 13995 27572 14037 27581
rect 13995 27532 13996 27572
rect 14036 27532 14037 27572
rect 13995 27523 14037 27532
rect 17059 27572 17117 27573
rect 17059 27532 17068 27572
rect 17108 27532 17117 27572
rect 17059 27531 17117 27532
rect 17443 27572 17501 27573
rect 17443 27532 17452 27572
rect 17492 27532 17501 27572
rect 17443 27531 17501 27532
rect 19459 27572 19517 27573
rect 19459 27532 19468 27572
rect 19508 27532 19517 27572
rect 19459 27531 19517 27532
rect 19843 27572 19901 27573
rect 19843 27532 19852 27572
rect 19892 27532 19901 27572
rect 19843 27531 19901 27532
rect 3435 27488 3477 27497
rect 3435 27448 3436 27488
rect 3476 27448 3477 27488
rect 3435 27439 3477 27448
rect 5731 27488 5789 27489
rect 5731 27448 5740 27488
rect 5780 27448 5789 27488
rect 5731 27447 5789 27448
rect 13131 27488 13173 27497
rect 13131 27448 13132 27488
rect 13172 27448 13173 27488
rect 13131 27439 13173 27448
rect 17259 27488 17301 27497
rect 17259 27448 17260 27488
rect 17300 27448 17301 27488
rect 17259 27439 17301 27448
rect 17643 27488 17685 27497
rect 17643 27448 17644 27488
rect 17684 27448 17685 27488
rect 17643 27439 17685 27448
rect 1611 27404 1653 27413
rect 1611 27364 1612 27404
rect 1652 27364 1653 27404
rect 1611 27355 1653 27364
rect 3243 27404 3285 27413
rect 3243 27364 3244 27404
rect 3284 27364 3285 27404
rect 3243 27355 3285 27364
rect 11595 27404 11637 27413
rect 11595 27364 11596 27404
rect 11636 27364 11637 27404
rect 11595 27355 11637 27364
rect 19659 27404 19701 27413
rect 19659 27364 19660 27404
rect 19700 27364 19701 27404
rect 19659 27355 19701 27364
rect 20043 27404 20085 27413
rect 20043 27364 20044 27404
rect 20084 27364 20085 27404
rect 20043 27355 20085 27364
rect 1152 27236 20352 27260
rect 1152 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 20352 27236
rect 1152 27172 20352 27196
rect 8715 27068 8757 27077
rect 8715 27028 8716 27068
rect 8756 27028 8757 27068
rect 8715 27019 8757 27028
rect 9195 27068 9237 27077
rect 9195 27028 9196 27068
rect 9236 27028 9237 27068
rect 9195 27019 9237 27028
rect 13419 27068 13461 27077
rect 13419 27028 13420 27068
rect 13460 27028 13461 27068
rect 13419 27019 13461 27028
rect 15531 27068 15573 27077
rect 15531 27028 15532 27068
rect 15572 27028 15573 27068
rect 15531 27019 15573 27028
rect 6411 26984 6453 26993
rect 6411 26944 6412 26984
rect 6452 26944 6453 26984
rect 6411 26935 6453 26944
rect 9771 26984 9813 26993
rect 9771 26944 9772 26984
rect 9812 26944 9813 26984
rect 9771 26935 9813 26944
rect 17163 26984 17205 26993
rect 17163 26944 17164 26984
rect 17204 26944 17205 26984
rect 17163 26935 17205 26944
rect 10539 26900 10581 26909
rect 10539 26860 10540 26900
rect 10580 26860 10581 26900
rect 10539 26851 10581 26860
rect 10635 26900 10677 26909
rect 10635 26860 10636 26900
rect 10676 26860 10677 26900
rect 10635 26851 10677 26860
rect 15331 26900 15389 26901
rect 15331 26860 15340 26900
rect 15380 26860 15389 26900
rect 15331 26859 15389 26860
rect 19363 26900 19421 26901
rect 19363 26860 19372 26900
rect 19412 26860 19421 26900
rect 19363 26859 19421 26860
rect 19747 26900 19805 26901
rect 19747 26860 19756 26900
rect 19796 26860 19805 26900
rect 19747 26859 19805 26860
rect 3387 26825 3429 26834
rect 8235 26830 8277 26839
rect 1227 26816 1269 26825
rect 1227 26776 1228 26816
rect 1268 26776 1269 26816
rect 1227 26767 1269 26776
rect 1323 26816 1365 26825
rect 1323 26776 1324 26816
rect 1364 26776 1365 26816
rect 1323 26767 1365 26776
rect 1803 26816 1845 26825
rect 1803 26776 1804 26816
rect 1844 26776 1845 26816
rect 1803 26767 1845 26776
rect 1899 26816 1941 26825
rect 1899 26776 1900 26816
rect 1940 26776 1941 26816
rect 1899 26767 1941 26776
rect 2283 26816 2325 26825
rect 2283 26776 2284 26816
rect 2324 26776 2325 26816
rect 2283 26767 2325 26776
rect 2379 26816 2421 26825
rect 2379 26776 2380 26816
rect 2420 26776 2421 26816
rect 2379 26767 2421 26776
rect 2851 26816 2909 26817
rect 2851 26776 2860 26816
rect 2900 26776 2909 26816
rect 3387 26785 3388 26825
rect 3428 26785 3429 26825
rect 3387 26776 3429 26785
rect 4011 26816 4053 26825
rect 4011 26776 4012 26816
rect 4052 26776 4053 26816
rect 2851 26775 2909 26776
rect 4011 26767 4053 26776
rect 4107 26816 4149 26825
rect 4107 26776 4108 26816
rect 4148 26776 4149 26816
rect 4107 26767 4149 26776
rect 4203 26816 4245 26825
rect 4203 26776 4204 26816
rect 4244 26776 4245 26816
rect 4203 26767 4245 26776
rect 4299 26816 4341 26825
rect 4299 26776 4300 26816
rect 4340 26776 4341 26816
rect 4299 26767 4341 26776
rect 4675 26816 4733 26817
rect 4675 26776 4684 26816
rect 4724 26776 4733 26816
rect 4675 26775 4733 26776
rect 5923 26816 5981 26817
rect 5923 26776 5932 26816
rect 5972 26776 5981 26816
rect 5923 26775 5981 26776
rect 6699 26816 6741 26825
rect 6699 26776 6700 26816
rect 6740 26776 6741 26816
rect 6699 26767 6741 26776
rect 6795 26816 6837 26825
rect 6795 26776 6796 26816
rect 6836 26776 6837 26816
rect 6795 26767 6837 26776
rect 7179 26816 7221 26825
rect 7179 26776 7180 26816
rect 7220 26776 7221 26816
rect 7179 26767 7221 26776
rect 7275 26816 7317 26825
rect 7275 26776 7276 26816
rect 7316 26776 7317 26816
rect 7275 26767 7317 26776
rect 7747 26816 7805 26817
rect 7747 26776 7756 26816
rect 7796 26776 7805 26816
rect 8235 26790 8236 26830
rect 8276 26790 8277 26830
rect 11595 26830 11637 26839
rect 8235 26781 8277 26790
rect 8715 26816 8757 26825
rect 7747 26775 7805 26776
rect 8715 26776 8716 26816
rect 8756 26776 8757 26816
rect 8715 26767 8757 26776
rect 9003 26816 9045 26825
rect 9003 26776 9004 26816
rect 9044 26776 9045 26816
rect 9003 26767 9045 26776
rect 9195 26816 9237 26825
rect 9195 26776 9196 26816
rect 9236 26776 9237 26816
rect 9195 26767 9237 26776
rect 9387 26816 9429 26825
rect 9387 26776 9388 26816
rect 9428 26776 9429 26816
rect 9387 26767 9429 26776
rect 9475 26816 9533 26817
rect 9475 26776 9484 26816
rect 9524 26776 9533 26816
rect 9475 26775 9533 26776
rect 9667 26816 9725 26817
rect 9667 26776 9676 26816
rect 9716 26776 9725 26816
rect 9667 26775 9725 26776
rect 10059 26816 10101 26825
rect 10059 26776 10060 26816
rect 10100 26776 10101 26816
rect 10059 26767 10101 26776
rect 10155 26816 10197 26825
rect 10155 26776 10156 26816
rect 10196 26776 10197 26816
rect 10155 26767 10197 26776
rect 11107 26816 11165 26817
rect 11107 26776 11116 26816
rect 11156 26776 11165 26816
rect 11595 26790 11596 26830
rect 11636 26790 11637 26830
rect 19035 26825 19077 26834
rect 11595 26781 11637 26790
rect 11971 26816 12029 26817
rect 11107 26775 11165 26776
rect 11971 26776 11980 26816
rect 12020 26776 12029 26816
rect 11971 26775 12029 26776
rect 13219 26816 13277 26817
rect 13219 26776 13228 26816
rect 13268 26776 13277 26816
rect 13219 26775 13277 26776
rect 13603 26816 13661 26817
rect 13603 26776 13612 26816
rect 13652 26776 13661 26816
rect 13603 26775 13661 26776
rect 14851 26816 14909 26817
rect 14851 26776 14860 26816
rect 14900 26776 14909 26816
rect 14851 26775 14909 26776
rect 15715 26816 15773 26817
rect 15715 26776 15724 26816
rect 15764 26776 15773 26816
rect 15715 26775 15773 26776
rect 16963 26816 17021 26817
rect 16963 26776 16972 26816
rect 17012 26776 17021 26816
rect 16963 26775 17021 26776
rect 17451 26816 17493 26825
rect 17451 26776 17452 26816
rect 17492 26776 17493 26816
rect 17451 26767 17493 26776
rect 17547 26816 17589 26825
rect 17547 26776 17548 26816
rect 17588 26776 17589 26816
rect 17547 26767 17589 26776
rect 17931 26816 17973 26825
rect 17931 26776 17932 26816
rect 17972 26776 17973 26816
rect 17931 26767 17973 26776
rect 18027 26816 18069 26825
rect 18027 26776 18028 26816
rect 18068 26776 18069 26816
rect 18027 26767 18069 26776
rect 18499 26816 18557 26817
rect 18499 26776 18508 26816
rect 18548 26776 18557 26816
rect 19035 26785 19036 26825
rect 19076 26785 19077 26825
rect 19035 26776 19077 26785
rect 18499 26775 18557 26776
rect 3531 26732 3573 26741
rect 3531 26692 3532 26732
rect 3572 26692 3573 26732
rect 3531 26683 3573 26692
rect 11787 26732 11829 26741
rect 11787 26692 11788 26732
rect 11828 26692 11829 26732
rect 11787 26683 11829 26692
rect 1507 26648 1565 26649
rect 1507 26608 1516 26648
rect 1556 26608 1565 26648
rect 1507 26607 1565 26608
rect 3819 26648 3861 26657
rect 3819 26608 3820 26648
rect 3860 26608 3861 26648
rect 3819 26599 3861 26608
rect 6123 26648 6165 26657
rect 6123 26608 6124 26648
rect 6164 26608 6165 26648
rect 6123 26599 6165 26608
rect 8427 26648 8469 26657
rect 8427 26608 8428 26648
rect 8468 26608 8469 26648
rect 8427 26599 8469 26608
rect 15051 26648 15093 26657
rect 15051 26608 15052 26648
rect 15092 26608 15093 26648
rect 15051 26599 15093 26608
rect 19179 26648 19221 26657
rect 19179 26608 19180 26648
rect 19220 26608 19221 26648
rect 19179 26599 19221 26608
rect 19563 26648 19605 26657
rect 19563 26608 19564 26648
rect 19604 26608 19605 26648
rect 19563 26599 19605 26608
rect 19947 26648 19989 26657
rect 19947 26608 19948 26648
rect 19988 26608 19989 26648
rect 19947 26599 19989 26608
rect 1152 26480 20452 26504
rect 1152 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20452 26480
rect 1152 26416 20452 26440
rect 1419 26312 1461 26321
rect 1419 26272 1420 26312
rect 1460 26272 1461 26312
rect 1419 26263 1461 26272
rect 4491 26312 4533 26321
rect 4491 26272 4492 26312
rect 4532 26272 4533 26312
rect 4491 26263 4533 26272
rect 10923 26312 10965 26321
rect 10923 26272 10924 26312
rect 10964 26272 10965 26312
rect 10923 26263 10965 26272
rect 14571 26312 14613 26321
rect 14571 26272 14572 26312
rect 14612 26272 14613 26312
rect 14571 26263 14613 26272
rect 19563 26312 19605 26321
rect 19563 26272 19564 26312
rect 19604 26272 19605 26312
rect 19563 26263 19605 26272
rect 3531 26228 3573 26237
rect 3531 26188 3532 26228
rect 3572 26188 3573 26228
rect 3531 26179 3573 26188
rect 5355 26228 5397 26237
rect 5355 26188 5356 26228
rect 5396 26188 5397 26228
rect 5355 26179 5397 26188
rect 7275 26228 7317 26237
rect 7275 26188 7276 26228
rect 7316 26188 7317 26228
rect 7275 26179 7317 26188
rect 12555 26228 12597 26237
rect 12555 26188 12556 26228
rect 12596 26188 12597 26228
rect 12555 26179 12597 26188
rect 1227 26144 1269 26153
rect 1227 26104 1228 26144
rect 1268 26104 1269 26144
rect 1227 26095 1269 26104
rect 1323 26144 1365 26153
rect 1323 26104 1324 26144
rect 1364 26104 1365 26144
rect 1323 26095 1365 26104
rect 1515 26144 1557 26153
rect 1515 26104 1516 26144
rect 1556 26104 1557 26144
rect 1515 26095 1557 26104
rect 1803 26144 1845 26153
rect 1803 26104 1804 26144
rect 1844 26104 1845 26144
rect 1803 26095 1845 26104
rect 1899 26144 1941 26153
rect 1899 26104 1900 26144
rect 1940 26104 1941 26144
rect 1899 26095 1941 26104
rect 2283 26144 2325 26153
rect 2283 26104 2284 26144
rect 2324 26104 2325 26144
rect 2283 26095 2325 26104
rect 2851 26144 2909 26145
rect 2851 26104 2860 26144
rect 2900 26104 2909 26144
rect 2851 26103 2909 26104
rect 3339 26139 3381 26148
rect 3339 26099 3340 26139
rect 3380 26099 3381 26139
rect 4963 26144 5021 26145
rect 4963 26104 4972 26144
rect 5012 26104 5021 26144
rect 4963 26103 5021 26104
rect 5259 26144 5301 26153
rect 5259 26104 5260 26144
rect 5300 26104 5301 26144
rect 3339 26090 3381 26099
rect 5259 26095 5301 26104
rect 5827 26144 5885 26145
rect 5827 26104 5836 26144
rect 5876 26104 5885 26144
rect 5827 26103 5885 26104
rect 7075 26144 7133 26145
rect 7075 26104 7084 26144
rect 7124 26104 7133 26144
rect 7075 26103 7133 26104
rect 7459 26144 7517 26145
rect 7459 26104 7468 26144
rect 7508 26104 7517 26144
rect 7459 26103 7517 26104
rect 8707 26144 8765 26145
rect 8707 26104 8716 26144
rect 8756 26104 8765 26144
rect 8707 26103 8765 26104
rect 9195 26144 9237 26153
rect 9195 26104 9196 26144
rect 9236 26104 9237 26144
rect 9195 26095 9237 26104
rect 9291 26144 9333 26153
rect 9291 26104 9292 26144
rect 9332 26104 9333 26144
rect 9291 26095 9333 26104
rect 9675 26144 9717 26153
rect 9675 26104 9676 26144
rect 9716 26104 9717 26144
rect 9675 26095 9717 26104
rect 10243 26144 10301 26145
rect 10243 26104 10252 26144
rect 10292 26104 10301 26144
rect 10243 26103 10301 26104
rect 10731 26139 10773 26148
rect 10731 26099 10732 26139
rect 10772 26099 10773 26139
rect 11107 26144 11165 26145
rect 11107 26104 11116 26144
rect 11156 26104 11165 26144
rect 11107 26103 11165 26104
rect 12355 26144 12413 26145
rect 12355 26104 12364 26144
rect 12404 26104 12413 26144
rect 12355 26103 12413 26104
rect 12843 26144 12885 26153
rect 12843 26104 12844 26144
rect 12884 26104 12885 26144
rect 10731 26090 10773 26099
rect 12843 26095 12885 26104
rect 12939 26144 12981 26153
rect 12939 26104 12940 26144
rect 12980 26104 12981 26144
rect 12939 26095 12981 26104
rect 13323 26144 13365 26153
rect 13323 26104 13324 26144
rect 13364 26104 13365 26144
rect 13323 26095 13365 26104
rect 13419 26144 13461 26153
rect 13419 26104 13420 26144
rect 13460 26104 13461 26144
rect 13419 26095 13461 26104
rect 13891 26144 13949 26145
rect 13891 26104 13900 26144
rect 13940 26104 13949 26144
rect 14947 26144 15005 26145
rect 13891 26103 13949 26104
rect 14379 26130 14421 26139
rect 14379 26090 14380 26130
rect 14420 26090 14421 26130
rect 14947 26104 14956 26144
rect 14996 26104 15005 26144
rect 14947 26103 15005 26104
rect 16195 26144 16253 26145
rect 16195 26104 16204 26144
rect 16244 26104 16253 26144
rect 16195 26103 16253 26104
rect 16387 26144 16445 26145
rect 16387 26104 16396 26144
rect 16436 26104 16445 26144
rect 16387 26103 16445 26104
rect 17635 26144 17693 26145
rect 17635 26104 17644 26144
rect 17684 26104 17693 26144
rect 17635 26103 17693 26104
rect 18115 26144 18173 26145
rect 18115 26104 18124 26144
rect 18164 26104 18173 26144
rect 18115 26103 18173 26104
rect 19363 26144 19421 26145
rect 19363 26104 19372 26144
rect 19412 26104 19421 26144
rect 19363 26103 19421 26104
rect 14379 26081 14421 26090
rect 2379 26060 2421 26069
rect 2379 26020 2380 26060
rect 2420 26020 2421 26060
rect 2379 26011 2421 26020
rect 4195 26060 4253 26061
rect 4195 26020 4204 26060
rect 4244 26020 4253 26060
rect 4195 26019 4253 26020
rect 4675 26060 4733 26061
rect 4675 26020 4684 26060
rect 4724 26020 4733 26060
rect 4675 26019 4733 26020
rect 9771 26060 9813 26069
rect 9771 26020 9772 26060
rect 9812 26020 9813 26060
rect 9771 26011 9813 26020
rect 19747 26060 19805 26061
rect 19747 26020 19756 26060
rect 19796 26020 19805 26060
rect 19747 26019 19805 26020
rect 3819 25976 3861 25985
rect 3819 25936 3820 25976
rect 3860 25936 3861 25976
rect 3819 25927 3861 25936
rect 5635 25976 5693 25977
rect 5635 25936 5644 25976
rect 5684 25936 5693 25976
rect 5635 25935 5693 25936
rect 4011 25892 4053 25901
rect 4011 25852 4012 25892
rect 4052 25852 4053 25892
rect 4011 25843 4053 25852
rect 8907 25892 8949 25901
rect 8907 25852 8908 25892
rect 8948 25852 8949 25892
rect 8907 25843 8949 25852
rect 14763 25892 14805 25901
rect 14763 25852 14764 25892
rect 14804 25852 14805 25892
rect 14763 25843 14805 25852
rect 17835 25892 17877 25901
rect 17835 25852 17836 25892
rect 17876 25852 17877 25892
rect 17835 25843 17877 25852
rect 19947 25892 19989 25901
rect 19947 25852 19948 25892
rect 19988 25852 19989 25892
rect 19947 25843 19989 25852
rect 1152 25724 20352 25748
rect 1152 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 20352 25724
rect 1152 25660 20352 25684
rect 2859 25556 2901 25565
rect 2859 25516 2860 25556
rect 2900 25516 2901 25556
rect 2859 25507 2901 25516
rect 6219 25556 6261 25565
rect 6219 25516 6220 25556
rect 6260 25516 6261 25556
rect 6219 25507 6261 25516
rect 10539 25556 10581 25565
rect 10539 25516 10540 25556
rect 10580 25516 10581 25556
rect 10539 25507 10581 25516
rect 12555 25556 12597 25565
rect 12555 25516 12556 25556
rect 12596 25516 12597 25556
rect 12555 25507 12597 25516
rect 14667 25556 14709 25565
rect 14667 25516 14668 25556
rect 14708 25516 14709 25556
rect 14667 25507 14709 25516
rect 3043 25388 3101 25389
rect 3043 25348 3052 25388
rect 3092 25348 3101 25388
rect 3043 25347 3101 25348
rect 4683 25388 4725 25397
rect 4683 25348 4684 25388
rect 4724 25348 4725 25388
rect 4683 25339 4725 25348
rect 6019 25388 6077 25389
rect 6019 25348 6028 25388
rect 6068 25348 6077 25388
rect 6019 25347 6077 25348
rect 10339 25388 10397 25389
rect 10339 25348 10348 25388
rect 10388 25348 10397 25388
rect 10339 25347 10397 25348
rect 12355 25388 12413 25389
rect 12355 25348 12364 25388
rect 12404 25348 12413 25388
rect 12355 25347 12413 25348
rect 14467 25388 14525 25389
rect 14467 25348 14476 25388
rect 14516 25348 14525 25388
rect 14467 25347 14525 25348
rect 15531 25388 15573 25397
rect 15531 25348 15532 25388
rect 15572 25348 15573 25388
rect 15531 25339 15573 25348
rect 19363 25388 19421 25389
rect 19363 25348 19372 25388
rect 19412 25348 19421 25388
rect 19363 25347 19421 25348
rect 19747 25388 19805 25389
rect 19747 25348 19756 25388
rect 19796 25348 19805 25388
rect 19747 25347 19805 25348
rect 3627 25309 3669 25318
rect 16539 25313 16581 25322
rect 1219 25304 1277 25305
rect 1219 25264 1228 25304
rect 1268 25264 1277 25304
rect 1219 25263 1277 25264
rect 2467 25304 2525 25305
rect 2467 25264 2476 25304
rect 2516 25264 2525 25304
rect 2467 25263 2525 25264
rect 3627 25269 3628 25309
rect 3668 25269 3669 25309
rect 3627 25260 3669 25269
rect 4099 25304 4157 25305
rect 4099 25264 4108 25304
rect 4148 25264 4157 25304
rect 4099 25263 4157 25264
rect 4587 25304 4629 25313
rect 4587 25264 4588 25304
rect 4628 25264 4629 25304
rect 4587 25255 4629 25264
rect 5067 25304 5109 25313
rect 5067 25264 5068 25304
rect 5108 25264 5109 25304
rect 5067 25255 5109 25264
rect 5163 25304 5205 25313
rect 5163 25264 5164 25304
rect 5204 25264 5205 25304
rect 5163 25255 5205 25264
rect 5547 25304 5589 25313
rect 5547 25264 5548 25304
rect 5588 25264 5589 25304
rect 5547 25255 5589 25264
rect 5643 25304 5685 25313
rect 5643 25264 5644 25304
rect 5684 25264 5685 25304
rect 5643 25255 5685 25264
rect 6403 25304 6461 25305
rect 6403 25264 6412 25304
rect 6452 25264 6461 25304
rect 6403 25263 6461 25264
rect 7651 25304 7709 25305
rect 7651 25264 7660 25304
rect 7700 25264 7709 25304
rect 7651 25263 7709 25264
rect 8035 25304 8093 25305
rect 8035 25264 8044 25304
rect 8084 25264 8093 25304
rect 8035 25263 8093 25264
rect 9283 25304 9341 25305
rect 9283 25264 9292 25304
rect 9332 25264 9341 25304
rect 9283 25263 9341 25264
rect 10723 25304 10781 25305
rect 10723 25264 10732 25304
rect 10772 25264 10781 25304
rect 10723 25263 10781 25264
rect 11971 25304 12029 25305
rect 11971 25264 11980 25304
rect 12020 25264 12029 25304
rect 11971 25263 12029 25264
rect 12739 25304 12797 25305
rect 12739 25264 12748 25304
rect 12788 25264 12797 25304
rect 12739 25263 12797 25264
rect 13987 25304 14045 25305
rect 13987 25264 13996 25304
rect 14036 25264 14045 25304
rect 13987 25263 14045 25264
rect 14955 25304 14997 25313
rect 14955 25264 14956 25304
rect 14996 25264 14997 25304
rect 14955 25255 14997 25264
rect 15051 25304 15093 25313
rect 15051 25264 15052 25304
rect 15092 25264 15093 25304
rect 15051 25255 15093 25264
rect 15435 25304 15477 25313
rect 15435 25264 15436 25304
rect 15476 25264 15477 25304
rect 15435 25255 15477 25264
rect 16003 25304 16061 25305
rect 16003 25264 16012 25304
rect 16052 25264 16061 25304
rect 16539 25273 16540 25313
rect 16580 25273 16581 25313
rect 16539 25264 16581 25273
rect 17259 25304 17301 25313
rect 17259 25264 17260 25304
rect 17300 25264 17301 25304
rect 16003 25263 16061 25264
rect 17259 25255 17301 25264
rect 17355 25304 17397 25313
rect 17355 25264 17356 25304
rect 17396 25264 17397 25304
rect 17355 25255 17397 25264
rect 17739 25304 17781 25313
rect 17739 25264 17740 25304
rect 17780 25264 17781 25304
rect 17739 25255 17781 25264
rect 17835 25304 17877 25313
rect 18795 25309 18837 25318
rect 17835 25264 17836 25304
rect 17876 25264 17877 25304
rect 17835 25255 17877 25264
rect 18307 25304 18365 25305
rect 18307 25264 18316 25304
rect 18356 25264 18365 25304
rect 18307 25263 18365 25264
rect 18795 25269 18796 25309
rect 18836 25269 18837 25309
rect 18795 25260 18837 25269
rect 3435 25220 3477 25229
rect 3435 25180 3436 25220
rect 3476 25180 3477 25220
rect 3435 25171 3477 25180
rect 16683 25220 16725 25229
rect 16683 25180 16684 25220
rect 16724 25180 16725 25220
rect 16683 25171 16725 25180
rect 18987 25220 19029 25229
rect 18987 25180 18988 25220
rect 19028 25180 19029 25220
rect 18987 25171 19029 25180
rect 2667 25136 2709 25145
rect 2667 25096 2668 25136
rect 2708 25096 2709 25136
rect 2667 25087 2709 25096
rect 5827 25136 5885 25137
rect 5827 25096 5836 25136
rect 5876 25096 5885 25136
rect 5827 25095 5885 25096
rect 7851 25136 7893 25145
rect 7851 25096 7852 25136
rect 7892 25096 7893 25136
rect 7851 25087 7893 25096
rect 9483 25136 9525 25145
rect 9483 25096 9484 25136
rect 9524 25096 9525 25136
rect 9483 25087 9525 25096
rect 12171 25136 12213 25145
rect 12171 25096 12172 25136
rect 12212 25096 12213 25136
rect 12171 25087 12213 25096
rect 14187 25136 14229 25145
rect 14187 25096 14188 25136
rect 14228 25096 14229 25136
rect 14187 25087 14229 25096
rect 19563 25136 19605 25145
rect 19563 25096 19564 25136
rect 19604 25096 19605 25136
rect 19563 25087 19605 25096
rect 19947 25136 19989 25145
rect 19947 25096 19948 25136
rect 19988 25096 19989 25136
rect 19947 25087 19989 25096
rect 1152 24968 20452 24992
rect 1152 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20452 24968
rect 1152 24904 20452 24928
rect 12171 24800 12213 24809
rect 12171 24760 12172 24800
rect 12212 24760 12213 24800
rect 12171 24751 12213 24760
rect 14475 24800 14517 24809
rect 14475 24760 14476 24800
rect 14516 24760 14517 24800
rect 14475 24751 14517 24760
rect 14955 24800 14997 24809
rect 14955 24760 14956 24800
rect 14996 24760 14997 24800
rect 14955 24751 14997 24760
rect 16587 24800 16629 24809
rect 16587 24760 16588 24800
rect 16628 24760 16629 24800
rect 16587 24751 16629 24760
rect 17259 24800 17301 24809
rect 17259 24760 17260 24800
rect 17300 24760 17301 24800
rect 17259 24751 17301 24760
rect 19275 24800 19317 24809
rect 19275 24760 19276 24800
rect 19316 24760 19317 24800
rect 19275 24751 19317 24760
rect 8139 24716 8181 24725
rect 8139 24676 8140 24716
rect 8180 24676 8181 24716
rect 8139 24667 8181 24676
rect 1219 24632 1277 24633
rect 1219 24592 1228 24632
rect 1268 24592 1277 24632
rect 1219 24591 1277 24592
rect 2467 24632 2525 24633
rect 2467 24592 2476 24632
rect 2516 24592 2525 24632
rect 2467 24591 2525 24592
rect 3043 24632 3101 24633
rect 3043 24592 3052 24632
rect 3092 24592 3101 24632
rect 3043 24591 3101 24592
rect 4291 24632 4349 24633
rect 4291 24592 4300 24632
rect 4340 24592 4349 24632
rect 4291 24591 4349 24592
rect 4675 24632 4733 24633
rect 4675 24592 4684 24632
rect 4724 24592 4733 24632
rect 4675 24591 4733 24592
rect 5923 24632 5981 24633
rect 5923 24592 5932 24632
rect 5972 24592 5981 24632
rect 5923 24591 5981 24592
rect 6411 24632 6453 24641
rect 6411 24592 6412 24632
rect 6452 24592 6453 24632
rect 6411 24583 6453 24592
rect 6507 24632 6549 24641
rect 6507 24592 6508 24632
rect 6548 24592 6549 24632
rect 6507 24583 6549 24592
rect 6891 24632 6933 24641
rect 6891 24592 6892 24632
rect 6932 24592 6933 24632
rect 6891 24583 6933 24592
rect 7459 24632 7517 24633
rect 7459 24592 7468 24632
rect 7508 24592 7517 24632
rect 7459 24591 7517 24592
rect 7947 24627 7989 24636
rect 7947 24587 7948 24627
rect 7988 24587 7989 24627
rect 8707 24632 8765 24633
rect 8707 24592 8716 24632
rect 8756 24592 8765 24632
rect 8707 24591 8765 24592
rect 9955 24632 10013 24633
rect 9955 24592 9964 24632
rect 10004 24592 10013 24632
rect 9955 24591 10013 24592
rect 10443 24632 10485 24641
rect 10443 24592 10444 24632
rect 10484 24592 10485 24632
rect 7947 24578 7989 24587
rect 10443 24583 10485 24592
rect 10539 24632 10581 24641
rect 10539 24592 10540 24632
rect 10580 24592 10581 24632
rect 10539 24583 10581 24592
rect 11491 24632 11549 24633
rect 11491 24592 11500 24632
rect 11540 24592 11549 24632
rect 12451 24632 12509 24633
rect 11491 24591 11549 24592
rect 12027 24590 12069 24599
rect 12451 24592 12460 24632
rect 12500 24592 12509 24632
rect 12451 24591 12509 24592
rect 12747 24632 12789 24641
rect 12747 24592 12748 24632
rect 12788 24592 12789 24632
rect 6987 24548 7029 24557
rect 6987 24508 6988 24548
rect 7028 24508 7029 24548
rect 6987 24499 7029 24508
rect 10923 24548 10965 24557
rect 10923 24508 10924 24548
rect 10964 24508 10965 24548
rect 10923 24499 10965 24508
rect 11019 24548 11061 24557
rect 11019 24508 11020 24548
rect 11060 24508 11061 24548
rect 12027 24550 12028 24590
rect 12068 24550 12069 24590
rect 12747 24583 12789 24592
rect 12843 24632 12885 24641
rect 12843 24592 12844 24632
rect 12884 24592 12885 24632
rect 12843 24583 12885 24592
rect 13795 24632 13853 24633
rect 13795 24592 13804 24632
rect 13844 24592 13853 24632
rect 13795 24591 13853 24592
rect 14283 24627 14325 24636
rect 14283 24587 14284 24627
rect 14324 24587 14325 24627
rect 15139 24632 15197 24633
rect 15139 24592 15148 24632
rect 15188 24592 15197 24632
rect 15139 24591 15197 24592
rect 16387 24632 16445 24633
rect 16387 24592 16396 24632
rect 16436 24592 16445 24632
rect 16387 24591 16445 24592
rect 17827 24632 17885 24633
rect 17827 24592 17836 24632
rect 17876 24592 17885 24632
rect 17827 24591 17885 24592
rect 19075 24632 19133 24633
rect 19075 24592 19084 24632
rect 19124 24592 19133 24632
rect 19075 24591 19133 24592
rect 19851 24632 19893 24641
rect 19851 24592 19852 24632
rect 19892 24592 19893 24632
rect 14283 24578 14325 24587
rect 19851 24583 19893 24592
rect 20043 24632 20085 24641
rect 20043 24592 20044 24632
rect 20084 24592 20085 24632
rect 20043 24583 20085 24592
rect 12027 24541 12069 24550
rect 12363 24548 12405 24557
rect 11019 24499 11061 24508
rect 12363 24508 12364 24548
rect 12404 24508 12405 24548
rect 12363 24499 12405 24508
rect 13227 24548 13269 24557
rect 13227 24508 13228 24548
rect 13268 24508 13269 24548
rect 13227 24499 13269 24508
rect 13323 24548 13365 24557
rect 13323 24508 13324 24548
rect 13364 24508 13365 24548
rect 13323 24499 13365 24508
rect 14755 24548 14813 24549
rect 14755 24508 14764 24548
rect 14804 24508 14813 24548
rect 14755 24507 14813 24508
rect 17059 24548 17117 24549
rect 17059 24508 17068 24548
rect 17108 24508 17117 24548
rect 17059 24507 17117 24508
rect 17443 24548 17501 24549
rect 17443 24508 17452 24548
rect 17492 24508 17501 24548
rect 17443 24507 17501 24508
rect 19459 24548 19517 24549
rect 19459 24508 19468 24548
rect 19508 24508 19517 24548
rect 19459 24507 19517 24508
rect 17643 24464 17685 24473
rect 17643 24424 17644 24464
rect 17684 24424 17685 24464
rect 17643 24415 17685 24424
rect 2667 24380 2709 24389
rect 2667 24340 2668 24380
rect 2708 24340 2709 24380
rect 2667 24331 2709 24340
rect 4491 24380 4533 24389
rect 4491 24340 4492 24380
rect 4532 24340 4533 24380
rect 4491 24331 4533 24340
rect 6123 24380 6165 24389
rect 6123 24340 6124 24380
rect 6164 24340 6165 24380
rect 6123 24331 6165 24340
rect 10155 24380 10197 24389
rect 10155 24340 10156 24380
rect 10196 24340 10197 24380
rect 10155 24331 10197 24340
rect 19659 24380 19701 24389
rect 19659 24340 19660 24380
rect 19700 24340 19701 24380
rect 19659 24331 19701 24340
rect 19851 24380 19893 24389
rect 19851 24340 19852 24380
rect 19892 24340 19893 24380
rect 19851 24331 19893 24340
rect 1152 24212 20352 24236
rect 1152 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 20352 24212
rect 1152 24148 20352 24172
rect 12747 24044 12789 24053
rect 12747 24004 12748 24044
rect 12788 24004 12789 24044
rect 12747 23995 12789 24004
rect 13227 24044 13269 24053
rect 13227 24004 13228 24044
rect 13268 24004 13269 24044
rect 13227 23995 13269 24004
rect 13611 24044 13653 24053
rect 13611 24004 13612 24044
rect 13652 24004 13653 24044
rect 13611 23995 13653 24004
rect 19755 24044 19797 24053
rect 19755 24004 19756 24044
rect 19796 24004 19797 24044
rect 19755 23995 19797 24004
rect 13995 23960 14037 23969
rect 13995 23920 13996 23960
rect 14036 23920 14037 23960
rect 13995 23911 14037 23920
rect 14379 23960 14421 23969
rect 14379 23920 14380 23960
rect 14420 23920 14421 23960
rect 14379 23911 14421 23920
rect 14763 23960 14805 23969
rect 14763 23920 14764 23960
rect 14804 23920 14805 23960
rect 14763 23911 14805 23920
rect 19371 23960 19413 23969
rect 19371 23920 19372 23960
rect 19412 23920 19413 23960
rect 19371 23911 19413 23920
rect 6699 23876 6741 23885
rect 6699 23836 6700 23876
rect 6740 23836 6741 23876
rect 6699 23827 6741 23836
rect 9771 23876 9813 23885
rect 9771 23836 9772 23876
rect 9812 23836 9813 23876
rect 9771 23827 9813 23836
rect 13027 23876 13085 23877
rect 13027 23836 13036 23876
rect 13076 23836 13085 23876
rect 13027 23835 13085 23836
rect 13411 23876 13469 23877
rect 13411 23836 13420 23876
rect 13460 23836 13469 23876
rect 13411 23835 13469 23836
rect 13795 23876 13853 23877
rect 13795 23836 13804 23876
rect 13844 23836 13853 23876
rect 13795 23835 13853 23836
rect 14179 23876 14237 23877
rect 14179 23836 14188 23876
rect 14228 23836 14237 23876
rect 14179 23835 14237 23836
rect 14563 23876 14621 23877
rect 14563 23836 14572 23876
rect 14612 23836 14621 23876
rect 14563 23835 14621 23836
rect 15531 23876 15573 23885
rect 15531 23836 15532 23876
rect 15572 23836 15573 23876
rect 15531 23827 15573 23836
rect 19939 23876 19997 23877
rect 19939 23836 19948 23876
rect 19988 23836 19997 23876
rect 19939 23835 19997 23836
rect 7659 23806 7701 23815
rect 1419 23792 1461 23801
rect 1419 23752 1420 23792
rect 1460 23752 1461 23792
rect 1419 23743 1461 23752
rect 1515 23792 1557 23801
rect 1515 23752 1516 23792
rect 1556 23752 1557 23792
rect 1515 23743 1557 23752
rect 1611 23792 1653 23801
rect 1611 23752 1612 23792
rect 1652 23752 1653 23792
rect 1611 23743 1653 23752
rect 1899 23792 1941 23801
rect 1899 23752 1900 23792
rect 1940 23752 1941 23792
rect 1899 23743 1941 23752
rect 1995 23792 2037 23801
rect 1995 23752 1996 23792
rect 2036 23752 2037 23792
rect 1995 23743 2037 23752
rect 2091 23792 2133 23801
rect 2091 23752 2092 23792
rect 2132 23752 2133 23792
rect 2091 23743 2133 23752
rect 2275 23792 2333 23793
rect 2275 23752 2284 23792
rect 2324 23752 2333 23792
rect 2275 23751 2333 23752
rect 3523 23792 3581 23793
rect 3523 23752 3532 23792
rect 3572 23752 3581 23792
rect 3523 23751 3581 23752
rect 4291 23792 4349 23793
rect 4291 23752 4300 23792
rect 4340 23752 4349 23792
rect 4291 23751 4349 23752
rect 5539 23792 5597 23793
rect 5539 23752 5548 23792
rect 5588 23752 5597 23792
rect 5539 23751 5597 23752
rect 6123 23792 6165 23801
rect 6123 23752 6124 23792
rect 6164 23752 6165 23792
rect 6123 23743 6165 23752
rect 6219 23792 6261 23801
rect 6219 23752 6220 23792
rect 6260 23752 6261 23792
rect 6219 23743 6261 23752
rect 6603 23792 6645 23801
rect 6603 23752 6604 23792
rect 6644 23752 6645 23792
rect 6603 23743 6645 23752
rect 7171 23792 7229 23793
rect 7171 23752 7180 23792
rect 7220 23752 7229 23792
rect 7659 23766 7660 23806
rect 7700 23766 7701 23806
rect 10827 23806 10869 23815
rect 7659 23757 7701 23766
rect 9291 23792 9333 23801
rect 7171 23751 7229 23752
rect 9291 23752 9292 23792
rect 9332 23752 9333 23792
rect 9291 23743 9333 23752
rect 9387 23792 9429 23801
rect 9387 23752 9388 23792
rect 9428 23752 9429 23792
rect 9387 23743 9429 23752
rect 9867 23792 9909 23801
rect 9867 23752 9868 23792
rect 9908 23752 9909 23792
rect 9867 23743 9909 23752
rect 10339 23792 10397 23793
rect 10339 23752 10348 23792
rect 10388 23752 10397 23792
rect 10827 23766 10828 23806
rect 10868 23766 10869 23806
rect 16635 23801 16677 23810
rect 10827 23757 10869 23766
rect 11299 23792 11357 23793
rect 10339 23751 10397 23752
rect 11299 23752 11308 23792
rect 11348 23752 11357 23792
rect 11299 23751 11357 23752
rect 12547 23792 12605 23793
rect 12547 23752 12556 23792
rect 12596 23752 12605 23792
rect 12547 23751 12605 23752
rect 15051 23792 15093 23801
rect 15051 23752 15052 23792
rect 15092 23752 15093 23792
rect 15051 23743 15093 23752
rect 15147 23792 15189 23801
rect 15147 23752 15148 23792
rect 15188 23752 15189 23792
rect 15147 23743 15189 23752
rect 15627 23792 15669 23801
rect 15627 23752 15628 23792
rect 15668 23752 15669 23792
rect 15627 23743 15669 23752
rect 16099 23792 16157 23793
rect 16099 23752 16108 23792
rect 16148 23752 16157 23792
rect 16635 23761 16636 23801
rect 16676 23761 16677 23801
rect 16635 23752 16677 23761
rect 17259 23797 17301 23806
rect 17259 23757 17260 23797
rect 17300 23757 17301 23797
rect 16099 23751 16157 23752
rect 17259 23748 17301 23757
rect 17731 23792 17789 23793
rect 17731 23752 17740 23792
rect 17780 23752 17789 23792
rect 17731 23751 17789 23752
rect 18219 23792 18261 23801
rect 18219 23752 18220 23792
rect 18260 23752 18261 23792
rect 18219 23743 18261 23752
rect 18315 23792 18357 23801
rect 18315 23752 18316 23792
rect 18356 23752 18357 23792
rect 18315 23743 18357 23752
rect 18699 23792 18741 23801
rect 18699 23752 18700 23792
rect 18740 23752 18741 23792
rect 18699 23743 18741 23752
rect 18795 23792 18837 23801
rect 18795 23752 18796 23792
rect 18836 23752 18837 23792
rect 18795 23743 18837 23752
rect 19075 23792 19133 23793
rect 19075 23752 19084 23792
rect 19124 23752 19133 23792
rect 19075 23751 19133 23752
rect 19179 23792 19221 23801
rect 19179 23752 19180 23792
rect 19220 23752 19221 23792
rect 19179 23743 19221 23752
rect 19371 23792 19413 23801
rect 19371 23752 19372 23792
rect 19412 23752 19413 23792
rect 19371 23743 19413 23752
rect 19563 23792 19605 23801
rect 19563 23752 19564 23792
rect 19604 23752 19605 23792
rect 19563 23743 19605 23752
rect 19755 23792 19797 23801
rect 19755 23752 19756 23792
rect 19796 23752 19797 23792
rect 19755 23743 19797 23752
rect 11019 23708 11061 23717
rect 11019 23668 11020 23708
rect 11060 23668 11061 23708
rect 11019 23659 11061 23668
rect 16779 23708 16821 23717
rect 16779 23668 16780 23708
rect 16820 23668 16821 23708
rect 16779 23659 16821 23668
rect 1315 23624 1373 23625
rect 1315 23584 1324 23624
rect 1364 23584 1373 23624
rect 1315 23583 1373 23584
rect 1795 23624 1853 23625
rect 1795 23584 1804 23624
rect 1844 23584 1853 23624
rect 1795 23583 1853 23584
rect 3723 23624 3765 23633
rect 3723 23584 3724 23624
rect 3764 23584 3765 23624
rect 3723 23575 3765 23584
rect 4011 23624 4053 23633
rect 4011 23584 4012 23624
rect 4052 23584 4053 23624
rect 4011 23575 4053 23584
rect 5739 23624 5781 23633
rect 5739 23584 5740 23624
rect 5780 23584 5781 23624
rect 5739 23575 5781 23584
rect 7851 23624 7893 23633
rect 7851 23584 7852 23624
rect 7892 23584 7893 23624
rect 7851 23575 7893 23584
rect 17067 23624 17109 23633
rect 17067 23584 17068 23624
rect 17108 23584 17109 23624
rect 17067 23575 17109 23584
rect 20139 23624 20181 23633
rect 20139 23584 20140 23624
rect 20180 23584 20181 23624
rect 20139 23575 20181 23584
rect 1152 23456 20452 23480
rect 1152 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20452 23456
rect 1152 23392 20452 23416
rect 1515 23288 1557 23297
rect 1515 23248 1516 23288
rect 1556 23248 1557 23288
rect 1515 23239 1557 23248
rect 3619 23288 3677 23289
rect 3619 23248 3628 23288
rect 3668 23248 3677 23288
rect 3619 23247 3677 23248
rect 6603 23288 6645 23297
rect 6603 23248 6604 23288
rect 6644 23248 6645 23288
rect 6603 23239 6645 23248
rect 13323 23288 13365 23297
rect 13323 23248 13324 23288
rect 13364 23248 13365 23288
rect 13323 23239 13365 23248
rect 14955 23288 14997 23297
rect 14955 23248 14956 23288
rect 14996 23248 14997 23288
rect 14955 23239 14997 23248
rect 16683 23288 16725 23297
rect 16683 23248 16684 23288
rect 16724 23248 16725 23288
rect 16683 23239 16725 23248
rect 17067 23288 17109 23297
rect 17067 23248 17068 23288
rect 17108 23248 17109 23288
rect 17067 23239 17109 23248
rect 19459 23288 19517 23289
rect 19459 23248 19468 23288
rect 19508 23248 19517 23288
rect 19459 23247 19517 23248
rect 5835 23204 5877 23213
rect 5835 23164 5836 23204
rect 5876 23164 5877 23204
rect 5835 23155 5877 23164
rect 1699 23120 1757 23121
rect 1699 23080 1708 23120
rect 1748 23080 1757 23120
rect 1699 23079 1757 23080
rect 2947 23120 3005 23121
rect 2947 23080 2956 23120
rect 2996 23080 3005 23120
rect 2947 23079 3005 23080
rect 3339 23120 3381 23129
rect 3339 23080 3340 23120
rect 3380 23080 3381 23120
rect 3339 23071 3381 23080
rect 3435 23120 3477 23129
rect 3435 23080 3436 23120
rect 3476 23080 3477 23120
rect 3435 23071 3477 23080
rect 4107 23120 4149 23129
rect 4107 23080 4108 23120
rect 4148 23080 4149 23120
rect 4107 23071 4149 23080
rect 4203 23120 4245 23129
rect 4203 23080 4204 23120
rect 4244 23080 4245 23120
rect 4203 23071 4245 23080
rect 4683 23120 4725 23129
rect 4683 23080 4684 23120
rect 4724 23080 4725 23120
rect 4683 23071 4725 23080
rect 5155 23120 5213 23121
rect 5155 23080 5164 23120
rect 5204 23080 5213 23120
rect 7075 23120 7133 23121
rect 5155 23079 5213 23080
rect 5691 23110 5733 23119
rect 5691 23070 5692 23110
rect 5732 23070 5733 23110
rect 7075 23080 7084 23120
rect 7124 23080 7133 23120
rect 7075 23079 7133 23080
rect 8323 23120 8381 23121
rect 8323 23080 8332 23120
rect 8372 23080 8381 23120
rect 8323 23079 8381 23080
rect 9475 23120 9533 23121
rect 9475 23080 9484 23120
rect 9524 23080 9533 23120
rect 9475 23079 9533 23080
rect 10723 23120 10781 23121
rect 10723 23080 10732 23120
rect 10772 23080 10781 23120
rect 10723 23079 10781 23080
rect 11395 23120 11453 23121
rect 11395 23080 11404 23120
rect 11444 23080 11453 23120
rect 11395 23079 11453 23080
rect 12643 23120 12701 23121
rect 12643 23080 12652 23120
rect 12692 23080 12701 23120
rect 12643 23079 12701 23080
rect 13507 23120 13565 23121
rect 13507 23080 13516 23120
rect 13556 23080 13565 23120
rect 13507 23079 13565 23080
rect 14755 23120 14813 23121
rect 14755 23080 14764 23120
rect 14804 23080 14813 23120
rect 14755 23079 14813 23080
rect 15235 23120 15293 23121
rect 15235 23080 15244 23120
rect 15284 23080 15293 23120
rect 15235 23079 15293 23080
rect 16483 23120 16541 23121
rect 16483 23080 16492 23120
rect 16532 23080 16541 23120
rect 16483 23079 16541 23080
rect 16971 23120 17013 23129
rect 16971 23080 16972 23120
rect 17012 23080 17013 23120
rect 16971 23071 17013 23080
rect 17163 23120 17205 23129
rect 17163 23080 17164 23120
rect 17204 23080 17205 23120
rect 17163 23071 17205 23080
rect 17347 23120 17405 23121
rect 17347 23080 17356 23120
rect 17396 23080 17405 23120
rect 17347 23079 17405 23080
rect 18595 23120 18653 23121
rect 18595 23080 18604 23120
rect 18644 23080 18653 23120
rect 18595 23079 18653 23080
rect 18987 23120 19029 23129
rect 18987 23080 18988 23120
rect 19028 23080 19029 23120
rect 18987 23071 19029 23080
rect 19179 23120 19221 23129
rect 19179 23080 19180 23120
rect 19220 23080 19221 23120
rect 19179 23071 19221 23080
rect 19275 23120 19317 23129
rect 19275 23080 19276 23120
rect 19316 23080 19317 23120
rect 19275 23071 19317 23080
rect 19563 23120 19605 23129
rect 19563 23080 19564 23120
rect 19604 23080 19605 23120
rect 19563 23071 19605 23080
rect 19659 23120 19701 23129
rect 19659 23080 19660 23120
rect 19700 23080 19701 23120
rect 19659 23071 19701 23080
rect 19755 23120 19797 23129
rect 19755 23080 19756 23120
rect 19796 23080 19797 23120
rect 20139 23120 20181 23129
rect 19755 23071 19797 23080
rect 19947 23109 19989 23118
rect 5691 23061 5733 23070
rect 19947 23069 19948 23109
rect 19988 23069 19989 23109
rect 20139 23080 20140 23120
rect 20180 23080 20181 23120
rect 20139 23071 20181 23080
rect 20227 23120 20285 23121
rect 20227 23080 20236 23120
rect 20276 23080 20285 23120
rect 20227 23079 20285 23080
rect 19947 23060 19989 23069
rect 1315 23036 1373 23037
rect 1315 22996 1324 23036
rect 1364 22996 1373 23036
rect 1315 22995 1373 22996
rect 4587 23036 4629 23045
rect 4587 22996 4588 23036
rect 4628 22996 4629 23036
rect 4587 22987 4629 22996
rect 6019 23036 6077 23037
rect 6019 22996 6028 23036
rect 6068 22996 6077 23036
rect 6019 22995 6077 22996
rect 6403 23036 6461 23037
rect 6403 22996 6412 23036
rect 6452 22996 6461 23036
rect 6403 22995 6461 22996
rect 13123 23036 13181 23037
rect 13123 22996 13132 23036
rect 13172 22996 13181 23036
rect 13123 22995 13181 22996
rect 3147 22868 3189 22877
rect 3147 22828 3148 22868
rect 3188 22828 3189 22868
rect 3147 22819 3189 22828
rect 6219 22868 6261 22877
rect 6219 22828 6220 22868
rect 6260 22828 6261 22868
rect 6219 22819 6261 22828
rect 8523 22868 8565 22877
rect 8523 22828 8524 22868
rect 8564 22828 8565 22868
rect 8523 22819 8565 22828
rect 10923 22868 10965 22877
rect 10923 22828 10924 22868
rect 10964 22828 10965 22868
rect 10923 22819 10965 22828
rect 12843 22868 12885 22877
rect 12843 22828 12844 22868
rect 12884 22828 12885 22868
rect 12843 22819 12885 22828
rect 18795 22868 18837 22877
rect 18795 22828 18796 22868
rect 18836 22828 18837 22868
rect 18795 22819 18837 22828
rect 19947 22868 19989 22877
rect 19947 22828 19948 22868
rect 19988 22828 19989 22868
rect 19947 22819 19989 22828
rect 1152 22700 20352 22724
rect 1152 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 20352 22700
rect 1152 22636 20352 22660
rect 1515 22532 1557 22541
rect 1515 22492 1516 22532
rect 1556 22492 1557 22532
rect 1515 22483 1557 22492
rect 1707 22532 1749 22541
rect 1707 22492 1708 22532
rect 1748 22492 1749 22532
rect 1707 22483 1749 22492
rect 4491 22532 4533 22541
rect 4491 22492 4492 22532
rect 4532 22492 4533 22532
rect 4491 22483 4533 22492
rect 13515 22532 13557 22541
rect 13515 22492 13516 22532
rect 13556 22492 13557 22532
rect 13515 22483 13557 22492
rect 19275 22532 19317 22541
rect 19275 22492 19276 22532
rect 19316 22492 19317 22532
rect 19275 22483 19317 22492
rect 4107 22448 4149 22457
rect 4107 22408 4108 22448
rect 4148 22408 4149 22448
rect 4107 22399 4149 22408
rect 4683 22448 4725 22457
rect 4683 22408 4684 22448
rect 4724 22408 4725 22448
rect 4683 22399 4725 22408
rect 1315 22364 1373 22365
rect 1315 22324 1324 22364
rect 1364 22324 1373 22364
rect 1315 22323 1373 22324
rect 1891 22364 1949 22365
rect 1891 22324 1900 22364
rect 1940 22324 1949 22364
rect 1891 22323 1949 22324
rect 4291 22364 4349 22365
rect 4291 22324 4300 22364
rect 4340 22324 4349 22364
rect 4291 22323 4349 22324
rect 7275 22364 7317 22373
rect 7275 22324 7276 22364
rect 7316 22324 7317 22364
rect 9675 22364 9717 22373
rect 2371 22322 2429 22323
rect 2371 22282 2380 22322
rect 2420 22282 2429 22322
rect 7275 22315 7317 22324
rect 8283 22322 8325 22331
rect 2371 22281 2429 22282
rect 3619 22280 3677 22281
rect 3619 22240 3628 22280
rect 3668 22240 3677 22280
rect 3619 22239 3677 22240
rect 4963 22280 5021 22281
rect 4963 22240 4972 22280
rect 5012 22240 5021 22280
rect 4963 22239 5021 22240
rect 6211 22280 6269 22281
rect 6211 22240 6220 22280
rect 6260 22240 6269 22280
rect 6211 22239 6269 22240
rect 6699 22280 6741 22289
rect 6699 22240 6700 22280
rect 6740 22240 6741 22280
rect 6699 22231 6741 22240
rect 6795 22280 6837 22289
rect 6795 22240 6796 22280
rect 6836 22240 6837 22280
rect 6795 22231 6837 22240
rect 7179 22280 7221 22289
rect 8283 22282 8284 22322
rect 8324 22282 8325 22322
rect 9675 22324 9676 22364
rect 9716 22324 9717 22364
rect 9675 22315 9717 22324
rect 13315 22364 13373 22365
rect 13315 22324 13324 22364
rect 13364 22324 13373 22364
rect 13315 22323 13373 22324
rect 19939 22364 19997 22365
rect 19939 22324 19948 22364
rect 19988 22324 19997 22364
rect 19939 22323 19997 22324
rect 10779 22289 10821 22298
rect 12747 22294 12789 22303
rect 7179 22240 7180 22280
rect 7220 22240 7221 22280
rect 7179 22231 7221 22240
rect 7747 22280 7805 22281
rect 7747 22240 7756 22280
rect 7796 22240 7805 22280
rect 8283 22273 8325 22282
rect 9195 22280 9237 22289
rect 7747 22239 7805 22240
rect 9195 22240 9196 22280
rect 9236 22240 9237 22280
rect 9195 22231 9237 22240
rect 9291 22280 9333 22289
rect 9291 22240 9292 22280
rect 9332 22240 9333 22280
rect 9291 22231 9333 22240
rect 9771 22280 9813 22289
rect 9771 22240 9772 22280
rect 9812 22240 9813 22280
rect 9771 22231 9813 22240
rect 10243 22280 10301 22281
rect 10243 22240 10252 22280
rect 10292 22240 10301 22280
rect 10779 22249 10780 22289
rect 10820 22249 10821 22289
rect 10779 22240 10821 22249
rect 11211 22280 11253 22289
rect 11211 22240 11212 22280
rect 11252 22240 11253 22280
rect 10243 22239 10301 22240
rect 11211 22231 11253 22240
rect 11307 22280 11349 22289
rect 11307 22240 11308 22280
rect 11348 22240 11349 22280
rect 11307 22231 11349 22240
rect 11691 22280 11733 22289
rect 11691 22240 11692 22280
rect 11732 22240 11733 22280
rect 11691 22231 11733 22240
rect 11787 22280 11829 22289
rect 11787 22240 11788 22280
rect 11828 22240 11829 22280
rect 11787 22231 11829 22240
rect 12259 22280 12317 22281
rect 12259 22240 12268 22280
rect 12308 22240 12317 22280
rect 12747 22254 12748 22294
rect 12788 22254 12789 22294
rect 12747 22245 12789 22254
rect 13803 22280 13845 22289
rect 12259 22239 12317 22240
rect 13803 22240 13804 22280
rect 13844 22240 13845 22280
rect 13803 22231 13845 22240
rect 13899 22280 13941 22289
rect 13899 22240 13900 22280
rect 13940 22240 13941 22280
rect 13899 22231 13941 22240
rect 14283 22280 14325 22289
rect 14283 22240 14284 22280
rect 14324 22240 14325 22280
rect 14283 22231 14325 22240
rect 14379 22280 14421 22289
rect 15339 22285 15381 22294
rect 14379 22240 14380 22280
rect 14420 22240 14421 22280
rect 14379 22231 14421 22240
rect 14851 22280 14909 22281
rect 14851 22240 14860 22280
rect 14900 22240 14909 22280
rect 14851 22239 14909 22240
rect 15339 22245 15340 22285
rect 15380 22245 15381 22285
rect 15339 22236 15381 22245
rect 15907 22280 15965 22281
rect 15907 22240 15916 22280
rect 15956 22240 15965 22280
rect 15907 22239 15965 22240
rect 17155 22280 17213 22281
rect 17155 22240 17164 22280
rect 17204 22240 17213 22280
rect 17155 22239 17213 22240
rect 17539 22280 17597 22281
rect 17539 22240 17548 22280
rect 17588 22240 17597 22280
rect 17539 22239 17597 22240
rect 17827 22280 17885 22281
rect 17827 22240 17836 22280
rect 17876 22240 17885 22280
rect 17827 22239 17885 22240
rect 19075 22280 19133 22281
rect 19075 22240 19084 22280
rect 19124 22240 19133 22280
rect 19075 22239 19133 22240
rect 19467 22280 19509 22289
rect 19467 22240 19468 22280
rect 19508 22240 19509 22280
rect 19467 22231 19509 22240
rect 19563 22280 19605 22289
rect 19563 22240 19564 22280
rect 19604 22240 19605 22280
rect 19563 22231 19605 22240
rect 19659 22280 19701 22289
rect 19659 22240 19660 22280
rect 19700 22240 19701 22280
rect 19659 22231 19701 22240
rect 19755 22280 19797 22289
rect 19755 22240 19756 22280
rect 19796 22240 19797 22280
rect 19755 22231 19797 22240
rect 2187 22196 2229 22205
rect 2187 22156 2188 22196
rect 2228 22156 2229 22196
rect 2187 22147 2229 22156
rect 15531 22196 15573 22205
rect 15531 22156 15532 22196
rect 15572 22156 15573 22196
rect 15531 22147 15573 22156
rect 17355 22196 17397 22205
rect 17355 22156 17356 22196
rect 17396 22156 17397 22196
rect 17355 22147 17397 22156
rect 3819 22112 3861 22121
rect 3819 22072 3820 22112
rect 3860 22072 3861 22112
rect 3819 22063 3861 22072
rect 6411 22112 6453 22121
rect 6411 22072 6412 22112
rect 6452 22072 6453 22112
rect 6411 22063 6453 22072
rect 8427 22112 8469 22121
rect 8427 22072 8428 22112
rect 8468 22072 8469 22112
rect 8427 22063 8469 22072
rect 10923 22112 10965 22121
rect 10923 22072 10924 22112
rect 10964 22072 10965 22112
rect 10923 22063 10965 22072
rect 12939 22112 12981 22121
rect 12939 22072 12940 22112
rect 12980 22072 12981 22112
rect 12939 22063 12981 22072
rect 17643 22112 17685 22121
rect 17643 22072 17644 22112
rect 17684 22072 17685 22112
rect 17643 22063 17685 22072
rect 20139 22112 20181 22121
rect 20139 22072 20140 22112
rect 20180 22072 20181 22112
rect 20139 22063 20181 22072
rect 1152 21944 20452 21968
rect 1152 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20452 21944
rect 1152 21880 20452 21904
rect 1515 21776 1557 21785
rect 1515 21736 1516 21776
rect 1556 21736 1557 21776
rect 1515 21727 1557 21736
rect 1899 21776 1941 21785
rect 1899 21736 1900 21776
rect 1940 21736 1941 21776
rect 1899 21727 1941 21736
rect 2283 21776 2325 21785
rect 2283 21736 2284 21776
rect 2324 21736 2325 21776
rect 2283 21727 2325 21736
rect 4299 21776 4341 21785
rect 4299 21736 4300 21776
rect 4340 21736 4341 21776
rect 4299 21727 4341 21736
rect 9483 21776 9525 21785
rect 9483 21736 9484 21776
rect 9524 21736 9525 21776
rect 9483 21727 9525 21736
rect 11115 21776 11157 21785
rect 11115 21736 11116 21776
rect 11156 21736 11157 21776
rect 11115 21727 11157 21736
rect 13707 21776 13749 21785
rect 13707 21736 13708 21776
rect 13748 21736 13749 21776
rect 13707 21727 13749 21736
rect 15339 21776 15381 21785
rect 15339 21736 15340 21776
rect 15380 21736 15381 21776
rect 15339 21727 15381 21736
rect 7851 21692 7893 21701
rect 7851 21652 7852 21692
rect 7892 21652 7893 21692
rect 7851 21643 7893 21652
rect 18603 21692 18645 21701
rect 18603 21652 18604 21692
rect 18644 21652 18645 21692
rect 18603 21643 18645 21652
rect 2571 21608 2613 21617
rect 2571 21568 2572 21608
rect 2612 21568 2613 21608
rect 2571 21559 2613 21568
rect 2667 21608 2709 21617
rect 2667 21568 2668 21608
rect 2708 21568 2709 21608
rect 2667 21559 2709 21568
rect 3051 21608 3093 21617
rect 3051 21568 3052 21608
rect 3092 21568 3093 21608
rect 3051 21559 3093 21568
rect 3147 21608 3189 21617
rect 3147 21568 3148 21608
rect 3188 21568 3189 21608
rect 3147 21559 3189 21568
rect 3619 21608 3677 21609
rect 3619 21568 3628 21608
rect 3668 21568 3677 21608
rect 3619 21567 3677 21568
rect 4107 21603 4149 21612
rect 4107 21563 4108 21603
rect 4148 21563 4149 21603
rect 4579 21608 4637 21609
rect 4579 21568 4588 21608
rect 4628 21568 4637 21608
rect 4579 21567 4637 21568
rect 4875 21608 4917 21617
rect 4875 21568 4876 21608
rect 4916 21568 4917 21608
rect 4107 21554 4149 21563
rect 4875 21559 4917 21568
rect 4971 21608 5013 21617
rect 4971 21568 4972 21608
rect 5012 21568 5013 21608
rect 4971 21559 5013 21568
rect 6123 21608 6165 21617
rect 6123 21568 6124 21608
rect 6164 21568 6165 21608
rect 6123 21559 6165 21568
rect 6219 21608 6261 21617
rect 6219 21568 6220 21608
rect 6260 21568 6261 21608
rect 6219 21559 6261 21568
rect 6603 21608 6645 21617
rect 6603 21568 6604 21608
rect 6644 21568 6645 21608
rect 6603 21559 6645 21568
rect 7171 21608 7229 21609
rect 7171 21568 7180 21608
rect 7220 21568 7229 21608
rect 7171 21567 7229 21568
rect 7659 21603 7701 21612
rect 7659 21563 7660 21603
rect 7700 21563 7701 21603
rect 8035 21608 8093 21609
rect 8035 21568 8044 21608
rect 8084 21568 8093 21608
rect 8035 21567 8093 21568
rect 9283 21608 9341 21609
rect 9283 21568 9292 21608
rect 9332 21568 9341 21608
rect 9283 21567 9341 21568
rect 9667 21608 9725 21609
rect 9667 21568 9676 21608
rect 9716 21568 9725 21608
rect 9667 21567 9725 21568
rect 10915 21608 10973 21609
rect 10915 21568 10924 21608
rect 10964 21568 10973 21608
rect 10915 21567 10973 21568
rect 12259 21608 12317 21609
rect 12259 21568 12268 21608
rect 12308 21568 12317 21608
rect 12259 21567 12317 21568
rect 13507 21608 13565 21609
rect 13507 21568 13516 21608
rect 13556 21568 13565 21608
rect 13507 21567 13565 21568
rect 13891 21608 13949 21609
rect 13891 21568 13900 21608
rect 13940 21568 13949 21608
rect 13891 21567 13949 21568
rect 15139 21608 15197 21609
rect 15139 21568 15148 21608
rect 15188 21568 15197 21608
rect 15139 21567 15197 21568
rect 15523 21608 15581 21609
rect 15523 21568 15532 21608
rect 15572 21568 15581 21608
rect 15523 21567 15581 21568
rect 16771 21608 16829 21609
rect 16771 21568 16780 21608
rect 16820 21568 16829 21608
rect 16771 21567 16829 21568
rect 17155 21608 17213 21609
rect 17155 21568 17164 21608
rect 17204 21568 17213 21608
rect 17155 21567 17213 21568
rect 18403 21608 18461 21609
rect 18403 21568 18412 21608
rect 18452 21568 18461 21608
rect 18403 21567 18461 21568
rect 18795 21608 18837 21617
rect 18795 21568 18796 21608
rect 18836 21568 18837 21608
rect 7659 21554 7701 21563
rect 18795 21559 18837 21568
rect 19083 21615 19125 21624
rect 19083 21575 19084 21615
rect 19124 21575 19125 21615
rect 19083 21566 19125 21575
rect 19275 21608 19317 21617
rect 19275 21568 19276 21608
rect 19316 21568 19317 21608
rect 19275 21559 19317 21568
rect 19371 21608 19413 21617
rect 19371 21568 19372 21608
rect 19412 21568 19413 21608
rect 19371 21559 19413 21568
rect 19467 21608 19509 21617
rect 19467 21568 19468 21608
rect 19508 21568 19509 21608
rect 19467 21559 19509 21568
rect 19563 21608 19605 21617
rect 19563 21568 19564 21608
rect 19604 21568 19605 21608
rect 19563 21559 19605 21568
rect 19755 21608 19797 21617
rect 19755 21568 19756 21608
rect 19796 21568 19797 21608
rect 19755 21559 19797 21568
rect 19947 21608 19989 21617
rect 19947 21568 19948 21608
rect 19988 21568 19989 21608
rect 19947 21559 19989 21568
rect 20035 21608 20093 21609
rect 20035 21568 20044 21608
rect 20084 21568 20093 21608
rect 20035 21567 20093 21568
rect 1315 21524 1373 21525
rect 1315 21484 1324 21524
rect 1364 21484 1373 21524
rect 1315 21483 1373 21484
rect 1699 21524 1757 21525
rect 1699 21484 1708 21524
rect 1748 21484 1757 21524
rect 1699 21483 1757 21484
rect 2083 21524 2141 21525
rect 2083 21484 2092 21524
rect 2132 21484 2141 21524
rect 2083 21483 2141 21484
rect 6699 21524 6741 21533
rect 6699 21484 6700 21524
rect 6740 21484 6741 21524
rect 6699 21475 6741 21484
rect 5251 21440 5309 21441
rect 5251 21400 5260 21440
rect 5300 21400 5309 21440
rect 5251 21399 5309 21400
rect 19755 21440 19797 21449
rect 19755 21400 19756 21440
rect 19796 21400 19797 21440
rect 19755 21391 19797 21400
rect 16971 21356 17013 21365
rect 16971 21316 16972 21356
rect 17012 21316 17013 21356
rect 16971 21307 17013 21316
rect 19083 21356 19125 21365
rect 19083 21316 19084 21356
rect 19124 21316 19125 21356
rect 19083 21307 19125 21316
rect 1152 21188 20352 21212
rect 1152 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 20352 21188
rect 1152 21124 20352 21148
rect 1515 21020 1557 21029
rect 1515 20980 1516 21020
rect 1556 20980 1557 21020
rect 1515 20971 1557 20980
rect 6795 21020 6837 21029
rect 6795 20980 6796 21020
rect 6836 20980 6837 21020
rect 6795 20971 6837 20980
rect 15339 21020 15381 21029
rect 15339 20980 15340 21020
rect 15380 20980 15381 21020
rect 15339 20971 15381 20980
rect 4491 20936 4533 20945
rect 4491 20896 4492 20936
rect 4532 20896 4533 20936
rect 4491 20887 4533 20896
rect 5163 20936 5205 20945
rect 5163 20896 5164 20936
rect 5204 20896 5205 20936
rect 5163 20887 5205 20896
rect 15723 20936 15765 20945
rect 15723 20896 15724 20936
rect 15764 20896 15765 20936
rect 15723 20887 15765 20896
rect 19275 20936 19317 20945
rect 19275 20896 19276 20936
rect 19316 20896 19317 20936
rect 19275 20887 19317 20896
rect 20043 20936 20085 20945
rect 20043 20896 20044 20936
rect 20084 20896 20085 20936
rect 20043 20887 20085 20896
rect 1315 20852 1373 20853
rect 1315 20812 1324 20852
rect 1364 20812 1373 20852
rect 1315 20811 1373 20812
rect 2859 20852 2901 20861
rect 2859 20812 2860 20852
rect 2900 20812 2901 20852
rect 2859 20803 2901 20812
rect 2955 20852 2997 20861
rect 2955 20812 2956 20852
rect 2996 20812 2997 20852
rect 4291 20852 4349 20853
rect 2955 20803 2997 20812
rect 3963 20810 4005 20819
rect 4291 20812 4300 20852
rect 4340 20812 4349 20852
rect 4291 20811 4349 20812
rect 13515 20852 13557 20861
rect 13515 20812 13516 20852
rect 13556 20812 13557 20852
rect 2379 20768 2421 20777
rect 2379 20728 2380 20768
rect 2420 20728 2421 20768
rect 2379 20719 2421 20728
rect 2475 20768 2517 20777
rect 3963 20770 3964 20810
rect 4004 20770 4005 20810
rect 13515 20803 13557 20812
rect 15139 20852 15197 20853
rect 15139 20812 15148 20852
rect 15188 20812 15197 20852
rect 15139 20811 15197 20812
rect 16971 20852 17013 20861
rect 16971 20812 16972 20852
rect 17012 20812 17013 20852
rect 16971 20803 17013 20812
rect 17067 20852 17109 20861
rect 17067 20812 17068 20852
rect 17108 20812 17109 20852
rect 17067 20803 17109 20812
rect 19179 20852 19221 20861
rect 19179 20812 19180 20852
rect 19220 20812 19221 20852
rect 19179 20803 19221 20812
rect 19371 20852 19413 20861
rect 19371 20812 19372 20852
rect 19412 20812 19413 20852
rect 19371 20803 19413 20812
rect 14619 20777 14661 20786
rect 18027 20782 18069 20791
rect 2475 20728 2476 20768
rect 2516 20728 2517 20768
rect 2475 20719 2517 20728
rect 3427 20768 3485 20769
rect 3427 20728 3436 20768
rect 3476 20728 3485 20768
rect 3963 20761 4005 20770
rect 5347 20768 5405 20769
rect 3427 20727 3485 20728
rect 5347 20728 5356 20768
rect 5396 20728 5405 20768
rect 5347 20727 5405 20728
rect 6595 20768 6653 20769
rect 6595 20728 6604 20768
rect 6644 20728 6653 20768
rect 6595 20727 6653 20728
rect 8035 20768 8093 20769
rect 8035 20728 8044 20768
rect 8084 20728 8093 20768
rect 8035 20727 8093 20728
rect 9283 20768 9341 20769
rect 9283 20728 9292 20768
rect 9332 20728 9341 20768
rect 9283 20727 9341 20728
rect 9667 20768 9725 20769
rect 9667 20728 9676 20768
rect 9716 20728 9725 20768
rect 9667 20727 9725 20728
rect 10915 20768 10973 20769
rect 10915 20728 10924 20768
rect 10964 20728 10973 20768
rect 10915 20727 10973 20728
rect 11299 20768 11357 20769
rect 11299 20728 11308 20768
rect 11348 20728 11357 20768
rect 11299 20727 11357 20728
rect 12547 20768 12605 20769
rect 12547 20728 12556 20768
rect 12596 20728 12605 20768
rect 12547 20727 12605 20728
rect 13035 20768 13077 20777
rect 13035 20728 13036 20768
rect 13076 20728 13077 20768
rect 13035 20719 13077 20728
rect 13131 20768 13173 20777
rect 13131 20728 13132 20768
rect 13172 20728 13173 20768
rect 13131 20719 13173 20728
rect 13611 20768 13653 20777
rect 13611 20728 13612 20768
rect 13652 20728 13653 20768
rect 13611 20719 13653 20728
rect 14083 20768 14141 20769
rect 14083 20728 14092 20768
rect 14132 20728 14141 20768
rect 14619 20737 14620 20777
rect 14660 20737 14661 20777
rect 14619 20728 14661 20737
rect 15531 20768 15573 20777
rect 15531 20728 15532 20768
rect 15572 20728 15573 20768
rect 14083 20727 14141 20728
rect 15531 20719 15573 20728
rect 15723 20768 15765 20777
rect 15723 20728 15724 20768
rect 15764 20728 15765 20768
rect 15723 20719 15765 20728
rect 15907 20768 15965 20769
rect 15907 20728 15916 20768
rect 15956 20728 15965 20768
rect 15907 20727 15965 20728
rect 16011 20768 16053 20777
rect 16011 20728 16012 20768
rect 16052 20728 16053 20768
rect 16011 20719 16053 20728
rect 16195 20768 16253 20769
rect 16195 20728 16204 20768
rect 16244 20728 16253 20768
rect 16195 20727 16253 20728
rect 16491 20768 16533 20777
rect 16491 20728 16492 20768
rect 16532 20728 16533 20768
rect 16491 20719 16533 20728
rect 16587 20768 16629 20777
rect 16587 20728 16588 20768
rect 16628 20728 16629 20768
rect 16587 20719 16629 20728
rect 17539 20768 17597 20769
rect 17539 20728 17548 20768
rect 17588 20728 17597 20768
rect 18027 20742 18028 20782
rect 18068 20742 18069 20782
rect 18027 20733 18069 20742
rect 18507 20768 18549 20777
rect 17539 20727 17597 20728
rect 18507 20728 18508 20768
rect 18548 20728 18549 20768
rect 18507 20719 18549 20728
rect 18603 20768 18645 20777
rect 18603 20728 18604 20768
rect 18644 20728 18645 20768
rect 18603 20719 18645 20728
rect 18699 20768 18741 20777
rect 18699 20728 18700 20768
rect 18740 20728 18741 20768
rect 18699 20719 18741 20728
rect 19075 20768 19133 20769
rect 19075 20728 19084 20768
rect 19124 20728 19133 20768
rect 19075 20727 19133 20728
rect 19467 20768 19509 20777
rect 19467 20728 19468 20768
rect 19508 20728 19509 20768
rect 19467 20719 19509 20728
rect 19659 20768 19701 20777
rect 19659 20728 19660 20768
rect 19700 20728 19701 20768
rect 19659 20719 19701 20728
rect 19851 20768 19893 20777
rect 19851 20728 19852 20768
rect 19892 20728 19893 20768
rect 19851 20719 19893 20728
rect 20043 20768 20085 20777
rect 20043 20728 20044 20768
rect 20084 20728 20085 20768
rect 20043 20719 20085 20728
rect 20235 20768 20277 20777
rect 20235 20728 20236 20768
rect 20276 20728 20277 20768
rect 20235 20719 20277 20728
rect 4107 20684 4149 20693
rect 4107 20644 4108 20684
rect 4148 20644 4149 20684
rect 4107 20635 4149 20644
rect 12747 20684 12789 20693
rect 12747 20644 12748 20684
rect 12788 20644 12789 20684
rect 12747 20635 12789 20644
rect 18219 20684 18261 20693
rect 18219 20644 18220 20684
rect 18260 20644 18261 20684
rect 18219 20635 18261 20644
rect 1699 20600 1757 20601
rect 1699 20560 1708 20600
rect 1748 20560 1757 20600
rect 1699 20559 1757 20560
rect 9483 20600 9525 20609
rect 9483 20560 9484 20600
rect 9524 20560 9525 20600
rect 9483 20551 9525 20560
rect 11115 20600 11157 20609
rect 11115 20560 11116 20600
rect 11156 20560 11157 20600
rect 11115 20551 11157 20560
rect 14763 20600 14805 20609
rect 14763 20560 14764 20600
rect 14804 20560 14805 20600
rect 14763 20551 14805 20560
rect 16203 20600 16245 20609
rect 16203 20560 16204 20600
rect 16244 20560 16245 20600
rect 16203 20551 16245 20560
rect 18403 20600 18461 20601
rect 18403 20560 18412 20600
rect 18452 20560 18461 20600
rect 18403 20559 18461 20560
rect 19755 20600 19797 20609
rect 19755 20560 19756 20600
rect 19796 20560 19797 20600
rect 19755 20551 19797 20560
rect 1152 20432 20452 20456
rect 1152 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20452 20432
rect 1152 20368 20452 20392
rect 12643 20264 12701 20265
rect 12643 20224 12652 20264
rect 12692 20224 12701 20264
rect 12643 20223 12701 20224
rect 18019 20264 18077 20265
rect 18019 20224 18028 20264
rect 18068 20224 18077 20264
rect 18019 20223 18077 20224
rect 2955 20180 2997 20189
rect 2955 20140 2956 20180
rect 2996 20140 2997 20180
rect 2955 20131 2997 20140
rect 6891 20180 6933 20189
rect 6891 20140 6892 20180
rect 6932 20140 6933 20180
rect 6891 20131 6933 20140
rect 7083 20180 7125 20189
rect 7083 20140 7084 20180
rect 7124 20140 7125 20180
rect 7083 20131 7125 20140
rect 11691 20180 11733 20189
rect 11691 20140 11692 20180
rect 11732 20140 11733 20180
rect 11691 20131 11733 20140
rect 14763 20180 14805 20189
rect 14763 20140 14764 20180
rect 14804 20140 14805 20180
rect 14763 20131 14805 20140
rect 17451 20180 17493 20189
rect 17451 20140 17452 20180
rect 17492 20140 17493 20180
rect 17451 20131 17493 20140
rect 1507 20096 1565 20097
rect 1507 20056 1516 20096
rect 1556 20056 1565 20096
rect 1507 20055 1565 20056
rect 2755 20096 2813 20097
rect 2755 20056 2764 20096
rect 2804 20056 2813 20096
rect 2755 20055 2813 20056
rect 3139 20096 3197 20097
rect 3139 20056 3148 20096
rect 3188 20056 3197 20096
rect 3139 20055 3197 20056
rect 4387 20096 4445 20097
rect 4387 20056 4396 20096
rect 4436 20056 4445 20096
rect 4387 20055 4445 20056
rect 5163 20096 5205 20105
rect 5163 20056 5164 20096
rect 5204 20056 5205 20096
rect 5163 20047 5205 20056
rect 5259 20096 5301 20105
rect 5259 20056 5260 20096
rect 5300 20056 5301 20096
rect 5259 20047 5301 20056
rect 6211 20096 6269 20097
rect 6211 20056 6220 20096
rect 6260 20056 6269 20096
rect 7747 20096 7805 20097
rect 6211 20055 6269 20056
rect 6699 20082 6741 20091
rect 6699 20042 6700 20082
rect 6740 20042 6741 20082
rect 6699 20033 6741 20042
rect 7275 20082 7317 20091
rect 7275 20042 7276 20082
rect 7316 20042 7317 20082
rect 7747 20056 7756 20096
rect 7796 20056 7805 20096
rect 7747 20055 7805 20056
rect 8715 20096 8757 20105
rect 8715 20056 8716 20096
rect 8756 20056 8757 20096
rect 8715 20047 8757 20056
rect 8811 20096 8853 20105
rect 8811 20056 8812 20096
rect 8852 20056 8853 20096
rect 8811 20047 8853 20056
rect 9963 20096 10005 20105
rect 9963 20056 9964 20096
rect 10004 20056 10005 20096
rect 9963 20047 10005 20056
rect 10059 20096 10101 20105
rect 10059 20056 10060 20096
rect 10100 20056 10101 20096
rect 10059 20047 10101 20056
rect 11011 20096 11069 20097
rect 11011 20056 11020 20096
rect 11060 20056 11069 20096
rect 11011 20055 11069 20056
rect 11499 20091 11541 20100
rect 11499 20051 11500 20091
rect 11540 20051 11541 20091
rect 12163 20096 12221 20097
rect 12163 20056 12172 20096
rect 12212 20056 12221 20096
rect 12163 20055 12221 20056
rect 12259 20096 12317 20097
rect 12259 20056 12268 20096
rect 12308 20056 12317 20096
rect 12259 20055 12317 20056
rect 12459 20096 12501 20105
rect 12459 20056 12460 20096
rect 12500 20056 12501 20096
rect 11499 20042 11541 20051
rect 12459 20047 12501 20056
rect 12555 20096 12597 20105
rect 12555 20056 12556 20096
rect 12596 20056 12597 20096
rect 13035 20096 13077 20105
rect 12555 20047 12597 20056
rect 12712 20081 12754 20090
rect 7275 20033 7317 20042
rect 12712 20041 12713 20081
rect 12753 20041 12754 20081
rect 13035 20056 13036 20096
rect 13076 20056 13077 20096
rect 13035 20047 13077 20056
rect 13131 20096 13173 20105
rect 13131 20056 13132 20096
rect 13172 20056 13173 20096
rect 13131 20047 13173 20056
rect 14083 20096 14141 20097
rect 14083 20056 14092 20096
rect 14132 20056 14141 20096
rect 14955 20096 14997 20105
rect 14083 20055 14141 20056
rect 14619 20054 14661 20063
rect 12712 20032 12754 20041
rect 4875 20012 4917 20021
rect 4875 19972 4876 20012
rect 4916 19972 4917 20012
rect 4875 19963 4917 19972
rect 5643 20012 5685 20021
rect 5643 19972 5644 20012
rect 5684 19972 5685 20012
rect 5643 19963 5685 19972
rect 5739 20012 5781 20021
rect 5739 19972 5740 20012
rect 5780 19972 5781 20012
rect 5739 19963 5781 19972
rect 8235 20012 8277 20021
rect 8235 19972 8236 20012
rect 8276 19972 8277 20012
rect 8235 19963 8277 19972
rect 8331 20012 8373 20021
rect 8331 19972 8332 20012
rect 8372 19972 8373 20012
rect 8331 19963 8373 19972
rect 10443 20012 10485 20021
rect 10443 19972 10444 20012
rect 10484 19972 10485 20012
rect 10443 19963 10485 19972
rect 10539 20012 10581 20021
rect 10539 19972 10540 20012
rect 10580 19972 10581 20012
rect 10539 19963 10581 19972
rect 13515 20012 13557 20021
rect 13515 19972 13516 20012
rect 13556 19972 13557 20012
rect 13515 19963 13557 19972
rect 13611 20012 13653 20021
rect 13611 19972 13612 20012
rect 13652 19972 13653 20012
rect 14619 20014 14620 20054
rect 14660 20014 14661 20054
rect 14955 20056 14956 20096
rect 14996 20056 14997 20096
rect 14955 20047 14997 20056
rect 15147 20096 15189 20105
rect 15147 20056 15148 20096
rect 15188 20056 15189 20096
rect 15147 20047 15189 20056
rect 15427 20096 15485 20097
rect 15427 20056 15436 20096
rect 15476 20056 15485 20096
rect 15427 20055 15485 20056
rect 15819 20096 15861 20105
rect 15819 20056 15820 20096
rect 15860 20056 15861 20096
rect 15819 20047 15861 20056
rect 16003 20096 16061 20097
rect 16003 20056 16012 20096
rect 16052 20056 16061 20096
rect 16003 20055 16061 20056
rect 17251 20096 17309 20097
rect 17251 20056 17260 20096
rect 17300 20056 17309 20096
rect 17251 20055 17309 20056
rect 17827 20096 17885 20097
rect 17827 20056 17836 20096
rect 17876 20056 17885 20096
rect 17827 20055 17885 20056
rect 17931 20096 17973 20105
rect 17931 20056 17932 20096
rect 17972 20056 17973 20096
rect 17931 20047 17973 20056
rect 18123 20096 18165 20105
rect 18123 20056 18124 20096
rect 18164 20056 18165 20096
rect 18123 20047 18165 20056
rect 18699 20096 18741 20105
rect 18699 20056 18700 20096
rect 18740 20056 18741 20096
rect 18307 20054 18365 20055
rect 14619 20005 14661 20014
rect 15531 20012 15573 20021
rect 13611 19963 13653 19972
rect 15531 19972 15532 20012
rect 15572 19972 15573 20012
rect 15531 19963 15573 19972
rect 15723 20012 15765 20021
rect 18307 20014 18316 20054
rect 18356 20014 18365 20054
rect 18699 20047 18741 20056
rect 19179 20096 19221 20105
rect 19179 20056 19180 20096
rect 19220 20056 19221 20096
rect 19179 20047 19221 20056
rect 19275 20096 19317 20105
rect 19275 20056 19276 20096
rect 19316 20056 19317 20096
rect 19275 20047 19317 20056
rect 19555 20096 19613 20097
rect 19555 20056 19564 20096
rect 19604 20056 19613 20096
rect 19555 20055 19613 20056
rect 19843 20096 19901 20097
rect 19843 20056 19852 20096
rect 19892 20056 19901 20096
rect 19843 20055 19901 20056
rect 19947 20096 19989 20105
rect 19947 20056 19948 20096
rect 19988 20056 19989 20096
rect 19947 20047 19989 20056
rect 20131 20054 20189 20055
rect 18307 20013 18365 20014
rect 15723 19972 15724 20012
rect 15764 19972 15765 20012
rect 15723 19963 15765 19972
rect 18411 20012 18453 20021
rect 18411 19972 18412 20012
rect 18452 19972 18453 20012
rect 18411 19963 18453 19972
rect 18603 20012 18645 20021
rect 20131 20014 20140 20054
rect 20180 20014 20189 20054
rect 20131 20013 20189 20014
rect 18603 19972 18604 20012
rect 18644 19972 18645 20012
rect 18603 19963 18645 19972
rect 1323 19928 1365 19937
rect 1323 19888 1324 19928
rect 1364 19888 1365 19928
rect 1323 19879 1365 19888
rect 4587 19928 4629 19937
rect 4587 19888 4588 19928
rect 4628 19888 4629 19928
rect 4587 19879 4629 19888
rect 15627 19928 15669 19937
rect 15627 19888 15628 19928
rect 15668 19888 15669 19928
rect 18883 19928 18941 19929
rect 15627 19879 15669 19888
rect 18507 19886 18549 19895
rect 18883 19888 18892 19928
rect 18932 19888 18941 19928
rect 18883 19887 18941 19888
rect 15147 19844 15189 19853
rect 15147 19804 15148 19844
rect 15188 19804 15189 19844
rect 18507 19846 18508 19886
rect 18548 19846 18549 19886
rect 18507 19837 18549 19846
rect 19947 19844 19989 19853
rect 15147 19795 15189 19804
rect 19947 19804 19948 19844
rect 19988 19804 19989 19844
rect 19947 19795 19989 19804
rect 1152 19676 20352 19700
rect 1152 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 20352 19676
rect 1152 19612 20352 19636
rect 1707 19508 1749 19517
rect 1707 19468 1708 19508
rect 1748 19468 1749 19508
rect 1707 19459 1749 19468
rect 7371 19508 7413 19517
rect 7371 19468 7372 19508
rect 7412 19468 7413 19508
rect 7371 19459 7413 19468
rect 13035 19508 13077 19517
rect 13035 19468 13036 19508
rect 13076 19468 13077 19508
rect 13035 19459 13077 19468
rect 14763 19508 14805 19517
rect 14763 19468 14764 19508
rect 14804 19468 14805 19508
rect 14763 19459 14805 19468
rect 16395 19508 16437 19517
rect 16395 19468 16396 19508
rect 16436 19468 16437 19508
rect 16395 19459 16437 19468
rect 17547 19508 17589 19517
rect 17547 19468 17548 19508
rect 17588 19468 17589 19508
rect 17547 19459 17589 19468
rect 5163 19424 5205 19433
rect 5163 19384 5164 19424
rect 5204 19384 5205 19424
rect 5163 19375 5205 19384
rect 1323 19340 1365 19349
rect 1323 19300 1324 19340
rect 1364 19300 1365 19340
rect 1323 19291 1365 19300
rect 1507 19340 1565 19341
rect 1507 19300 1516 19340
rect 1556 19300 1565 19340
rect 1507 19299 1565 19300
rect 3243 19340 3285 19349
rect 3243 19300 3244 19340
rect 3284 19300 3285 19340
rect 3243 19291 3285 19300
rect 2763 19256 2805 19265
rect 2763 19216 2764 19256
rect 2804 19216 2805 19256
rect 2763 19207 2805 19216
rect 2859 19256 2901 19265
rect 2859 19216 2860 19256
rect 2900 19216 2901 19256
rect 2859 19207 2901 19216
rect 3339 19256 3381 19265
rect 4299 19261 4341 19270
rect 3339 19216 3340 19256
rect 3380 19216 3381 19256
rect 3339 19207 3381 19216
rect 3811 19256 3869 19257
rect 3811 19216 3820 19256
rect 3860 19216 3869 19256
rect 3811 19215 3869 19216
rect 4299 19221 4300 19261
rect 4340 19221 4341 19261
rect 4299 19212 4341 19221
rect 5731 19256 5789 19257
rect 5731 19216 5740 19256
rect 5780 19216 5789 19256
rect 5731 19215 5789 19216
rect 6979 19256 7037 19257
rect 6979 19216 6988 19256
rect 7028 19216 7037 19256
rect 6979 19215 7037 19216
rect 7555 19256 7613 19257
rect 7555 19216 7564 19256
rect 7604 19216 7613 19256
rect 7555 19215 7613 19216
rect 8803 19256 8861 19257
rect 8803 19216 8812 19256
rect 8852 19216 8861 19256
rect 8803 19215 8861 19216
rect 9675 19256 9717 19265
rect 9675 19216 9676 19256
rect 9716 19216 9717 19256
rect 9675 19207 9717 19216
rect 9771 19256 9813 19265
rect 9771 19216 9772 19256
rect 9812 19216 9813 19256
rect 9771 19207 9813 19216
rect 10155 19256 10197 19265
rect 10155 19216 10156 19256
rect 10196 19216 10197 19256
rect 10155 19207 10197 19216
rect 10251 19256 10293 19265
rect 11211 19261 11253 19270
rect 10251 19216 10252 19256
rect 10292 19216 10293 19256
rect 10251 19207 10293 19216
rect 10723 19256 10781 19257
rect 10723 19216 10732 19256
rect 10772 19216 10781 19256
rect 10723 19215 10781 19216
rect 11211 19221 11212 19261
rect 11252 19221 11253 19261
rect 11211 19212 11253 19221
rect 11587 19256 11645 19257
rect 11587 19216 11596 19256
rect 11636 19216 11645 19256
rect 11587 19215 11645 19216
rect 12835 19256 12893 19257
rect 12835 19216 12844 19256
rect 12884 19216 12893 19256
rect 12835 19215 12893 19216
rect 13315 19256 13373 19257
rect 13315 19216 13324 19256
rect 13364 19216 13373 19256
rect 13315 19215 13373 19216
rect 14563 19256 14621 19257
rect 14563 19216 14572 19256
rect 14612 19216 14621 19256
rect 14563 19215 14621 19216
rect 14947 19256 15005 19257
rect 14947 19216 14956 19256
rect 14996 19216 15005 19256
rect 14947 19215 15005 19216
rect 16195 19256 16253 19257
rect 16195 19216 16204 19256
rect 16244 19216 16253 19256
rect 16195 19215 16253 19216
rect 16579 19256 16637 19257
rect 16579 19216 16588 19256
rect 16628 19216 16637 19256
rect 16579 19215 16637 19216
rect 16675 19256 16733 19257
rect 16675 19216 16684 19256
rect 16724 19216 16733 19256
rect 16675 19215 16733 19216
rect 16875 19256 16917 19265
rect 16875 19216 16876 19256
rect 16916 19216 16917 19256
rect 16875 19207 16917 19216
rect 16971 19256 17013 19265
rect 16971 19216 16972 19256
rect 17012 19216 17013 19256
rect 16971 19207 17013 19216
rect 17118 19256 17176 19257
rect 17118 19216 17127 19256
rect 17167 19216 17176 19256
rect 17118 19215 17176 19216
rect 17355 19256 17397 19265
rect 17355 19216 17356 19256
rect 17396 19216 17397 19256
rect 17355 19207 17397 19216
rect 17547 19256 17589 19265
rect 17547 19216 17548 19256
rect 17588 19216 17589 19256
rect 17547 19207 17589 19216
rect 17731 19256 17789 19257
rect 17731 19216 17740 19256
rect 17780 19216 17789 19256
rect 17731 19215 17789 19216
rect 18979 19256 19037 19257
rect 18979 19216 18988 19256
rect 19028 19216 19037 19256
rect 18979 19215 19037 19216
rect 19459 19256 19517 19257
rect 19459 19216 19468 19256
rect 19508 19216 19517 19256
rect 19459 19215 19517 19216
rect 19755 19256 19797 19265
rect 19755 19216 19756 19256
rect 19796 19216 19797 19256
rect 19755 19207 19797 19216
rect 11403 19172 11445 19181
rect 11403 19132 11404 19172
rect 11444 19132 11445 19172
rect 11403 19123 11445 19132
rect 19179 19172 19221 19181
rect 19179 19132 19180 19172
rect 19220 19132 19221 19172
rect 19179 19123 19221 19132
rect 19851 19172 19893 19181
rect 19851 19132 19852 19172
rect 19892 19132 19893 19172
rect 19851 19123 19893 19132
rect 4491 19088 4533 19097
rect 4491 19048 4492 19088
rect 4532 19048 4533 19088
rect 4491 19039 4533 19048
rect 7179 19088 7221 19097
rect 7179 19048 7180 19088
rect 7220 19048 7221 19088
rect 7179 19039 7221 19048
rect 16395 19088 16437 19097
rect 16395 19048 16396 19088
rect 16436 19048 16437 19088
rect 16395 19039 16437 19048
rect 16963 19088 17021 19089
rect 16963 19048 16972 19088
rect 17012 19048 17021 19088
rect 16963 19047 17021 19048
rect 20139 19046 20181 19055
rect 20139 19006 20140 19046
rect 20180 19006 20181 19046
rect 20139 18997 20181 19006
rect 1152 18920 20452 18944
rect 1152 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20452 18920
rect 1152 18856 20452 18880
rect 6987 18752 7029 18761
rect 6987 18712 6988 18752
rect 7028 18712 7029 18752
rect 6987 18703 7029 18712
rect 9483 18752 9525 18761
rect 9483 18712 9484 18752
rect 9524 18712 9525 18752
rect 9483 18703 9525 18712
rect 11115 18752 11157 18761
rect 11115 18712 11116 18752
rect 11156 18712 11157 18752
rect 11115 18703 11157 18712
rect 13227 18752 13269 18761
rect 13227 18712 13228 18752
rect 13268 18712 13269 18752
rect 13227 18703 13269 18712
rect 14859 18752 14901 18761
rect 14859 18712 14860 18752
rect 14900 18712 14901 18752
rect 14859 18703 14901 18712
rect 19179 18752 19221 18761
rect 19179 18712 19180 18752
rect 19220 18712 19221 18752
rect 19179 18703 19221 18712
rect 19555 18752 19613 18753
rect 19555 18712 19564 18752
rect 19604 18712 19613 18752
rect 19555 18711 19613 18712
rect 4395 18668 4437 18677
rect 4395 18628 4396 18668
rect 4436 18628 4437 18668
rect 4395 18619 4437 18628
rect 5067 18668 5109 18677
rect 5067 18628 5068 18668
rect 5108 18628 5109 18668
rect 5067 18619 5109 18628
rect 15043 18626 15101 18627
rect 2083 18584 2141 18585
rect 2083 18544 2092 18584
rect 2132 18544 2141 18584
rect 2083 18543 2141 18544
rect 2667 18584 2709 18593
rect 2667 18544 2668 18584
rect 2708 18544 2709 18584
rect 2667 18535 2709 18544
rect 2763 18584 2805 18593
rect 2763 18544 2764 18584
rect 2804 18544 2805 18584
rect 2763 18535 2805 18544
rect 3715 18584 3773 18585
rect 3715 18544 3724 18584
rect 3764 18544 3773 18584
rect 4675 18584 4733 18585
rect 3715 18543 3773 18544
rect 4203 18570 4245 18579
rect 4203 18530 4204 18570
rect 4244 18530 4245 18570
rect 4675 18544 4684 18584
rect 4724 18544 4733 18584
rect 4675 18543 4733 18544
rect 4971 18584 5013 18593
rect 4971 18544 4972 18584
rect 5012 18544 5013 18584
rect 4971 18535 5013 18544
rect 5539 18584 5597 18585
rect 5539 18544 5548 18584
rect 5588 18544 5597 18584
rect 5539 18543 5597 18544
rect 6787 18584 6845 18585
rect 6787 18544 6796 18584
rect 6836 18544 6845 18584
rect 6787 18543 6845 18544
rect 8035 18584 8093 18585
rect 8035 18544 8044 18584
rect 8084 18544 8093 18584
rect 8035 18543 8093 18544
rect 9283 18584 9341 18585
rect 9283 18544 9292 18584
rect 9332 18544 9341 18584
rect 9283 18543 9341 18544
rect 9667 18584 9725 18585
rect 9667 18544 9676 18584
rect 9716 18544 9725 18584
rect 9667 18543 9725 18544
rect 10915 18584 10973 18585
rect 10915 18544 10924 18584
rect 10964 18544 10973 18584
rect 10915 18543 10973 18544
rect 11299 18584 11357 18585
rect 11299 18544 11308 18584
rect 11348 18544 11357 18584
rect 11299 18543 11357 18544
rect 11403 18584 11445 18593
rect 15043 18586 15052 18626
rect 15092 18586 15101 18626
rect 15043 18585 15101 18586
rect 11403 18544 11404 18584
rect 11444 18544 11445 18584
rect 11403 18535 11445 18544
rect 11587 18584 11645 18585
rect 11587 18544 11596 18584
rect 11636 18544 11645 18584
rect 11587 18543 11645 18544
rect 11779 18584 11837 18585
rect 11779 18544 11788 18584
rect 11828 18544 11837 18584
rect 11779 18543 11837 18544
rect 13027 18584 13085 18585
rect 13027 18544 13036 18584
rect 13076 18544 13085 18584
rect 13027 18543 13085 18544
rect 13411 18584 13469 18585
rect 13411 18544 13420 18584
rect 13460 18544 13469 18584
rect 13411 18543 13469 18544
rect 14659 18584 14717 18585
rect 14659 18544 14668 18584
rect 14708 18544 14717 18584
rect 14659 18543 14717 18544
rect 16291 18584 16349 18585
rect 16291 18544 16300 18584
rect 16340 18544 16349 18584
rect 16291 18543 16349 18544
rect 16771 18584 16829 18585
rect 16771 18544 16780 18584
rect 16820 18544 16829 18584
rect 16771 18543 16829 18544
rect 17067 18584 17109 18593
rect 17067 18544 17068 18584
rect 17108 18544 17109 18584
rect 17067 18535 17109 18544
rect 17163 18584 17205 18593
rect 17163 18544 17164 18584
rect 17204 18544 17205 18584
rect 17163 18535 17205 18544
rect 17731 18584 17789 18585
rect 17731 18544 17740 18584
rect 17780 18544 17789 18584
rect 17731 18543 17789 18544
rect 18979 18584 19037 18585
rect 18979 18544 18988 18584
rect 19028 18544 19037 18584
rect 18979 18543 19037 18544
rect 19363 18584 19421 18585
rect 19363 18544 19372 18584
rect 19412 18544 19421 18584
rect 19363 18543 19421 18544
rect 19459 18584 19517 18585
rect 19459 18544 19468 18584
rect 19508 18544 19517 18584
rect 19459 18543 19517 18544
rect 19659 18584 19701 18593
rect 19659 18544 19660 18584
rect 19700 18544 19701 18584
rect 19659 18535 19701 18544
rect 19755 18584 19797 18593
rect 19755 18544 19756 18584
rect 19796 18544 19797 18584
rect 19755 18535 19797 18544
rect 19902 18584 19960 18585
rect 19902 18544 19911 18584
rect 19951 18544 19960 18584
rect 19902 18543 19960 18544
rect 20131 18584 20189 18585
rect 20131 18544 20140 18584
rect 20180 18544 20189 18584
rect 20131 18543 20189 18544
rect 4203 18521 4245 18530
rect 3147 18500 3189 18509
rect 3147 18460 3148 18500
rect 3188 18460 3189 18500
rect 3147 18451 3189 18460
rect 3243 18500 3285 18509
rect 3243 18460 3244 18500
rect 3284 18460 3285 18500
rect 3243 18451 3285 18460
rect 1515 18416 1557 18425
rect 1515 18376 1516 18416
rect 1556 18376 1557 18416
rect 1515 18367 1557 18376
rect 1803 18416 1845 18425
rect 1803 18376 1804 18416
rect 1844 18376 1845 18416
rect 1803 18367 1845 18376
rect 16491 18416 16533 18425
rect 16491 18376 16492 18416
rect 16532 18376 16533 18416
rect 16491 18367 16533 18376
rect 17443 18416 17501 18417
rect 17443 18376 17452 18416
rect 17492 18376 17501 18416
rect 17443 18375 17501 18376
rect 1995 18332 2037 18341
rect 1995 18292 1996 18332
rect 2036 18292 2037 18332
rect 1995 18283 2037 18292
rect 5347 18332 5405 18333
rect 5347 18292 5356 18332
rect 5396 18292 5405 18332
rect 5347 18291 5405 18292
rect 11595 18332 11637 18341
rect 11595 18292 11596 18332
rect 11636 18292 11637 18332
rect 11595 18283 11637 18292
rect 20235 18332 20277 18341
rect 20235 18292 20236 18332
rect 20276 18292 20277 18332
rect 20235 18283 20277 18292
rect 1152 18164 20352 18188
rect 1152 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 20352 18164
rect 1152 18100 20352 18124
rect 2667 17996 2709 18005
rect 2667 17956 2668 17996
rect 2708 17956 2709 17996
rect 2667 17947 2709 17956
rect 4299 17996 4341 18005
rect 4299 17956 4300 17996
rect 4340 17956 4341 17996
rect 4299 17947 4341 17956
rect 13131 17996 13173 18005
rect 13131 17956 13132 17996
rect 13172 17956 13173 17996
rect 13131 17947 13173 17956
rect 13315 17996 13373 17997
rect 13315 17956 13324 17996
rect 13364 17956 13373 17996
rect 16299 17996 16341 18005
rect 13315 17955 13373 17956
rect 14475 17954 14517 17963
rect 14475 17914 14476 17954
rect 14516 17914 14517 17954
rect 16299 17956 16300 17996
rect 16340 17956 16341 17996
rect 16299 17947 16341 17956
rect 16483 17996 16541 17997
rect 16483 17956 16492 17996
rect 16532 17956 16541 17996
rect 16483 17955 16541 17956
rect 17547 17996 17589 18005
rect 17547 17956 17548 17996
rect 17588 17956 17589 17996
rect 17547 17947 17589 17956
rect 19179 17996 19221 18005
rect 19179 17956 19180 17996
rect 19220 17956 19221 17996
rect 19179 17947 19221 17956
rect 19947 17996 19989 18005
rect 19947 17956 19948 17996
rect 19988 17956 19989 17996
rect 19947 17947 19989 17956
rect 8899 17912 8957 17913
rect 8899 17872 8908 17912
rect 8948 17872 8957 17912
rect 14475 17905 14517 17914
rect 8899 17871 8957 17872
rect 14379 17870 14421 17879
rect 6699 17828 6741 17837
rect 6699 17788 6700 17828
rect 6740 17788 6741 17828
rect 6699 17779 6741 17788
rect 6795 17828 6837 17837
rect 6795 17788 6796 17828
rect 6836 17788 6837 17828
rect 14379 17830 14380 17870
rect 14420 17830 14421 17870
rect 14379 17821 14421 17830
rect 14571 17828 14613 17837
rect 6795 17779 6837 17788
rect 14283 17786 14325 17795
rect 1219 17744 1277 17745
rect 1219 17704 1228 17744
rect 1268 17704 1277 17744
rect 1219 17703 1277 17704
rect 2467 17744 2525 17745
rect 2467 17704 2476 17744
rect 2516 17704 2525 17744
rect 2467 17703 2525 17704
rect 2851 17744 2909 17745
rect 2851 17704 2860 17744
rect 2900 17704 2909 17744
rect 2851 17703 2909 17704
rect 4099 17744 4157 17745
rect 4099 17704 4108 17744
rect 4148 17704 4157 17744
rect 4099 17703 4157 17704
rect 4483 17744 4541 17745
rect 4483 17704 4492 17744
rect 4532 17704 4541 17744
rect 4483 17703 4541 17704
rect 5731 17744 5789 17745
rect 5731 17704 5740 17744
rect 5780 17704 5789 17744
rect 5731 17703 5789 17704
rect 6219 17744 6261 17753
rect 6219 17704 6220 17744
rect 6260 17704 6261 17744
rect 6219 17695 6261 17704
rect 6315 17744 6357 17753
rect 7755 17749 7797 17758
rect 6315 17704 6316 17744
rect 6356 17704 6357 17744
rect 6315 17695 6357 17704
rect 7267 17744 7325 17745
rect 7267 17704 7276 17744
rect 7316 17704 7325 17744
rect 7267 17703 7325 17704
rect 7755 17709 7756 17749
rect 7796 17709 7797 17749
rect 7755 17700 7797 17709
rect 8227 17744 8285 17745
rect 8227 17704 8236 17744
rect 8276 17704 8285 17744
rect 8227 17703 8285 17704
rect 8523 17744 8565 17753
rect 8523 17704 8524 17744
rect 8564 17704 8565 17744
rect 8523 17695 8565 17704
rect 9187 17744 9245 17745
rect 9187 17704 9196 17744
rect 9236 17704 9245 17744
rect 9187 17703 9245 17704
rect 9571 17744 9629 17745
rect 9571 17704 9580 17744
rect 9620 17704 9629 17744
rect 9571 17703 9629 17704
rect 10819 17744 10877 17745
rect 10819 17704 10828 17744
rect 10868 17704 10877 17744
rect 10819 17703 10877 17704
rect 11395 17744 11453 17745
rect 11395 17704 11404 17744
rect 11444 17704 11453 17744
rect 11395 17703 11453 17704
rect 12643 17744 12701 17745
rect 12643 17704 12652 17744
rect 12692 17704 12701 17744
rect 12643 17703 12701 17704
rect 13027 17744 13085 17745
rect 13027 17704 13036 17744
rect 13076 17704 13085 17744
rect 13027 17703 13085 17704
rect 13707 17744 13749 17753
rect 14283 17746 14284 17786
rect 14324 17746 14325 17786
rect 14571 17788 14572 17828
rect 14612 17788 14613 17828
rect 14571 17779 14613 17788
rect 19363 17828 19421 17829
rect 19363 17788 19372 17828
rect 19412 17788 19421 17828
rect 19363 17787 19421 17788
rect 19747 17828 19805 17829
rect 19747 17788 19756 17828
rect 19796 17788 19805 17828
rect 19747 17787 19805 17788
rect 14659 17786 14717 17787
rect 13707 17704 13708 17744
rect 13748 17704 13749 17744
rect 13707 17695 13749 17704
rect 13987 17744 14045 17745
rect 13987 17704 13996 17744
rect 14036 17704 14045 17744
rect 14283 17737 14325 17746
rect 14659 17746 14668 17786
rect 14708 17746 14717 17786
rect 14659 17745 14717 17746
rect 14851 17744 14909 17745
rect 13987 17703 14045 17704
rect 14851 17704 14860 17744
rect 14900 17704 14909 17744
rect 14851 17703 14909 17704
rect 16099 17744 16157 17745
rect 16099 17704 16108 17744
rect 16148 17704 16157 17744
rect 16099 17703 16157 17704
rect 16875 17744 16917 17753
rect 16875 17704 16876 17744
rect 16916 17704 16917 17744
rect 16875 17695 16917 17704
rect 17155 17744 17213 17745
rect 17155 17704 17164 17744
rect 17204 17704 17213 17744
rect 17155 17703 17213 17704
rect 17443 17744 17501 17745
rect 17443 17704 17452 17744
rect 17492 17704 17501 17744
rect 17443 17703 17501 17704
rect 17731 17744 17789 17745
rect 17731 17704 17740 17744
rect 17780 17704 17789 17744
rect 17731 17703 17789 17704
rect 18979 17744 19037 17745
rect 18979 17704 18988 17744
rect 19028 17704 19037 17744
rect 18979 17703 19037 17704
rect 5931 17660 5973 17669
rect 5931 17620 5932 17660
rect 5972 17620 5973 17660
rect 5931 17611 5973 17620
rect 7947 17660 7989 17669
rect 7947 17620 7948 17660
rect 7988 17620 7989 17660
rect 7947 17611 7989 17620
rect 8619 17660 8661 17669
rect 8619 17620 8620 17660
rect 8660 17620 8661 17660
rect 8619 17611 8661 17620
rect 12843 17660 12885 17669
rect 12843 17620 12844 17660
rect 12884 17620 12885 17660
rect 12843 17611 12885 17620
rect 13611 17660 13653 17669
rect 13611 17620 13612 17660
rect 13652 17620 13653 17660
rect 13611 17611 13653 17620
rect 16779 17660 16821 17669
rect 16779 17620 16780 17660
rect 16820 17620 16821 17660
rect 16779 17611 16821 17620
rect 9099 17576 9141 17585
rect 9099 17536 9100 17576
rect 9140 17536 9141 17576
rect 9099 17527 9141 17536
rect 11019 17576 11061 17585
rect 11019 17536 11020 17576
rect 11060 17536 11061 17576
rect 11019 17527 11061 17536
rect 19563 17576 19605 17585
rect 19563 17536 19564 17576
rect 19604 17536 19605 17576
rect 19563 17527 19605 17536
rect 1152 17408 20452 17432
rect 1152 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20452 17408
rect 1152 17344 20452 17368
rect 5931 17240 5973 17249
rect 5931 17200 5932 17240
rect 5972 17200 5973 17240
rect 5931 17191 5973 17200
rect 7947 17240 7989 17249
rect 7947 17200 7948 17240
rect 7988 17200 7989 17240
rect 7947 17191 7989 17200
rect 12843 17240 12885 17249
rect 12843 17200 12844 17240
rect 12884 17200 12885 17240
rect 12843 17191 12885 17200
rect 1419 17156 1461 17165
rect 1419 17116 1420 17156
rect 1460 17116 1461 17156
rect 1419 17107 1461 17116
rect 4107 17156 4149 17165
rect 4107 17116 4108 17156
rect 4148 17116 4149 17156
rect 4107 17107 4149 17116
rect 9579 17156 9621 17165
rect 9579 17116 9580 17156
rect 9620 17116 9621 17156
rect 9579 17107 9621 17116
rect 18795 17156 18837 17165
rect 18795 17116 18796 17156
rect 18836 17116 18837 17156
rect 18795 17107 18837 17116
rect 20126 17083 20168 17092
rect 1323 17072 1365 17081
rect 1323 17032 1324 17072
rect 1364 17032 1365 17072
rect 1323 17023 1365 17032
rect 1515 17072 1557 17081
rect 1515 17032 1516 17072
rect 1556 17032 1557 17072
rect 1515 17023 1557 17032
rect 1603 17072 1661 17073
rect 1603 17032 1612 17072
rect 1652 17032 1661 17072
rect 1603 17031 1661 17032
rect 1803 17072 1845 17081
rect 1803 17032 1804 17072
rect 1844 17032 1845 17072
rect 1803 17023 1845 17032
rect 1899 17072 1941 17081
rect 1899 17032 1900 17072
rect 1940 17032 1941 17072
rect 1899 17023 1941 17032
rect 1995 17072 2037 17081
rect 1995 17032 1996 17072
rect 2036 17032 2037 17072
rect 1995 17023 2037 17032
rect 2091 17072 2133 17081
rect 2091 17032 2092 17072
rect 2132 17032 2133 17072
rect 2091 17023 2133 17032
rect 2379 17072 2421 17081
rect 2379 17032 2380 17072
rect 2420 17032 2421 17072
rect 2379 17023 2421 17032
rect 2475 17072 2517 17081
rect 2475 17032 2476 17072
rect 2516 17032 2517 17072
rect 2475 17023 2517 17032
rect 2955 17072 2997 17081
rect 2955 17032 2956 17072
rect 2996 17032 2997 17072
rect 2955 17023 2997 17032
rect 3427 17072 3485 17073
rect 3427 17032 3436 17072
rect 3476 17032 3485 17072
rect 3427 17031 3485 17032
rect 3915 17067 3957 17076
rect 3915 17027 3916 17067
rect 3956 17027 3957 17067
rect 4483 17072 4541 17073
rect 4483 17032 4492 17072
rect 4532 17032 4541 17072
rect 4483 17031 4541 17032
rect 5731 17072 5789 17073
rect 5731 17032 5740 17072
rect 5780 17032 5789 17072
rect 5731 17031 5789 17032
rect 6219 17072 6261 17081
rect 6219 17032 6220 17072
rect 6260 17032 6261 17072
rect 3915 17018 3957 17027
rect 6219 17023 6261 17032
rect 6315 17072 6357 17081
rect 6315 17032 6316 17072
rect 6356 17032 6357 17072
rect 6315 17023 6357 17032
rect 7267 17072 7325 17073
rect 7267 17032 7276 17072
rect 7316 17032 7325 17072
rect 7267 17031 7325 17032
rect 7755 17067 7797 17076
rect 7755 17027 7756 17067
rect 7796 17027 7797 17067
rect 8227 17072 8285 17073
rect 8227 17032 8236 17072
rect 8276 17032 8285 17072
rect 8227 17031 8285 17032
rect 8707 17072 8765 17073
rect 8707 17032 8716 17072
rect 8756 17032 8765 17072
rect 8707 17031 8765 17032
rect 9003 17072 9045 17081
rect 9003 17032 9004 17072
rect 9044 17032 9045 17072
rect 7755 17018 7797 17027
rect 9003 17023 9045 17032
rect 9099 17072 9141 17081
rect 9099 17032 9100 17072
rect 9140 17032 9141 17072
rect 9099 17023 9141 17032
rect 9763 17072 9821 17073
rect 9763 17032 9772 17072
rect 9812 17032 9821 17072
rect 9763 17031 9821 17032
rect 11011 17072 11069 17073
rect 11011 17032 11020 17072
rect 11060 17032 11069 17072
rect 11011 17031 11069 17032
rect 11395 17072 11453 17073
rect 11395 17032 11404 17072
rect 11444 17032 11453 17072
rect 11395 17031 11453 17032
rect 12643 17072 12701 17073
rect 12643 17032 12652 17072
rect 12692 17032 12701 17072
rect 12643 17031 12701 17032
rect 13411 17072 13469 17073
rect 13411 17032 13420 17072
rect 13460 17032 13469 17072
rect 13411 17031 13469 17032
rect 13707 17072 13749 17081
rect 13707 17032 13708 17072
rect 13748 17032 13749 17072
rect 13707 17023 13749 17032
rect 13803 17072 13845 17081
rect 13803 17032 13804 17072
rect 13844 17032 13845 17072
rect 13803 17023 13845 17032
rect 14467 17072 14525 17073
rect 14467 17032 14476 17072
rect 14516 17032 14525 17072
rect 14467 17031 14525 17032
rect 15715 17072 15773 17073
rect 15715 17032 15724 17072
rect 15764 17032 15773 17072
rect 15715 17031 15773 17032
rect 16107 17072 16149 17081
rect 16107 17032 16108 17072
rect 16148 17032 16149 17072
rect 16107 17023 16149 17032
rect 16483 17072 16541 17073
rect 16483 17032 16492 17072
rect 16532 17032 16541 17072
rect 16483 17031 16541 17032
rect 16675 17072 16733 17073
rect 16675 17032 16684 17072
rect 16724 17032 16733 17072
rect 16675 17031 16733 17032
rect 17067 17072 17109 17081
rect 17067 17032 17068 17072
rect 17108 17032 17109 17072
rect 17067 17023 17109 17032
rect 17347 17072 17405 17073
rect 17347 17032 17356 17072
rect 17396 17032 17405 17072
rect 17347 17031 17405 17032
rect 18595 17072 18653 17073
rect 18595 17032 18604 17072
rect 18644 17032 18653 17072
rect 18595 17031 18653 17032
rect 18979 17072 19037 17073
rect 18979 17032 18988 17072
rect 19028 17032 19037 17072
rect 18979 17031 19037 17032
rect 19371 17072 19413 17081
rect 19371 17032 19372 17072
rect 19412 17032 19413 17072
rect 19371 17023 19413 17032
rect 19563 17072 19605 17081
rect 19563 17032 19564 17072
rect 19604 17032 19605 17072
rect 19563 17023 19605 17032
rect 19939 17072 19997 17073
rect 19939 17032 19948 17072
rect 19988 17032 19997 17072
rect 20126 17043 20127 17083
rect 20167 17043 20168 17083
rect 20126 17034 20168 17043
rect 19939 17031 19997 17032
rect 2859 16988 2901 16997
rect 2859 16948 2860 16988
rect 2900 16948 2901 16988
rect 2859 16939 2901 16948
rect 6699 16988 6741 16997
rect 6699 16948 6700 16988
rect 6740 16948 6741 16988
rect 6699 16939 6741 16948
rect 6795 16988 6837 16997
rect 6795 16948 6796 16988
rect 6836 16948 6837 16988
rect 6795 16939 6837 16948
rect 16203 16988 16245 16997
rect 16203 16948 16204 16988
rect 16244 16948 16245 16988
rect 16203 16939 16245 16948
rect 16395 16988 16437 16997
rect 16395 16948 16396 16988
rect 16436 16948 16437 16988
rect 16395 16939 16437 16948
rect 16779 16988 16821 16997
rect 16779 16948 16780 16988
rect 16820 16948 16821 16988
rect 16779 16939 16821 16948
rect 16971 16988 17013 16997
rect 16971 16948 16972 16988
rect 17012 16948 17013 16988
rect 16971 16939 17013 16948
rect 19083 16988 19125 16997
rect 19083 16948 19084 16988
rect 19124 16948 19125 16988
rect 19083 16939 19125 16948
rect 19275 16988 19317 16997
rect 19275 16948 19276 16988
rect 19316 16948 19317 16988
rect 19275 16939 19317 16948
rect 19659 16988 19701 16997
rect 19659 16948 19660 16988
rect 19700 16948 19701 16988
rect 19659 16939 19701 16948
rect 19851 16988 19893 16997
rect 19851 16948 19852 16988
rect 19892 16948 19893 16988
rect 19851 16939 19893 16948
rect 20235 16988 20277 16997
rect 20235 16948 20236 16988
rect 20276 16948 20277 16988
rect 20235 16939 20277 16948
rect 14083 16904 14141 16905
rect 14083 16864 14092 16904
rect 14132 16864 14141 16904
rect 14083 16863 14141 16864
rect 16299 16904 16341 16913
rect 16299 16864 16300 16904
rect 16340 16864 16341 16904
rect 16299 16855 16341 16864
rect 16875 16904 16917 16913
rect 16875 16864 16876 16904
rect 16916 16864 16917 16904
rect 16875 16855 16917 16864
rect 19179 16904 19221 16913
rect 19179 16864 19180 16904
rect 19220 16864 19221 16904
rect 19179 16855 19221 16864
rect 19755 16904 19797 16913
rect 19755 16864 19756 16904
rect 19796 16864 19797 16904
rect 19755 16855 19797 16864
rect 8139 16820 8181 16829
rect 8139 16780 8140 16820
rect 8180 16780 8181 16820
rect 8139 16771 8181 16780
rect 9379 16820 9437 16821
rect 9379 16780 9388 16820
rect 9428 16780 9437 16820
rect 9379 16779 9437 16780
rect 15915 16820 15957 16829
rect 15915 16780 15916 16820
rect 15956 16780 15957 16820
rect 15915 16771 15957 16780
rect 1152 16652 20352 16676
rect 1152 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 20352 16652
rect 1152 16588 20352 16612
rect 19947 16484 19989 16493
rect 19947 16444 19948 16484
rect 19988 16444 19989 16484
rect 19947 16435 19989 16444
rect 8523 16400 8565 16409
rect 8523 16360 8524 16400
rect 8564 16360 8565 16400
rect 8523 16351 8565 16360
rect 18891 16400 18933 16409
rect 18891 16360 18892 16400
rect 18932 16360 18933 16400
rect 18891 16351 18933 16360
rect 2859 16316 2901 16325
rect 2859 16276 2860 16316
rect 2900 16276 2901 16316
rect 2859 16267 2901 16276
rect 9675 16316 9717 16325
rect 9675 16276 9676 16316
rect 9716 16276 9717 16316
rect 9675 16267 9717 16276
rect 15723 16316 15765 16325
rect 15723 16276 15724 16316
rect 15764 16276 15765 16316
rect 15723 16267 15765 16276
rect 15819 16316 15861 16325
rect 15819 16276 15820 16316
rect 15860 16276 15861 16316
rect 15819 16267 15861 16276
rect 20139 16274 20181 16283
rect 10731 16246 10773 16255
rect 1219 16232 1277 16233
rect 1219 16192 1228 16232
rect 1268 16192 1277 16232
rect 1219 16191 1277 16192
rect 1323 16232 1365 16241
rect 1323 16192 1324 16232
rect 1364 16192 1365 16232
rect 1323 16183 1365 16192
rect 1515 16232 1557 16241
rect 1515 16192 1516 16232
rect 1556 16192 1557 16232
rect 1515 16183 1557 16192
rect 1707 16232 1749 16241
rect 1707 16192 1708 16232
rect 1748 16192 1749 16232
rect 1707 16183 1749 16192
rect 1899 16232 1941 16241
rect 1899 16192 1900 16232
rect 1940 16192 1941 16232
rect 1899 16183 1941 16192
rect 1987 16232 2045 16233
rect 1987 16192 1996 16232
rect 2036 16192 2045 16232
rect 1987 16191 2045 16192
rect 2283 16232 2325 16241
rect 2283 16192 2284 16232
rect 2324 16192 2325 16232
rect 2283 16183 2325 16192
rect 2379 16232 2421 16241
rect 2379 16192 2380 16232
rect 2420 16192 2421 16232
rect 2379 16183 2421 16192
rect 2763 16232 2805 16241
rect 3819 16237 3861 16246
rect 2763 16192 2764 16232
rect 2804 16192 2805 16232
rect 2763 16183 2805 16192
rect 3331 16232 3389 16233
rect 3331 16192 3340 16232
rect 3380 16192 3389 16232
rect 3331 16191 3389 16192
rect 3819 16197 3820 16237
rect 3860 16197 3861 16237
rect 3819 16188 3861 16197
rect 4195 16232 4253 16233
rect 4195 16192 4204 16232
rect 4244 16192 4253 16232
rect 4195 16191 4253 16192
rect 4299 16232 4341 16241
rect 4299 16192 4300 16232
rect 4340 16192 4341 16232
rect 4299 16183 4341 16192
rect 4579 16232 4637 16233
rect 4579 16192 4588 16232
rect 4628 16192 4637 16232
rect 4579 16191 4637 16192
rect 5827 16232 5885 16233
rect 5827 16192 5836 16232
rect 5876 16192 5885 16232
rect 5827 16191 5885 16192
rect 6302 16232 6360 16233
rect 6302 16192 6311 16232
rect 6351 16192 6360 16232
rect 6302 16191 6360 16192
rect 6411 16232 6453 16241
rect 6411 16192 6412 16232
rect 6452 16192 6453 16232
rect 6411 16183 6453 16192
rect 6507 16232 6549 16241
rect 6507 16192 6508 16232
rect 6548 16192 6549 16232
rect 6507 16183 6549 16192
rect 6691 16232 6749 16233
rect 6691 16192 6700 16232
rect 6740 16192 6749 16232
rect 6691 16191 6749 16192
rect 6787 16232 6845 16233
rect 6787 16192 6796 16232
rect 6836 16192 6845 16232
rect 6787 16191 6845 16192
rect 7075 16232 7133 16233
rect 7075 16192 7084 16232
rect 7124 16192 7133 16232
rect 7075 16191 7133 16192
rect 8323 16232 8381 16233
rect 8323 16192 8332 16232
rect 8372 16192 8381 16232
rect 8323 16191 8381 16192
rect 8715 16232 8757 16241
rect 8715 16192 8716 16232
rect 8756 16192 8757 16232
rect 8715 16183 8757 16192
rect 8907 16232 8949 16241
rect 8907 16192 8908 16232
rect 8948 16192 8949 16232
rect 8907 16183 8949 16192
rect 9195 16232 9237 16241
rect 9195 16192 9196 16232
rect 9236 16192 9237 16232
rect 9195 16183 9237 16192
rect 9291 16232 9333 16241
rect 9291 16192 9292 16232
rect 9332 16192 9333 16232
rect 9291 16183 9333 16192
rect 9771 16232 9813 16241
rect 9771 16192 9772 16232
rect 9812 16192 9813 16232
rect 9771 16183 9813 16192
rect 10243 16232 10301 16233
rect 10243 16192 10252 16232
rect 10292 16192 10301 16232
rect 10731 16206 10732 16246
rect 10772 16206 10773 16246
rect 10731 16197 10773 16206
rect 11587 16232 11645 16233
rect 10243 16191 10301 16192
rect 11587 16192 11596 16232
rect 11636 16192 11645 16232
rect 11587 16191 11645 16192
rect 12835 16232 12893 16233
rect 12835 16192 12844 16232
rect 12884 16192 12893 16232
rect 12835 16191 12893 16192
rect 13507 16232 13565 16233
rect 13507 16192 13516 16232
rect 13556 16192 13565 16232
rect 13507 16191 13565 16192
rect 14755 16232 14813 16233
rect 14755 16192 14764 16232
rect 14804 16192 14813 16232
rect 14755 16191 14813 16192
rect 15243 16232 15285 16241
rect 15243 16192 15244 16232
rect 15284 16192 15285 16232
rect 15243 16183 15285 16192
rect 15339 16232 15381 16241
rect 16779 16237 16821 16246
rect 15339 16192 15340 16232
rect 15380 16192 15381 16232
rect 15339 16183 15381 16192
rect 16291 16232 16349 16233
rect 16291 16192 16300 16232
rect 16340 16192 16349 16232
rect 16291 16191 16349 16192
rect 16779 16197 16780 16237
rect 16820 16197 16821 16237
rect 16779 16188 16821 16197
rect 17251 16232 17309 16233
rect 17251 16192 17260 16232
rect 17300 16192 17309 16232
rect 17251 16191 17309 16192
rect 17443 16232 17501 16233
rect 17443 16192 17452 16232
rect 17492 16192 17501 16232
rect 17443 16191 17501 16192
rect 18691 16232 18749 16233
rect 18691 16192 18700 16232
rect 18740 16192 18749 16232
rect 18691 16191 18749 16192
rect 19171 16232 19229 16233
rect 19171 16192 19180 16232
rect 19220 16192 19229 16232
rect 19171 16191 19229 16192
rect 19267 16232 19325 16233
rect 19267 16192 19276 16232
rect 19316 16192 19325 16232
rect 19267 16191 19325 16192
rect 19467 16232 19509 16241
rect 19467 16192 19468 16232
rect 19508 16192 19509 16232
rect 19467 16183 19509 16192
rect 19563 16232 19605 16241
rect 19563 16192 19564 16232
rect 19604 16192 19605 16232
rect 19563 16183 19605 16192
rect 19720 16239 19762 16248
rect 19720 16199 19721 16239
rect 19761 16199 19762 16239
rect 20139 16234 20140 16274
rect 20180 16234 20181 16274
rect 19720 16190 19762 16199
rect 19939 16232 19997 16233
rect 19939 16192 19948 16232
rect 19988 16192 19997 16232
rect 20139 16225 20181 16234
rect 20227 16232 20285 16233
rect 19939 16191 19997 16192
rect 20227 16192 20236 16232
rect 20276 16192 20285 16232
rect 20227 16191 20285 16192
rect 10923 16148 10965 16157
rect 10923 16108 10924 16148
rect 10964 16108 10965 16148
rect 10923 16099 10965 16108
rect 1411 16064 1469 16065
rect 1411 16024 1420 16064
rect 1460 16024 1469 16064
rect 1411 16023 1469 16024
rect 1795 16064 1853 16065
rect 1795 16024 1804 16064
rect 1844 16024 1853 16064
rect 1795 16023 1853 16024
rect 4011 16064 4053 16073
rect 4011 16024 4012 16064
rect 4052 16024 4053 16064
rect 4011 16015 4053 16024
rect 6027 16064 6069 16073
rect 6027 16024 6028 16064
rect 6068 16024 6069 16064
rect 6027 16015 6069 16024
rect 6307 16064 6365 16065
rect 6307 16024 6316 16064
rect 6356 16024 6365 16064
rect 6307 16023 6365 16024
rect 8811 16064 8853 16073
rect 8811 16024 8812 16064
rect 8852 16024 8853 16064
rect 8811 16015 8853 16024
rect 13035 16064 13077 16073
rect 13035 16024 13036 16064
rect 13076 16024 13077 16064
rect 13035 16015 13077 16024
rect 14955 16064 14997 16073
rect 14955 16024 14956 16064
rect 14996 16024 14997 16064
rect 14955 16015 14997 16024
rect 16971 16064 17013 16073
rect 16971 16024 16972 16064
rect 17012 16024 17013 16064
rect 16971 16015 17013 16024
rect 17163 16064 17205 16073
rect 17163 16024 17164 16064
rect 17204 16024 17205 16064
rect 17163 16015 17205 16024
rect 19363 16064 19421 16065
rect 19363 16024 19372 16064
rect 19412 16024 19421 16064
rect 19363 16023 19421 16024
rect 1152 15896 20452 15920
rect 1152 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20452 15896
rect 1152 15832 20452 15856
rect 2667 15728 2709 15737
rect 2667 15688 2668 15728
rect 2708 15688 2709 15728
rect 2667 15679 2709 15688
rect 10923 15728 10965 15737
rect 10923 15688 10924 15728
rect 10964 15688 10965 15728
rect 10923 15679 10965 15688
rect 14947 15728 15005 15729
rect 14947 15688 14956 15728
rect 14996 15688 15005 15728
rect 14947 15687 15005 15688
rect 3339 15644 3381 15653
rect 3339 15604 3340 15644
rect 3380 15604 3381 15644
rect 3339 15595 3381 15604
rect 6891 15644 6933 15653
rect 6891 15604 6892 15644
rect 6932 15604 6933 15644
rect 6891 15595 6933 15604
rect 8907 15644 8949 15653
rect 8907 15604 8908 15644
rect 8948 15604 8949 15644
rect 8907 15595 8949 15604
rect 13419 15644 13461 15653
rect 13419 15604 13420 15644
rect 13460 15604 13461 15644
rect 13419 15595 13461 15604
rect 17451 15644 17493 15653
rect 17451 15604 17452 15644
rect 17492 15604 17493 15644
rect 17451 15595 17493 15604
rect 1219 15560 1277 15561
rect 1219 15520 1228 15560
rect 1268 15520 1277 15560
rect 1219 15519 1277 15520
rect 2467 15560 2525 15561
rect 2467 15520 2476 15560
rect 2516 15520 2525 15560
rect 2467 15519 2525 15520
rect 2947 15560 3005 15561
rect 2947 15520 2956 15560
rect 2996 15520 3005 15560
rect 2947 15519 3005 15520
rect 3243 15560 3285 15569
rect 3243 15520 3244 15560
rect 3284 15520 3285 15560
rect 3243 15511 3285 15520
rect 3811 15560 3869 15561
rect 3811 15520 3820 15560
rect 3860 15520 3869 15560
rect 3811 15519 3869 15520
rect 5059 15560 5117 15561
rect 5059 15520 5068 15560
rect 5108 15520 5117 15560
rect 5059 15519 5117 15520
rect 5443 15560 5501 15561
rect 5443 15520 5452 15560
rect 5492 15520 5501 15560
rect 5443 15519 5501 15520
rect 6691 15560 6749 15561
rect 6691 15520 6700 15560
rect 6740 15520 6749 15560
rect 6691 15519 6749 15520
rect 7179 15560 7221 15569
rect 7179 15520 7180 15560
rect 7220 15520 7221 15560
rect 7179 15511 7221 15520
rect 7275 15560 7317 15569
rect 7275 15520 7276 15560
rect 7316 15520 7317 15560
rect 7275 15511 7317 15520
rect 8227 15560 8285 15561
rect 8227 15520 8236 15560
rect 8276 15520 8285 15560
rect 9195 15560 9237 15569
rect 8227 15519 8285 15520
rect 8715 15546 8757 15555
rect 8715 15506 8716 15546
rect 8756 15506 8757 15546
rect 9195 15520 9196 15560
rect 9236 15520 9237 15560
rect 9195 15511 9237 15520
rect 9291 15560 9333 15569
rect 9291 15520 9292 15560
rect 9332 15520 9333 15560
rect 9291 15511 9333 15520
rect 9675 15560 9717 15569
rect 9675 15520 9676 15560
rect 9716 15520 9717 15560
rect 9675 15511 9717 15520
rect 9771 15560 9813 15569
rect 9771 15520 9772 15560
rect 9812 15520 9813 15560
rect 9771 15511 9813 15520
rect 10243 15560 10301 15561
rect 10243 15520 10252 15560
rect 10292 15520 10301 15560
rect 10243 15519 10301 15520
rect 10731 15555 10773 15564
rect 10731 15515 10732 15555
rect 10772 15515 10773 15555
rect 11395 15560 11453 15561
rect 10731 15506 10773 15515
rect 11107 15547 11165 15548
rect 11107 15507 11116 15547
rect 11156 15507 11165 15547
rect 11395 15520 11404 15560
rect 11444 15520 11453 15560
rect 11395 15519 11453 15520
rect 11787 15560 11829 15569
rect 11787 15520 11788 15560
rect 11828 15520 11829 15560
rect 11787 15511 11829 15520
rect 11971 15560 12029 15561
rect 11971 15520 11980 15560
rect 12020 15520 12029 15560
rect 11971 15519 12029 15520
rect 13219 15560 13277 15561
rect 13219 15520 13228 15560
rect 13268 15520 13277 15560
rect 13219 15519 13277 15520
rect 13899 15560 13941 15569
rect 13899 15520 13900 15560
rect 13940 15520 13941 15560
rect 13899 15511 13941 15520
rect 13995 15560 14037 15569
rect 13995 15520 13996 15560
rect 14036 15520 14037 15560
rect 13995 15511 14037 15520
rect 14275 15560 14333 15561
rect 14275 15520 14284 15560
rect 14324 15520 14333 15560
rect 14763 15560 14805 15569
rect 14275 15519 14333 15520
rect 14605 15545 14647 15554
rect 11107 15506 11165 15507
rect 8715 15497 8757 15506
rect 14605 15505 14606 15545
rect 14646 15505 14647 15545
rect 14763 15520 14764 15560
rect 14804 15520 14805 15560
rect 14763 15511 14805 15520
rect 14859 15560 14901 15569
rect 14859 15520 14860 15560
rect 14900 15520 14901 15560
rect 14859 15511 14901 15520
rect 15043 15560 15101 15561
rect 15043 15520 15052 15560
rect 15092 15520 15101 15560
rect 15043 15519 15101 15520
rect 15139 15560 15197 15561
rect 15139 15520 15148 15560
rect 15188 15520 15197 15560
rect 15139 15519 15197 15520
rect 15723 15560 15765 15569
rect 15723 15520 15724 15560
rect 15764 15520 15765 15560
rect 15723 15511 15765 15520
rect 15819 15560 15861 15569
rect 15819 15520 15820 15560
rect 15860 15520 15861 15560
rect 15819 15511 15861 15520
rect 16203 15560 16245 15569
rect 16203 15520 16204 15560
rect 16244 15520 16245 15560
rect 16203 15511 16245 15520
rect 16771 15560 16829 15561
rect 16771 15520 16780 15560
rect 16820 15520 16829 15560
rect 16771 15519 16829 15520
rect 17259 15555 17301 15564
rect 17259 15515 17260 15555
rect 17300 15515 17301 15555
rect 17635 15560 17693 15561
rect 17635 15520 17644 15560
rect 17684 15520 17693 15560
rect 17635 15519 17693 15520
rect 18883 15560 18941 15561
rect 18883 15520 18892 15560
rect 18932 15520 18941 15560
rect 18883 15519 18941 15520
rect 19363 15560 19421 15561
rect 19363 15520 19372 15560
rect 19412 15520 19421 15560
rect 19363 15519 19421 15520
rect 19659 15560 19701 15569
rect 19659 15520 19660 15560
rect 19700 15520 19701 15560
rect 17259 15506 17301 15515
rect 19659 15511 19701 15520
rect 19755 15560 19797 15569
rect 19755 15520 19756 15560
rect 19796 15520 19797 15560
rect 19755 15511 19797 15520
rect 14605 15496 14647 15505
rect 7659 15476 7701 15485
rect 7659 15436 7660 15476
rect 7700 15436 7701 15476
rect 7659 15427 7701 15436
rect 7755 15476 7797 15485
rect 7755 15436 7756 15476
rect 7796 15436 7797 15476
rect 7755 15427 7797 15436
rect 11499 15476 11541 15485
rect 11499 15436 11500 15476
rect 11540 15436 11541 15476
rect 11499 15427 11541 15436
rect 11691 15476 11733 15485
rect 11691 15436 11692 15476
rect 11732 15436 11733 15476
rect 11691 15427 11733 15436
rect 16299 15476 16341 15485
rect 16299 15436 16300 15476
rect 16340 15436 16341 15476
rect 16299 15427 16341 15436
rect 5259 15392 5301 15401
rect 5259 15352 5260 15392
rect 5300 15352 5301 15392
rect 5259 15343 5301 15352
rect 11595 15392 11637 15401
rect 11595 15352 11596 15392
rect 11636 15352 11637 15392
rect 11595 15343 11637 15352
rect 13603 15392 13661 15393
rect 13603 15352 13612 15392
rect 13652 15352 13661 15392
rect 13603 15351 13661 15352
rect 20035 15392 20093 15393
rect 20035 15352 20044 15392
rect 20084 15352 20093 15392
rect 20035 15351 20093 15352
rect 3619 15308 3677 15309
rect 3619 15268 3628 15308
rect 3668 15268 3677 15308
rect 3619 15267 3677 15268
rect 11211 15308 11253 15317
rect 11211 15268 11212 15308
rect 11252 15268 11253 15308
rect 11211 15259 11253 15268
rect 19083 15308 19125 15317
rect 19083 15268 19084 15308
rect 19124 15268 19125 15308
rect 19083 15259 19125 15268
rect 1152 15140 20352 15164
rect 1152 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 20352 15140
rect 1152 15076 20352 15100
rect 3339 14972 3381 14981
rect 3339 14932 3340 14972
rect 3380 14932 3381 14972
rect 3339 14923 3381 14932
rect 3531 14972 3573 14981
rect 3531 14932 3532 14972
rect 3572 14932 3573 14972
rect 3531 14923 3573 14932
rect 9003 14972 9045 14981
rect 9003 14932 9004 14972
rect 9044 14932 9045 14972
rect 9003 14923 9045 14932
rect 13323 14972 13365 14981
rect 13323 14932 13324 14972
rect 13364 14932 13365 14972
rect 13323 14923 13365 14932
rect 14275 14972 14333 14973
rect 14275 14932 14284 14972
rect 14324 14932 14333 14972
rect 14275 14931 14333 14932
rect 16963 14972 17021 14973
rect 16963 14932 16972 14972
rect 17012 14932 17021 14972
rect 16963 14931 17021 14932
rect 18315 14972 18357 14981
rect 18315 14932 18316 14972
rect 18356 14932 18357 14972
rect 18315 14923 18357 14932
rect 19843 14972 19901 14973
rect 19843 14932 19852 14972
rect 19892 14932 19901 14972
rect 19843 14931 19901 14932
rect 20235 14972 20277 14981
rect 20235 14932 20236 14972
rect 20276 14932 20277 14972
rect 20235 14923 20277 14932
rect 1515 14888 1557 14897
rect 1515 14848 1516 14888
rect 1556 14848 1557 14888
rect 1515 14839 1557 14848
rect 5155 14888 5213 14889
rect 5155 14848 5164 14888
rect 5204 14848 5213 14888
rect 5155 14847 5213 14848
rect 6315 14888 6357 14897
rect 6315 14848 6316 14888
rect 6356 14848 6357 14888
rect 6315 14839 6357 14848
rect 6891 14888 6933 14897
rect 6891 14848 6892 14888
rect 6932 14848 6933 14888
rect 6891 14839 6933 14848
rect 10827 14888 10869 14897
rect 10827 14848 10828 14888
rect 10868 14848 10869 14888
rect 10827 14839 10869 14848
rect 14667 14888 14709 14897
rect 14667 14848 14668 14888
rect 14708 14848 14709 14888
rect 14667 14839 14709 14848
rect 1419 14804 1461 14813
rect 1419 14764 1420 14804
rect 1460 14764 1461 14804
rect 1419 14755 1461 14764
rect 1611 14804 1653 14813
rect 1611 14764 1612 14804
rect 1652 14764 1653 14804
rect 1611 14755 1653 14764
rect 6219 14804 6261 14813
rect 6219 14764 6220 14804
rect 6260 14764 6261 14804
rect 6219 14755 6261 14764
rect 6411 14804 6453 14813
rect 6411 14764 6412 14804
rect 6452 14764 6453 14804
rect 6411 14755 6453 14764
rect 10731 14804 10773 14813
rect 10731 14764 10732 14804
rect 10772 14764 10773 14804
rect 10731 14755 10773 14764
rect 10923 14804 10965 14813
rect 10923 14764 10924 14804
rect 10964 14764 10965 14804
rect 10923 14755 10965 14764
rect 14571 14804 14613 14813
rect 14571 14764 14572 14804
rect 14612 14764 14613 14804
rect 14571 14755 14613 14764
rect 14763 14804 14805 14813
rect 14763 14764 14764 14804
rect 14804 14764 14805 14804
rect 14763 14755 14805 14764
rect 18115 14804 18173 14805
rect 18115 14764 18124 14804
rect 18164 14764 18173 14804
rect 18115 14763 18173 14764
rect 17251 14762 17309 14763
rect 1323 14720 1365 14729
rect 1323 14680 1324 14720
rect 1364 14680 1365 14720
rect 1323 14671 1365 14680
rect 1699 14720 1757 14721
rect 1699 14680 1708 14720
rect 1748 14680 1757 14720
rect 1699 14679 1757 14680
rect 1891 14720 1949 14721
rect 1891 14680 1900 14720
rect 1940 14680 1949 14720
rect 1891 14679 1949 14680
rect 3139 14720 3197 14721
rect 3139 14680 3148 14720
rect 3188 14680 3197 14720
rect 3139 14679 3197 14680
rect 3715 14720 3773 14721
rect 3715 14680 3724 14720
rect 3764 14680 3773 14720
rect 3715 14679 3773 14680
rect 4963 14720 5021 14721
rect 4963 14680 4972 14720
rect 5012 14680 5021 14720
rect 4963 14679 5021 14680
rect 5451 14720 5493 14729
rect 5451 14680 5452 14720
rect 5492 14680 5493 14720
rect 5451 14671 5493 14680
rect 5547 14720 5589 14729
rect 5547 14680 5548 14720
rect 5588 14680 5589 14720
rect 5547 14671 5589 14680
rect 5827 14720 5885 14721
rect 5827 14680 5836 14720
rect 5876 14680 5885 14720
rect 5827 14679 5885 14680
rect 6123 14720 6165 14729
rect 6123 14680 6124 14720
rect 6164 14680 6165 14720
rect 6123 14671 6165 14680
rect 6499 14720 6557 14721
rect 6499 14680 6508 14720
rect 6548 14680 6557 14720
rect 6499 14679 6557 14680
rect 6795 14720 6837 14729
rect 6795 14680 6796 14720
rect 6836 14680 6837 14720
rect 6795 14671 6837 14680
rect 6987 14720 7029 14729
rect 6987 14680 6988 14720
rect 7028 14680 7029 14720
rect 6987 14671 7029 14680
rect 7083 14720 7125 14729
rect 7083 14680 7084 14720
rect 7124 14680 7125 14720
rect 7083 14671 7125 14680
rect 7555 14720 7613 14721
rect 7555 14680 7564 14720
rect 7604 14680 7613 14720
rect 7555 14679 7613 14680
rect 8803 14720 8861 14721
rect 8803 14680 8812 14720
rect 8852 14680 8861 14720
rect 8803 14679 8861 14680
rect 9195 14720 9237 14729
rect 9195 14680 9196 14720
rect 9236 14680 9237 14720
rect 9195 14671 9237 14680
rect 9291 14720 9333 14729
rect 9291 14680 9292 14720
rect 9332 14680 9333 14720
rect 9291 14671 9333 14680
rect 9675 14720 9717 14729
rect 9675 14680 9676 14720
rect 9716 14680 9717 14720
rect 9675 14671 9717 14680
rect 9771 14720 9813 14729
rect 9771 14680 9772 14720
rect 9812 14680 9813 14720
rect 9771 14671 9813 14680
rect 9867 14720 9909 14729
rect 9867 14680 9868 14720
rect 9908 14680 9909 14720
rect 9867 14671 9909 14680
rect 9963 14720 10005 14729
rect 9963 14680 9964 14720
rect 10004 14680 10005 14720
rect 9963 14671 10005 14680
rect 10155 14720 10197 14729
rect 10155 14680 10156 14720
rect 10196 14680 10197 14720
rect 10155 14671 10197 14680
rect 10347 14720 10389 14729
rect 10347 14680 10348 14720
rect 10388 14680 10389 14720
rect 10347 14671 10389 14680
rect 10443 14720 10485 14729
rect 10443 14680 10444 14720
rect 10484 14680 10485 14720
rect 10443 14671 10485 14680
rect 10635 14720 10677 14729
rect 10635 14680 10636 14720
rect 10676 14680 10677 14720
rect 10635 14671 10677 14680
rect 11011 14720 11069 14721
rect 11011 14680 11020 14720
rect 11060 14680 11069 14720
rect 11011 14679 11069 14680
rect 11211 14720 11253 14729
rect 11211 14680 11212 14720
rect 11252 14680 11253 14720
rect 11211 14671 11253 14680
rect 11403 14720 11445 14729
rect 11403 14680 11404 14720
rect 11444 14680 11445 14720
rect 11403 14671 11445 14680
rect 11587 14720 11645 14721
rect 11587 14680 11596 14720
rect 11636 14680 11645 14720
rect 11587 14679 11645 14680
rect 12835 14720 12893 14721
rect 12835 14680 12844 14720
rect 12884 14680 12893 14720
rect 12835 14679 12893 14680
rect 13219 14720 13277 14721
rect 13219 14680 13228 14720
rect 13268 14680 13277 14720
rect 13219 14679 13277 14680
rect 13603 14720 13661 14721
rect 13603 14680 13612 14720
rect 13652 14680 13661 14720
rect 13603 14679 13661 14680
rect 13899 14720 13941 14729
rect 13899 14680 13900 14720
rect 13940 14680 13941 14720
rect 13899 14671 13941 14680
rect 14467 14720 14525 14721
rect 14467 14680 14476 14720
rect 14516 14680 14525 14720
rect 14467 14679 14525 14680
rect 14859 14720 14901 14729
rect 17251 14722 17260 14762
rect 17300 14722 17309 14762
rect 17251 14721 17309 14722
rect 14859 14680 14860 14720
rect 14900 14680 14901 14720
rect 14859 14671 14901 14680
rect 15331 14720 15389 14721
rect 15331 14680 15340 14720
rect 15380 14680 15389 14720
rect 15331 14679 15389 14680
rect 16579 14720 16637 14721
rect 16579 14680 16588 14720
rect 16628 14680 16637 14720
rect 16579 14679 16637 14680
rect 17355 14720 17397 14729
rect 17355 14680 17356 14720
rect 17396 14680 17397 14720
rect 17355 14671 17397 14680
rect 17635 14720 17693 14721
rect 17635 14680 17644 14720
rect 17684 14680 17693 14720
rect 17635 14679 17693 14680
rect 18499 14720 18557 14721
rect 18499 14680 18508 14720
rect 18548 14680 18557 14720
rect 18499 14679 18557 14680
rect 18603 14720 18645 14729
rect 18603 14680 18604 14720
rect 18644 14680 18645 14720
rect 18603 14671 18645 14680
rect 18787 14720 18845 14721
rect 18787 14680 18796 14720
rect 18836 14680 18845 14720
rect 18787 14679 18845 14680
rect 19171 14720 19229 14721
rect 19171 14680 19180 14720
rect 19220 14680 19229 14720
rect 19171 14679 19229 14680
rect 19467 14720 19509 14729
rect 19467 14680 19468 14720
rect 19508 14680 19509 14720
rect 19467 14671 19509 14680
rect 20043 14720 20085 14729
rect 20043 14680 20044 14720
rect 20084 14680 20085 14720
rect 20043 14671 20085 14680
rect 20235 14720 20277 14729
rect 20235 14680 20236 14720
rect 20276 14680 20277 14720
rect 20235 14671 20277 14680
rect 11307 14636 11349 14645
rect 11307 14596 11308 14636
rect 11348 14596 11349 14636
rect 11307 14587 11349 14596
rect 13995 14636 14037 14645
rect 13995 14596 13996 14636
rect 14036 14596 14037 14636
rect 13995 14587 14037 14596
rect 16779 14636 16821 14645
rect 16779 14596 16780 14636
rect 16820 14596 16821 14636
rect 16779 14587 16821 14596
rect 19563 14636 19605 14645
rect 19563 14596 19564 14636
rect 19604 14596 19605 14636
rect 19563 14587 19605 14596
rect 3531 14552 3573 14561
rect 3531 14512 3532 14552
rect 3572 14512 3573 14552
rect 3531 14503 3573 14512
rect 9475 14552 9533 14553
rect 9475 14512 9484 14552
rect 9524 14512 9533 14552
rect 9475 14511 9533 14512
rect 10251 14552 10293 14561
rect 10251 14512 10252 14552
rect 10292 14512 10293 14552
rect 10251 14503 10293 14512
rect 13035 14552 13077 14561
rect 13035 14512 13036 14552
rect 13076 14512 13077 14552
rect 13035 14503 13077 14512
rect 18795 14552 18837 14561
rect 18795 14512 18796 14552
rect 18836 14512 18837 14552
rect 18795 14503 18837 14512
rect 1152 14384 20452 14408
rect 1152 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20452 14384
rect 1152 14320 20452 14344
rect 2667 14216 2709 14225
rect 2667 14176 2668 14216
rect 2708 14176 2709 14216
rect 2667 14167 2709 14176
rect 4299 14216 4341 14225
rect 4299 14176 4300 14216
rect 4340 14176 4341 14216
rect 4299 14167 4341 14176
rect 12267 14216 12309 14225
rect 12267 14176 12268 14216
rect 12308 14176 12309 14216
rect 12267 14167 12309 14176
rect 12843 14216 12885 14225
rect 12843 14176 12844 14216
rect 12884 14176 12885 14216
rect 12843 14167 12885 14176
rect 16203 14216 16245 14225
rect 16203 14176 16204 14216
rect 16244 14176 16245 14216
rect 16203 14167 16245 14176
rect 16587 14216 16629 14225
rect 16587 14176 16588 14216
rect 16628 14176 16629 14216
rect 16587 14167 16629 14176
rect 17067 14216 17109 14225
rect 17067 14176 17068 14216
rect 17108 14176 17109 14216
rect 17067 14167 17109 14176
rect 20235 14216 20277 14225
rect 20235 14176 20236 14216
rect 20276 14176 20277 14216
rect 20235 14167 20277 14176
rect 4779 14132 4821 14141
rect 4779 14092 4780 14132
rect 4820 14092 4821 14132
rect 4779 14083 4821 14092
rect 8907 14132 8949 14141
rect 8907 14092 8908 14132
rect 8948 14092 8949 14132
rect 8907 14083 8949 14092
rect 11787 14132 11829 14141
rect 11787 14092 11788 14132
rect 11828 14092 11829 14132
rect 11787 14083 11829 14092
rect 14475 14132 14517 14141
rect 14475 14092 14476 14132
rect 14516 14092 14517 14132
rect 14475 14083 14517 14092
rect 14955 14132 14997 14141
rect 14955 14092 14956 14132
rect 14996 14092 14997 14132
rect 14955 14083 14997 14092
rect 1219 14048 1277 14049
rect 1219 14008 1228 14048
rect 1268 14008 1277 14048
rect 1219 14007 1277 14008
rect 2467 14048 2525 14049
rect 2467 14008 2476 14048
rect 2516 14008 2525 14048
rect 2467 14007 2525 14008
rect 2851 14048 2909 14049
rect 2851 14008 2860 14048
rect 2900 14008 2909 14048
rect 2851 14007 2909 14008
rect 4099 14048 4157 14049
rect 4099 14008 4108 14048
rect 4148 14008 4157 14048
rect 4099 14007 4157 14008
rect 4875 14048 4917 14057
rect 4875 14008 4876 14048
rect 4916 14008 4917 14048
rect 4875 13999 4917 14008
rect 5155 14048 5213 14049
rect 5155 14008 5164 14048
rect 5204 14008 5213 14048
rect 5155 14007 5213 14008
rect 5539 14048 5597 14049
rect 5539 14008 5548 14048
rect 5588 14008 5597 14048
rect 5539 14007 5597 14008
rect 5923 14048 5981 14049
rect 5923 14008 5932 14048
rect 5972 14008 5981 14048
rect 5923 14007 5981 14008
rect 7171 14048 7229 14049
rect 7171 14008 7180 14048
rect 7220 14008 7229 14048
rect 7171 14007 7229 14008
rect 7459 14048 7517 14049
rect 7459 14008 7468 14048
rect 7508 14008 7517 14048
rect 7459 14007 7517 14008
rect 8707 14048 8765 14049
rect 8707 14008 8716 14048
rect 8756 14008 8765 14048
rect 8707 14007 8765 14008
rect 10339 14048 10397 14049
rect 10339 14008 10348 14048
rect 10388 14008 10397 14048
rect 10339 14007 10397 14008
rect 10819 14048 10877 14049
rect 10819 14008 10828 14048
rect 10868 14008 10877 14048
rect 10819 14007 10877 14008
rect 11115 14048 11157 14057
rect 11115 14008 11116 14048
rect 11156 14008 11157 14048
rect 9091 14006 9149 14007
rect 9091 13966 9100 14006
rect 9140 13966 9149 14006
rect 11115 13999 11157 14008
rect 11211 14048 11253 14057
rect 11211 14008 11212 14048
rect 11252 14008 11253 14048
rect 11211 13999 11253 14008
rect 11691 14048 11733 14057
rect 11691 14008 11692 14048
rect 11732 14008 11733 14048
rect 11691 13999 11733 14008
rect 11883 14048 11925 14057
rect 11883 14008 11884 14048
rect 11924 14008 11925 14048
rect 11883 13999 11925 14008
rect 11971 14048 12029 14049
rect 11971 14008 11980 14048
rect 12020 14008 12029 14048
rect 11971 14007 12029 14008
rect 12171 14048 12213 14057
rect 12171 14008 12172 14048
rect 12212 14008 12213 14048
rect 12171 13999 12213 14008
rect 12363 14048 12405 14057
rect 12363 14008 12364 14048
rect 12404 14008 12405 14048
rect 12363 13999 12405 14008
rect 12547 14048 12605 14049
rect 12547 14008 12556 14048
rect 12596 14008 12605 14048
rect 12547 14007 12605 14008
rect 12651 14048 12693 14057
rect 12651 14008 12652 14048
rect 12692 14008 12693 14048
rect 12651 13999 12693 14008
rect 12835 14048 12893 14049
rect 12835 14008 12844 14048
rect 12884 14008 12893 14048
rect 12835 14007 12893 14008
rect 13027 14048 13085 14049
rect 13027 14008 13036 14048
rect 13076 14008 13085 14048
rect 13027 14007 13085 14008
rect 14275 14048 14333 14049
rect 14275 14008 14284 14048
rect 14324 14008 14333 14048
rect 14275 14007 14333 14008
rect 14667 14048 14709 14057
rect 14667 14008 14668 14048
rect 14708 14008 14709 14048
rect 14667 13999 14709 14008
rect 14763 14048 14805 14057
rect 14763 14008 14764 14048
rect 14804 14008 14805 14048
rect 14763 13999 14805 14008
rect 14859 14048 14901 14057
rect 14859 14008 14860 14048
rect 14900 14008 14901 14048
rect 14859 13999 14901 14008
rect 15147 14048 15189 14057
rect 15147 14008 15148 14048
rect 15188 14008 15189 14048
rect 15147 13999 15189 14008
rect 15339 14048 15381 14057
rect 15339 14008 15340 14048
rect 15380 14008 15381 14048
rect 15339 13999 15381 14008
rect 15427 14048 15485 14049
rect 15427 14008 15436 14048
rect 15476 14008 15485 14048
rect 15427 14007 15485 14008
rect 15627 14048 15669 14057
rect 15627 14008 15628 14048
rect 15668 14008 15669 14048
rect 15627 13999 15669 14008
rect 15723 14048 15765 14057
rect 15723 14008 15724 14048
rect 15764 14008 15765 14048
rect 15723 13999 15765 14008
rect 15819 14048 15861 14057
rect 15819 14008 15820 14048
rect 15860 14008 15861 14048
rect 15819 13999 15861 14008
rect 15915 14048 15957 14057
rect 15915 14008 15916 14048
rect 15956 14008 15957 14048
rect 15915 13999 15957 14008
rect 16107 14048 16149 14057
rect 16107 14008 16108 14048
rect 16148 14008 16149 14048
rect 16107 13999 16149 14008
rect 16299 14048 16341 14057
rect 16299 14008 16300 14048
rect 16340 14008 16341 14048
rect 16299 13999 16341 14008
rect 16491 14048 16533 14057
rect 16491 14008 16492 14048
rect 16532 14008 16533 14048
rect 16491 13999 16533 14008
rect 16683 14048 16725 14057
rect 16683 14008 16684 14048
rect 16724 14008 16725 14048
rect 16683 13999 16725 14008
rect 17251 14048 17309 14049
rect 17251 14008 17260 14048
rect 17300 14008 17309 14048
rect 17251 14007 17309 14008
rect 18499 14048 18557 14049
rect 18499 14008 18508 14048
rect 18548 14008 18557 14048
rect 18499 14007 18557 14008
rect 18883 14048 18941 14049
rect 18883 14008 18892 14048
rect 18932 14008 18941 14048
rect 18883 14007 18941 14008
rect 19275 14048 19317 14057
rect 19275 14008 19276 14048
rect 19316 14008 19317 14048
rect 19275 13999 19317 14008
rect 19459 14048 19517 14049
rect 19459 14008 19468 14048
rect 19508 14008 19517 14048
rect 19459 14007 19517 14008
rect 19851 14048 19893 14057
rect 19851 14008 19852 14048
rect 19892 14008 19893 14048
rect 19851 13999 19893 14008
rect 9091 13965 9149 13966
rect 16867 13964 16925 13965
rect 16867 13924 16876 13964
rect 16916 13924 16925 13964
rect 16867 13923 16925 13924
rect 18987 13964 19029 13973
rect 18987 13924 18988 13964
rect 19028 13924 19029 13964
rect 18987 13915 19029 13924
rect 19179 13964 19221 13973
rect 19179 13924 19180 13964
rect 19220 13924 19221 13964
rect 19179 13915 19221 13924
rect 19563 13964 19605 13973
rect 19563 13924 19564 13964
rect 19604 13924 19605 13964
rect 19563 13915 19605 13924
rect 19755 13964 19797 13973
rect 19755 13924 19756 13964
rect 19796 13924 19797 13964
rect 19755 13915 19797 13924
rect 20035 13964 20093 13965
rect 20035 13924 20044 13964
rect 20084 13924 20093 13964
rect 20035 13923 20093 13924
rect 4483 13880 4541 13881
rect 4483 13840 4492 13880
rect 4532 13840 4541 13880
rect 4483 13839 4541 13840
rect 10539 13880 10581 13889
rect 10539 13840 10540 13880
rect 10580 13840 10581 13880
rect 10539 13831 10581 13840
rect 11491 13880 11549 13881
rect 11491 13840 11500 13880
rect 11540 13840 11549 13880
rect 11491 13839 11549 13840
rect 18699 13880 18741 13889
rect 18699 13840 18700 13880
rect 18740 13840 18741 13880
rect 18699 13831 18741 13840
rect 19083 13880 19125 13889
rect 19083 13840 19084 13880
rect 19124 13840 19125 13880
rect 19083 13831 19125 13840
rect 19659 13880 19701 13889
rect 19659 13840 19660 13880
rect 19700 13840 19701 13880
rect 19659 13831 19701 13840
rect 4299 13796 4341 13805
rect 4299 13756 4300 13796
rect 4340 13756 4341 13796
rect 4299 13747 4341 13756
rect 5451 13796 5493 13805
rect 5451 13756 5452 13796
rect 5492 13756 5493 13796
rect 5451 13747 5493 13756
rect 5739 13796 5781 13805
rect 5739 13756 5740 13796
rect 5780 13756 5781 13796
rect 5739 13747 5781 13756
rect 15147 13796 15189 13805
rect 15147 13756 15148 13796
rect 15188 13756 15189 13796
rect 15147 13747 15189 13756
rect 1152 13628 20352 13652
rect 1152 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 20352 13628
rect 1152 13564 20352 13588
rect 2667 13460 2709 13469
rect 2667 13420 2668 13460
rect 2708 13420 2709 13460
rect 2667 13411 2709 13420
rect 9963 13460 10005 13469
rect 9963 13420 9964 13460
rect 10004 13420 10005 13460
rect 9963 13411 10005 13420
rect 10827 13460 10869 13469
rect 10827 13420 10828 13460
rect 10868 13420 10869 13460
rect 10827 13411 10869 13420
rect 16875 13460 16917 13469
rect 16875 13420 16876 13460
rect 16916 13420 16917 13460
rect 16875 13411 16917 13420
rect 18507 13460 18549 13469
rect 18507 13420 18508 13460
rect 18548 13420 18549 13460
rect 18507 13411 18549 13420
rect 19459 13460 19517 13461
rect 19459 13420 19468 13460
rect 19508 13420 19517 13460
rect 19459 13419 19517 13420
rect 19659 13460 19701 13469
rect 19659 13420 19660 13460
rect 19700 13420 19701 13460
rect 19659 13411 19701 13420
rect 7179 13292 7221 13301
rect 7179 13252 7180 13292
rect 7220 13252 7221 13292
rect 7179 13243 7221 13252
rect 10443 13292 10485 13301
rect 10443 13252 10444 13292
rect 10484 13252 10485 13292
rect 9763 13250 9821 13251
rect 8187 13217 8229 13226
rect 1219 13208 1277 13209
rect 1219 13168 1228 13208
rect 1268 13168 1277 13208
rect 1219 13167 1277 13168
rect 2467 13208 2525 13209
rect 2467 13168 2476 13208
rect 2516 13168 2525 13208
rect 2467 13167 2525 13168
rect 3043 13208 3101 13209
rect 3043 13168 3052 13208
rect 3092 13168 3101 13208
rect 3043 13167 3101 13168
rect 4291 13208 4349 13209
rect 4291 13168 4300 13208
rect 4340 13168 4349 13208
rect 4291 13167 4349 13168
rect 4867 13208 4925 13209
rect 4867 13168 4876 13208
rect 4916 13168 4925 13208
rect 4867 13167 4925 13168
rect 6115 13208 6173 13209
rect 6115 13168 6124 13208
rect 6164 13168 6173 13208
rect 6115 13167 6173 13168
rect 6603 13208 6645 13217
rect 6603 13168 6604 13208
rect 6644 13168 6645 13208
rect 6603 13159 6645 13168
rect 6699 13208 6741 13217
rect 6699 13168 6700 13208
rect 6740 13168 6741 13208
rect 6699 13159 6741 13168
rect 7083 13208 7125 13217
rect 7083 13168 7084 13208
rect 7124 13168 7125 13208
rect 7083 13159 7125 13168
rect 7651 13208 7709 13209
rect 7651 13168 7660 13208
rect 7700 13168 7709 13208
rect 8187 13177 8188 13217
rect 8228 13177 8229 13217
rect 9763 13210 9772 13250
rect 9812 13210 9821 13250
rect 10443 13243 10485 13252
rect 13611 13292 13653 13301
rect 13611 13252 13612 13292
rect 13652 13252 13653 13292
rect 13611 13243 13653 13252
rect 13707 13292 13749 13301
rect 13707 13252 13708 13292
rect 13748 13252 13749 13292
rect 13707 13243 13749 13252
rect 14715 13217 14757 13226
rect 9763 13209 9821 13210
rect 8187 13168 8229 13177
rect 8515 13208 8573 13209
rect 8515 13168 8524 13208
rect 8564 13168 8573 13208
rect 7651 13167 7709 13168
rect 8515 13167 8573 13168
rect 10347 13208 10389 13217
rect 10347 13168 10348 13208
rect 10388 13168 10389 13208
rect 10347 13159 10389 13168
rect 10635 13208 10677 13217
rect 10635 13168 10636 13208
rect 10676 13168 10677 13208
rect 10635 13159 10677 13168
rect 11115 13208 11157 13217
rect 11115 13168 11116 13208
rect 11156 13168 11157 13208
rect 11115 13159 11157 13168
rect 11203 13208 11261 13209
rect 11203 13168 11212 13208
rect 11252 13168 11261 13208
rect 11203 13167 11261 13168
rect 11499 13208 11541 13217
rect 11499 13168 11500 13208
rect 11540 13168 11541 13208
rect 11499 13159 11541 13168
rect 11691 13208 11733 13217
rect 11691 13168 11692 13208
rect 11732 13168 11733 13208
rect 11691 13159 11733 13168
rect 11779 13208 11837 13209
rect 11779 13168 11788 13208
rect 11828 13168 11837 13208
rect 11779 13167 11837 13168
rect 12075 13208 12117 13217
rect 12075 13168 12076 13208
rect 12116 13168 12117 13208
rect 12075 13159 12117 13168
rect 12171 13208 12213 13217
rect 12171 13168 12172 13208
rect 12212 13168 12213 13208
rect 12171 13159 12213 13168
rect 12267 13208 12309 13217
rect 12267 13168 12268 13208
rect 12308 13168 12309 13208
rect 12267 13159 12309 13168
rect 12555 13208 12597 13217
rect 12555 13168 12556 13208
rect 12596 13168 12597 13208
rect 12555 13159 12597 13168
rect 12843 13208 12885 13217
rect 12843 13168 12844 13208
rect 12884 13168 12885 13208
rect 12843 13159 12885 13168
rect 13131 13208 13173 13217
rect 13131 13168 13132 13208
rect 13172 13168 13173 13208
rect 13131 13159 13173 13168
rect 13227 13208 13269 13217
rect 13227 13168 13228 13208
rect 13268 13168 13269 13208
rect 13227 13159 13269 13168
rect 14179 13208 14237 13209
rect 14179 13168 14188 13208
rect 14228 13168 14237 13208
rect 14715 13177 14716 13217
rect 14756 13177 14757 13217
rect 14715 13168 14757 13177
rect 15051 13208 15093 13217
rect 15051 13168 15052 13208
rect 15092 13168 15093 13208
rect 14179 13167 14237 13168
rect 15051 13159 15093 13168
rect 15243 13208 15285 13217
rect 15243 13168 15244 13208
rect 15284 13168 15285 13208
rect 15243 13159 15285 13168
rect 15427 13208 15485 13209
rect 15427 13168 15436 13208
rect 15476 13168 15485 13208
rect 15427 13167 15485 13168
rect 16675 13208 16733 13209
rect 16675 13168 16684 13208
rect 16724 13168 16733 13208
rect 16675 13167 16733 13168
rect 17059 13208 17117 13209
rect 17059 13168 17068 13208
rect 17108 13168 17117 13208
rect 17059 13167 17117 13168
rect 18307 13208 18365 13209
rect 18307 13168 18316 13208
rect 18356 13168 18365 13208
rect 18307 13167 18365 13168
rect 18787 13208 18845 13209
rect 18787 13168 18796 13208
rect 18836 13168 18845 13208
rect 18787 13167 18845 13168
rect 19083 13208 19125 13217
rect 19083 13168 19084 13208
rect 19124 13168 19125 13208
rect 19083 13159 19125 13168
rect 19179 13208 19221 13217
rect 19179 13168 19180 13208
rect 19220 13168 19221 13208
rect 19179 13159 19221 13168
rect 19651 13208 19709 13209
rect 19651 13168 19660 13208
rect 19700 13168 19709 13208
rect 19651 13167 19709 13168
rect 19747 13208 19805 13209
rect 19747 13168 19756 13208
rect 19796 13168 19805 13208
rect 19747 13167 19805 13168
rect 19947 13208 19989 13217
rect 19947 13168 19948 13208
rect 19988 13168 19989 13208
rect 19947 13159 19989 13168
rect 20043 13208 20085 13217
rect 20043 13168 20044 13208
rect 20084 13168 20085 13208
rect 20043 13159 20085 13168
rect 20136 13208 20194 13209
rect 20136 13168 20145 13208
rect 20185 13168 20194 13208
rect 20136 13167 20194 13168
rect 8331 13124 8373 13133
rect 8331 13084 8332 13124
rect 8372 13084 8373 13124
rect 8331 13075 8373 13084
rect 12747 13124 12789 13133
rect 12747 13084 12748 13124
rect 12788 13084 12789 13124
rect 12747 13075 12789 13084
rect 2859 13040 2901 13049
rect 2859 13000 2860 13040
rect 2900 13000 2901 13040
rect 2859 12991 2901 13000
rect 4483 13040 4541 13041
rect 4483 13000 4492 13040
rect 4532 13000 4541 13040
rect 4483 12999 4541 13000
rect 6315 13040 6357 13049
rect 6315 13000 6316 13040
rect 6356 13000 6357 13040
rect 6315 12991 6357 13000
rect 9963 13040 10005 13049
rect 9963 13000 9964 13040
rect 10004 13000 10005 13040
rect 9963 12991 10005 13000
rect 11587 13040 11645 13041
rect 11587 13000 11596 13040
rect 11636 13000 11645 13040
rect 11587 12999 11645 13000
rect 12355 13040 12413 13041
rect 12355 13000 12364 13040
rect 12404 13000 12413 13040
rect 12355 12999 12413 13000
rect 14859 13040 14901 13049
rect 14859 13000 14860 13040
rect 14900 13000 14901 13040
rect 14859 12991 14901 13000
rect 15147 13040 15189 13049
rect 15147 13000 15148 13040
rect 15188 13000 15189 13040
rect 15147 12991 15189 13000
rect 11307 12982 11349 12991
rect 11307 12942 11308 12982
rect 11348 12942 11349 12982
rect 11307 12933 11349 12942
rect 1152 12872 20452 12896
rect 1152 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20452 12872
rect 1152 12808 20452 12832
rect 2667 12704 2709 12713
rect 2667 12664 2668 12704
rect 2708 12664 2709 12704
rect 2667 12655 2709 12664
rect 5835 12704 5877 12713
rect 5835 12664 5836 12704
rect 5876 12664 5877 12704
rect 5835 12655 5877 12664
rect 9771 12704 9813 12713
rect 9771 12664 9772 12704
rect 9812 12664 9813 12704
rect 9771 12655 9813 12664
rect 10627 12704 10685 12705
rect 10627 12664 10636 12704
rect 10676 12664 10685 12704
rect 10627 12663 10685 12664
rect 18699 12704 18741 12713
rect 18699 12664 18700 12704
rect 18740 12664 18741 12704
rect 18699 12655 18741 12664
rect 5643 12620 5685 12629
rect 5643 12580 5644 12620
rect 5684 12580 5685 12620
rect 5643 12571 5685 12580
rect 13611 12620 13653 12629
rect 13611 12580 13612 12620
rect 13652 12580 13653 12620
rect 13611 12571 13653 12580
rect 13899 12620 13941 12629
rect 13899 12580 13900 12620
rect 13940 12580 13941 12620
rect 13899 12571 13941 12580
rect 15723 12620 15765 12629
rect 15723 12580 15724 12620
rect 15764 12580 15765 12620
rect 15723 12571 15765 12580
rect 1219 12536 1277 12537
rect 1219 12496 1228 12536
rect 1268 12496 1277 12536
rect 1219 12495 1277 12496
rect 2467 12536 2525 12537
rect 2467 12496 2476 12536
rect 2516 12496 2525 12536
rect 2467 12495 2525 12496
rect 2947 12536 3005 12537
rect 2947 12496 2956 12536
rect 2996 12496 3005 12536
rect 2947 12495 3005 12496
rect 3531 12536 3573 12545
rect 3531 12496 3532 12536
rect 3572 12496 3573 12536
rect 3531 12487 3573 12496
rect 3627 12536 3669 12545
rect 3627 12496 3628 12536
rect 3668 12496 3669 12536
rect 3627 12487 3669 12496
rect 3907 12536 3965 12537
rect 3907 12496 3916 12536
rect 3956 12496 3965 12536
rect 3907 12495 3965 12496
rect 4195 12536 4253 12537
rect 4195 12496 4204 12536
rect 4244 12496 4253 12536
rect 4195 12495 4253 12496
rect 5443 12536 5501 12537
rect 5443 12496 5452 12536
rect 5492 12496 5501 12536
rect 6499 12536 6557 12537
rect 5443 12495 5501 12496
rect 5979 12526 6021 12535
rect 5979 12486 5980 12526
rect 6020 12486 6021 12526
rect 6499 12496 6508 12536
rect 6548 12496 6557 12536
rect 6499 12495 6557 12496
rect 6987 12536 7029 12545
rect 6987 12496 6988 12536
rect 7028 12496 7029 12536
rect 6987 12487 7029 12496
rect 7467 12536 7509 12545
rect 7467 12496 7468 12536
rect 7508 12496 7509 12536
rect 7467 12487 7509 12496
rect 7563 12536 7605 12545
rect 7563 12496 7564 12536
rect 7604 12496 7605 12536
rect 7563 12487 7605 12496
rect 7851 12536 7893 12545
rect 7851 12496 7852 12536
rect 7892 12496 7893 12536
rect 7851 12487 7893 12496
rect 8043 12536 8085 12545
rect 8043 12496 8044 12536
rect 8084 12496 8085 12536
rect 8043 12487 8085 12496
rect 8131 12536 8189 12537
rect 8131 12496 8140 12536
rect 8180 12496 8189 12536
rect 8131 12495 8189 12496
rect 8323 12536 8381 12537
rect 8323 12496 8332 12536
rect 8372 12496 8381 12536
rect 8323 12495 8381 12496
rect 9571 12536 9629 12537
rect 9571 12496 9580 12536
rect 9620 12496 9629 12536
rect 9571 12495 9629 12496
rect 9963 12536 10005 12545
rect 9963 12496 9964 12536
rect 10004 12496 10005 12536
rect 9963 12487 10005 12496
rect 10155 12536 10197 12545
rect 10155 12496 10156 12536
rect 10196 12496 10197 12536
rect 10155 12487 10197 12496
rect 10243 12536 10301 12537
rect 10243 12496 10252 12536
rect 10292 12496 10301 12536
rect 10243 12495 10301 12496
rect 10731 12536 10773 12545
rect 10731 12496 10732 12536
rect 10772 12496 10773 12536
rect 10731 12487 10773 12496
rect 10827 12536 10869 12545
rect 10827 12496 10828 12536
rect 10868 12496 10869 12536
rect 10827 12487 10869 12496
rect 10923 12536 10965 12545
rect 10923 12496 10924 12536
rect 10964 12496 10965 12536
rect 11307 12536 11349 12545
rect 10923 12487 10965 12496
rect 11211 12491 11253 12500
rect 5979 12477 6021 12486
rect 7083 12452 7125 12461
rect 7083 12412 7084 12452
rect 7124 12412 7125 12452
rect 11211 12451 11212 12491
rect 11252 12451 11253 12491
rect 11307 12496 11308 12536
rect 11348 12496 11349 12536
rect 11307 12487 11349 12496
rect 11403 12536 11445 12545
rect 11403 12496 11404 12536
rect 11444 12496 11445 12536
rect 11403 12487 11445 12496
rect 11499 12536 11541 12545
rect 11499 12496 11500 12536
rect 11540 12496 11541 12536
rect 11499 12487 11541 12496
rect 11691 12536 11733 12545
rect 11691 12496 11692 12536
rect 11732 12496 11733 12536
rect 11691 12487 11733 12496
rect 11883 12536 11925 12545
rect 11883 12496 11884 12536
rect 11924 12496 11925 12536
rect 11883 12487 11925 12496
rect 11971 12536 12029 12537
rect 11971 12496 11980 12536
rect 12020 12496 12029 12536
rect 11971 12495 12029 12496
rect 12163 12536 12221 12537
rect 12163 12496 12172 12536
rect 12212 12496 12221 12536
rect 12163 12495 12221 12496
rect 13411 12536 13469 12537
rect 13411 12496 13420 12536
rect 13460 12496 13469 12536
rect 13411 12495 13469 12496
rect 13803 12536 13845 12545
rect 13803 12496 13804 12536
rect 13844 12496 13845 12536
rect 13803 12487 13845 12496
rect 13995 12536 14037 12545
rect 13995 12496 13996 12536
rect 14036 12496 14037 12536
rect 13995 12487 14037 12496
rect 14083 12536 14141 12537
rect 14083 12496 14092 12536
rect 14132 12496 14141 12536
rect 14083 12495 14141 12496
rect 14275 12536 14333 12537
rect 14275 12496 14284 12536
rect 14324 12496 14333 12536
rect 14275 12495 14333 12496
rect 15523 12536 15581 12537
rect 15523 12496 15532 12536
rect 15572 12496 15581 12536
rect 15523 12495 15581 12496
rect 15915 12536 15957 12545
rect 15915 12496 15916 12536
rect 15956 12496 15957 12536
rect 15915 12487 15957 12496
rect 16107 12536 16149 12545
rect 16107 12496 16108 12536
rect 16148 12496 16149 12536
rect 16107 12487 16149 12496
rect 16291 12536 16349 12537
rect 16291 12496 16300 12536
rect 16340 12496 16349 12536
rect 16291 12495 16349 12496
rect 16683 12536 16725 12545
rect 16683 12496 16684 12536
rect 16724 12496 16725 12536
rect 16683 12487 16725 12496
rect 17251 12536 17309 12537
rect 17251 12496 17260 12536
rect 17300 12496 17309 12536
rect 17251 12495 17309 12496
rect 18499 12536 18557 12537
rect 18499 12496 18508 12536
rect 18548 12496 18557 12536
rect 18499 12495 18557 12496
rect 19171 12536 19229 12537
rect 19171 12496 19180 12536
rect 19220 12496 19229 12536
rect 19171 12495 19229 12496
rect 19467 12536 19509 12545
rect 19467 12496 19468 12536
rect 19508 12496 19509 12536
rect 19467 12487 19509 12496
rect 19563 12536 19605 12545
rect 19563 12496 19564 12536
rect 19604 12496 19605 12536
rect 19563 12487 19605 12496
rect 11211 12442 11253 12451
rect 16395 12452 16437 12461
rect 7083 12403 7125 12412
rect 16395 12412 16396 12452
rect 16436 12412 16437 12452
rect 16395 12403 16437 12412
rect 16587 12452 16629 12461
rect 16587 12412 16588 12452
rect 16628 12412 16629 12452
rect 16587 12403 16629 12412
rect 16867 12452 16925 12453
rect 16867 12412 16876 12452
rect 16916 12412 16925 12452
rect 16867 12411 16925 12412
rect 20035 12452 20093 12453
rect 20035 12412 20044 12452
rect 20084 12412 20093 12452
rect 20035 12411 20093 12412
rect 3235 12368 3293 12369
rect 3235 12328 3244 12368
rect 3284 12328 3293 12368
rect 3235 12327 3293 12328
rect 9963 12368 10005 12377
rect 9963 12328 9964 12368
rect 10004 12328 10005 12368
rect 9963 12319 10005 12328
rect 16107 12368 16149 12377
rect 16107 12328 16108 12368
rect 16148 12328 16149 12368
rect 16107 12319 16149 12328
rect 16491 12368 16533 12377
rect 16491 12328 16492 12368
rect 16532 12328 16533 12368
rect 16491 12319 16533 12328
rect 17067 12368 17109 12377
rect 17067 12328 17068 12368
rect 17108 12328 17109 12368
rect 17067 12319 17109 12328
rect 19843 12368 19901 12369
rect 19843 12328 19852 12368
rect 19892 12328 19901 12368
rect 19843 12327 19901 12328
rect 20235 12368 20277 12377
rect 20235 12328 20236 12368
rect 20276 12328 20277 12368
rect 20235 12319 20277 12328
rect 3051 12284 3093 12293
rect 3051 12244 3052 12284
rect 3092 12244 3093 12284
rect 3051 12235 3093 12244
rect 7851 12284 7893 12293
rect 7851 12244 7852 12284
rect 7892 12244 7893 12284
rect 7851 12235 7893 12244
rect 11691 12284 11733 12293
rect 11691 12244 11692 12284
rect 11732 12244 11733 12284
rect 11691 12235 11733 12244
rect 1152 12116 20352 12140
rect 1152 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 20352 12116
rect 1152 12052 20352 12076
rect 1515 11948 1557 11957
rect 1515 11908 1516 11948
rect 1556 11908 1557 11948
rect 1515 11899 1557 11908
rect 8323 11948 8381 11949
rect 8323 11908 8332 11948
rect 8372 11908 8381 11948
rect 8323 11907 8381 11908
rect 11403 11948 11445 11957
rect 11403 11908 11404 11948
rect 11444 11908 11445 11948
rect 11403 11899 11445 11908
rect 13035 11948 13077 11957
rect 13035 11908 13036 11948
rect 13076 11908 13077 11948
rect 13035 11899 13077 11908
rect 16587 11948 16629 11957
rect 16587 11908 16588 11948
rect 16628 11908 16629 11948
rect 16587 11899 16629 11908
rect 17643 11948 17685 11957
rect 17643 11908 17644 11948
rect 17684 11908 17685 11948
rect 17643 11899 17685 11908
rect 17835 11948 17877 11957
rect 17835 11908 17836 11948
rect 17876 11908 17877 11948
rect 17835 11899 17877 11908
rect 20043 11948 20085 11957
rect 20043 11908 20044 11948
rect 20084 11908 20085 11948
rect 20043 11899 20085 11908
rect 8139 11864 8181 11873
rect 8139 11824 8140 11864
rect 8180 11824 8181 11864
rect 8139 11815 8181 11824
rect 9579 11864 9621 11873
rect 9579 11824 9580 11864
rect 9620 11824 9621 11864
rect 9579 11815 9621 11824
rect 9483 11780 9525 11789
rect 9483 11740 9484 11780
rect 9524 11740 9525 11780
rect 2947 11738 3005 11739
rect 2947 11698 2956 11738
rect 2996 11698 3005 11738
rect 9483 11731 9525 11740
rect 9675 11780 9717 11789
rect 9675 11740 9676 11780
rect 9716 11740 9717 11780
rect 9675 11731 9717 11740
rect 17443 11780 17501 11781
rect 17443 11740 17452 11780
rect 17492 11740 17501 11780
rect 17443 11739 17501 11740
rect 19843 11780 19901 11781
rect 19843 11740 19852 11780
rect 19892 11740 19901 11780
rect 19843 11739 19901 11740
rect 2947 11697 3005 11698
rect 1315 11696 1373 11697
rect 1315 11656 1324 11696
rect 1364 11656 1373 11696
rect 1315 11655 1373 11656
rect 1699 11696 1757 11697
rect 1699 11656 1708 11696
rect 1748 11656 1757 11696
rect 1699 11655 1757 11656
rect 3139 11696 3197 11697
rect 3139 11656 3148 11696
rect 3188 11656 3197 11696
rect 3139 11655 3197 11656
rect 4387 11696 4445 11697
rect 4387 11656 4396 11696
rect 4436 11656 4445 11696
rect 4387 11655 4445 11656
rect 4867 11696 4925 11697
rect 4867 11656 4876 11696
rect 4916 11656 4925 11696
rect 4867 11655 4925 11656
rect 5251 11696 5309 11697
rect 5251 11656 5260 11696
rect 5300 11656 5309 11696
rect 5251 11655 5309 11656
rect 6499 11696 6557 11697
rect 6499 11656 6508 11696
rect 6548 11656 6557 11696
rect 6499 11655 6557 11656
rect 6691 11696 6749 11697
rect 6691 11656 6700 11696
rect 6740 11656 6749 11696
rect 6691 11655 6749 11656
rect 7939 11696 7997 11697
rect 7939 11656 7948 11696
rect 7988 11656 7997 11696
rect 7939 11655 7997 11656
rect 8619 11696 8661 11705
rect 8619 11656 8620 11696
rect 8660 11656 8661 11696
rect 8619 11647 8661 11656
rect 8715 11696 8757 11705
rect 8715 11656 8716 11696
rect 8756 11656 8757 11696
rect 8715 11647 8757 11656
rect 8995 11696 9053 11697
rect 8995 11656 9004 11696
rect 9044 11656 9053 11696
rect 8995 11655 9053 11656
rect 9387 11696 9429 11705
rect 9387 11656 9388 11696
rect 9428 11656 9429 11696
rect 9387 11647 9429 11656
rect 9763 11696 9821 11697
rect 9763 11656 9772 11696
rect 9812 11656 9821 11696
rect 9763 11655 9821 11656
rect 9955 11696 10013 11697
rect 9955 11656 9964 11696
rect 10004 11656 10013 11696
rect 9955 11655 10013 11656
rect 11203 11696 11261 11697
rect 11203 11656 11212 11696
rect 11252 11656 11261 11696
rect 11203 11655 11261 11656
rect 11587 11696 11645 11697
rect 11587 11656 11596 11696
rect 11636 11656 11645 11696
rect 11587 11655 11645 11656
rect 12835 11696 12893 11697
rect 12835 11656 12844 11696
rect 12884 11656 12893 11696
rect 12835 11655 12893 11656
rect 13411 11696 13469 11697
rect 13411 11656 13420 11696
rect 13460 11656 13469 11696
rect 13411 11655 13469 11656
rect 14659 11696 14717 11697
rect 14659 11656 14668 11696
rect 14708 11656 14717 11696
rect 14659 11655 14717 11656
rect 15043 11696 15101 11697
rect 15043 11656 15052 11696
rect 15092 11656 15101 11696
rect 15043 11655 15101 11656
rect 16291 11696 16349 11697
rect 16291 11656 16300 11696
rect 16340 11656 16349 11696
rect 16291 11655 16349 11656
rect 16579 11696 16637 11697
rect 16579 11656 16588 11696
rect 16628 11656 16637 11696
rect 16579 11655 16637 11656
rect 16675 11696 16733 11697
rect 16675 11656 16684 11696
rect 16724 11656 16733 11696
rect 16675 11655 16733 11656
rect 16875 11696 16917 11705
rect 16875 11656 16876 11696
rect 16916 11656 16917 11696
rect 16875 11647 16917 11656
rect 16971 11696 17013 11705
rect 16971 11656 16972 11696
rect 17012 11656 17013 11696
rect 16971 11647 17013 11656
rect 17118 11696 17176 11697
rect 17118 11656 17127 11696
rect 17167 11656 17176 11696
rect 17118 11655 17176 11656
rect 17835 11696 17877 11705
rect 17835 11656 17836 11696
rect 17876 11656 17877 11696
rect 17835 11647 17877 11656
rect 18027 11696 18069 11705
rect 18027 11656 18028 11696
rect 18068 11656 18069 11696
rect 18027 11647 18069 11656
rect 18211 11696 18269 11697
rect 18211 11656 18220 11696
rect 18260 11656 18269 11696
rect 18211 11655 18269 11656
rect 19459 11696 19517 11697
rect 19459 11656 19468 11696
rect 19508 11656 19517 11696
rect 19459 11655 19517 11656
rect 4779 11612 4821 11621
rect 4779 11572 4780 11612
rect 4820 11572 4821 11612
rect 4779 11563 4821 11572
rect 1227 11528 1269 11537
rect 1227 11488 1228 11528
rect 1268 11488 1269 11528
rect 1227 11479 1269 11488
rect 1515 11528 1557 11537
rect 1515 11488 1516 11528
rect 1556 11488 1557 11528
rect 1515 11479 1557 11488
rect 4587 11528 4629 11537
rect 4587 11488 4588 11528
rect 4628 11488 4629 11528
rect 4587 11479 4629 11488
rect 5067 11528 5109 11537
rect 5067 11488 5068 11528
rect 5108 11488 5109 11528
rect 5067 11479 5109 11488
rect 11403 11528 11445 11537
rect 11403 11488 11404 11528
rect 11444 11488 11445 11528
rect 11403 11479 11445 11488
rect 13035 11528 13077 11537
rect 13035 11488 13036 11528
rect 13076 11488 13077 11528
rect 13035 11479 13077 11488
rect 13227 11528 13269 11537
rect 13227 11488 13228 11528
rect 13268 11488 13269 11528
rect 13227 11479 13269 11488
rect 14859 11528 14901 11537
rect 14859 11488 14860 11528
rect 14900 11488 14901 11528
rect 14859 11479 14901 11488
rect 19659 11528 19701 11537
rect 19659 11488 19660 11528
rect 19700 11488 19701 11528
rect 19659 11479 19701 11488
rect 1152 11360 20452 11384
rect 1152 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20452 11360
rect 1152 11296 20452 11320
rect 1323 11192 1365 11201
rect 1323 11152 1324 11192
rect 1364 11152 1365 11192
rect 1323 11143 1365 11152
rect 2947 11192 3005 11193
rect 2947 11152 2956 11192
rect 2996 11152 3005 11192
rect 2947 11151 3005 11152
rect 18123 11192 18165 11201
rect 18123 11152 18124 11192
rect 18164 11152 18165 11192
rect 18123 11143 18165 11152
rect 20235 11192 20277 11201
rect 20235 11152 20236 11192
rect 20276 11152 20277 11192
rect 20235 11143 20277 11152
rect 6603 11108 6645 11117
rect 6603 11068 6604 11108
rect 6644 11068 6645 11108
rect 6603 11059 6645 11068
rect 6795 11108 6837 11117
rect 6795 11068 6796 11108
rect 6836 11068 6837 11108
rect 6795 11059 6837 11068
rect 9291 11108 9333 11117
rect 9291 11068 9292 11108
rect 9332 11068 9333 11108
rect 9291 11059 9333 11068
rect 12747 11108 12789 11117
rect 12747 11068 12748 11108
rect 12788 11068 12789 11108
rect 12747 11059 12789 11068
rect 1507 11024 1565 11025
rect 1507 10984 1516 11024
rect 1556 10984 1565 11024
rect 1507 10983 1565 10984
rect 2755 11024 2813 11025
rect 2755 10984 2764 11024
rect 2804 10984 2813 11024
rect 2755 10983 2813 10984
rect 3147 11024 3189 11033
rect 3147 10984 3148 11024
rect 3188 10984 3189 11024
rect 3715 11024 3773 11025
rect 3147 10975 3189 10984
rect 3240 11014 3298 11015
rect 3240 10974 3249 11014
rect 3289 10974 3298 11014
rect 3715 10984 3724 11024
rect 3764 10984 3773 11024
rect 3715 10983 3773 10984
rect 4963 11024 5021 11025
rect 4963 10984 4972 11024
rect 5012 10984 5021 11024
rect 4963 10983 5021 10984
rect 5155 11024 5213 11025
rect 5155 10984 5164 11024
rect 5204 10984 5213 11024
rect 5155 10983 5213 10984
rect 6403 11024 6461 11025
rect 6403 10984 6412 11024
rect 6452 10984 6461 11024
rect 6403 10983 6461 10984
rect 6987 11019 7029 11028
rect 3240 10973 3298 10974
rect 6987 10979 6988 11019
rect 7028 10979 7029 11019
rect 7459 11024 7517 11025
rect 7459 10984 7468 11024
rect 7508 10984 7517 11024
rect 7459 10983 7517 10984
rect 7947 11024 7989 11033
rect 7947 10984 7948 11024
rect 7988 10984 7989 11024
rect 6987 10970 7029 10979
rect 7947 10975 7989 10984
rect 8427 11024 8469 11033
rect 8427 10984 8428 11024
rect 8468 10984 8469 11024
rect 8427 10975 8469 10984
rect 8523 11024 8565 11033
rect 8523 10984 8524 11024
rect 8564 10984 8565 11024
rect 8523 10975 8565 10984
rect 8811 11024 8853 11033
rect 8811 10984 8812 11024
rect 8852 10984 8853 11024
rect 8811 10975 8853 10984
rect 9099 11024 9141 11033
rect 9099 10984 9100 11024
rect 9140 10984 9141 11024
rect 9099 10975 9141 10984
rect 9475 11024 9533 11025
rect 9475 10984 9484 11024
rect 9524 10984 9533 11024
rect 9475 10983 9533 10984
rect 10723 11024 10781 11025
rect 10723 10984 10732 11024
rect 10772 10984 10781 11024
rect 10723 10983 10781 10984
rect 11019 11024 11061 11033
rect 11019 10984 11020 11024
rect 11060 10984 11061 11024
rect 11019 10975 11061 10984
rect 11115 11024 11157 11033
rect 11115 10984 11116 11024
rect 11156 10984 11157 11024
rect 11115 10975 11157 10984
rect 12067 11024 12125 11025
rect 12067 10984 12076 11024
rect 12116 10984 12125 11024
rect 12067 10983 12125 10984
rect 12555 11019 12597 11028
rect 12555 10979 12556 11019
rect 12596 10979 12597 11019
rect 13027 11024 13085 11025
rect 13027 10984 13036 11024
rect 13076 10984 13085 11024
rect 13027 10983 13085 10984
rect 14275 11024 14333 11025
rect 14275 10984 14284 11024
rect 14324 10984 14333 11024
rect 14275 10983 14333 10984
rect 14851 11024 14909 11025
rect 14851 10984 14860 11024
rect 14900 10984 14909 11024
rect 14851 10983 14909 10984
rect 15043 11024 15101 11025
rect 15043 10984 15052 11024
rect 15092 10984 15101 11024
rect 15043 10983 15101 10984
rect 16291 11024 16349 11025
rect 16291 10984 16300 11024
rect 16340 10984 16349 11024
rect 16291 10983 16349 10984
rect 16771 11024 16829 11025
rect 16771 10984 16780 11024
rect 16820 10984 16829 11024
rect 16771 10983 16829 10984
rect 17067 11024 17109 11033
rect 17067 10984 17068 11024
rect 17108 10984 17109 11024
rect 12555 10970 12597 10979
rect 17067 10975 17109 10984
rect 17163 11024 17205 11033
rect 17163 10984 17164 11024
rect 17204 10984 17205 11024
rect 17163 10975 17205 10984
rect 17643 11024 17685 11033
rect 17643 10984 17644 11024
rect 17684 10984 17685 11024
rect 17643 10975 17685 10984
rect 17835 11024 17877 11033
rect 17835 10984 17836 11024
rect 17876 10984 17877 11024
rect 17835 10975 17877 10984
rect 18027 11024 18069 11033
rect 18027 10984 18028 11024
rect 18068 10984 18069 11024
rect 18027 10975 18069 10984
rect 18219 11024 18261 11033
rect 18219 10984 18220 11024
rect 18260 10984 18261 11024
rect 18219 10975 18261 10984
rect 18403 11024 18461 11025
rect 18403 10984 18412 11024
rect 18452 10984 18461 11024
rect 18403 10983 18461 10984
rect 19651 11024 19709 11025
rect 19651 10984 19660 11024
rect 19700 10984 19709 11024
rect 19651 10983 19709 10984
rect 8043 10940 8085 10949
rect 8043 10900 8044 10940
rect 8084 10900 8085 10940
rect 8043 10891 8085 10900
rect 11499 10940 11541 10949
rect 11499 10900 11500 10940
rect 11540 10900 11541 10940
rect 11499 10891 11541 10900
rect 11595 10940 11637 10949
rect 11595 10900 11596 10940
rect 11636 10900 11637 10940
rect 11595 10891 11637 10900
rect 20035 10940 20093 10941
rect 20035 10900 20044 10940
rect 20084 10900 20093 10940
rect 20035 10899 20093 10900
rect 17443 10856 17501 10857
rect 17443 10816 17452 10856
rect 17492 10816 17501 10856
rect 17443 10815 17501 10816
rect 3531 10772 3573 10781
rect 3531 10732 3532 10772
rect 3572 10732 3573 10772
rect 3531 10723 3573 10732
rect 9099 10772 9141 10781
rect 9099 10732 9100 10772
rect 9140 10732 9141 10772
rect 9099 10723 9141 10732
rect 14475 10772 14517 10781
rect 14475 10732 14476 10772
rect 14516 10732 14517 10772
rect 14475 10723 14517 10732
rect 14763 10772 14805 10781
rect 14763 10732 14764 10772
rect 14804 10732 14805 10772
rect 14763 10723 14805 10732
rect 16491 10772 16533 10781
rect 16491 10732 16492 10772
rect 16532 10732 16533 10772
rect 16491 10723 16533 10732
rect 17643 10772 17685 10781
rect 17643 10732 17644 10772
rect 17684 10732 17685 10772
rect 17643 10723 17685 10732
rect 19851 10772 19893 10781
rect 19851 10732 19852 10772
rect 19892 10732 19893 10772
rect 19851 10723 19893 10732
rect 1152 10604 20352 10628
rect 1152 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 20352 10604
rect 1152 10540 20352 10564
rect 2667 10436 2709 10445
rect 2667 10396 2668 10436
rect 2708 10396 2709 10436
rect 2667 10387 2709 10396
rect 2851 10436 2909 10437
rect 2851 10396 2860 10436
rect 2900 10396 2909 10436
rect 2851 10395 2909 10396
rect 9859 10436 9917 10437
rect 9859 10396 9868 10436
rect 9908 10396 9917 10436
rect 9859 10395 9917 10396
rect 15819 10436 15861 10445
rect 15819 10396 15820 10436
rect 15860 10396 15861 10436
rect 15819 10387 15861 10396
rect 11403 10352 11445 10361
rect 11403 10312 11404 10352
rect 11444 10312 11445 10352
rect 11403 10303 11445 10312
rect 11979 10352 12021 10361
rect 11979 10312 11980 10352
rect 12020 10312 12021 10352
rect 11979 10303 12021 10312
rect 16203 10352 16245 10361
rect 16203 10312 16204 10352
rect 16244 10312 16245 10352
rect 16203 10303 16245 10312
rect 16579 10352 16637 10353
rect 16579 10312 16588 10352
rect 16628 10312 16637 10352
rect 16579 10311 16637 10312
rect 17739 10352 17781 10361
rect 17739 10312 17740 10352
rect 17780 10312 17781 10352
rect 17739 10303 17781 10312
rect 5067 10268 5109 10277
rect 5067 10228 5068 10268
rect 5108 10228 5109 10268
rect 5067 10219 5109 10228
rect 10923 10268 10965 10277
rect 10923 10228 10924 10268
rect 10964 10228 10965 10268
rect 10923 10219 10965 10228
rect 11307 10268 11349 10277
rect 11307 10228 11308 10268
rect 11348 10228 11349 10268
rect 11307 10219 11349 10228
rect 11499 10268 11541 10277
rect 11499 10228 11500 10268
rect 11540 10228 11541 10268
rect 11499 10219 11541 10228
rect 11883 10268 11925 10277
rect 11883 10228 11884 10268
rect 11924 10228 11925 10268
rect 11883 10219 11925 10228
rect 12075 10268 12117 10277
rect 12075 10228 12076 10268
rect 12116 10228 12117 10268
rect 12075 10219 12117 10228
rect 13707 10268 13749 10277
rect 13707 10228 13708 10268
rect 13748 10228 13749 10268
rect 12355 10226 12413 10227
rect 4011 10198 4053 10207
rect 1219 10184 1277 10185
rect 1219 10144 1228 10184
rect 1268 10144 1277 10184
rect 1219 10143 1277 10144
rect 2467 10184 2525 10185
rect 2467 10144 2476 10184
rect 2516 10144 2525 10184
rect 2467 10143 2525 10144
rect 3243 10184 3285 10193
rect 3243 10144 3244 10184
rect 3284 10144 3285 10184
rect 3243 10135 3285 10144
rect 3523 10184 3581 10185
rect 3523 10144 3532 10184
rect 3572 10144 3581 10184
rect 4011 10158 4012 10198
rect 4052 10158 4053 10198
rect 4011 10149 4053 10158
rect 4483 10184 4541 10185
rect 3523 10143 3581 10144
rect 4483 10144 4492 10184
rect 4532 10144 4541 10184
rect 4483 10143 4541 10144
rect 4971 10184 5013 10193
rect 4971 10144 4972 10184
rect 5012 10144 5013 10184
rect 4971 10135 5013 10144
rect 5451 10184 5493 10193
rect 5451 10144 5452 10184
rect 5492 10144 5493 10184
rect 5451 10135 5493 10144
rect 5547 10184 5589 10193
rect 5547 10144 5548 10184
rect 5588 10144 5589 10184
rect 5547 10135 5589 10144
rect 5923 10184 5981 10185
rect 5923 10144 5932 10184
rect 5972 10144 5981 10184
rect 5923 10143 5981 10144
rect 7171 10184 7229 10185
rect 7171 10144 7180 10184
rect 7220 10144 7229 10184
rect 7171 10143 7229 10144
rect 7755 10184 7797 10193
rect 7755 10144 7756 10184
rect 7796 10144 7797 10184
rect 7755 10135 7797 10144
rect 7851 10184 7893 10193
rect 7851 10144 7852 10184
rect 7892 10144 7893 10184
rect 7851 10135 7893 10144
rect 7947 10184 7989 10193
rect 7947 10144 7948 10184
rect 7988 10144 7989 10184
rect 7947 10135 7989 10144
rect 8043 10184 8085 10193
rect 8043 10144 8044 10184
rect 8084 10144 8085 10184
rect 8043 10135 8085 10144
rect 8227 10184 8285 10185
rect 8227 10144 8236 10184
rect 8276 10144 8285 10184
rect 8227 10143 8285 10144
rect 9475 10184 9533 10185
rect 9475 10144 9484 10184
rect 9524 10144 9533 10184
rect 9475 10143 9533 10144
rect 10155 10184 10197 10193
rect 10155 10144 10156 10184
rect 10196 10144 10197 10184
rect 10155 10135 10197 10144
rect 10251 10184 10293 10193
rect 10251 10144 10252 10184
rect 10292 10144 10293 10184
rect 10251 10135 10293 10144
rect 10531 10184 10589 10185
rect 10531 10144 10540 10184
rect 10580 10144 10589 10184
rect 10531 10143 10589 10144
rect 10827 10184 10869 10193
rect 10827 10144 10828 10184
rect 10868 10144 10869 10184
rect 10827 10135 10869 10144
rect 11019 10184 11061 10193
rect 11019 10144 11020 10184
rect 11060 10144 11061 10184
rect 11019 10135 11061 10144
rect 11203 10184 11261 10185
rect 11203 10144 11212 10184
rect 11252 10144 11261 10184
rect 11203 10143 11261 10144
rect 11595 10184 11637 10193
rect 11595 10144 11596 10184
rect 11636 10144 11637 10184
rect 11595 10135 11637 10144
rect 11779 10184 11837 10185
rect 11779 10144 11788 10184
rect 11828 10144 11837 10184
rect 11779 10143 11837 10144
rect 12171 10184 12213 10193
rect 12355 10186 12364 10226
rect 12404 10186 12413 10226
rect 13707 10219 13749 10228
rect 13803 10268 13845 10277
rect 13803 10228 13804 10268
rect 13844 10228 13845 10268
rect 13803 10219 13845 10228
rect 16107 10268 16149 10277
rect 16107 10228 16108 10268
rect 16148 10228 16149 10268
rect 16107 10219 16149 10228
rect 16299 10268 16341 10277
rect 16299 10228 16300 10268
rect 16340 10228 16341 10268
rect 16299 10219 16341 10228
rect 19843 10226 19901 10227
rect 14763 10198 14805 10207
rect 12355 10185 12413 10186
rect 12171 10144 12172 10184
rect 12212 10144 12213 10184
rect 12171 10135 12213 10144
rect 12555 10184 12597 10193
rect 12555 10144 12556 10184
rect 12596 10144 12597 10184
rect 12555 10135 12597 10144
rect 12643 10184 12701 10185
rect 12643 10144 12652 10184
rect 12692 10144 12701 10184
rect 12643 10143 12701 10144
rect 12835 10184 12893 10185
rect 12835 10144 12844 10184
rect 12884 10144 12893 10184
rect 12835 10143 12893 10144
rect 13227 10184 13269 10193
rect 13227 10144 13228 10184
rect 13268 10144 13269 10184
rect 13227 10135 13269 10144
rect 13323 10184 13365 10193
rect 13323 10144 13324 10184
rect 13364 10144 13365 10184
rect 13323 10135 13365 10144
rect 14275 10184 14333 10185
rect 14275 10144 14284 10184
rect 14324 10144 14333 10184
rect 14763 10158 14764 10198
rect 14804 10158 14805 10198
rect 14763 10149 14805 10158
rect 15235 10184 15293 10185
rect 14275 10143 14333 10144
rect 15235 10144 15244 10184
rect 15284 10144 15293 10184
rect 15235 10143 15293 10144
rect 15523 10184 15581 10185
rect 15523 10144 15532 10184
rect 15572 10144 15581 10184
rect 15523 10143 15581 10144
rect 15627 10184 15669 10193
rect 15627 10144 15628 10184
rect 15668 10144 15669 10184
rect 15627 10135 15669 10144
rect 15811 10184 15869 10185
rect 15811 10144 15820 10184
rect 15860 10144 15869 10184
rect 15811 10143 15869 10144
rect 16003 10184 16061 10185
rect 16003 10144 16012 10184
rect 16052 10144 16061 10184
rect 16003 10143 16061 10144
rect 16395 10184 16437 10193
rect 16395 10144 16396 10184
rect 16436 10144 16437 10184
rect 16395 10135 16437 10144
rect 16875 10184 16917 10193
rect 16875 10144 16876 10184
rect 16916 10144 16917 10184
rect 16875 10135 16917 10144
rect 16971 10184 17013 10193
rect 16971 10144 16972 10184
rect 17012 10144 17013 10184
rect 16971 10135 17013 10144
rect 17251 10184 17309 10185
rect 17251 10144 17260 10184
rect 17300 10144 17309 10184
rect 17251 10143 17309 10144
rect 17739 10184 17781 10193
rect 17739 10144 17740 10184
rect 17780 10144 17781 10184
rect 17739 10135 17781 10144
rect 18115 10184 18173 10185
rect 18115 10144 18124 10184
rect 18164 10144 18173 10184
rect 18115 10143 18173 10144
rect 19363 10184 19421 10185
rect 19363 10144 19372 10184
rect 19412 10144 19421 10184
rect 19363 10143 19421 10144
rect 19755 10184 19797 10193
rect 19843 10186 19852 10226
rect 19892 10186 19901 10226
rect 19843 10185 19901 10186
rect 19755 10144 19756 10184
rect 19796 10144 19797 10184
rect 19755 10135 19797 10144
rect 19947 10184 19989 10193
rect 19947 10144 19948 10184
rect 19988 10144 19989 10184
rect 19947 10135 19989 10144
rect 3147 10100 3189 10109
rect 3147 10060 3148 10100
rect 3188 10060 3189 10100
rect 3147 10051 3189 10060
rect 3819 10100 3861 10109
rect 3819 10060 3820 10100
rect 3860 10060 3861 10100
rect 3819 10051 3861 10060
rect 7371 10100 7413 10109
rect 7371 10060 7372 10100
rect 7412 10060 7413 10100
rect 7371 10051 7413 10060
rect 9675 10016 9717 10025
rect 9675 9976 9676 10016
rect 9716 9976 9717 10016
rect 9675 9967 9717 9976
rect 12363 10016 12405 10025
rect 12363 9976 12364 10016
rect 12404 9976 12405 10016
rect 12363 9967 12405 9976
rect 12939 10016 12981 10025
rect 12939 9976 12940 10016
rect 12980 9976 12981 10016
rect 12939 9967 12981 9976
rect 14955 10016 14997 10025
rect 14955 9976 14956 10016
rect 14996 9976 14997 10016
rect 14955 9967 14997 9976
rect 15339 10016 15381 10025
rect 15339 9976 15340 10016
rect 15380 9976 15381 10016
rect 15339 9967 15381 9976
rect 17931 10016 17973 10025
rect 17931 9976 17932 10016
rect 17972 9976 17973 10016
rect 17931 9967 17973 9976
rect 19563 10016 19605 10025
rect 19563 9976 19564 10016
rect 19604 9976 19605 10016
rect 19563 9967 19605 9976
rect 20035 10016 20093 10017
rect 20035 9976 20044 10016
rect 20084 9976 20093 10016
rect 20035 9975 20093 9976
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 3243 9680 3285 9689
rect 3243 9640 3244 9680
rect 3284 9640 3285 9680
rect 3243 9631 3285 9640
rect 4483 9680 4541 9681
rect 4483 9640 4492 9680
rect 4532 9640 4541 9680
rect 4483 9639 4541 9640
rect 9955 9680 10013 9681
rect 9955 9640 9964 9680
rect 10004 9640 10013 9680
rect 9955 9639 10013 9640
rect 12075 9680 12117 9689
rect 12075 9640 12076 9680
rect 12116 9640 12117 9680
rect 12075 9631 12117 9640
rect 12643 9680 12701 9681
rect 12643 9640 12652 9680
rect 12692 9640 12701 9680
rect 12643 9639 12701 9640
rect 17923 9680 17981 9681
rect 17923 9640 17932 9680
rect 17972 9640 17981 9680
rect 17923 9639 17981 9640
rect 3723 9596 3765 9605
rect 3723 9556 3724 9596
rect 3764 9556 3765 9596
rect 3723 9547 3765 9556
rect 13515 9596 13557 9605
rect 13515 9556 13516 9596
rect 13556 9556 13557 9596
rect 13515 9547 13557 9556
rect 17067 9596 17109 9605
rect 17067 9556 17068 9596
rect 17108 9556 17109 9596
rect 17067 9547 17109 9556
rect 20126 9523 20168 9532
rect 1323 9512 1365 9521
rect 1323 9472 1324 9512
rect 1364 9472 1365 9512
rect 1323 9463 1365 9472
rect 1515 9512 1557 9521
rect 1515 9472 1516 9512
rect 1556 9472 1557 9512
rect 1515 9463 1557 9472
rect 1603 9512 1661 9513
rect 1603 9472 1612 9512
rect 1652 9472 1661 9512
rect 1603 9471 1661 9472
rect 1795 9512 1853 9513
rect 1795 9472 1804 9512
rect 1844 9472 1853 9512
rect 1795 9471 1853 9472
rect 3043 9512 3101 9513
rect 3043 9472 3052 9512
rect 3092 9472 3101 9512
rect 3043 9471 3101 9472
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 4099 9512 4157 9513
rect 4099 9472 4108 9512
rect 4148 9472 4157 9512
rect 4099 9471 4157 9472
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4587 9512 4629 9521
rect 4587 9472 4588 9512
rect 4628 9472 4629 9512
rect 4587 9463 4629 9472
rect 4675 9512 4733 9513
rect 4675 9472 4684 9512
rect 4724 9472 4733 9512
rect 4675 9471 4733 9472
rect 4867 9512 4925 9513
rect 4867 9472 4876 9512
rect 4916 9472 4925 9512
rect 4867 9471 4925 9472
rect 6115 9512 6173 9513
rect 6115 9472 6124 9512
rect 6164 9472 6173 9512
rect 6115 9471 6173 9472
rect 6499 9512 6557 9513
rect 6499 9472 6508 9512
rect 6548 9472 6557 9512
rect 6499 9471 6557 9472
rect 7747 9512 7805 9513
rect 7747 9472 7756 9512
rect 7796 9472 7805 9512
rect 7747 9471 7805 9472
rect 8323 9512 8381 9513
rect 8323 9472 8332 9512
rect 8372 9472 8381 9512
rect 8323 9471 8381 9472
rect 9571 9512 9629 9513
rect 9571 9472 9580 9512
rect 9620 9472 9629 9512
rect 9571 9471 9629 9472
rect 9763 9512 9821 9513
rect 9763 9472 9772 9512
rect 9812 9472 9821 9512
rect 9763 9471 9821 9472
rect 9859 9512 9917 9513
rect 9859 9472 9868 9512
rect 9908 9472 9917 9512
rect 9859 9471 9917 9472
rect 10059 9512 10101 9521
rect 10059 9472 10060 9512
rect 10100 9472 10101 9512
rect 10059 9463 10101 9472
rect 10155 9512 10197 9521
rect 10155 9472 10156 9512
rect 10196 9472 10197 9512
rect 10155 9463 10197 9472
rect 10248 9512 10306 9513
rect 10248 9472 10257 9512
rect 10297 9472 10306 9512
rect 10248 9471 10306 9472
rect 10627 9512 10685 9513
rect 10627 9472 10636 9512
rect 10676 9472 10685 9512
rect 10627 9471 10685 9472
rect 11875 9512 11933 9513
rect 11875 9472 11884 9512
rect 11924 9472 11933 9512
rect 11875 9471 11933 9472
rect 12259 9512 12317 9513
rect 12259 9472 12268 9512
rect 12308 9472 12317 9512
rect 12555 9512 12597 9521
rect 12259 9471 12317 9472
rect 12403 9489 12461 9490
rect 12403 9449 12412 9489
rect 12452 9449 12461 9489
rect 12555 9472 12556 9512
rect 12596 9472 12597 9512
rect 13035 9512 13077 9521
rect 12808 9497 12850 9506
rect 12555 9463 12597 9472
rect 12643 9483 12701 9484
rect 12403 9448 12461 9449
rect 12643 9443 12652 9483
rect 12692 9443 12701 9483
rect 12808 9457 12809 9497
rect 12849 9457 12850 9497
rect 13035 9472 13036 9512
rect 13076 9472 13077 9512
rect 13035 9463 13077 9472
rect 13227 9512 13269 9521
rect 13227 9472 13228 9512
rect 13268 9472 13269 9512
rect 13227 9463 13269 9472
rect 13707 9507 13749 9516
rect 13707 9467 13708 9507
rect 13748 9467 13749 9507
rect 14179 9512 14237 9513
rect 14179 9472 14188 9512
rect 14228 9472 14237 9512
rect 14179 9471 14237 9472
rect 14763 9512 14805 9521
rect 14763 9472 14764 9512
rect 14804 9472 14805 9512
rect 13707 9458 13749 9467
rect 14763 9463 14805 9472
rect 15147 9512 15189 9521
rect 15147 9472 15148 9512
rect 15188 9472 15189 9512
rect 15147 9463 15189 9472
rect 15243 9512 15285 9521
rect 15243 9472 15244 9512
rect 15284 9472 15285 9512
rect 15243 9463 15285 9472
rect 15619 9512 15677 9513
rect 15619 9472 15628 9512
rect 15668 9472 15677 9512
rect 15619 9471 15677 9472
rect 16011 9512 16053 9521
rect 16011 9472 16012 9512
rect 16052 9472 16053 9512
rect 16011 9463 16053 9472
rect 16195 9512 16253 9513
rect 16195 9472 16204 9512
rect 16244 9472 16253 9512
rect 16195 9471 16253 9472
rect 16587 9512 16629 9521
rect 16587 9472 16588 9512
rect 16628 9472 16629 9512
rect 16587 9463 16629 9472
rect 17163 9512 17205 9521
rect 17163 9472 17164 9512
rect 17204 9472 17205 9512
rect 17163 9463 17205 9472
rect 17443 9512 17501 9513
rect 17443 9472 17452 9512
rect 17492 9472 17501 9512
rect 17443 9471 17501 9472
rect 17731 9512 17789 9513
rect 17731 9472 17740 9512
rect 17780 9472 17789 9512
rect 17731 9471 17789 9472
rect 17827 9512 17885 9513
rect 17827 9472 17836 9512
rect 17876 9472 17885 9512
rect 17827 9471 17885 9472
rect 18027 9512 18069 9521
rect 18027 9472 18028 9512
rect 18068 9472 18069 9512
rect 18027 9463 18069 9472
rect 18123 9512 18165 9521
rect 18123 9472 18124 9512
rect 18164 9472 18165 9512
rect 18123 9463 18165 9472
rect 18216 9512 18274 9513
rect 18216 9472 18225 9512
rect 18265 9472 18274 9512
rect 18216 9471 18274 9472
rect 18787 9512 18845 9513
rect 18787 9472 18796 9512
rect 18836 9472 18845 9512
rect 18787 9471 18845 9472
rect 19083 9512 19125 9521
rect 19083 9472 19084 9512
rect 19124 9472 19125 9512
rect 19083 9463 19125 9472
rect 19179 9512 19221 9521
rect 19179 9472 19180 9512
rect 19220 9472 19221 9512
rect 19179 9463 19221 9472
rect 19651 9512 19709 9513
rect 19651 9472 19660 9512
rect 19700 9472 19709 9512
rect 19651 9471 19709 9472
rect 19755 9512 19797 9521
rect 19755 9472 19756 9512
rect 19796 9472 19797 9512
rect 19755 9463 19797 9472
rect 19947 9512 19989 9521
rect 19947 9472 19948 9512
rect 19988 9472 19989 9512
rect 20126 9483 20127 9523
rect 20167 9483 20168 9523
rect 20126 9474 20168 9483
rect 19947 9463 19989 9472
rect 12808 9448 12850 9457
rect 12643 9442 12701 9443
rect 14667 9428 14709 9437
rect 14667 9388 14668 9428
rect 14708 9388 14709 9428
rect 14667 9379 14709 9388
rect 15723 9428 15765 9437
rect 15723 9388 15724 9428
rect 15764 9388 15765 9428
rect 15723 9379 15765 9388
rect 15915 9428 15957 9437
rect 15915 9388 15916 9428
rect 15956 9388 15957 9428
rect 15915 9379 15957 9388
rect 16299 9428 16341 9437
rect 16299 9388 16300 9428
rect 16340 9388 16341 9428
rect 16299 9379 16341 9388
rect 16491 9428 16533 9437
rect 16491 9388 16492 9428
rect 16532 9388 16533 9428
rect 16491 9379 16533 9388
rect 20235 9428 20277 9437
rect 20235 9388 20236 9428
rect 20276 9388 20277 9428
rect 20235 9379 20277 9388
rect 8139 9344 8181 9353
rect 8139 9304 8140 9344
rect 8180 9304 8181 9344
rect 8139 9295 8181 9304
rect 13035 9344 13077 9353
rect 13035 9304 13036 9344
rect 13076 9304 13077 9344
rect 13035 9295 13077 9304
rect 15819 9344 15861 9353
rect 15819 9304 15820 9344
rect 15860 9304 15861 9344
rect 15819 9295 15861 9304
rect 16395 9344 16437 9353
rect 16395 9304 16396 9344
rect 16436 9304 16437 9344
rect 16395 9295 16437 9304
rect 19459 9344 19517 9345
rect 19459 9304 19468 9344
rect 19508 9304 19517 9344
rect 19459 9303 19517 9304
rect 19947 9344 19989 9353
rect 19947 9304 19948 9344
rect 19988 9304 19989 9344
rect 19947 9295 19989 9304
rect 1323 9260 1365 9269
rect 1323 9220 1324 9260
rect 1364 9220 1365 9260
rect 1323 9211 1365 9220
rect 3427 9260 3485 9261
rect 3427 9220 3436 9260
rect 3476 9220 3485 9260
rect 3427 9219 3485 9220
rect 6315 9260 6357 9269
rect 6315 9220 6316 9260
rect 6356 9220 6357 9260
rect 6315 9211 6357 9220
rect 7947 9260 7989 9269
rect 7947 9220 7948 9260
rect 7988 9220 7989 9260
rect 7947 9211 7989 9220
rect 16771 9260 16829 9261
rect 16771 9220 16780 9260
rect 16820 9220 16829 9260
rect 16771 9219 16829 9220
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 3235 8924 3293 8925
rect 3235 8884 3244 8924
rect 3284 8884 3293 8924
rect 3235 8883 3293 8884
rect 10147 8924 10205 8925
rect 10147 8884 10156 8924
rect 10196 8884 10205 8924
rect 10147 8883 10205 8884
rect 11395 8924 11453 8925
rect 11395 8884 11404 8924
rect 11444 8884 11453 8924
rect 11395 8883 11453 8884
rect 13123 8924 13181 8925
rect 13123 8884 13132 8924
rect 13172 8884 13181 8924
rect 13123 8883 13181 8884
rect 16779 8924 16821 8933
rect 16779 8884 16780 8924
rect 16820 8884 16821 8924
rect 16779 8875 16821 8884
rect 17827 8924 17885 8925
rect 17827 8884 17836 8924
rect 17876 8884 17885 8924
rect 17827 8883 17885 8884
rect 6219 8840 6261 8849
rect 6219 8800 6220 8840
rect 6260 8800 6261 8840
rect 6219 8791 6261 8800
rect 2851 8756 2909 8757
rect 2851 8716 2860 8756
rect 2900 8716 2909 8756
rect 2851 8715 2909 8716
rect 18123 8756 18165 8765
rect 18123 8716 18124 8756
rect 18164 8716 18165 8756
rect 14659 8714 14717 8715
rect 8139 8686 8181 8695
rect 1219 8672 1277 8673
rect 1219 8632 1228 8672
rect 1268 8632 1277 8672
rect 1219 8631 1277 8632
rect 2467 8672 2525 8673
rect 2467 8632 2476 8672
rect 2516 8632 2525 8672
rect 2467 8631 2525 8632
rect 3531 8672 3573 8681
rect 3531 8632 3532 8672
rect 3572 8632 3573 8672
rect 3531 8623 3573 8632
rect 3627 8672 3669 8681
rect 3627 8632 3628 8672
rect 3668 8632 3669 8672
rect 3627 8623 3669 8632
rect 3907 8672 3965 8673
rect 3907 8632 3916 8672
rect 3956 8632 3965 8672
rect 3907 8631 3965 8632
rect 4299 8672 4341 8681
rect 4299 8632 4300 8672
rect 4340 8632 4341 8672
rect 4299 8623 4341 8632
rect 4395 8672 4437 8681
rect 4395 8632 4396 8672
rect 4436 8632 4437 8672
rect 4395 8623 4437 8632
rect 4779 8672 4821 8681
rect 4779 8632 4780 8672
rect 4820 8632 4821 8672
rect 4779 8623 4821 8632
rect 4875 8672 4917 8681
rect 5835 8677 5877 8686
rect 4875 8632 4876 8672
rect 4916 8632 4917 8672
rect 4875 8623 4917 8632
rect 5347 8672 5405 8673
rect 5347 8632 5356 8672
rect 5396 8632 5405 8672
rect 5347 8631 5405 8632
rect 5835 8637 5836 8677
rect 5876 8637 5877 8677
rect 5835 8628 5877 8637
rect 6603 8672 6645 8681
rect 6603 8632 6604 8672
rect 6644 8632 6645 8672
rect 6603 8623 6645 8632
rect 6699 8672 6741 8681
rect 6699 8632 6700 8672
rect 6740 8632 6741 8672
rect 6699 8623 6741 8632
rect 7083 8672 7125 8681
rect 7083 8632 7084 8672
rect 7124 8632 7125 8672
rect 7083 8623 7125 8632
rect 7179 8672 7221 8681
rect 7179 8632 7180 8672
rect 7220 8632 7221 8672
rect 7179 8623 7221 8632
rect 7651 8672 7709 8673
rect 7651 8632 7660 8672
rect 7700 8632 7709 8672
rect 8139 8646 8140 8686
rect 8180 8646 8181 8686
rect 8139 8637 8181 8646
rect 8515 8672 8573 8673
rect 7651 8631 7709 8632
rect 8515 8632 8524 8672
rect 8564 8632 8573 8672
rect 8515 8631 8573 8632
rect 9763 8672 9821 8673
rect 9763 8632 9772 8672
rect 9812 8632 9821 8672
rect 9763 8631 9821 8632
rect 10443 8672 10485 8681
rect 10443 8632 10444 8672
rect 10484 8632 10485 8672
rect 10443 8623 10485 8632
rect 10539 8672 10581 8681
rect 10539 8632 10540 8672
rect 10580 8632 10581 8672
rect 10539 8623 10581 8632
rect 10819 8672 10877 8673
rect 10819 8632 10828 8672
rect 10868 8632 10877 8672
rect 10819 8631 10877 8632
rect 11115 8672 11157 8681
rect 11115 8632 11116 8672
rect 11156 8632 11157 8672
rect 11115 8623 11157 8632
rect 11203 8672 11261 8673
rect 11203 8632 11212 8672
rect 11252 8632 11261 8672
rect 11203 8631 11261 8632
rect 11787 8672 11829 8681
rect 11787 8632 11788 8672
rect 11828 8632 11829 8672
rect 11787 8623 11829 8632
rect 12067 8672 12125 8673
rect 12067 8632 12076 8672
rect 12116 8632 12125 8672
rect 12067 8631 12125 8632
rect 12451 8672 12509 8673
rect 12451 8632 12460 8672
rect 12500 8632 12509 8672
rect 12451 8631 12509 8632
rect 12747 8672 12789 8681
rect 14659 8674 14668 8714
rect 14708 8674 14717 8714
rect 18123 8707 18165 8716
rect 18411 8691 18453 8700
rect 14659 8673 14717 8674
rect 12747 8632 12748 8672
rect 12788 8632 12789 8672
rect 12747 8623 12789 8632
rect 13411 8672 13469 8673
rect 13411 8632 13420 8672
rect 13460 8632 13469 8672
rect 13411 8631 13469 8632
rect 15043 8672 15101 8673
rect 15043 8632 15052 8672
rect 15092 8632 15101 8672
rect 15043 8631 15101 8632
rect 15331 8672 15389 8673
rect 15331 8632 15340 8672
rect 15380 8632 15389 8672
rect 15331 8631 15389 8632
rect 16579 8672 16637 8673
rect 16579 8632 16588 8672
rect 16628 8632 16637 8672
rect 16579 8631 16637 8632
rect 17155 8672 17213 8673
rect 17155 8632 17164 8672
rect 17204 8632 17213 8672
rect 17155 8631 17213 8632
rect 17451 8672 17493 8681
rect 17451 8632 17452 8672
rect 17492 8632 17493 8672
rect 17451 8623 17493 8632
rect 18019 8672 18077 8673
rect 18019 8632 18028 8672
rect 18068 8632 18077 8672
rect 18411 8651 18412 8691
rect 18452 8651 18453 8691
rect 18411 8642 18453 8651
rect 18507 8691 18549 8700
rect 18507 8651 18508 8691
rect 18548 8651 18549 8691
rect 19947 8686 19989 8695
rect 18507 8642 18549 8651
rect 18891 8672 18933 8681
rect 18019 8631 18077 8632
rect 18891 8632 18892 8672
rect 18932 8632 18933 8672
rect 18891 8623 18933 8632
rect 18987 8672 19029 8681
rect 18987 8632 18988 8672
rect 19028 8632 19029 8672
rect 18987 8623 19029 8632
rect 19459 8672 19517 8673
rect 19459 8632 19468 8672
rect 19508 8632 19517 8672
rect 19947 8646 19948 8686
rect 19988 8646 19989 8686
rect 19947 8637 19989 8646
rect 19459 8631 19517 8632
rect 6027 8588 6069 8597
rect 6027 8548 6028 8588
rect 6068 8548 6069 8588
rect 6027 8539 6069 8548
rect 9963 8588 10005 8597
rect 9963 8548 9964 8588
rect 10004 8548 10005 8588
rect 9963 8539 10005 8548
rect 11691 8588 11733 8597
rect 11691 8548 11692 8588
rect 11732 8548 11733 8588
rect 11691 8539 11733 8548
rect 12843 8588 12885 8597
rect 12843 8548 12844 8588
rect 12884 8548 12885 8588
rect 12843 8539 12885 8548
rect 17547 8588 17589 8597
rect 17547 8548 17548 8588
rect 17588 8548 17589 8588
rect 17547 8539 17589 8548
rect 2667 8504 2709 8513
rect 2667 8464 2668 8504
rect 2708 8464 2709 8504
rect 2667 8455 2709 8464
rect 3051 8504 3093 8513
rect 3051 8464 3052 8504
rect 3092 8464 3093 8504
rect 3051 8455 3093 8464
rect 8331 8504 8373 8513
rect 8331 8464 8332 8504
rect 8372 8464 8373 8504
rect 8331 8455 8373 8464
rect 14859 8504 14901 8513
rect 14859 8464 14860 8504
rect 14900 8464 14901 8504
rect 14859 8455 14901 8464
rect 15147 8504 15189 8513
rect 15147 8464 15148 8504
rect 15188 8464 15189 8504
rect 15147 8455 15189 8464
rect 20139 8504 20181 8513
rect 20139 8464 20140 8504
rect 20180 8464 20181 8504
rect 20139 8455 20181 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 2955 8168 2997 8177
rect 2955 8128 2956 8168
rect 2996 8128 2997 8168
rect 2955 8119 2997 8128
rect 5155 8168 5213 8169
rect 5155 8128 5164 8168
rect 5204 8128 5213 8168
rect 12747 8168 12789 8177
rect 5155 8127 5213 8128
rect 5835 8126 5877 8135
rect 2667 8084 2709 8093
rect 2667 8044 2668 8084
rect 2708 8044 2709 8084
rect 5835 8086 5836 8126
rect 5876 8086 5877 8126
rect 12747 8128 12748 8168
rect 12788 8128 12789 8168
rect 12747 8119 12789 8128
rect 14091 8168 14133 8177
rect 14091 8128 14092 8168
rect 14132 8128 14133 8168
rect 14091 8119 14133 8128
rect 17643 8168 17685 8177
rect 17643 8128 17644 8168
rect 17684 8128 17685 8168
rect 17643 8119 17685 8128
rect 18403 8168 18461 8169
rect 18403 8128 18412 8168
rect 18452 8128 18461 8168
rect 18403 8127 18461 8128
rect 5835 8077 5877 8086
rect 11883 8084 11925 8093
rect 2667 8035 2709 8044
rect 11883 8044 11884 8084
rect 11924 8044 11925 8084
rect 9667 8042 9725 8043
rect 1219 8000 1277 8001
rect 1219 7960 1228 8000
rect 1268 7960 1277 8000
rect 1219 7959 1277 7960
rect 2467 8000 2525 8001
rect 2467 7960 2476 8000
rect 2516 7960 2525 8000
rect 3619 8000 3677 8001
rect 2467 7959 2525 7960
rect 3099 7990 3141 7999
rect 3099 7950 3100 7990
rect 3140 7950 3141 7990
rect 3619 7960 3628 8000
rect 3668 7960 3677 8000
rect 3619 7959 3677 7960
rect 4587 8000 4629 8009
rect 4587 7960 4588 8000
rect 4628 7960 4629 8000
rect 4587 7951 4629 7960
rect 4683 8000 4725 8009
rect 4683 7960 4684 8000
rect 4724 7960 4725 8000
rect 4683 7951 4725 7960
rect 4963 8000 5021 8001
rect 4963 7960 4972 8000
rect 5012 7960 5021 8000
rect 4963 7959 5021 7960
rect 5059 8000 5117 8001
rect 5059 7960 5068 8000
rect 5108 7960 5117 8000
rect 5059 7959 5117 7960
rect 5259 8000 5301 8009
rect 5259 7960 5260 8000
rect 5300 7960 5301 8000
rect 5259 7951 5301 7960
rect 5355 8000 5397 8009
rect 5355 7960 5356 8000
rect 5396 7960 5397 8000
rect 5355 7951 5397 7960
rect 5448 8000 5506 8001
rect 5448 7960 5457 8000
rect 5497 7960 5506 8000
rect 6499 8000 6557 8001
rect 5448 7959 5506 7960
rect 5979 7990 6021 7999
rect 3099 7941 3141 7950
rect 5979 7950 5980 7990
rect 6020 7950 6021 7990
rect 6499 7960 6508 8000
rect 6548 7960 6557 8000
rect 6499 7959 6557 7960
rect 6987 8000 7029 8009
rect 6987 7960 6988 8000
rect 7028 7960 7029 8000
rect 6987 7951 7029 7960
rect 7083 8000 7125 8009
rect 7083 7960 7084 8000
rect 7124 7960 7125 8000
rect 7083 7951 7125 7960
rect 7467 8000 7509 8009
rect 7467 7960 7468 8000
rect 7508 7960 7509 8000
rect 7467 7951 7509 7960
rect 7563 8000 7605 8009
rect 9667 8002 9676 8042
rect 9716 8002 9725 8042
rect 11883 8035 11925 8044
rect 14955 8084 14997 8093
rect 14955 8044 14956 8084
rect 14996 8044 14997 8084
rect 14955 8035 14997 8044
rect 16875 8084 16917 8093
rect 16875 8044 16876 8084
rect 16916 8044 16917 8084
rect 16875 8035 16917 8044
rect 9667 8001 9725 8002
rect 7563 7960 7564 8000
rect 7604 7960 7605 8000
rect 7563 7951 7605 7960
rect 8035 8000 8093 8001
rect 8035 7960 8044 8000
rect 8084 7960 8093 8000
rect 8035 7959 8093 7960
rect 9283 8000 9341 8001
rect 9283 7960 9292 8000
rect 9332 7960 9341 8000
rect 9283 7959 9341 7960
rect 10059 8000 10101 8009
rect 10059 7960 10060 8000
rect 10100 7960 10101 8000
rect 10059 7951 10101 7960
rect 10435 8000 10493 8001
rect 10435 7960 10444 8000
rect 10484 7960 10493 8000
rect 10435 7959 10493 7960
rect 11683 8000 11741 8001
rect 11683 7960 11692 8000
rect 11732 7960 11741 8000
rect 11683 7959 11741 7960
rect 12067 8000 12125 8001
rect 12067 7960 12076 8000
rect 12116 7960 12125 8000
rect 12067 7959 12125 7960
rect 12267 8000 12309 8009
rect 12267 7960 12268 8000
rect 12308 7960 12309 8000
rect 12267 7951 12309 7960
rect 12355 8000 12413 8001
rect 12355 7960 12364 8000
rect 12404 7960 12413 8000
rect 12355 7959 12413 7960
rect 12651 8000 12693 8009
rect 12651 7960 12652 8000
rect 12692 7960 12693 8000
rect 12651 7951 12693 7960
rect 12843 8000 12885 8009
rect 12843 7960 12844 8000
rect 12884 7960 12885 8000
rect 12843 7951 12885 7960
rect 13035 8000 13077 8009
rect 13035 7960 13036 8000
rect 13076 7960 13077 8000
rect 13035 7951 13077 7960
rect 13323 8000 13365 8009
rect 13323 7960 13324 8000
rect 13364 7960 13365 8000
rect 13323 7951 13365 7960
rect 13515 8000 13557 8009
rect 13515 7960 13516 8000
rect 13556 7960 13557 8000
rect 13515 7951 13557 7960
rect 13611 8000 13653 8009
rect 13611 7960 13612 8000
rect 13652 7960 13653 8000
rect 13611 7951 13653 7960
rect 13707 8000 13749 8009
rect 13707 7960 13708 8000
rect 13748 7960 13749 8000
rect 13707 7951 13749 7960
rect 13803 8000 13845 8009
rect 13803 7960 13804 8000
rect 13844 7960 13845 8000
rect 13803 7951 13845 7960
rect 13995 8000 14037 8009
rect 13995 7960 13996 8000
rect 14036 7960 14037 8000
rect 13995 7951 14037 7960
rect 14187 8000 14229 8009
rect 14187 7960 14188 8000
rect 14228 7960 14229 8000
rect 14187 7951 14229 7960
rect 14563 8000 14621 8001
rect 14563 7960 14572 8000
rect 14612 7960 14621 8000
rect 14563 7959 14621 7960
rect 14859 8000 14901 8009
rect 14859 7960 14860 8000
rect 14900 7960 14901 8000
rect 14859 7951 14901 7960
rect 15427 8000 15485 8001
rect 15427 7960 15436 8000
rect 15476 7960 15485 8000
rect 15427 7959 15485 7960
rect 16675 8000 16733 8001
rect 16675 7960 16684 8000
rect 16724 7960 16733 8000
rect 16675 7959 16733 7960
rect 17059 8000 17117 8001
rect 17059 7960 17068 8000
rect 17108 7960 17117 8000
rect 17059 7959 17117 7960
rect 17163 8000 17205 8009
rect 17163 7960 17164 8000
rect 17204 7960 17205 8000
rect 17163 7951 17205 7960
rect 17347 8000 17405 8001
rect 17347 7960 17356 8000
rect 17396 7960 17405 8000
rect 17347 7959 17405 7960
rect 17547 8000 17589 8009
rect 17547 7960 17548 8000
rect 17588 7960 17589 8000
rect 17547 7951 17589 7960
rect 17739 8000 17781 8009
rect 17739 7960 17740 8000
rect 17780 7960 17781 8000
rect 17739 7951 17781 7960
rect 18507 8000 18549 8009
rect 18507 7960 18508 8000
rect 18548 7960 18549 8000
rect 18507 7951 18549 7960
rect 18603 8000 18645 8009
rect 18603 7960 18604 8000
rect 18644 7960 18645 8000
rect 18603 7951 18645 7960
rect 18699 8000 18741 8009
rect 18699 7960 18700 8000
rect 18740 7960 18741 8000
rect 18699 7951 18741 7960
rect 18883 8000 18941 8001
rect 18883 7960 18892 8000
rect 18932 7960 18941 8000
rect 18883 7959 18941 7960
rect 19275 8000 19317 8009
rect 19275 7960 19276 8000
rect 19316 7960 19317 8000
rect 19275 7951 19317 7960
rect 19459 8000 19517 8001
rect 19459 7960 19468 8000
rect 19508 7960 19517 8000
rect 19459 7959 19517 7960
rect 19851 8000 19893 8009
rect 19851 7960 19852 8000
rect 19892 7960 19893 8000
rect 19851 7951 19893 7960
rect 20043 8000 20085 8009
rect 20043 7960 20044 8000
rect 20084 7960 20085 8000
rect 20043 7951 20085 7960
rect 20235 8000 20277 8009
rect 20235 7960 20236 8000
rect 20276 7960 20277 8000
rect 20235 7951 20277 7960
rect 5979 7941 6021 7950
rect 4107 7916 4149 7925
rect 4107 7876 4108 7916
rect 4148 7876 4149 7916
rect 4107 7867 4149 7876
rect 4203 7916 4245 7925
rect 4203 7876 4204 7916
rect 4244 7876 4245 7916
rect 4203 7867 4245 7876
rect 9771 7916 9813 7925
rect 9771 7876 9772 7916
rect 9812 7876 9813 7916
rect 9771 7867 9813 7876
rect 9963 7916 10005 7925
rect 9963 7876 9964 7916
rect 10004 7876 10005 7916
rect 9963 7867 10005 7876
rect 18019 7916 18077 7917
rect 18019 7876 18028 7916
rect 18068 7876 18077 7916
rect 18019 7875 18077 7876
rect 18987 7916 19029 7925
rect 18987 7876 18988 7916
rect 19028 7876 19029 7916
rect 18987 7867 19029 7876
rect 19179 7916 19221 7925
rect 19179 7876 19180 7916
rect 19220 7876 19221 7916
rect 19179 7867 19221 7876
rect 19563 7916 19605 7925
rect 19563 7876 19564 7916
rect 19604 7876 19605 7916
rect 19563 7867 19605 7876
rect 19755 7916 19797 7925
rect 19755 7876 19756 7916
rect 19796 7876 19797 7916
rect 19755 7867 19797 7876
rect 9483 7832 9525 7841
rect 9483 7792 9484 7832
rect 9524 7792 9525 7832
rect 9483 7783 9525 7792
rect 9867 7832 9909 7841
rect 9867 7792 9868 7832
rect 9908 7792 9909 7832
rect 9867 7783 9909 7792
rect 12259 7832 12317 7833
rect 12259 7792 12268 7832
rect 12308 7792 12317 7832
rect 12259 7791 12317 7792
rect 17155 7832 17213 7833
rect 17155 7792 17164 7832
rect 17204 7792 17213 7832
rect 17155 7791 17213 7792
rect 19083 7832 19125 7841
rect 19083 7792 19084 7832
rect 19124 7792 19125 7832
rect 19083 7783 19125 7792
rect 19659 7832 19701 7841
rect 19659 7792 19660 7832
rect 19700 7792 19701 7832
rect 19659 7783 19701 7792
rect 20235 7832 20277 7841
rect 20235 7792 20236 7832
rect 20276 7792 20277 7832
rect 20235 7783 20277 7792
rect 13323 7748 13365 7757
rect 13323 7708 13324 7748
rect 13364 7708 13365 7748
rect 13323 7699 13365 7708
rect 15235 7748 15293 7749
rect 15235 7708 15244 7748
rect 15284 7708 15293 7748
rect 15235 7707 15293 7708
rect 18219 7748 18261 7757
rect 18219 7708 18220 7748
rect 18260 7708 18261 7748
rect 18219 7699 18261 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 3627 7412 3669 7421
rect 3627 7372 3628 7412
rect 3668 7372 3669 7412
rect 3627 7363 3669 7372
rect 5643 7412 5685 7421
rect 5643 7372 5644 7412
rect 5684 7372 5685 7412
rect 5643 7363 5685 7372
rect 5835 7412 5877 7421
rect 5835 7372 5836 7412
rect 5876 7372 5877 7412
rect 5835 7363 5877 7372
rect 13995 7412 14037 7421
rect 13995 7372 13996 7412
rect 14036 7372 14037 7412
rect 13995 7363 14037 7372
rect 14667 7412 14709 7421
rect 14667 7372 14668 7412
rect 14708 7372 14709 7412
rect 14667 7363 14709 7372
rect 17451 7412 17493 7421
rect 17451 7372 17452 7412
rect 17492 7372 17493 7412
rect 17451 7363 17493 7372
rect 19275 7412 19317 7421
rect 19275 7372 19276 7412
rect 19316 7372 19317 7412
rect 19275 7363 19317 7372
rect 8139 7328 8181 7337
rect 8139 7288 8140 7328
rect 8180 7288 8181 7328
rect 15043 7328 15101 7329
rect 8139 7279 8181 7288
rect 8331 7302 8373 7311
rect 8331 7262 8332 7302
rect 8372 7262 8373 7302
rect 15043 7288 15052 7328
rect 15092 7288 15101 7328
rect 15043 7287 15101 7288
rect 15627 7328 15669 7337
rect 15627 7288 15628 7328
rect 15668 7288 15669 7328
rect 15627 7279 15669 7288
rect 8331 7253 8373 7262
rect 9483 7244 9525 7253
rect 9483 7204 9484 7244
rect 9524 7204 9525 7244
rect 9483 7195 9525 7204
rect 9579 7244 9621 7253
rect 9579 7204 9580 7244
rect 9620 7204 9621 7244
rect 9579 7195 9621 7204
rect 11107 7244 11165 7245
rect 11107 7204 11116 7244
rect 11156 7204 11165 7244
rect 11107 7203 11165 7204
rect 11491 7244 11549 7245
rect 11491 7204 11500 7244
rect 11540 7204 11549 7244
rect 11491 7203 11549 7204
rect 15531 7244 15573 7253
rect 15531 7204 15532 7244
rect 15572 7204 15573 7244
rect 15531 7195 15573 7204
rect 15723 7244 15765 7253
rect 15723 7204 15724 7244
rect 15764 7204 15765 7244
rect 15723 7195 15765 7204
rect 1227 7160 1269 7169
rect 1227 7120 1228 7160
rect 1268 7120 1269 7160
rect 1227 7111 1269 7120
rect 1419 7160 1461 7169
rect 1419 7120 1420 7160
rect 1460 7120 1461 7160
rect 1419 7111 1461 7120
rect 1507 7160 1565 7161
rect 1507 7120 1516 7160
rect 1556 7120 1565 7160
rect 1507 7119 1565 7120
rect 1707 7160 1749 7169
rect 1707 7120 1708 7160
rect 1748 7120 1749 7160
rect 1707 7111 1749 7120
rect 1803 7160 1845 7169
rect 1803 7120 1804 7160
rect 1844 7120 1845 7160
rect 1803 7111 1845 7120
rect 1899 7160 1941 7169
rect 1899 7120 1900 7160
rect 1940 7120 1941 7160
rect 1899 7111 1941 7120
rect 1995 7160 2037 7169
rect 1995 7120 1996 7160
rect 2036 7120 2037 7160
rect 1995 7111 2037 7120
rect 2179 7160 2237 7161
rect 2179 7120 2188 7160
rect 2228 7120 2237 7160
rect 2179 7119 2237 7120
rect 3427 7160 3485 7161
rect 3427 7120 3436 7160
rect 3476 7120 3485 7160
rect 3427 7119 3485 7120
rect 3819 7160 3861 7169
rect 3819 7120 3820 7160
rect 3860 7120 3861 7160
rect 3819 7111 3861 7120
rect 4011 7160 4053 7169
rect 4011 7120 4012 7160
rect 4052 7120 4053 7160
rect 4011 7111 4053 7120
rect 4195 7160 4253 7161
rect 4195 7120 4204 7160
rect 4244 7120 4253 7160
rect 4195 7119 4253 7120
rect 5443 7160 5501 7161
rect 5443 7120 5452 7160
rect 5492 7120 5501 7160
rect 5443 7119 5501 7120
rect 6019 7160 6077 7161
rect 6019 7120 6028 7160
rect 6068 7120 6077 7160
rect 6019 7119 6077 7120
rect 7267 7160 7325 7161
rect 7267 7120 7276 7160
rect 7316 7120 7325 7160
rect 7267 7119 7325 7120
rect 7659 7160 7701 7169
rect 7659 7120 7660 7160
rect 7700 7120 7701 7160
rect 7659 7111 7701 7120
rect 7755 7160 7797 7169
rect 7755 7120 7756 7160
rect 7796 7120 7797 7160
rect 7755 7111 7797 7120
rect 7851 7160 7893 7169
rect 7851 7120 7852 7160
rect 7892 7120 7893 7160
rect 7851 7111 7893 7120
rect 7947 7160 7989 7169
rect 7947 7120 7948 7160
rect 7988 7120 7989 7160
rect 7947 7111 7989 7120
rect 8331 7152 8373 7161
rect 8331 7112 8332 7152
rect 8372 7112 8373 7152
rect 8707 7160 8765 7161
rect 8707 7120 8716 7160
rect 8756 7120 8765 7160
rect 8707 7119 8765 7120
rect 9003 7160 9045 7169
rect 9003 7120 9004 7160
rect 9044 7120 9045 7160
rect 8331 7103 8373 7112
rect 9003 7111 9045 7120
rect 9099 7160 9141 7169
rect 10539 7165 10581 7174
rect 9099 7120 9100 7160
rect 9140 7120 9141 7160
rect 9099 7111 9141 7120
rect 10051 7160 10109 7161
rect 10051 7120 10060 7160
rect 10100 7120 10109 7160
rect 10051 7119 10109 7120
rect 10539 7125 10540 7165
rect 10580 7125 10581 7165
rect 10539 7116 10581 7125
rect 11779 7160 11837 7161
rect 11779 7120 11788 7160
rect 11828 7120 11837 7160
rect 11779 7119 11837 7120
rect 12075 7160 12117 7169
rect 12075 7120 12076 7160
rect 12116 7120 12117 7160
rect 12075 7111 12117 7120
rect 12171 7160 12213 7169
rect 12171 7120 12172 7160
rect 12212 7120 12213 7160
rect 12171 7111 12213 7120
rect 12555 7160 12597 7169
rect 12555 7120 12556 7160
rect 12596 7120 12597 7160
rect 12555 7111 12597 7120
rect 12651 7160 12693 7169
rect 13611 7165 13653 7174
rect 12651 7120 12652 7160
rect 12692 7120 12693 7160
rect 12651 7111 12693 7120
rect 13123 7160 13181 7161
rect 13123 7120 13132 7160
rect 13172 7120 13181 7160
rect 13123 7119 13181 7120
rect 13611 7125 13612 7165
rect 13652 7125 13653 7165
rect 13611 7116 13653 7125
rect 13995 7160 14037 7169
rect 13995 7120 13996 7160
rect 14036 7120 14037 7160
rect 13995 7111 14037 7120
rect 14187 7160 14229 7169
rect 14187 7120 14188 7160
rect 14228 7120 14229 7160
rect 14187 7111 14229 7120
rect 14275 7160 14333 7161
rect 14275 7120 14284 7160
rect 14324 7120 14333 7160
rect 14275 7119 14333 7120
rect 14475 7160 14517 7169
rect 14475 7120 14476 7160
rect 14516 7120 14517 7160
rect 14475 7111 14517 7120
rect 14667 7160 14709 7169
rect 14667 7120 14668 7160
rect 14708 7120 14709 7160
rect 14667 7111 14709 7120
rect 14947 7160 15005 7161
rect 14947 7120 14956 7160
rect 14996 7120 15005 7160
rect 14947 7119 15005 7120
rect 15051 7160 15093 7169
rect 15051 7120 15052 7160
rect 15092 7120 15093 7160
rect 15051 7111 15093 7120
rect 15235 7160 15293 7161
rect 15235 7120 15244 7160
rect 15284 7120 15293 7160
rect 15235 7119 15293 7120
rect 15427 7160 15485 7161
rect 15427 7120 15436 7160
rect 15476 7120 15485 7160
rect 15427 7119 15485 7120
rect 15819 7160 15861 7169
rect 15819 7120 15820 7160
rect 15860 7120 15861 7160
rect 15819 7111 15861 7120
rect 16003 7160 16061 7161
rect 16003 7120 16012 7160
rect 16052 7120 16061 7160
rect 16003 7119 16061 7120
rect 17251 7160 17309 7161
rect 17251 7120 17260 7160
rect 17300 7120 17309 7160
rect 17251 7119 17309 7120
rect 17827 7160 17885 7161
rect 17827 7120 17836 7160
rect 17876 7120 17885 7160
rect 17827 7119 17885 7120
rect 19075 7160 19133 7161
rect 19075 7120 19084 7160
rect 19124 7120 19133 7160
rect 19075 7119 19133 7120
rect 19459 7160 19517 7161
rect 19459 7120 19468 7160
rect 19508 7120 19517 7160
rect 19459 7119 19517 7120
rect 19555 7160 19613 7161
rect 19555 7120 19564 7160
rect 19604 7120 19613 7160
rect 19555 7119 19613 7120
rect 19755 7160 19797 7169
rect 19755 7120 19756 7160
rect 19796 7120 19797 7160
rect 19755 7111 19797 7120
rect 19851 7160 19893 7169
rect 19851 7120 19852 7160
rect 19892 7120 19893 7160
rect 19851 7111 19893 7120
rect 19944 7160 20002 7161
rect 19944 7120 19953 7160
rect 19993 7120 20002 7160
rect 19944 7119 20002 7120
rect 1323 7076 1365 7085
rect 1323 7036 1324 7076
rect 1364 7036 1365 7076
rect 1323 7027 1365 7036
rect 8619 7076 8661 7085
rect 8619 7036 8620 7076
rect 8660 7036 8661 7076
rect 8619 7027 8661 7036
rect 3915 6992 3957 7001
rect 3915 6952 3916 6992
rect 3956 6952 3957 6992
rect 3915 6943 3957 6952
rect 10731 6992 10773 7001
rect 10731 6952 10732 6992
rect 10772 6952 10773 6992
rect 10731 6943 10773 6952
rect 10923 6992 10965 7001
rect 10923 6952 10924 6992
rect 10964 6952 10965 6992
rect 10923 6943 10965 6952
rect 11307 6992 11349 7001
rect 11307 6952 11308 6992
rect 11348 6952 11349 6992
rect 11307 6943 11349 6952
rect 11691 6992 11733 7001
rect 11691 6952 11692 6992
rect 11732 6952 11733 6992
rect 11691 6943 11733 6952
rect 13803 6992 13845 7001
rect 13803 6952 13804 6992
rect 13844 6952 13845 6992
rect 13803 6943 13845 6952
rect 19651 6992 19709 6993
rect 19651 6952 19660 6992
rect 19700 6952 19709 6992
rect 19651 6951 19709 6952
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 1603 6656 1661 6657
rect 1603 6616 1612 6656
rect 1652 6616 1661 6656
rect 1603 6615 1661 6616
rect 2371 6656 2429 6657
rect 2371 6616 2380 6656
rect 2420 6616 2429 6656
rect 2371 6615 2429 6616
rect 2571 6656 2613 6665
rect 2571 6616 2572 6656
rect 2612 6616 2613 6656
rect 2571 6607 2613 6616
rect 6027 6656 6069 6665
rect 6027 6616 6028 6656
rect 6068 6616 6069 6656
rect 6027 6607 6069 6616
rect 10251 6656 10293 6665
rect 10251 6616 10252 6656
rect 10292 6616 10293 6656
rect 10251 6607 10293 6616
rect 11883 6656 11925 6665
rect 11883 6616 11884 6656
rect 11924 6616 11925 6656
rect 11883 6607 11925 6616
rect 13515 6656 13557 6665
rect 13515 6616 13516 6656
rect 13556 6616 13557 6656
rect 13515 6607 13557 6616
rect 14379 6656 14421 6665
rect 14379 6616 14380 6656
rect 14420 6616 14421 6656
rect 14379 6607 14421 6616
rect 16107 6656 16149 6665
rect 16107 6616 16108 6656
rect 16148 6616 16149 6656
rect 16107 6607 16149 6616
rect 17259 6614 17301 6623
rect 6411 6572 6453 6581
rect 6411 6532 6412 6572
rect 6452 6532 6453 6572
rect 17259 6574 17260 6614
rect 17300 6574 17301 6614
rect 17259 6565 17301 6574
rect 6411 6523 6453 6532
rect 1896 6497 1954 6498
rect 1227 6488 1269 6497
rect 1227 6448 1228 6488
rect 1268 6448 1269 6488
rect 1227 6439 1269 6448
rect 1419 6488 1461 6497
rect 1419 6448 1420 6488
rect 1460 6448 1461 6488
rect 1419 6439 1461 6448
rect 1803 6488 1845 6497
rect 1803 6448 1804 6488
rect 1844 6448 1845 6488
rect 1896 6457 1905 6497
rect 1945 6457 1954 6497
rect 1896 6456 1954 6457
rect 2091 6488 2133 6497
rect 1803 6439 1845 6448
rect 2091 6448 2092 6488
rect 2132 6448 2133 6488
rect 2091 6439 2133 6448
rect 2187 6488 2229 6497
rect 2187 6448 2188 6488
rect 2228 6448 2229 6488
rect 2187 6439 2229 6448
rect 2763 6483 2805 6492
rect 2763 6443 2764 6483
rect 2804 6443 2805 6483
rect 3235 6488 3293 6489
rect 3235 6448 3244 6488
rect 3284 6448 3293 6488
rect 3235 6447 3293 6448
rect 3723 6488 3765 6497
rect 3723 6448 3724 6488
rect 3764 6448 3765 6488
rect 2763 6434 2805 6443
rect 3723 6439 3765 6448
rect 3819 6488 3861 6497
rect 3819 6448 3820 6488
rect 3860 6448 3861 6488
rect 3819 6439 3861 6448
rect 4203 6488 4245 6497
rect 4203 6448 4204 6488
rect 4244 6448 4245 6488
rect 4203 6439 4245 6448
rect 4299 6488 4341 6497
rect 4299 6448 4300 6488
rect 4340 6448 4341 6488
rect 4299 6439 4341 6448
rect 4579 6488 4637 6489
rect 4579 6448 4588 6488
rect 4628 6448 4637 6488
rect 4579 6447 4637 6448
rect 5827 6488 5885 6489
rect 5827 6448 5836 6488
rect 5876 6448 5885 6488
rect 7075 6488 7133 6489
rect 5827 6447 5885 6448
rect 6603 6474 6645 6483
rect 6603 6434 6604 6474
rect 6644 6434 6645 6474
rect 7075 6448 7084 6488
rect 7124 6448 7133 6488
rect 7075 6447 7133 6448
rect 7563 6488 7605 6497
rect 7563 6448 7564 6488
rect 7604 6448 7605 6488
rect 7563 6439 7605 6448
rect 8043 6488 8085 6497
rect 8043 6448 8044 6488
rect 8084 6448 8085 6488
rect 8043 6439 8085 6448
rect 8139 6488 8181 6497
rect 8139 6448 8140 6488
rect 8180 6448 8181 6488
rect 8139 6439 8181 6448
rect 8427 6488 8469 6497
rect 8427 6448 8428 6488
rect 8468 6448 8469 6488
rect 8427 6439 8469 6448
rect 8619 6488 8661 6497
rect 8619 6448 8620 6488
rect 8660 6448 8661 6488
rect 8619 6439 8661 6448
rect 8803 6488 8861 6489
rect 8803 6448 8812 6488
rect 8852 6448 8861 6488
rect 8803 6447 8861 6448
rect 10051 6488 10109 6489
rect 10051 6448 10060 6488
rect 10100 6448 10109 6488
rect 10051 6447 10109 6448
rect 10435 6488 10493 6489
rect 10435 6448 10444 6488
rect 10484 6448 10493 6488
rect 10435 6447 10493 6448
rect 11683 6488 11741 6489
rect 11683 6448 11692 6488
rect 11732 6448 11741 6488
rect 11683 6447 11741 6448
rect 13315 6488 13373 6489
rect 13315 6448 13324 6488
rect 13364 6448 13373 6488
rect 13315 6447 13373 6448
rect 13707 6488 13749 6497
rect 13707 6448 13708 6488
rect 13748 6448 13749 6488
rect 12067 6446 12125 6447
rect 6603 6425 6645 6434
rect 7659 6404 7701 6413
rect 12067 6406 12076 6446
rect 12116 6406 12125 6446
rect 13707 6439 13749 6448
rect 13899 6488 13941 6497
rect 13899 6448 13900 6488
rect 13940 6448 13941 6488
rect 13899 6439 13941 6448
rect 13987 6488 14045 6489
rect 13987 6448 13996 6488
rect 14036 6448 14045 6488
rect 13987 6447 14045 6448
rect 14283 6488 14325 6497
rect 14283 6448 14284 6488
rect 14324 6448 14325 6488
rect 14283 6439 14325 6448
rect 14475 6488 14517 6497
rect 14475 6448 14476 6488
rect 14516 6448 14517 6488
rect 14475 6439 14517 6448
rect 14659 6488 14717 6489
rect 14659 6448 14668 6488
rect 14708 6448 14717 6488
rect 14659 6447 14717 6448
rect 15907 6488 15965 6489
rect 15907 6448 15916 6488
rect 15956 6448 15965 6488
rect 15907 6447 15965 6448
rect 16291 6488 16349 6489
rect 16291 6448 16300 6488
rect 16340 6448 16349 6488
rect 16291 6447 16349 6448
rect 16387 6488 16445 6489
rect 16387 6448 16396 6488
rect 16436 6448 16445 6488
rect 16387 6447 16445 6448
rect 16587 6488 16629 6497
rect 16587 6448 16588 6488
rect 16628 6448 16629 6488
rect 16587 6439 16629 6448
rect 16683 6488 16725 6497
rect 17067 6488 17109 6497
rect 16683 6448 16684 6488
rect 16724 6448 16725 6488
rect 16683 6439 16725 6448
rect 16819 6487 16877 6488
rect 16819 6447 16828 6487
rect 16868 6447 16877 6487
rect 16819 6446 16877 6447
rect 17067 6448 17068 6488
rect 17108 6448 17109 6488
rect 17067 6439 17109 6448
rect 17443 6488 17501 6489
rect 17443 6448 17452 6488
rect 17492 6448 17501 6488
rect 17443 6447 17501 6448
rect 17731 6488 17789 6489
rect 17731 6448 17740 6488
rect 17780 6448 17789 6488
rect 17731 6447 17789 6448
rect 18979 6488 19037 6489
rect 18979 6448 18988 6488
rect 19028 6448 19037 6488
rect 18979 6447 19037 6448
rect 19659 6488 19701 6497
rect 19659 6448 19660 6488
rect 19700 6448 19701 6488
rect 19659 6439 19701 6448
rect 19755 6488 19797 6497
rect 19755 6448 19756 6488
rect 19796 6448 19797 6488
rect 19755 6439 19797 6448
rect 20035 6488 20093 6489
rect 20035 6448 20044 6488
rect 20084 6448 20093 6488
rect 20035 6447 20093 6448
rect 12067 6405 12125 6406
rect 7659 6364 7660 6404
rect 7700 6364 7701 6404
rect 7659 6355 7701 6364
rect 17163 6404 17205 6413
rect 17163 6364 17164 6404
rect 17204 6364 17205 6404
rect 17163 6355 17205 6364
rect 17355 6404 17397 6413
rect 17355 6364 17356 6404
rect 17396 6364 17397 6404
rect 17355 6355 17397 6364
rect 8619 6320 8661 6329
rect 8619 6280 8620 6320
rect 8660 6280 8661 6320
rect 8619 6271 8661 6280
rect 19363 6320 19421 6321
rect 19363 6280 19372 6320
rect 19412 6280 19421 6320
rect 19363 6279 19421 6280
rect 1419 6236 1461 6245
rect 1419 6196 1420 6236
rect 1460 6196 1461 6236
rect 1419 6187 1461 6196
rect 13707 6236 13749 6245
rect 13707 6196 13708 6236
rect 13748 6196 13749 6236
rect 13707 6187 13749 6196
rect 16299 6236 16341 6245
rect 16299 6196 16300 6236
rect 16340 6196 16341 6236
rect 16299 6187 16341 6196
rect 19179 6236 19221 6245
rect 19179 6196 19180 6236
rect 19220 6196 19221 6236
rect 19179 6187 19221 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 2763 5900 2805 5909
rect 2763 5860 2764 5900
rect 2804 5860 2805 5900
rect 2763 5851 2805 5860
rect 5931 5900 5973 5909
rect 5931 5860 5932 5900
rect 5972 5860 5973 5900
rect 5931 5851 5973 5860
rect 7563 5900 7605 5909
rect 7563 5860 7564 5900
rect 7604 5860 7605 5900
rect 7563 5851 7605 5860
rect 11883 5900 11925 5909
rect 11883 5860 11884 5900
rect 11924 5860 11925 5900
rect 11883 5851 11925 5860
rect 15531 5900 15573 5909
rect 15531 5860 15532 5900
rect 15572 5860 15573 5900
rect 15531 5851 15573 5860
rect 16867 5900 16925 5901
rect 16867 5860 16876 5900
rect 16916 5860 16925 5900
rect 16867 5859 16925 5860
rect 19843 5900 19901 5901
rect 19843 5860 19852 5900
rect 19892 5860 19901 5900
rect 19843 5859 19901 5860
rect 20235 5900 20277 5909
rect 20235 5860 20236 5900
rect 20276 5860 20277 5900
rect 20235 5851 20277 5860
rect 1803 5816 1845 5825
rect 1803 5776 1804 5816
rect 1844 5776 1845 5816
rect 1803 5767 1845 5776
rect 2379 5816 2421 5825
rect 2379 5776 2380 5816
rect 2420 5776 2421 5816
rect 2379 5767 2421 5776
rect 9867 5816 9909 5825
rect 9867 5776 9868 5816
rect 9908 5776 9909 5816
rect 9867 5767 9909 5776
rect 2283 5732 2325 5741
rect 2283 5692 2284 5732
rect 2324 5692 2325 5732
rect 2283 5683 2325 5692
rect 2475 5732 2517 5741
rect 2475 5692 2476 5732
rect 2516 5692 2517 5732
rect 2475 5683 2517 5692
rect 8907 5732 8949 5741
rect 8907 5692 8908 5732
rect 8948 5692 8949 5732
rect 8907 5683 8949 5692
rect 9003 5732 9045 5741
rect 9003 5692 9004 5732
rect 9044 5692 9045 5732
rect 9003 5683 9045 5692
rect 10051 5732 10109 5733
rect 10051 5692 10060 5732
rect 10100 5692 10109 5732
rect 10051 5691 10109 5692
rect 13515 5732 13557 5741
rect 13515 5692 13516 5732
rect 13556 5692 13557 5732
rect 13515 5683 13557 5692
rect 17163 5732 17205 5741
rect 17163 5692 17164 5732
rect 17204 5692 17205 5732
rect 17163 5683 17205 5692
rect 1219 5648 1277 5649
rect 1219 5608 1228 5648
rect 1268 5608 1277 5648
rect 1219 5607 1277 5608
rect 1323 5648 1365 5657
rect 1323 5608 1324 5648
rect 1364 5608 1365 5648
rect 1323 5599 1365 5608
rect 1515 5648 1557 5657
rect 1515 5608 1516 5648
rect 1556 5608 1557 5648
rect 1515 5599 1557 5608
rect 1707 5648 1749 5657
rect 1707 5608 1708 5648
rect 1748 5608 1749 5648
rect 1707 5599 1749 5608
rect 1899 5648 1941 5657
rect 1899 5608 1900 5648
rect 1940 5608 1941 5648
rect 1899 5599 1941 5608
rect 1995 5648 2037 5657
rect 1995 5608 1996 5648
rect 2036 5608 2037 5648
rect 1995 5599 2037 5608
rect 2187 5648 2229 5657
rect 7947 5653 7989 5662
rect 2187 5608 2188 5648
rect 2228 5608 2229 5648
rect 2187 5599 2229 5608
rect 2563 5648 2621 5649
rect 2563 5608 2572 5648
rect 2612 5608 2621 5648
rect 2563 5607 2621 5608
rect 2947 5648 3005 5649
rect 2947 5608 2956 5648
rect 2996 5608 3005 5648
rect 2947 5607 3005 5608
rect 4195 5648 4253 5649
rect 4195 5608 4204 5648
rect 4244 5608 4253 5648
rect 4195 5607 4253 5608
rect 4483 5648 4541 5649
rect 4483 5608 4492 5648
rect 4532 5608 4541 5648
rect 4483 5607 4541 5608
rect 5731 5648 5789 5649
rect 5731 5608 5740 5648
rect 5780 5608 5789 5648
rect 5731 5607 5789 5608
rect 6115 5648 6173 5649
rect 6115 5608 6124 5648
rect 6164 5608 6173 5648
rect 6115 5607 6173 5608
rect 7363 5648 7421 5649
rect 7363 5608 7372 5648
rect 7412 5608 7421 5648
rect 7363 5607 7421 5608
rect 7947 5613 7948 5653
rect 7988 5613 7989 5653
rect 7947 5604 7989 5613
rect 8419 5648 8477 5649
rect 8419 5608 8428 5648
rect 8468 5608 8477 5648
rect 8419 5607 8477 5608
rect 9387 5648 9429 5657
rect 9387 5608 9388 5648
rect 9428 5608 9429 5648
rect 9387 5599 9429 5608
rect 9483 5648 9525 5657
rect 9483 5608 9484 5648
rect 9524 5608 9525 5648
rect 9483 5599 9525 5608
rect 10435 5648 10493 5649
rect 10435 5608 10444 5648
rect 10484 5608 10493 5648
rect 10435 5607 10493 5608
rect 11683 5648 11741 5649
rect 11683 5608 11692 5648
rect 11732 5608 11741 5648
rect 11683 5607 11741 5608
rect 12363 5648 12405 5657
rect 12363 5608 12364 5648
rect 12404 5608 12405 5648
rect 12363 5599 12405 5608
rect 12459 5648 12501 5657
rect 12459 5608 12460 5648
rect 12500 5608 12501 5648
rect 12459 5599 12501 5608
rect 12555 5648 12597 5657
rect 12555 5608 12556 5648
rect 12596 5608 12597 5648
rect 12555 5599 12597 5608
rect 12939 5648 12981 5657
rect 12939 5608 12940 5648
rect 12980 5608 12981 5648
rect 12939 5599 12981 5608
rect 13035 5648 13077 5657
rect 13035 5608 13036 5648
rect 13076 5608 13077 5648
rect 13035 5599 13077 5608
rect 13131 5648 13173 5657
rect 13131 5608 13132 5648
rect 13172 5608 13173 5648
rect 13131 5599 13173 5608
rect 13227 5648 13269 5657
rect 13227 5608 13228 5648
rect 13268 5608 13269 5648
rect 13227 5599 13269 5608
rect 13419 5648 13461 5657
rect 13419 5608 13420 5648
rect 13460 5608 13461 5648
rect 13419 5599 13461 5608
rect 13611 5648 13653 5657
rect 13611 5608 13612 5648
rect 13652 5608 13653 5648
rect 13611 5599 13653 5608
rect 13891 5648 13949 5649
rect 13891 5608 13900 5648
rect 13940 5608 13949 5648
rect 13891 5607 13949 5608
rect 14083 5648 14141 5649
rect 14083 5608 14092 5648
rect 14132 5608 14141 5648
rect 14083 5607 14141 5608
rect 15331 5648 15389 5649
rect 15331 5608 15340 5648
rect 15380 5608 15389 5648
rect 15331 5607 15389 5608
rect 15723 5648 15765 5657
rect 15723 5608 15724 5648
rect 15764 5608 15765 5648
rect 15723 5599 15765 5608
rect 15915 5648 15957 5657
rect 15915 5608 15916 5648
rect 15956 5608 15957 5648
rect 15915 5599 15957 5608
rect 16195 5648 16253 5649
rect 16195 5608 16204 5648
rect 16244 5608 16253 5648
rect 16195 5607 16253 5608
rect 16491 5648 16533 5657
rect 16491 5608 16492 5648
rect 16532 5608 16533 5648
rect 16491 5599 16533 5608
rect 16587 5648 16629 5657
rect 16587 5608 16588 5648
rect 16628 5608 16629 5648
rect 16587 5599 16629 5608
rect 17067 5648 17109 5657
rect 17067 5608 17068 5648
rect 17108 5608 17109 5648
rect 17067 5599 17109 5608
rect 17259 5648 17301 5657
rect 17259 5608 17260 5648
rect 17300 5608 17301 5648
rect 17259 5599 17301 5608
rect 17443 5648 17501 5649
rect 17443 5608 17452 5648
rect 17492 5608 17501 5648
rect 17443 5607 17501 5608
rect 18691 5648 18749 5649
rect 18691 5608 18700 5648
rect 18740 5608 18749 5648
rect 18691 5607 18749 5608
rect 19171 5648 19229 5649
rect 19171 5608 19180 5648
rect 19220 5608 19229 5648
rect 19171 5607 19229 5608
rect 19467 5648 19509 5657
rect 19467 5608 19468 5648
rect 19508 5608 19509 5648
rect 19467 5599 19509 5608
rect 19563 5648 19605 5657
rect 19563 5608 19564 5648
rect 19604 5608 19605 5648
rect 19563 5599 19605 5608
rect 20043 5648 20085 5657
rect 20043 5608 20044 5648
rect 20084 5608 20085 5648
rect 20043 5599 20085 5608
rect 20235 5648 20277 5657
rect 20235 5608 20236 5648
rect 20276 5608 20277 5648
rect 20235 5599 20277 5608
rect 1411 5480 1469 5481
rect 1411 5440 1420 5480
rect 1460 5440 1469 5480
rect 1411 5439 1469 5440
rect 7755 5480 7797 5489
rect 7755 5440 7756 5480
rect 7796 5440 7797 5480
rect 7755 5431 7797 5440
rect 9763 5480 9821 5481
rect 9763 5440 9772 5480
rect 9812 5440 9821 5480
rect 9763 5439 9821 5440
rect 10251 5480 10293 5489
rect 10251 5440 10252 5480
rect 10292 5440 10293 5480
rect 10251 5431 10293 5440
rect 12171 5480 12213 5489
rect 12171 5440 12172 5480
rect 12212 5440 12213 5480
rect 12171 5431 12213 5440
rect 12643 5480 12701 5481
rect 12643 5440 12652 5480
rect 12692 5440 12701 5480
rect 12643 5439 12701 5440
rect 13803 5480 13845 5489
rect 13803 5440 13804 5480
rect 13844 5440 13845 5480
rect 13803 5431 13845 5440
rect 15531 5480 15573 5489
rect 15531 5440 15532 5480
rect 15572 5440 15573 5480
rect 15531 5431 15573 5440
rect 15819 5480 15861 5489
rect 15819 5440 15820 5480
rect 15860 5440 15861 5480
rect 15819 5431 15861 5440
rect 18891 5480 18933 5489
rect 18891 5440 18892 5480
rect 18932 5440 18933 5480
rect 18891 5431 18933 5440
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 15627 5144 15669 5153
rect 15627 5104 15628 5144
rect 15668 5104 15669 5144
rect 15627 5095 15669 5104
rect 15915 5144 15957 5153
rect 15915 5104 15916 5144
rect 15956 5104 15957 5144
rect 15915 5095 15957 5104
rect 17347 5144 17405 5145
rect 17347 5104 17356 5144
rect 17396 5104 17405 5144
rect 17347 5103 17405 5104
rect 17731 5144 17789 5145
rect 17731 5104 17740 5144
rect 17780 5104 17789 5144
rect 17731 5103 17789 5104
rect 6315 5060 6357 5069
rect 6315 5020 6316 5060
rect 6356 5020 6357 5060
rect 6315 5011 6357 5020
rect 7371 5060 7413 5069
rect 7371 5020 7372 5060
rect 7412 5020 7413 5060
rect 7371 5011 7413 5020
rect 8331 5060 8373 5069
rect 8331 5020 8332 5060
rect 8372 5020 8373 5060
rect 8331 5011 8373 5020
rect 10347 5060 10389 5069
rect 10347 5020 10348 5060
rect 10388 5020 10389 5060
rect 10347 5011 10389 5020
rect 11115 5060 11157 5069
rect 11115 5020 11116 5060
rect 11156 5020 11157 5060
rect 11115 5011 11157 5020
rect 16587 5060 16629 5069
rect 16587 5020 16588 5060
rect 16628 5020 16629 5060
rect 16587 5011 16629 5020
rect 19179 5060 19221 5069
rect 19179 5020 19180 5060
rect 19220 5020 19221 5060
rect 19179 5011 19221 5020
rect 1227 4976 1269 4985
rect 1227 4936 1228 4976
rect 1268 4936 1269 4976
rect 1227 4927 1269 4936
rect 1411 4976 1469 4977
rect 1411 4936 1420 4976
rect 1460 4936 1469 4976
rect 1411 4935 1469 4936
rect 1603 4976 1661 4977
rect 1603 4936 1612 4976
rect 1652 4936 1661 4976
rect 1603 4935 1661 4936
rect 2851 4976 2909 4977
rect 2851 4936 2860 4976
rect 2900 4936 2909 4976
rect 2851 4935 2909 4936
rect 3235 4976 3293 4977
rect 3235 4936 3244 4976
rect 3284 4936 3293 4976
rect 3235 4935 3293 4936
rect 4483 4976 4541 4977
rect 4483 4936 4492 4976
rect 4532 4936 4541 4976
rect 4483 4935 4541 4936
rect 4867 4976 4925 4977
rect 4867 4936 4876 4976
rect 4916 4936 4925 4976
rect 4867 4935 4925 4936
rect 6115 4976 6173 4977
rect 6115 4936 6124 4976
rect 6164 4936 6173 4976
rect 6115 4935 6173 4936
rect 7651 4976 7709 4977
rect 7651 4936 7660 4976
rect 7700 4936 7709 4976
rect 7651 4935 7709 4936
rect 7755 4976 7797 4985
rect 7755 4936 7756 4976
rect 7796 4936 7797 4976
rect 7755 4927 7797 4936
rect 7939 4976 7997 4977
rect 7939 4936 7948 4976
rect 7988 4936 7997 4976
rect 8995 4976 9053 4977
rect 7939 4935 7997 4936
rect 8523 4962 8565 4971
rect 8523 4922 8524 4962
rect 8564 4922 8565 4962
rect 8995 4936 9004 4976
rect 9044 4936 9053 4976
rect 8995 4935 9053 4936
rect 9579 4976 9621 4985
rect 9579 4936 9580 4976
rect 9620 4936 9621 4976
rect 9579 4927 9621 4936
rect 9963 4976 10005 4985
rect 9963 4936 9964 4976
rect 10004 4936 10005 4976
rect 9963 4927 10005 4936
rect 10059 4976 10101 4985
rect 10059 4936 10060 4976
rect 10100 4936 10101 4976
rect 10059 4927 10101 4936
rect 10635 4976 10677 4985
rect 10635 4936 10636 4976
rect 10676 4936 10677 4976
rect 10635 4927 10677 4936
rect 10923 4976 10965 4985
rect 10923 4936 10924 4976
rect 10964 4936 10965 4976
rect 11779 4976 11837 4977
rect 10923 4927 10965 4936
rect 11307 4962 11349 4971
rect 8523 4913 8565 4922
rect 11307 4922 11308 4962
rect 11348 4922 11349 4962
rect 11779 4936 11788 4976
rect 11828 4936 11837 4976
rect 11779 4935 11837 4936
rect 12267 4976 12309 4985
rect 12267 4936 12268 4976
rect 12308 4936 12309 4976
rect 12267 4927 12309 4936
rect 12363 4976 12405 4985
rect 12363 4936 12364 4976
rect 12404 4936 12405 4976
rect 12363 4927 12405 4936
rect 12747 4976 12789 4985
rect 12747 4936 12748 4976
rect 12788 4936 12789 4976
rect 12747 4927 12789 4936
rect 12843 4976 12885 4985
rect 12843 4936 12844 4976
rect 12884 4936 12885 4976
rect 12843 4927 12885 4936
rect 13131 4976 13173 4985
rect 13131 4936 13132 4976
rect 13172 4936 13173 4976
rect 13131 4927 13173 4936
rect 13323 4976 13365 4985
rect 13323 4936 13324 4976
rect 13364 4936 13365 4976
rect 13323 4927 13365 4936
rect 13411 4976 13469 4977
rect 13411 4936 13420 4976
rect 13460 4936 13469 4976
rect 13411 4935 13469 4936
rect 13707 4976 13749 4985
rect 13707 4936 13708 4976
rect 13748 4936 13749 4976
rect 13707 4927 13749 4936
rect 13803 4976 13845 4985
rect 13803 4936 13804 4976
rect 13844 4936 13845 4976
rect 13803 4927 13845 4936
rect 13899 4976 13941 4985
rect 13899 4936 13900 4976
rect 13940 4936 13941 4976
rect 13899 4927 13941 4936
rect 13995 4976 14037 4985
rect 13995 4936 13996 4976
rect 14036 4936 14037 4976
rect 13995 4927 14037 4936
rect 14179 4976 14237 4977
rect 14179 4936 14188 4976
rect 14228 4936 14237 4976
rect 14179 4935 14237 4936
rect 15427 4976 15485 4977
rect 15427 4936 15436 4976
rect 15476 4936 15485 4976
rect 15427 4935 15485 4936
rect 15811 4976 15869 4977
rect 15811 4936 15820 4976
rect 15860 4936 15869 4976
rect 15811 4935 15869 4936
rect 16195 4976 16253 4977
rect 16195 4936 16204 4976
rect 16244 4936 16253 4976
rect 16195 4935 16253 4936
rect 16491 4976 16533 4985
rect 16491 4936 16492 4976
rect 16532 4936 16533 4976
rect 16491 4927 16533 4936
rect 17067 4976 17109 4985
rect 17067 4936 17068 4976
rect 17108 4936 17109 4976
rect 17067 4927 17109 4936
rect 17163 4976 17205 4985
rect 17163 4936 17164 4976
rect 17204 4936 17205 4976
rect 17163 4927 17205 4936
rect 17827 4976 17885 4977
rect 17827 4936 17836 4976
rect 17876 4936 17885 4976
rect 17827 4935 17885 4936
rect 18403 4976 18461 4977
rect 18403 4936 18412 4976
rect 18452 4936 18461 4976
rect 18403 4935 18461 4936
rect 18507 4976 18549 4985
rect 18507 4936 18508 4976
rect 18548 4936 18549 4976
rect 18507 4927 18549 4936
rect 18691 4976 18749 4977
rect 18691 4936 18700 4976
rect 18740 4936 18749 4976
rect 18691 4935 18749 4936
rect 19275 4976 19317 4985
rect 19275 4936 19276 4976
rect 19316 4936 19317 4976
rect 19275 4927 19317 4936
rect 19555 4976 19613 4977
rect 19555 4936 19564 4976
rect 19604 4936 19613 4976
rect 19555 4935 19613 4936
rect 11307 4913 11349 4922
rect 6507 4892 6549 4901
rect 6507 4852 6508 4892
rect 6548 4852 6549 4892
rect 6507 4843 6549 4852
rect 6979 4892 7037 4893
rect 6979 4852 6988 4892
rect 7028 4852 7037 4892
rect 6979 4851 7037 4852
rect 9483 4892 9525 4901
rect 9483 4852 9484 4892
rect 9524 4852 9525 4892
rect 9483 4843 9525 4852
rect 19843 4892 19901 4893
rect 19843 4852 19852 4892
rect 19892 4852 19901 4892
rect 19843 4851 19901 4852
rect 7747 4808 7805 4809
rect 7747 4768 7756 4808
rect 7796 4768 7805 4808
rect 7747 4767 7805 4768
rect 10923 4808 10965 4817
rect 10923 4768 10924 4808
rect 10964 4768 10965 4808
rect 10923 4759 10965 4768
rect 16867 4808 16925 4809
rect 16867 4768 16876 4808
rect 16916 4768 16925 4808
rect 16867 4767 16925 4768
rect 18499 4808 18557 4809
rect 18499 4768 18508 4808
rect 18548 4768 18557 4808
rect 18499 4767 18557 4768
rect 20043 4808 20085 4817
rect 20043 4768 20044 4808
rect 20084 4768 20085 4808
rect 20043 4759 20085 4768
rect 1323 4724 1365 4733
rect 1323 4684 1324 4724
rect 1364 4684 1365 4724
rect 1323 4675 1365 4684
rect 3051 4724 3093 4733
rect 3051 4684 3052 4724
rect 3092 4684 3093 4724
rect 3051 4675 3093 4684
rect 4683 4724 4725 4733
rect 4683 4684 4684 4724
rect 4724 4684 4725 4724
rect 4683 4675 4725 4684
rect 7179 4724 7221 4733
rect 7179 4684 7180 4724
rect 7220 4684 7221 4724
rect 7179 4675 7221 4684
rect 13131 4724 13173 4733
rect 13131 4684 13132 4724
rect 13172 4684 13173 4724
rect 13131 4675 13173 4684
rect 18019 4724 18077 4725
rect 18019 4684 18028 4724
rect 18068 4684 18077 4724
rect 18019 4683 18077 4684
rect 18883 4724 18941 4725
rect 18883 4684 18892 4724
rect 18932 4684 18941 4724
rect 18883 4683 18941 4684
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 3435 4388 3477 4397
rect 3435 4348 3436 4388
rect 3476 4348 3477 4388
rect 3435 4339 3477 4348
rect 6987 4388 7029 4397
rect 6987 4348 6988 4388
rect 7028 4348 7029 4388
rect 6987 4339 7029 4348
rect 10923 4388 10965 4397
rect 10923 4348 10924 4388
rect 10964 4348 10965 4388
rect 10923 4339 10965 4348
rect 13515 4388 13557 4397
rect 13515 4348 13516 4388
rect 13556 4348 13557 4388
rect 13515 4339 13557 4348
rect 18219 4388 18261 4397
rect 18219 4348 18220 4388
rect 18260 4348 18261 4388
rect 18219 4339 18261 4348
rect 5643 4304 5685 4313
rect 5643 4264 5644 4304
rect 5684 4264 5685 4304
rect 5643 4255 5685 4264
rect 5931 4304 5973 4313
rect 5931 4264 5932 4304
rect 5972 4264 5973 4304
rect 5931 4255 5973 4264
rect 6219 4304 6261 4313
rect 6219 4264 6220 4304
rect 6260 4264 6261 4304
rect 6219 4255 6261 4264
rect 9099 4304 9141 4313
rect 9099 4264 9100 4304
rect 9140 4264 9141 4304
rect 9099 4255 9141 4264
rect 9291 4304 9333 4313
rect 9291 4264 9292 4304
rect 9332 4264 9333 4304
rect 9291 4255 9333 4264
rect 18603 4304 18645 4313
rect 18603 4264 18604 4304
rect 18644 4264 18645 4304
rect 18603 4255 18645 4264
rect 19747 4304 19805 4305
rect 19747 4264 19756 4304
rect 19796 4264 19805 4304
rect 19747 4263 19805 4264
rect 9571 4231 9629 4232
rect 1227 4220 1269 4229
rect 1227 4180 1228 4220
rect 1268 4180 1269 4220
rect 1227 4171 1269 4180
rect 4779 4220 4821 4229
rect 4779 4180 4780 4220
rect 4820 4180 4821 4220
rect 4779 4171 4821 4180
rect 4875 4220 4917 4229
rect 4875 4180 4876 4220
rect 4916 4180 4917 4220
rect 9571 4191 9580 4231
rect 9620 4191 9629 4231
rect 9571 4190 9629 4191
rect 9955 4220 10013 4221
rect 4875 4171 4917 4180
rect 9955 4180 9964 4220
rect 10004 4180 10013 4220
rect 9955 4179 10013 4180
rect 10443 4220 10485 4229
rect 10443 4180 10444 4220
rect 10484 4180 10485 4220
rect 10443 4171 10485 4180
rect 11587 4220 11645 4221
rect 11587 4180 11596 4220
rect 11636 4180 11645 4220
rect 11587 4179 11645 4180
rect 16587 4220 16629 4229
rect 16587 4180 16588 4220
rect 16628 4180 16629 4220
rect 16587 4171 16629 4180
rect 18507 4220 18549 4229
rect 18507 4180 18508 4220
rect 18548 4180 18549 4220
rect 18507 4171 18549 4180
rect 18699 4220 18741 4229
rect 18699 4180 18700 4220
rect 18740 4180 18741 4220
rect 18699 4171 18741 4180
rect 1515 4136 1557 4145
rect 1515 4096 1516 4136
rect 1556 4096 1557 4136
rect 1515 4087 1557 4096
rect 1611 4136 1653 4145
rect 1611 4096 1612 4136
rect 1652 4096 1653 4136
rect 1611 4087 1653 4096
rect 1707 4136 1749 4145
rect 1707 4096 1708 4136
rect 1748 4096 1749 4136
rect 1707 4087 1749 4096
rect 1803 4136 1845 4145
rect 3819 4141 3861 4150
rect 1803 4096 1804 4136
rect 1844 4096 1845 4136
rect 1803 4087 1845 4096
rect 1987 4136 2045 4137
rect 1987 4096 1996 4136
rect 2036 4096 2045 4136
rect 1987 4095 2045 4096
rect 3235 4136 3293 4137
rect 3235 4096 3244 4136
rect 3284 4096 3293 4136
rect 3235 4095 3293 4096
rect 3819 4101 3820 4141
rect 3860 4101 3861 4141
rect 3819 4092 3861 4101
rect 4291 4136 4349 4137
rect 4291 4096 4300 4136
rect 4340 4096 4349 4136
rect 4291 4095 4349 4096
rect 5259 4136 5301 4145
rect 5259 4096 5260 4136
rect 5300 4096 5301 4136
rect 5259 4087 5301 4096
rect 5355 4136 5397 4145
rect 5355 4096 5356 4136
rect 5396 4096 5397 4136
rect 5355 4087 5397 4096
rect 6507 4136 6549 4145
rect 6507 4096 6508 4136
rect 6548 4096 6549 4136
rect 6507 4087 6549 4096
rect 6603 4136 6645 4145
rect 6603 4096 6604 4136
rect 6644 4096 6645 4136
rect 6795 4136 6837 4145
rect 6603 4087 6645 4096
rect 6699 4115 6741 4124
rect 6699 4075 6700 4115
rect 6740 4075 6741 4115
rect 6795 4096 6796 4136
rect 6836 4096 6837 4136
rect 6795 4087 6837 4096
rect 7075 4136 7133 4137
rect 7075 4096 7084 4136
rect 7124 4096 7133 4136
rect 7075 4095 7133 4096
rect 7275 4136 7317 4145
rect 7275 4096 7276 4136
rect 7316 4096 7317 4136
rect 7275 4087 7317 4096
rect 7467 4136 7509 4145
rect 7467 4096 7468 4136
rect 7508 4096 7509 4136
rect 7467 4087 7509 4096
rect 7651 4136 7709 4137
rect 7651 4096 7660 4136
rect 7700 4096 7709 4136
rect 7651 4095 7709 4096
rect 8899 4136 8957 4137
rect 8899 4096 8908 4136
rect 8948 4096 8957 4136
rect 8899 4095 8957 4096
rect 10347 4136 10389 4145
rect 10347 4096 10348 4136
rect 10388 4096 10389 4136
rect 10347 4087 10389 4096
rect 10539 4136 10581 4145
rect 10539 4096 10540 4136
rect 10580 4096 10581 4136
rect 10539 4087 10581 4096
rect 10731 4136 10773 4145
rect 10731 4096 10732 4136
rect 10772 4096 10773 4136
rect 10731 4087 10773 4096
rect 10923 4136 10965 4145
rect 10923 4096 10924 4136
rect 10964 4096 10965 4136
rect 10923 4087 10965 4096
rect 11115 4136 11157 4145
rect 11115 4096 11116 4136
rect 11156 4096 11157 4136
rect 11115 4087 11157 4096
rect 11307 4136 11349 4145
rect 11307 4096 11308 4136
rect 11348 4096 11349 4136
rect 11307 4087 11349 4096
rect 11395 4136 11453 4137
rect 11395 4096 11404 4136
rect 11444 4096 11453 4136
rect 11395 4095 11453 4096
rect 12067 4136 12125 4137
rect 12067 4096 12076 4136
rect 12116 4096 12125 4136
rect 12067 4095 12125 4096
rect 13315 4136 13373 4137
rect 13315 4096 13324 4136
rect 13364 4096 13373 4136
rect 13315 4095 13373 4096
rect 13707 4136 13749 4145
rect 13707 4096 13708 4136
rect 13748 4096 13749 4136
rect 13707 4087 13749 4096
rect 13803 4136 13845 4145
rect 13803 4096 13804 4136
rect 13844 4096 13845 4136
rect 13803 4087 13845 4096
rect 13899 4136 13941 4145
rect 13899 4096 13900 4136
rect 13940 4096 13941 4136
rect 13899 4087 13941 4096
rect 14275 4136 14333 4137
rect 14275 4096 14284 4136
rect 14324 4096 14333 4136
rect 14275 4095 14333 4096
rect 15523 4136 15581 4137
rect 15523 4096 15532 4136
rect 15572 4096 15581 4136
rect 15523 4095 15581 4096
rect 16011 4136 16053 4145
rect 16011 4096 16012 4136
rect 16052 4096 16053 4136
rect 16011 4087 16053 4096
rect 16107 4136 16149 4145
rect 16107 4096 16108 4136
rect 16148 4096 16149 4136
rect 16107 4087 16149 4096
rect 16491 4136 16533 4145
rect 17547 4141 17589 4150
rect 16491 4096 16492 4136
rect 16532 4096 16533 4136
rect 16491 4087 16533 4096
rect 17059 4136 17117 4137
rect 17059 4096 17068 4136
rect 17108 4096 17117 4136
rect 17059 4095 17117 4096
rect 17547 4101 17548 4141
rect 17588 4101 17589 4141
rect 17547 4092 17589 4101
rect 17923 4136 17981 4137
rect 17923 4096 17932 4136
rect 17972 4096 17981 4136
rect 17923 4095 17981 4096
rect 18027 4136 18069 4145
rect 18027 4096 18028 4136
rect 18068 4096 18069 4136
rect 18027 4087 18069 4096
rect 18219 4136 18261 4145
rect 18219 4096 18220 4136
rect 18260 4096 18261 4136
rect 18219 4087 18261 4096
rect 18411 4136 18453 4145
rect 18411 4096 18412 4136
rect 18452 4096 18453 4136
rect 18411 4087 18453 4096
rect 18787 4136 18845 4137
rect 18787 4096 18796 4136
rect 18836 4096 18845 4136
rect 18787 4095 18845 4096
rect 19075 4136 19133 4137
rect 19075 4096 19084 4136
rect 19124 4096 19133 4136
rect 19075 4095 19133 4096
rect 19371 4136 19413 4145
rect 19371 4096 19372 4136
rect 19412 4096 19413 4136
rect 19371 4087 19413 4096
rect 19467 4136 19509 4145
rect 19467 4096 19468 4136
rect 19508 4096 19509 4136
rect 19467 4087 19509 4096
rect 19947 4136 19989 4145
rect 19947 4096 19948 4136
rect 19988 4096 19989 4136
rect 19947 4087 19989 4096
rect 20121 4141 20163 4150
rect 20121 4101 20122 4141
rect 20162 4101 20163 4141
rect 20121 4092 20163 4101
rect 6699 4066 6741 4075
rect 3627 4052 3669 4061
rect 3627 4012 3628 4052
rect 3668 4012 3669 4052
rect 3627 4003 3669 4012
rect 15723 4052 15765 4061
rect 15723 4012 15724 4052
rect 15764 4012 15765 4052
rect 15723 4003 15765 4012
rect 7371 3968 7413 3977
rect 7371 3928 7372 3968
rect 7412 3928 7413 3968
rect 7371 3919 7413 3928
rect 9771 3968 9813 3977
rect 9771 3928 9772 3968
rect 9812 3928 9813 3968
rect 9771 3919 9813 3928
rect 10155 3968 10197 3977
rect 10155 3928 10156 3968
rect 10196 3928 10197 3968
rect 10155 3919 10197 3928
rect 11203 3968 11261 3969
rect 11203 3928 11212 3968
rect 11252 3928 11261 3968
rect 11203 3927 11261 3928
rect 11787 3968 11829 3977
rect 11787 3928 11788 3968
rect 11828 3928 11829 3968
rect 11787 3919 11829 3928
rect 13987 3968 14045 3969
rect 13987 3928 13996 3968
rect 14036 3928 14045 3968
rect 13987 3927 14045 3928
rect 17739 3968 17781 3977
rect 17739 3928 17740 3968
rect 17780 3928 17781 3968
rect 17739 3919 17781 3928
rect 20043 3968 20085 3977
rect 20043 3928 20044 3968
rect 20084 3928 20085 3968
rect 20043 3919 20085 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 1411 3632 1469 3633
rect 1411 3592 1420 3632
rect 1460 3592 1469 3632
rect 1411 3591 1469 3592
rect 3619 3632 3677 3633
rect 3619 3592 3628 3632
rect 3668 3592 3677 3632
rect 3619 3591 3677 3592
rect 6499 3632 6557 3633
rect 6499 3592 6508 3632
rect 6548 3592 6557 3632
rect 6499 3591 6557 3592
rect 8235 3632 8277 3641
rect 8235 3592 8236 3632
rect 8276 3592 8277 3632
rect 8235 3583 8277 3592
rect 12075 3632 12117 3641
rect 12075 3592 12076 3632
rect 12116 3592 12117 3632
rect 12075 3583 12117 3592
rect 17067 3632 17109 3641
rect 17067 3592 17068 3632
rect 17108 3592 17109 3632
rect 17067 3583 17109 3592
rect 3435 3548 3477 3557
rect 3435 3508 3436 3548
rect 3476 3508 3477 3548
rect 3435 3499 3477 3508
rect 6315 3548 6357 3557
rect 6315 3508 6316 3548
rect 6356 3508 6357 3548
rect 6315 3499 6357 3508
rect 8523 3548 8565 3557
rect 8523 3508 8524 3548
rect 8564 3508 8565 3548
rect 8523 3499 8565 3508
rect 15819 3548 15861 3557
rect 15819 3508 15820 3548
rect 15860 3508 15861 3548
rect 15819 3499 15861 3508
rect 20043 3548 20085 3557
rect 20043 3508 20044 3548
rect 20084 3508 20085 3548
rect 20043 3499 20085 3508
rect 1987 3464 2045 3465
rect 1987 3424 1996 3464
rect 2036 3424 2045 3464
rect 1987 3423 2045 3424
rect 3235 3464 3293 3465
rect 3235 3424 3244 3464
rect 3284 3424 3293 3464
rect 3235 3423 3293 3424
rect 3723 3464 3765 3473
rect 3723 3424 3724 3464
rect 3764 3424 3765 3464
rect 3723 3415 3765 3424
rect 3819 3464 3861 3473
rect 3819 3424 3820 3464
rect 3860 3424 3861 3464
rect 3819 3415 3861 3424
rect 3915 3464 3957 3473
rect 3915 3424 3916 3464
rect 3956 3424 3957 3464
rect 3915 3415 3957 3424
rect 4587 3464 4629 3473
rect 4587 3424 4588 3464
rect 4628 3424 4629 3464
rect 5635 3464 5693 3465
rect 4587 3415 4629 3424
rect 4683 3445 4725 3454
rect 4683 3405 4684 3445
rect 4724 3405 4725 3445
rect 5635 3424 5644 3464
rect 5684 3424 5693 3464
rect 6787 3464 6845 3465
rect 5635 3423 5693 3424
rect 6123 3450 6165 3459
rect 4683 3396 4725 3405
rect 6123 3410 6124 3450
rect 6164 3410 6165 3450
rect 6787 3424 6796 3464
rect 6836 3424 6845 3464
rect 6787 3423 6845 3424
rect 8035 3464 8093 3465
rect 8035 3424 8044 3464
rect 8084 3424 8093 3464
rect 9187 3464 9245 3465
rect 8035 3423 8093 3424
rect 6123 3401 6165 3410
rect 8667 3422 8709 3431
rect 9187 3424 9196 3464
rect 9236 3424 9245 3464
rect 9187 3423 9245 3424
rect 9675 3464 9717 3473
rect 9675 3424 9676 3464
rect 9716 3424 9717 3464
rect 5067 3380 5109 3389
rect 5067 3340 5068 3380
rect 5108 3340 5109 3380
rect 5067 3331 5109 3340
rect 5163 3380 5205 3389
rect 5163 3340 5164 3380
rect 5204 3340 5205 3380
rect 8667 3382 8668 3422
rect 8708 3382 8709 3422
rect 9675 3415 9717 3424
rect 10155 3464 10197 3473
rect 10155 3424 10156 3464
rect 10196 3424 10197 3464
rect 10155 3415 10197 3424
rect 10251 3464 10293 3473
rect 10251 3424 10252 3464
rect 10292 3424 10293 3464
rect 10251 3415 10293 3424
rect 11499 3464 11541 3473
rect 11499 3424 11500 3464
rect 11540 3424 11541 3464
rect 11499 3415 11541 3424
rect 11595 3464 11637 3473
rect 11595 3424 11596 3464
rect 11636 3424 11637 3464
rect 11595 3415 11637 3424
rect 11691 3464 11733 3473
rect 11691 3424 11692 3464
rect 11732 3424 11733 3464
rect 11691 3415 11733 3424
rect 11787 3464 11829 3473
rect 11787 3424 11788 3464
rect 11828 3424 11829 3464
rect 11787 3415 11829 3424
rect 12259 3464 12317 3465
rect 12259 3424 12268 3464
rect 12308 3424 12317 3464
rect 12259 3423 12317 3424
rect 13507 3464 13565 3465
rect 13507 3424 13516 3464
rect 13556 3424 13565 3464
rect 13507 3423 13565 3424
rect 13891 3464 13949 3465
rect 13891 3424 13900 3464
rect 13940 3424 13949 3464
rect 13891 3423 13949 3424
rect 15139 3464 15197 3465
rect 15139 3424 15148 3464
rect 15188 3424 15197 3464
rect 15139 3423 15197 3424
rect 15427 3464 15485 3465
rect 15427 3424 15436 3464
rect 15476 3424 15485 3464
rect 15427 3423 15485 3424
rect 15723 3464 15765 3473
rect 15723 3424 15724 3464
rect 15764 3424 15765 3464
rect 15723 3415 15765 3424
rect 16683 3464 16725 3473
rect 16683 3424 16684 3464
rect 16724 3424 16725 3464
rect 16683 3415 16725 3424
rect 16779 3464 16821 3473
rect 16779 3424 16780 3464
rect 16820 3424 16821 3464
rect 16779 3415 16821 3424
rect 16875 3464 16917 3473
rect 16875 3424 16876 3464
rect 16916 3424 16917 3464
rect 16875 3415 16917 3424
rect 17251 3464 17309 3465
rect 17251 3424 17260 3464
rect 17300 3424 17309 3464
rect 17251 3423 17309 3424
rect 17355 3464 17397 3473
rect 17355 3424 17356 3464
rect 17396 3424 17397 3464
rect 17355 3415 17397 3424
rect 17547 3464 17589 3473
rect 17547 3424 17548 3464
rect 17588 3424 17589 3464
rect 17547 3415 17589 3424
rect 17739 3464 17781 3473
rect 17739 3424 17740 3464
rect 17780 3424 17781 3464
rect 17739 3415 17781 3424
rect 17931 3464 17973 3473
rect 17931 3424 17932 3464
rect 17972 3424 17973 3464
rect 17931 3415 17973 3424
rect 18019 3464 18077 3465
rect 18019 3424 18028 3464
rect 18068 3424 18077 3464
rect 18019 3423 18077 3424
rect 18219 3464 18261 3473
rect 18219 3424 18220 3464
rect 18260 3424 18261 3464
rect 18219 3415 18261 3424
rect 18411 3464 18453 3473
rect 18411 3424 18412 3464
rect 18452 3424 18453 3464
rect 18411 3415 18453 3424
rect 18595 3464 18653 3465
rect 18595 3424 18604 3464
rect 18644 3424 18653 3464
rect 18595 3423 18653 3424
rect 18987 3464 19029 3473
rect 18987 3424 18988 3464
rect 19028 3424 19029 3464
rect 18987 3415 19029 3424
rect 19171 3464 19229 3465
rect 19171 3424 19180 3464
rect 19220 3424 19229 3464
rect 19171 3423 19229 3424
rect 19267 3464 19325 3465
rect 19267 3424 19276 3464
rect 19316 3424 19325 3464
rect 19267 3423 19325 3424
rect 19467 3464 19509 3473
rect 19467 3424 19468 3464
rect 19508 3424 19509 3464
rect 19467 3415 19509 3424
rect 19563 3464 19605 3473
rect 19563 3424 19564 3464
rect 19604 3424 19605 3464
rect 19563 3415 19605 3424
rect 19699 3464 19757 3465
rect 19699 3424 19708 3464
rect 19748 3424 19757 3464
rect 19699 3423 19757 3424
rect 19947 3464 19989 3473
rect 19947 3424 19948 3464
rect 19988 3424 19989 3464
rect 19947 3415 19989 3424
rect 20120 3451 20178 3452
rect 20120 3411 20129 3451
rect 20169 3411 20178 3451
rect 20120 3410 20178 3411
rect 8667 3373 8709 3382
rect 9771 3380 9813 3389
rect 5163 3331 5205 3340
rect 9771 3340 9772 3380
rect 9812 3340 9813 3380
rect 9771 3331 9813 3340
rect 10723 3380 10781 3381
rect 10723 3340 10732 3380
rect 10772 3340 10781 3380
rect 10723 3339 10781 3340
rect 11107 3380 11165 3381
rect 11107 3340 11116 3380
rect 11156 3340 11165 3380
rect 11107 3339 11165 3340
rect 18699 3380 18741 3389
rect 18699 3340 18700 3380
rect 18740 3340 18741 3380
rect 18699 3331 18741 3340
rect 18891 3380 18933 3389
rect 18891 3340 18892 3380
rect 18932 3340 18933 3380
rect 18891 3331 18933 3340
rect 1707 3296 1749 3305
rect 1707 3256 1708 3296
rect 1748 3256 1749 3296
rect 1707 3247 1749 3256
rect 4299 3296 4341 3305
rect 4299 3256 4300 3296
rect 4340 3256 4341 3296
rect 4299 3247 4341 3256
rect 16299 3296 16341 3305
rect 16299 3256 16300 3296
rect 16340 3256 16341 3296
rect 16299 3247 16341 3256
rect 17739 3296 17781 3305
rect 17739 3256 17740 3296
rect 17780 3256 17781 3296
rect 17739 3247 17781 3256
rect 18795 3296 18837 3305
rect 18795 3256 18796 3296
rect 18836 3256 18837 3296
rect 18795 3247 18837 3256
rect 10923 3212 10965 3221
rect 10923 3172 10924 3212
rect 10964 3172 10965 3212
rect 10923 3163 10965 3172
rect 11307 3212 11349 3221
rect 11307 3172 11308 3212
rect 11348 3172 11349 3212
rect 11307 3163 11349 3172
rect 13707 3212 13749 3221
rect 13707 3172 13708 3212
rect 13748 3172 13749 3212
rect 13707 3163 13749 3172
rect 16099 3212 16157 3213
rect 16099 3172 16108 3212
rect 16148 3172 16157 3212
rect 16099 3171 16157 3172
rect 17547 3212 17589 3221
rect 17547 3172 17548 3212
rect 17588 3172 17589 3212
rect 17547 3163 17589 3172
rect 18219 3212 18261 3221
rect 18219 3172 18220 3212
rect 18260 3172 18261 3212
rect 18219 3163 18261 3172
rect 19179 3212 19221 3221
rect 19179 3172 19180 3212
rect 19220 3172 19221 3212
rect 19179 3163 19221 3172
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 3627 2876 3669 2885
rect 3627 2836 3628 2876
rect 3668 2836 3669 2876
rect 3627 2827 3669 2836
rect 5739 2876 5781 2885
rect 5739 2836 5740 2876
rect 5780 2836 5781 2876
rect 5739 2827 5781 2836
rect 14091 2876 14133 2885
rect 14091 2836 14092 2876
rect 14132 2836 14133 2876
rect 14091 2827 14133 2836
rect 17355 2876 17397 2885
rect 17355 2836 17356 2876
rect 17396 2836 17397 2876
rect 17355 2827 17397 2836
rect 19467 2876 19509 2885
rect 19467 2836 19468 2876
rect 19508 2836 19509 2876
rect 19467 2827 19509 2836
rect 1611 2792 1653 2801
rect 1611 2752 1612 2792
rect 1652 2752 1653 2792
rect 1611 2743 1653 2752
rect 1899 2792 1941 2801
rect 1899 2752 1900 2792
rect 1940 2752 1941 2792
rect 1899 2743 1941 2752
rect 4875 2792 4917 2801
rect 4875 2752 4876 2792
rect 4916 2752 4917 2792
rect 4875 2743 4917 2752
rect 6123 2792 6165 2801
rect 6123 2752 6124 2792
rect 6164 2752 6165 2792
rect 6123 2743 6165 2752
rect 6507 2792 6549 2801
rect 6507 2752 6508 2792
rect 6548 2752 6549 2792
rect 6507 2743 6549 2752
rect 9291 2792 9333 2801
rect 9291 2752 9292 2792
rect 9332 2752 9333 2792
rect 9291 2743 9333 2752
rect 17547 2792 17589 2801
rect 17547 2752 17548 2792
rect 17588 2752 17589 2792
rect 17547 2743 17589 2752
rect 11203 2719 11261 2720
rect 5059 2708 5117 2709
rect 5059 2668 5068 2708
rect 5108 2668 5117 2708
rect 5059 2667 5117 2668
rect 6027 2708 6069 2717
rect 6027 2668 6028 2708
rect 6068 2668 6069 2708
rect 6027 2659 6069 2668
rect 6219 2708 6261 2717
rect 6219 2668 6220 2708
rect 6260 2668 6261 2708
rect 6219 2659 6261 2668
rect 7371 2708 7413 2717
rect 7371 2668 7372 2708
rect 7412 2668 7413 2708
rect 7371 2659 7413 2668
rect 7467 2708 7509 2717
rect 7467 2668 7468 2708
rect 7508 2668 7509 2708
rect 11203 2679 11212 2719
rect 11252 2679 11261 2719
rect 11203 2678 11261 2679
rect 11875 2708 11933 2709
rect 7467 2659 7509 2668
rect 11875 2668 11884 2708
rect 11924 2668 11933 2708
rect 11875 2667 11933 2668
rect 12171 2708 12213 2717
rect 12171 2668 12172 2708
rect 12212 2668 12213 2708
rect 12171 2659 12213 2668
rect 8427 2638 8469 2647
rect 1419 2624 1461 2633
rect 1419 2584 1420 2624
rect 1460 2584 1461 2624
rect 1419 2575 1461 2584
rect 2179 2624 2237 2625
rect 2179 2584 2188 2624
rect 2228 2584 2237 2624
rect 2179 2583 2237 2584
rect 3427 2624 3485 2625
rect 3427 2584 3436 2624
rect 3476 2584 3485 2624
rect 3427 2583 3485 2584
rect 4395 2624 4437 2633
rect 4395 2584 4396 2624
rect 4436 2584 4437 2624
rect 4395 2575 4437 2584
rect 4491 2624 4533 2633
rect 4491 2584 4492 2624
rect 4532 2584 4533 2624
rect 4491 2575 4533 2584
rect 5443 2624 5501 2625
rect 5443 2584 5452 2624
rect 5492 2584 5501 2624
rect 5443 2583 5501 2584
rect 5547 2624 5589 2633
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5547 2575 5589 2584
rect 5739 2624 5781 2633
rect 5739 2584 5740 2624
rect 5780 2584 5781 2624
rect 5739 2575 5781 2584
rect 5923 2624 5981 2625
rect 5923 2584 5932 2624
rect 5972 2584 5981 2624
rect 5923 2583 5981 2584
rect 6315 2624 6357 2633
rect 6315 2584 6316 2624
rect 6356 2584 6357 2624
rect 6315 2575 6357 2584
rect 6891 2624 6933 2633
rect 6891 2584 6892 2624
rect 6932 2584 6933 2624
rect 6891 2575 6933 2584
rect 6987 2624 7029 2633
rect 6987 2584 6988 2624
rect 7028 2584 7029 2624
rect 6987 2575 7029 2584
rect 7939 2624 7997 2625
rect 7939 2584 7948 2624
rect 7988 2584 7997 2624
rect 8427 2598 8428 2638
rect 8468 2598 8469 2638
rect 12075 2637 12117 2646
rect 8427 2589 8469 2598
rect 9003 2624 9045 2633
rect 7939 2583 7997 2584
rect 9003 2584 9004 2624
rect 9044 2584 9045 2624
rect 9003 2575 9045 2584
rect 9099 2624 9141 2633
rect 9099 2584 9100 2624
rect 9140 2584 9141 2624
rect 9099 2575 9141 2584
rect 9763 2624 9821 2625
rect 9763 2584 9772 2624
rect 9812 2584 9821 2624
rect 9763 2583 9821 2584
rect 11011 2624 11069 2625
rect 11011 2584 11020 2624
rect 11060 2584 11069 2624
rect 12075 2597 12076 2637
rect 12116 2597 12117 2637
rect 12075 2588 12117 2597
rect 12267 2624 12309 2633
rect 11011 2583 11069 2584
rect 12267 2584 12268 2624
rect 12308 2584 12309 2624
rect 12267 2575 12309 2584
rect 12643 2624 12701 2625
rect 12643 2584 12652 2624
rect 12692 2584 12701 2624
rect 12643 2583 12701 2584
rect 13891 2624 13949 2625
rect 13891 2584 13900 2624
rect 13940 2584 13949 2624
rect 13891 2583 13949 2584
rect 14275 2624 14333 2625
rect 14275 2584 14284 2624
rect 14324 2584 14333 2624
rect 14275 2583 14333 2584
rect 15523 2624 15581 2625
rect 15523 2584 15532 2624
rect 15572 2584 15581 2624
rect 15523 2583 15581 2584
rect 15715 2624 15773 2625
rect 15715 2584 15724 2624
rect 15764 2584 15773 2624
rect 15715 2583 15773 2584
rect 16963 2624 17021 2625
rect 16963 2584 16972 2624
rect 17012 2584 17021 2624
rect 16963 2583 17021 2584
rect 17547 2624 17589 2633
rect 17547 2584 17548 2624
rect 17588 2584 17589 2624
rect 17547 2575 17589 2584
rect 18019 2624 18077 2625
rect 18019 2584 18028 2624
rect 18068 2584 18077 2624
rect 18019 2583 18077 2584
rect 19267 2624 19325 2625
rect 19267 2584 19276 2624
rect 19316 2584 19325 2624
rect 19267 2583 19325 2584
rect 19651 2624 19709 2625
rect 19651 2584 19660 2624
rect 19700 2584 19709 2624
rect 19651 2583 19709 2584
rect 19755 2624 19797 2633
rect 19755 2584 19756 2624
rect 19796 2584 19797 2624
rect 19755 2575 19797 2584
rect 19947 2624 19989 2633
rect 19947 2584 19948 2624
rect 19988 2584 19989 2624
rect 19947 2575 19989 2584
rect 4011 2540 4053 2549
rect 4011 2500 4012 2540
rect 4052 2500 4053 2540
rect 4011 2491 4053 2500
rect 4779 2540 4821 2549
rect 4779 2500 4780 2540
rect 4820 2500 4821 2540
rect 4779 2491 4821 2500
rect 8619 2540 8661 2549
rect 8619 2500 8620 2540
rect 8660 2500 8661 2540
rect 8619 2491 8661 2500
rect 17163 2540 17205 2549
rect 17163 2500 17164 2540
rect 17204 2500 17205 2540
rect 17163 2491 17205 2500
rect 19851 2540 19893 2549
rect 19851 2500 19852 2540
rect 19892 2500 19893 2540
rect 19851 2491 19893 2500
rect 20139 2540 20181 2549
rect 20139 2500 20140 2540
rect 20180 2500 20181 2540
rect 20139 2491 20181 2500
rect 4195 2456 4253 2457
rect 4195 2416 4204 2456
rect 4244 2416 4253 2456
rect 4195 2415 4253 2416
rect 5259 2456 5301 2465
rect 5259 2416 5260 2456
rect 5300 2416 5301 2456
rect 5259 2407 5301 2416
rect 8803 2456 8861 2457
rect 8803 2416 8812 2456
rect 8852 2416 8861 2456
rect 8803 2415 8861 2416
rect 9579 2456 9621 2465
rect 9579 2416 9580 2456
rect 9620 2416 9621 2456
rect 9579 2407 9621 2416
rect 11403 2456 11445 2465
rect 11403 2416 11404 2456
rect 11444 2416 11445 2456
rect 11403 2407 11445 2416
rect 11691 2456 11733 2465
rect 11691 2416 11692 2456
rect 11732 2416 11733 2456
rect 11691 2407 11733 2416
rect 12459 2456 12501 2465
rect 12459 2416 12460 2456
rect 12500 2416 12501 2456
rect 12459 2407 12501 2416
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 1603 2120 1661 2121
rect 1603 2080 1612 2120
rect 1652 2080 1661 2120
rect 1603 2079 1661 2080
rect 1891 2120 1949 2121
rect 1891 2080 1900 2120
rect 1940 2080 1949 2120
rect 1891 2079 1949 2080
rect 5739 2120 5781 2129
rect 5739 2080 5740 2120
rect 5780 2080 5781 2120
rect 5739 2071 5781 2080
rect 8331 2120 8373 2129
rect 8331 2080 8332 2120
rect 8372 2080 8373 2120
rect 8331 2071 8373 2080
rect 9963 2120 10005 2129
rect 9963 2080 9964 2120
rect 10004 2080 10005 2120
rect 9963 2071 10005 2080
rect 11979 2120 12021 2129
rect 11979 2080 11980 2120
rect 12020 2080 12021 2120
rect 11979 2071 12021 2080
rect 17355 2120 17397 2129
rect 17355 2080 17356 2120
rect 17396 2080 17397 2120
rect 17355 2071 17397 2080
rect 19371 2120 19413 2129
rect 19371 2080 19372 2120
rect 19412 2080 19413 2120
rect 19371 2071 19413 2080
rect 19659 2120 19701 2129
rect 19659 2080 19660 2120
rect 19700 2080 19701 2120
rect 19659 2071 19701 2080
rect 20235 2120 20277 2129
rect 20235 2080 20236 2120
rect 20276 2080 20277 2120
rect 20235 2071 20277 2080
rect 8139 2036 8181 2045
rect 8139 1996 8140 2036
rect 8180 1996 8181 2036
rect 8139 1987 8181 1996
rect 15531 2036 15573 2045
rect 15531 1996 15532 2036
rect 15572 1996 15573 2036
rect 15531 1987 15573 1996
rect 2179 1952 2237 1953
rect 2179 1912 2188 1952
rect 2228 1912 2237 1952
rect 2179 1911 2237 1912
rect 3427 1952 3485 1953
rect 3427 1912 3436 1952
rect 3476 1912 3485 1952
rect 3427 1911 3485 1912
rect 4011 1952 4053 1961
rect 4011 1912 4012 1952
rect 4052 1912 4053 1952
rect 4011 1903 4053 1912
rect 4107 1952 4149 1961
rect 4107 1912 4108 1952
rect 4148 1912 4149 1952
rect 4107 1903 4149 1912
rect 4491 1952 4533 1961
rect 4491 1912 4492 1952
rect 4532 1912 4533 1952
rect 4491 1903 4533 1912
rect 5059 1952 5117 1953
rect 5059 1912 5068 1952
rect 5108 1912 5117 1952
rect 5059 1911 5117 1912
rect 5547 1947 5589 1956
rect 5547 1907 5548 1947
rect 5588 1907 5589 1947
rect 5547 1898 5589 1907
rect 6411 1952 6453 1961
rect 6411 1912 6412 1952
rect 6452 1912 6453 1952
rect 6411 1903 6453 1912
rect 6507 1952 6549 1961
rect 6507 1912 6508 1952
rect 6548 1912 6549 1952
rect 6507 1903 6549 1912
rect 6987 1952 7029 1961
rect 6987 1912 6988 1952
rect 7028 1912 7029 1952
rect 6987 1903 7029 1912
rect 7459 1952 7517 1953
rect 7459 1912 7468 1952
rect 7508 1912 7517 1952
rect 8515 1952 8573 1953
rect 7459 1911 7517 1912
rect 7947 1938 7989 1947
rect 7947 1898 7948 1938
rect 7988 1898 7989 1938
rect 8515 1912 8524 1952
rect 8564 1912 8573 1952
rect 8515 1911 8573 1912
rect 9763 1952 9821 1953
rect 9763 1912 9772 1952
rect 9812 1912 9821 1952
rect 9763 1911 9821 1912
rect 10147 1952 10205 1953
rect 10147 1912 10156 1952
rect 10196 1912 10205 1952
rect 10147 1911 10205 1912
rect 11395 1952 11453 1953
rect 11395 1912 11404 1952
rect 11444 1912 11453 1952
rect 11395 1911 11453 1912
rect 12163 1952 12221 1953
rect 12163 1912 12172 1952
rect 12212 1912 12221 1952
rect 12163 1911 12221 1912
rect 13411 1952 13469 1953
rect 13411 1912 13420 1952
rect 13460 1912 13469 1952
rect 13411 1911 13469 1912
rect 13603 1952 13661 1953
rect 13603 1912 13612 1952
rect 13652 1912 13661 1952
rect 13603 1911 13661 1912
rect 14851 1952 14909 1953
rect 14851 1912 14860 1952
rect 14900 1912 14909 1952
rect 14851 1911 14909 1912
rect 15243 1952 15285 1961
rect 15243 1912 15244 1952
rect 15284 1912 15285 1952
rect 15243 1903 15285 1912
rect 15339 1952 15381 1961
rect 15339 1912 15340 1952
rect 15380 1912 15381 1952
rect 15339 1903 15381 1912
rect 15435 1952 15477 1961
rect 15435 1912 15436 1952
rect 15476 1912 15477 1952
rect 15435 1903 15477 1912
rect 15907 1952 15965 1953
rect 15907 1912 15916 1952
rect 15956 1912 15965 1952
rect 15907 1911 15965 1912
rect 17155 1952 17213 1953
rect 17155 1912 17164 1952
rect 17204 1912 17213 1952
rect 17155 1911 17213 1912
rect 17923 1952 17981 1953
rect 17923 1912 17932 1952
rect 17972 1912 17981 1952
rect 17923 1911 17981 1912
rect 19171 1952 19229 1953
rect 19171 1912 19180 1952
rect 19220 1912 19229 1952
rect 19171 1911 19229 1912
rect 19651 1952 19709 1953
rect 19651 1912 19660 1952
rect 19700 1912 19709 1952
rect 19651 1911 19709 1912
rect 19851 1952 19893 1961
rect 19851 1912 19852 1952
rect 19892 1912 19893 1952
rect 19851 1903 19893 1912
rect 19939 1952 19997 1953
rect 19939 1912 19948 1952
rect 19988 1912 19997 1952
rect 19939 1911 19997 1912
rect 20126 1952 20168 1961
rect 20126 1912 20127 1952
rect 20167 1912 20168 1952
rect 20126 1903 20168 1912
rect 7947 1889 7989 1898
rect 1219 1868 1277 1869
rect 1219 1828 1228 1868
rect 1268 1828 1277 1868
rect 1219 1827 1277 1828
rect 4587 1868 4629 1877
rect 4587 1828 4588 1868
rect 4628 1828 4629 1868
rect 4587 1819 4629 1828
rect 5923 1868 5981 1869
rect 5923 1828 5932 1868
rect 5972 1828 5981 1868
rect 5923 1827 5981 1828
rect 6891 1868 6933 1877
rect 6891 1828 6892 1868
rect 6932 1828 6933 1868
rect 6891 1819 6933 1828
rect 11587 1868 11645 1869
rect 11587 1828 11596 1868
rect 11636 1828 11645 1868
rect 11587 1827 11645 1828
rect 17731 1868 17789 1869
rect 17731 1828 17740 1868
rect 17780 1828 17789 1868
rect 17731 1827 17789 1828
rect 1707 1784 1749 1793
rect 1707 1744 1708 1784
rect 1748 1744 1749 1784
rect 1707 1735 1749 1744
rect 3627 1784 3669 1793
rect 3627 1744 3628 1784
rect 3668 1744 3669 1784
rect 3627 1735 3669 1744
rect 1419 1700 1461 1709
rect 1419 1660 1420 1700
rect 1460 1660 1461 1700
rect 1419 1651 1461 1660
rect 6123 1700 6165 1709
rect 6123 1660 6124 1700
rect 6164 1660 6165 1700
rect 6123 1651 6165 1660
rect 11787 1700 11829 1709
rect 11787 1660 11788 1700
rect 11828 1660 11829 1700
rect 11787 1651 11829 1660
rect 15051 1700 15093 1709
rect 15051 1660 15052 1700
rect 15092 1660 15093 1700
rect 15051 1651 15093 1660
rect 17547 1700 17589 1709
rect 17547 1660 17548 1700
rect 17588 1660 17589 1700
rect 17547 1651 17589 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 9099 1364 9141 1373
rect 9099 1324 9100 1364
rect 9140 1324 9141 1364
rect 9099 1315 9141 1324
rect 11115 1364 11157 1373
rect 11115 1324 11116 1364
rect 11156 1324 11157 1364
rect 11115 1315 11157 1324
rect 12747 1364 12789 1373
rect 12747 1324 12748 1364
rect 12788 1324 12789 1364
rect 12747 1315 12789 1324
rect 19467 1364 19509 1373
rect 19467 1324 19468 1364
rect 19508 1324 19509 1364
rect 19467 1315 19509 1324
rect 1323 1280 1365 1289
rect 1323 1240 1324 1280
rect 1364 1240 1365 1280
rect 1323 1231 1365 1240
rect 3915 1280 3957 1289
rect 3915 1240 3916 1280
rect 3956 1240 3957 1280
rect 3915 1231 3957 1240
rect 4203 1280 4245 1289
rect 4203 1240 4204 1280
rect 4244 1240 4245 1280
rect 4203 1231 4245 1240
rect 4683 1280 4725 1289
rect 4683 1240 4684 1280
rect 4724 1240 4725 1280
rect 4683 1231 4725 1240
rect 7467 1280 7509 1289
rect 7467 1240 7468 1280
rect 7508 1240 7509 1280
rect 7467 1231 7509 1240
rect 12939 1280 12981 1289
rect 12939 1240 12940 1280
rect 12980 1240 12981 1280
rect 12939 1231 12981 1240
rect 1507 1196 1565 1197
rect 1507 1156 1516 1196
rect 1556 1156 1565 1196
rect 1507 1155 1565 1156
rect 2475 1196 2517 1205
rect 2475 1156 2476 1196
rect 2516 1156 2517 1196
rect 2475 1147 2517 1156
rect 2571 1196 2613 1205
rect 2571 1156 2572 1196
rect 2612 1156 2613 1196
rect 2571 1147 2613 1156
rect 4867 1196 4925 1197
rect 4867 1156 4876 1196
rect 4916 1156 4925 1196
rect 4867 1155 4925 1156
rect 5251 1196 5309 1197
rect 5251 1156 5260 1196
rect 5300 1156 5309 1196
rect 5251 1155 5309 1156
rect 5635 1196 5693 1197
rect 5635 1156 5644 1196
rect 5684 1156 5693 1196
rect 5635 1155 5693 1156
rect 9283 1196 9341 1197
rect 9283 1156 9292 1196
rect 9332 1156 9341 1196
rect 9283 1155 9341 1156
rect 13899 1196 13941 1205
rect 13899 1156 13900 1196
rect 13940 1156 13941 1196
rect 13899 1147 13941 1156
rect 19843 1196 19901 1197
rect 19843 1156 19852 1196
rect 19892 1156 19901 1196
rect 19843 1155 19901 1156
rect 20227 1196 20285 1197
rect 20227 1156 20236 1196
rect 20276 1156 20285 1196
rect 20227 1155 20285 1156
rect 1995 1112 2037 1121
rect 1995 1072 1996 1112
rect 2036 1072 2037 1112
rect 1995 1063 2037 1072
rect 2091 1112 2133 1121
rect 3531 1117 3573 1126
rect 2091 1072 2092 1112
rect 2132 1072 2133 1112
rect 2091 1063 2133 1072
rect 3043 1112 3101 1113
rect 3043 1072 3052 1112
rect 3092 1072 3101 1112
rect 3043 1071 3101 1072
rect 3531 1077 3532 1117
rect 3572 1077 3573 1117
rect 3531 1068 3573 1077
rect 6019 1112 6077 1113
rect 6019 1072 6028 1112
rect 6068 1072 6077 1112
rect 6019 1071 6077 1072
rect 7267 1112 7325 1113
rect 7267 1072 7276 1112
rect 7316 1072 7325 1112
rect 7267 1071 7325 1072
rect 7651 1112 7709 1113
rect 7651 1072 7660 1112
rect 7700 1072 7709 1112
rect 7651 1071 7709 1072
rect 8899 1112 8957 1113
rect 8899 1072 8908 1112
rect 8948 1072 8957 1112
rect 8899 1071 8957 1072
rect 9667 1112 9725 1113
rect 9667 1072 9676 1112
rect 9716 1072 9725 1112
rect 9667 1071 9725 1072
rect 10915 1112 10973 1113
rect 10915 1072 10924 1112
rect 10964 1072 10973 1112
rect 10915 1071 10973 1072
rect 11299 1112 11357 1113
rect 11299 1072 11308 1112
rect 11348 1072 11357 1112
rect 11299 1071 11357 1072
rect 12547 1112 12605 1113
rect 12547 1072 12556 1112
rect 12596 1072 12605 1112
rect 12547 1071 12605 1072
rect 12939 1112 12981 1121
rect 12939 1072 12940 1112
rect 12980 1072 12981 1112
rect 12939 1063 12981 1072
rect 13131 1112 13173 1121
rect 13131 1072 13132 1112
rect 13172 1072 13173 1112
rect 13131 1063 13173 1072
rect 13219 1112 13277 1113
rect 13219 1072 13228 1112
rect 13268 1072 13277 1112
rect 13219 1071 13277 1072
rect 13419 1112 13461 1121
rect 13419 1072 13420 1112
rect 13460 1072 13461 1112
rect 13419 1063 13461 1072
rect 13515 1112 13557 1121
rect 13515 1072 13516 1112
rect 13556 1072 13557 1112
rect 13515 1063 13557 1072
rect 13611 1112 13653 1121
rect 13611 1072 13612 1112
rect 13652 1072 13653 1112
rect 13611 1063 13653 1072
rect 13707 1112 13749 1121
rect 13707 1072 13708 1112
rect 13748 1072 13749 1112
rect 13707 1063 13749 1072
rect 14371 1112 14429 1113
rect 14371 1072 14380 1112
rect 14420 1072 14429 1112
rect 14371 1071 14429 1072
rect 15619 1112 15677 1113
rect 15619 1072 15628 1112
rect 15668 1072 15677 1112
rect 15619 1071 15677 1072
rect 16003 1112 16061 1113
rect 16003 1072 16012 1112
rect 16052 1072 16061 1112
rect 16003 1071 16061 1072
rect 17251 1112 17309 1113
rect 17251 1072 17260 1112
rect 17300 1072 17309 1112
rect 17251 1071 17309 1072
rect 17451 1112 17493 1121
rect 17451 1072 17452 1112
rect 17492 1072 17493 1112
rect 17451 1063 17493 1072
rect 17643 1112 17685 1121
rect 17643 1072 17644 1112
rect 17684 1072 17685 1112
rect 17643 1063 17685 1072
rect 17731 1112 17789 1113
rect 17731 1072 17740 1112
rect 17780 1072 17789 1112
rect 17731 1071 17789 1072
rect 18019 1112 18077 1113
rect 18019 1072 18028 1112
rect 18068 1072 18077 1112
rect 18019 1071 18077 1072
rect 19267 1112 19325 1113
rect 19267 1072 19276 1112
rect 19316 1072 19325 1112
rect 19267 1071 19325 1072
rect 3723 1028 3765 1037
rect 3723 988 3724 1028
rect 3764 988 3765 1028
rect 3723 979 3765 988
rect 17547 1028 17589 1037
rect 17547 988 17548 1028
rect 17588 988 17589 1028
rect 17547 979 17589 988
rect 1707 944 1749 953
rect 1707 904 1708 944
rect 1748 904 1749 944
rect 1707 895 1749 904
rect 5067 944 5109 953
rect 5067 904 5068 944
rect 5108 904 5109 944
rect 5067 895 5109 904
rect 5451 944 5493 953
rect 5451 904 5452 944
rect 5492 904 5493 944
rect 5451 895 5493 904
rect 5835 944 5877 953
rect 5835 904 5836 944
rect 5876 904 5877 944
rect 5835 895 5877 904
rect 9483 944 9525 953
rect 9483 904 9484 944
rect 9524 904 9525 944
rect 9483 895 9525 904
rect 14187 944 14229 953
rect 14187 904 14188 944
rect 14228 904 14229 944
rect 14187 895 14229 904
rect 15819 944 15861 953
rect 15819 904 15820 944
rect 15860 904 15861 944
rect 15819 895 15861 904
rect 19659 944 19701 953
rect 19659 904 19660 944
rect 19700 904 19701 944
rect 19659 895 19701 904
rect 20043 944 20085 953
rect 20043 904 20044 944
rect 20084 904 20085 944
rect 20043 895 20085 904
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 19468 41392 19508 41432
rect 19852 41392 19892 41432
rect 1612 41224 1652 41264
rect 2860 41224 2900 41264
rect 3244 41224 3284 41264
rect 4492 41224 4532 41264
rect 4972 41224 5012 41264
rect 5068 41224 5108 41264
rect 5260 41224 5300 41264
rect 5644 41224 5684 41264
rect 6892 41224 6932 41264
rect 7084 41224 7124 41264
rect 8332 41224 8372 41264
rect 8908 41224 8948 41264
rect 10156 41224 10196 41264
rect 10732 41224 10772 41264
rect 11980 41224 12020 41264
rect 12364 41224 12404 41264
rect 13612 41224 13652 41264
rect 13996 41224 14036 41264
rect 15244 41224 15284 41264
rect 15628 41224 15668 41264
rect 16876 41224 16916 41264
rect 17068 41224 17108 41264
rect 17260 41224 17300 41264
rect 17356 41224 17396 41264
rect 1228 41140 1268 41180
rect 17740 41140 17780 41180
rect 18124 41140 18164 41180
rect 18508 41140 18548 41180
rect 18892 41140 18932 41180
rect 19276 41140 19316 41180
rect 19660 41140 19700 41180
rect 20044 41140 20084 41180
rect 3052 41056 3092 41096
rect 17932 41056 17972 41096
rect 1420 40972 1460 41012
rect 4684 40972 4724 41012
rect 5260 40972 5300 41012
rect 5452 40972 5492 41012
rect 8524 40972 8564 41012
rect 10348 40972 10388 41012
rect 10540 40972 10580 41012
rect 12172 40972 12212 41012
rect 13804 40972 13844 41012
rect 15436 40972 15476 41012
rect 17068 40972 17108 41012
rect 17548 40972 17588 41012
rect 18316 40972 18356 41012
rect 18700 40972 18740 41012
rect 19084 40972 19124 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 6700 40636 6740 40676
rect 10348 40636 10388 40676
rect 12172 40636 12212 40676
rect 18508 40636 18548 40676
rect 19372 40636 19412 40676
rect 19756 40636 19796 40676
rect 13132 40552 13172 40592
rect 18124 40552 18164 40592
rect 18988 40552 19028 40592
rect 6508 40468 6548 40508
rect 10540 40468 10580 40508
rect 13324 40468 13364 40508
rect 17932 40468 17972 40508
rect 18316 40468 18356 40508
rect 18700 40468 18740 40508
rect 19180 40468 19220 40508
rect 19564 40468 19604 40508
rect 19948 40468 19988 40508
rect 1324 40384 1364 40424
rect 2572 40384 2612 40424
rect 2956 40384 2996 40424
rect 4204 40384 4244 40424
rect 4876 40384 4916 40424
rect 6124 40384 6164 40424
rect 6892 40384 6932 40424
rect 8140 40384 8180 40424
rect 8716 40384 8756 40424
rect 9964 40384 10004 40424
rect 10732 40384 10772 40424
rect 11980 40384 12020 40424
rect 12460 40384 12500 40424
rect 12748 40384 12788 40424
rect 13708 40384 13748 40424
rect 14956 40384 14996 40424
rect 15340 40384 15380 40424
rect 15436 40384 15476 40424
rect 15532 40384 15572 40424
rect 15628 40384 15668 40424
rect 15916 40384 15956 40424
rect 16012 40384 16052 40424
rect 16108 40363 16148 40403
rect 16396 40384 16436 40424
rect 16492 40384 16532 40424
rect 16588 40384 16628 40424
rect 16876 40384 16916 40424
rect 16972 40384 17012 40424
rect 17068 40384 17108 40424
rect 17260 40384 17300 40424
rect 17452 40384 17492 40424
rect 17548 40384 17588 40424
rect 20236 40384 20276 40424
rect 12844 40300 12884 40340
rect 20140 40300 20180 40340
rect 2764 40216 2804 40256
rect 4396 40216 4436 40256
rect 4684 40216 4724 40256
rect 6316 40216 6356 40256
rect 8332 40216 8372 40256
rect 10156 40216 10196 40256
rect 13516 40216 13556 40256
rect 15148 40216 15188 40256
rect 15820 40216 15860 40256
rect 16300 40216 16340 40256
rect 16780 40216 16820 40256
rect 17356 40216 17396 40256
rect 17740 40216 17780 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 7468 39880 7508 39920
rect 8236 39880 8276 39920
rect 18700 39880 18740 39920
rect 19180 39880 19220 39920
rect 19468 39880 19508 39920
rect 19852 39880 19892 39920
rect 6604 39796 6644 39836
rect 10444 39796 10484 39836
rect 12076 39796 12116 39836
rect 17740 39796 17780 39836
rect 1228 39712 1268 39752
rect 2476 39712 2516 39752
rect 3148 39712 3188 39752
rect 4396 39712 4436 39752
rect 4876 39712 4916 39752
rect 4972 39712 5012 39752
rect 5932 39712 5972 39752
rect 6412 39707 6452 39747
rect 8716 39712 8756 39752
rect 8812 39712 8852 39752
rect 9292 39712 9332 39752
rect 9772 39712 9812 39752
rect 10252 39707 10292 39747
rect 10636 39712 10676 39752
rect 11884 39712 11924 39752
rect 12364 39712 12404 39752
rect 12652 39712 12692 39752
rect 12748 39712 12788 39752
rect 13324 39712 13364 39752
rect 14572 39712 14612 39752
rect 14956 39712 14996 39752
rect 15052 39712 15092 39752
rect 15244 39712 15284 39752
rect 15532 39712 15572 39752
rect 15628 39712 15668 39752
rect 15820 39712 15860 39752
rect 16300 39712 16340 39752
rect 17548 39712 17588 39752
rect 19084 39712 19124 39752
rect 19276 39712 19316 39752
rect 5356 39628 5396 39668
rect 5452 39628 5492 39668
rect 6892 39628 6932 39668
rect 7084 39628 7124 39668
rect 7660 39628 7700 39668
rect 7852 39628 7892 39668
rect 8428 39628 8468 39668
rect 9196 39628 9236 39668
rect 16012 39628 16052 39668
rect 17932 39628 17972 39668
rect 18508 39628 18548 39668
rect 18892 39628 18932 39668
rect 19660 39628 19700 39668
rect 20044 39628 20084 39668
rect 2860 39544 2900 39584
rect 7276 39544 7316 39584
rect 13036 39544 13076 39584
rect 18124 39544 18164 39584
rect 2668 39460 2708 39500
rect 4588 39460 4628 39500
rect 8044 39460 8084 39500
rect 14764 39460 14804 39500
rect 15244 39460 15284 39500
rect 15820 39460 15860 39500
rect 18316 39460 18356 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 4972 39040 5012 39080
rect 6700 39040 6740 39080
rect 13900 39014 13940 39054
rect 15340 39040 15380 39080
rect 15532 39040 15572 39080
rect 15724 39040 15764 39080
rect 18412 39040 18452 39080
rect 18892 39040 18932 39080
rect 19852 39040 19892 39080
rect 1324 38956 1364 38996
rect 3340 38956 3380 38996
rect 4396 38956 4436 38996
rect 4780 38956 4820 38996
rect 9196 38956 9236 38996
rect 1708 38914 1748 38954
rect 16300 38956 16340 38996
rect 18316 38956 18356 38996
rect 18508 38956 18548 38996
rect 19084 38956 19124 38996
rect 19468 38956 19508 38996
rect 20044 38956 20084 38996
rect 2956 38872 2996 38912
rect 5260 38872 5300 38912
rect 6508 38872 6548 38912
rect 6892 38872 6932 38912
rect 8140 38872 8180 38912
rect 8620 38872 8660 38912
rect 8716 38872 8756 38912
rect 9100 38872 9140 38912
rect 9676 38872 9716 38912
rect 10156 38886 10196 38926
rect 10540 38872 10580 38912
rect 11788 38872 11828 38912
rect 12364 38872 12404 38912
rect 13612 38872 13652 38912
rect 13900 38864 13940 38904
rect 14284 38872 14324 38912
rect 14380 38872 14420 38912
rect 14476 38872 14516 38912
rect 14572 38872 14612 38912
rect 14764 38872 14804 38912
rect 14860 38872 14900 38912
rect 15052 38872 15092 38912
rect 15340 38872 15380 38912
rect 15724 38872 15764 38912
rect 15916 38872 15956 38912
rect 16012 38872 16052 38912
rect 16204 38872 16244 38912
rect 16396 38872 16436 38912
rect 16588 38872 16628 38912
rect 17836 38872 17876 38912
rect 18220 38872 18260 38912
rect 18604 38872 18644 38912
rect 18796 38872 18836 38912
rect 10348 38788 10388 38828
rect 11980 38788 12020 38828
rect 14956 38788 14996 38828
rect 1516 38704 1556 38744
rect 3148 38704 3188 38744
rect 3532 38704 3572 38744
rect 3820 38704 3860 38744
rect 4012 38704 4052 38744
rect 4588 38704 4628 38744
rect 8332 38704 8372 38744
rect 12172 38704 12212 38744
rect 14092 38704 14132 38744
rect 18028 38704 18068 38744
rect 19276 38704 19316 38744
rect 19660 38704 19700 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 1516 38368 1556 38408
rect 1900 38368 1940 38408
rect 4204 38368 4244 38408
rect 4396 38368 4436 38408
rect 14860 38368 14900 38408
rect 17836 38368 17876 38408
rect 5068 38284 5108 38324
rect 14380 38284 14420 38324
rect 2572 38200 2612 38240
rect 3820 38200 3860 38240
rect 4780 38200 4820 38240
rect 5260 38195 5300 38235
rect 5740 38200 5780 38240
rect 6700 38200 6740 38240
rect 6796 38200 6836 38240
rect 7660 38200 7700 38240
rect 8908 38200 8948 38240
rect 9292 38200 9332 38240
rect 10540 38200 10580 38240
rect 11116 38200 11156 38240
rect 12364 38200 12404 38240
rect 12556 38200 12596 38240
rect 12748 38200 12788 38240
rect 12940 38200 12980 38240
rect 14188 38200 14228 38240
rect 14572 38200 14612 38240
rect 14668 38200 14708 38240
rect 14764 38200 14804 38240
rect 15148 38200 15188 38240
rect 15436 38200 15476 38240
rect 15532 38200 15572 38240
rect 16396 38200 16436 38240
rect 17644 38200 17684 38240
rect 18220 38200 18260 38240
rect 18364 38190 18404 38230
rect 18508 38200 18548 38240
rect 18604 38200 18644 38240
rect 18705 38200 18745 38240
rect 18988 38200 19028 38240
rect 19372 38200 19412 38240
rect 1324 38116 1364 38156
rect 1708 38116 1748 38156
rect 2188 38116 2228 38156
rect 4012 38116 4052 38156
rect 4588 38116 4628 38156
rect 6220 38116 6260 38156
rect 6316 38116 6356 38156
rect 7276 38116 7316 38156
rect 16012 38116 16052 38156
rect 19084 38116 19124 38156
rect 19276 38116 19316 38156
rect 19564 38116 19604 38156
rect 19948 38116 19988 38156
rect 12748 38032 12788 38072
rect 15820 38032 15860 38072
rect 16204 38032 16244 38072
rect 19180 38032 19220 38072
rect 2380 37948 2420 37988
rect 7468 37948 7508 37988
rect 9100 37948 9140 37988
rect 10732 37948 10772 37988
rect 10924 37948 10964 37988
rect 18220 37948 18260 37988
rect 19756 37948 19796 37988
rect 20140 37948 20180 37988
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 1420 37612 1460 37652
rect 7180 37612 7220 37652
rect 9580 37612 9620 37652
rect 9964 37612 10004 37652
rect 13708 37612 13748 37652
rect 14380 37612 14420 37652
rect 14668 37612 14708 37652
rect 16108 37612 16148 37652
rect 17164 37612 17204 37652
rect 18316 37612 18356 37652
rect 18508 37612 18548 37652
rect 20236 37612 20276 37652
rect 4780 37528 4820 37568
rect 15724 37528 15764 37568
rect 1228 37444 1268 37484
rect 3628 37444 3668 37484
rect 4300 37444 4340 37484
rect 4972 37444 5012 37484
rect 6988 37444 7028 37484
rect 9388 37444 9428 37484
rect 9772 37444 9812 37484
rect 15628 37444 15668 37484
rect 15820 37444 15860 37484
rect 17356 37444 17396 37484
rect 1804 37374 1844 37414
rect 2284 37360 2324 37400
rect 2764 37360 2804 37400
rect 2860 37360 2900 37400
rect 3244 37340 3284 37380
rect 3340 37360 3380 37400
rect 5356 37360 5396 37400
rect 6604 37360 6644 37400
rect 7468 37360 7508 37400
rect 7564 37360 7604 37400
rect 7948 37360 7988 37400
rect 8044 37360 8084 37400
rect 8524 37360 8564 37400
rect 9004 37374 9044 37414
rect 10252 37360 10292 37400
rect 10444 37360 10484 37400
rect 11692 37360 11732 37400
rect 12268 37360 12308 37400
rect 13516 37360 13556 37400
rect 13708 37360 13748 37400
rect 13900 37360 13940 37400
rect 14092 37360 14132 37400
rect 14188 37360 14228 37400
rect 14380 37360 14420 37400
rect 14572 37360 14612 37400
rect 14860 37360 14900 37400
rect 14956 37360 14996 37400
rect 15052 37360 15092 37400
rect 15532 37360 15572 37400
rect 15916 37360 15956 37400
rect 16108 37360 16148 37400
rect 16684 37402 16724 37442
rect 19756 37444 19796 37484
rect 16300 37360 16340 37400
rect 16396 37360 16436 37400
rect 16780 37360 16820 37400
rect 16876 37360 16916 37400
rect 17932 37402 17972 37442
rect 17626 37345 17666 37385
rect 18892 37360 18932 37400
rect 19180 37360 19220 37400
rect 19468 37360 19508 37400
rect 20127 37349 20167 37389
rect 18028 37276 18068 37316
rect 18796 37276 18836 37316
rect 1612 37192 1652 37232
rect 3820 37192 3860 37232
rect 4108 37192 4148 37232
rect 4492 37192 4532 37232
rect 5164 37192 5204 37232
rect 6796 37192 6836 37232
rect 9196 37192 9236 37232
rect 10156 37192 10196 37232
rect 11884 37192 11924 37232
rect 12076 37192 12116 37232
rect 15148 37192 15188 37232
rect 16588 37192 16628 37232
rect 19564 37192 19604 37232
rect 19948 37192 19988 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 1516 36856 1556 36896
rect 5740 36856 5780 36896
rect 9388 36856 9428 36896
rect 15532 36856 15572 36896
rect 18124 36856 18164 36896
rect 19276 36856 19316 36896
rect 5164 36772 5204 36812
rect 11788 36772 11828 36812
rect 13804 36772 13844 36812
rect 15916 36772 15956 36812
rect 1708 36688 1748 36728
rect 2956 36667 2996 36707
rect 3436 36688 3476 36728
rect 3532 36708 3572 36748
rect 3916 36688 3956 36728
rect 4492 36688 4532 36728
rect 4972 36683 5012 36723
rect 5932 36688 5972 36728
rect 7180 36688 7220 36728
rect 7660 36688 7700 36728
rect 7756 36688 7796 36728
rect 8140 36688 8180 36728
rect 8716 36688 8756 36728
rect 9196 36683 9236 36723
rect 10060 36688 10100 36728
rect 10156 36688 10196 36728
rect 10540 36688 10580 36728
rect 10636 36688 10676 36728
rect 11116 36688 11156 36728
rect 11596 36674 11636 36714
rect 12076 36688 12116 36728
rect 12172 36688 12212 36728
rect 12556 36688 12596 36728
rect 13132 36688 13172 36728
rect 14092 36688 14132 36728
rect 15340 36688 15380 36728
rect 1324 36604 1364 36644
rect 4012 36604 4052 36644
rect 5548 36604 5588 36644
rect 8236 36604 8276 36644
rect 9580 36604 9620 36644
rect 12652 36604 12692 36644
rect 13660 36646 13700 36686
rect 15916 36665 15956 36705
rect 16012 36688 16052 36728
rect 16204 36673 16244 36713
rect 16300 36688 16340 36728
rect 16457 36673 16497 36713
rect 16684 36688 16724 36728
rect 17068 36688 17108 36728
rect 17260 36688 17300 36728
rect 17452 36688 17492 36728
rect 17836 36688 17876 36728
rect 17932 36688 17972 36728
rect 18124 36688 18164 36728
rect 18316 36688 18356 36728
rect 18508 36688 18548 36728
rect 16780 36604 16820 36644
rect 16972 36604 17012 36644
rect 17356 36604 17396 36644
rect 18412 36604 18452 36644
rect 18700 36604 18740 36644
rect 19084 36604 19124 36644
rect 19468 36604 19508 36644
rect 19852 36604 19892 36644
rect 9772 36520 9812 36560
rect 16876 36520 16916 36560
rect 18892 36520 18932 36560
rect 20044 36520 20084 36560
rect 3148 36436 3188 36476
rect 7372 36436 7412 36476
rect 19660 36436 19700 36476
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 1612 36100 1652 36140
rect 2572 36100 2612 36140
rect 11980 36100 12020 36140
rect 13804 36100 13844 36140
rect 16588 36142 16628 36182
rect 15436 36100 15476 36140
rect 16396 36016 16436 36056
rect 1420 35932 1460 35972
rect 1804 35932 1844 35972
rect 2380 35932 2420 35972
rect 3916 35932 3956 35972
rect 9196 35932 9236 35972
rect 19372 35932 19412 35972
rect 19756 35932 19796 35972
rect 2956 35862 2996 35902
rect 3436 35848 3476 35888
rect 4012 35848 4052 35888
rect 4396 35848 4436 35888
rect 4492 35848 4532 35888
rect 5068 35848 5108 35888
rect 5260 35848 5300 35888
rect 5356 35848 5396 35888
rect 5548 35848 5588 35888
rect 6796 35848 6836 35888
rect 7276 35848 7316 35888
rect 7372 35848 7412 35888
rect 7756 35848 7796 35888
rect 7852 35848 7892 35888
rect 8332 35848 8372 35888
rect 8812 35853 8852 35893
rect 9676 35848 9716 35888
rect 9772 35848 9812 35888
rect 9868 35848 9908 35888
rect 10060 35848 10100 35888
rect 10156 35848 10196 35888
rect 10252 35848 10292 35888
rect 10348 35848 10388 35888
rect 10540 35848 10580 35888
rect 11788 35848 11828 35888
rect 12364 35848 12404 35888
rect 13612 35848 13652 35888
rect 13996 35848 14036 35888
rect 15244 35848 15284 35888
rect 15724 35848 15764 35888
rect 16012 35848 16052 35888
rect 16972 35848 17012 35888
rect 17260 35848 17300 35888
rect 17740 35848 17780 35888
rect 18988 35848 19028 35888
rect 20127 35848 20167 35888
rect 2764 35764 2804 35804
rect 5164 35764 5204 35804
rect 6988 35764 7028 35804
rect 16108 35764 16148 35804
rect 16876 35764 16916 35804
rect 20236 35764 20276 35804
rect 1996 35680 2036 35720
rect 4780 35680 4820 35720
rect 9004 35680 9044 35720
rect 9388 35680 9428 35720
rect 9580 35680 9620 35720
rect 19180 35680 19220 35720
rect 19564 35680 19604 35720
rect 19948 35680 19988 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 9868 35344 9908 35384
rect 7660 35260 7700 35300
rect 12460 35260 12500 35300
rect 17164 35260 17204 35300
rect 19180 35260 19220 35300
rect 1900 35176 1940 35216
rect 3148 35176 3188 35216
rect 4204 35176 4244 35216
rect 5452 35176 5492 35216
rect 5932 35176 5972 35216
rect 6028 35176 6068 35216
rect 6988 35176 7028 35216
rect 7468 35162 7508 35202
rect 7852 35176 7892 35216
rect 8044 35176 8084 35216
rect 8236 35176 8276 35216
rect 9484 35176 9524 35216
rect 10060 35155 10100 35195
rect 11308 35176 11348 35216
rect 11596 35176 11636 35216
rect 12844 35176 12884 35216
rect 13132 35176 13172 35216
rect 13228 35176 13268 35216
rect 13708 35176 13748 35216
rect 14956 35176 14996 35216
rect 15340 35176 15380 35216
rect 15532 35176 15572 35216
rect 15724 35176 15764 35216
rect 16972 35176 17012 35216
rect 17452 35176 17492 35216
rect 17548 35176 17588 35216
rect 18508 35176 18548 35216
rect 19036 35166 19076 35206
rect 1516 35092 1556 35132
rect 3820 35092 3860 35132
rect 6412 35092 6452 35132
rect 6508 35092 6548 35132
rect 17932 35092 17972 35132
rect 18028 35092 18068 35132
rect 19660 35092 19700 35132
rect 19852 35092 19892 35132
rect 1324 35008 1364 35048
rect 1708 35008 1748 35048
rect 3532 35008 3572 35048
rect 4012 35008 4052 35048
rect 5644 35008 5684 35048
rect 19468 35008 19508 35048
rect 3340 34924 3380 34964
rect 7948 34924 7988 34964
rect 9676 34924 9716 34964
rect 13516 34924 13556 34964
rect 15148 34924 15188 34964
rect 15340 34924 15380 34964
rect 20044 34924 20084 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 3340 34588 3380 34628
rect 7180 34588 7220 34628
rect 14476 34588 14516 34628
rect 14668 34588 14708 34628
rect 3148 34407 3188 34447
rect 3676 34378 3716 34418
rect 4684 34420 4724 34460
rect 8428 34420 8468 34460
rect 8524 34420 8564 34460
rect 1324 34336 1364 34376
rect 1516 34336 1556 34376
rect 2764 34336 2804 34376
rect 4204 34336 4244 34376
rect 4780 34336 4820 34376
rect 5164 34336 5204 34376
rect 5260 34336 5300 34376
rect 5740 34336 5780 34376
rect 6988 34336 7028 34376
rect 7468 34315 7508 34355
rect 7564 34315 7604 34355
rect 7660 34336 7700 34376
rect 7948 34336 7988 34376
rect 9532 34378 9572 34418
rect 11500 34420 11540 34460
rect 8044 34336 8084 34376
rect 9004 34336 9044 34376
rect 9964 34336 10004 34376
rect 10060 34336 10100 34376
rect 10156 34336 10196 34376
rect 10348 34336 10388 34376
rect 10444 34336 10484 34376
rect 10540 34336 10580 34376
rect 10924 34336 10964 34376
rect 11020 34336 11060 34376
rect 11404 34336 11444 34376
rect 11980 34336 12020 34376
rect 12460 34341 12500 34381
rect 13036 34336 13076 34376
rect 14284 34336 14324 34376
rect 14668 34336 14708 34376
rect 14860 34336 14900 34376
rect 14956 34336 14996 34376
rect 16684 34336 16724 34376
rect 17068 34336 17108 34376
rect 18316 34336 18356 34376
rect 18700 34336 18740 34376
rect 19948 34357 19988 34397
rect 3532 34252 3572 34292
rect 15436 34294 15476 34334
rect 12652 34252 12692 34292
rect 1228 34168 1268 34208
rect 2956 34168 2996 34208
rect 7372 34168 7412 34208
rect 9676 34168 9716 34208
rect 9868 34168 9908 34208
rect 10636 34168 10676 34208
rect 15148 34168 15188 34208
rect 16876 34168 16916 34208
rect 18508 34168 18548 34208
rect 20140 34168 20180 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 3532 33832 3572 33872
rect 3820 33832 3860 33872
rect 4396 33832 4436 33872
rect 4684 33832 4724 33872
rect 11980 33832 12020 33872
rect 15436 33832 15476 33872
rect 19276 33832 19316 33872
rect 1324 33664 1364 33704
rect 1420 33664 1460 33704
rect 1612 33664 1652 33704
rect 1900 33664 1940 33704
rect 3148 33664 3188 33704
rect 4012 33664 4052 33704
rect 4108 33664 4148 33704
rect 4876 33664 4916 33704
rect 6124 33664 6164 33704
rect 6508 33664 6548 33704
rect 6604 33664 6644 33704
rect 6796 33664 6836 33704
rect 7276 33664 7316 33704
rect 8524 33664 8564 33704
rect 8908 33664 8948 33704
rect 10156 33664 10196 33704
rect 10540 33664 10580 33704
rect 11788 33643 11828 33683
rect 12364 33664 12404 33704
rect 13612 33664 13652 33704
rect 13996 33664 14036 33704
rect 15244 33664 15284 33704
rect 15628 33664 15668 33704
rect 16876 33664 16916 33704
rect 17548 33664 17588 33704
rect 17644 33664 17684 33704
rect 18604 33664 18644 33704
rect 19084 33659 19124 33699
rect 18028 33580 18068 33620
rect 18124 33580 18164 33620
rect 19468 33580 19508 33620
rect 19756 33580 19796 33620
rect 1420 33496 1460 33536
rect 20140 33496 20180 33536
rect 3340 33412 3380 33452
rect 6316 33412 6356 33452
rect 6796 33412 6836 33452
rect 7084 33412 7124 33452
rect 10348 33412 10388 33452
rect 13804 33412 13844 33452
rect 17068 33412 17108 33452
rect 19948 33412 19988 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 2380 33076 2420 33116
rect 10444 33076 10484 33116
rect 11308 33076 11348 33116
rect 16108 33076 16148 33116
rect 19084 33076 19124 33116
rect 4684 32992 4724 33032
rect 12364 32992 12404 33032
rect 20140 32992 20180 33032
rect 2188 32908 2228 32948
rect 3148 32908 3188 32948
rect 1420 32824 1460 32864
rect 1516 32824 1556 32864
rect 1708 32824 1748 32864
rect 1804 32824 1844 32864
rect 1961 32839 2001 32879
rect 2668 32824 2708 32864
rect 2764 32824 2804 32864
rect 3244 32824 3284 32864
rect 3724 32824 3764 32864
rect 4204 32838 4244 32878
rect 6652 32866 6692 32906
rect 14284 32908 14324 32948
rect 19372 32908 19412 32948
rect 19756 32908 19796 32948
rect 4876 32824 4916 32864
rect 6124 32824 6164 32864
rect 7180 32824 7220 32864
rect 7660 32824 7700 32864
rect 7756 32824 7796 32864
rect 8140 32824 8180 32864
rect 8236 32824 8276 32864
rect 8716 32824 8756 32864
rect 8812 32824 8852 32864
rect 9004 32824 9044 32864
rect 10252 32824 10292 32864
rect 10636 32824 10676 32864
rect 11596 32824 11636 32864
rect 11980 32824 12020 32864
rect 12076 32824 12116 32864
rect 12748 32824 12788 32864
rect 12844 32824 12884 32864
rect 13036 32824 13076 32864
rect 13324 32824 13364 32864
rect 13708 32824 13748 32864
rect 13804 32824 13844 32864
rect 14188 32824 14228 32864
rect 14764 32824 14804 32864
rect 15244 32838 15284 32878
rect 15628 32824 15668 32864
rect 15724 32824 15764 32864
rect 15820 32803 15860 32843
rect 15916 32824 15956 32864
rect 16108 32824 16148 32864
rect 16396 32824 16436 32864
rect 16972 32824 17012 32864
rect 4396 32740 4436 32780
rect 6316 32740 6356 32780
rect 13132 32740 13172 32780
rect 15436 32740 15476 32780
rect 16300 32782 16340 32822
rect 17068 32824 17108 32864
rect 17452 32824 17492 32864
rect 17548 32824 17588 32864
rect 18028 32824 18068 32864
rect 18508 32838 18548 32878
rect 18892 32824 18932 32864
rect 19084 32824 19124 32864
rect 18700 32740 18740 32780
rect 1900 32656 1940 32696
rect 8524 32656 8564 32696
rect 10444 32656 10484 32696
rect 6508 32614 6548 32654
rect 12556 32656 12596 32696
rect 19564 32656 19604 32696
rect 19948 32656 19988 32696
rect 11884 32598 11924 32638
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 2860 32320 2900 32360
rect 3244 32320 3284 32360
rect 10540 32320 10580 32360
rect 12268 32320 12308 32360
rect 13132 32320 13172 32360
rect 14476 32320 14516 32360
rect 19180 32320 19220 32360
rect 6700 32236 6740 32276
rect 6892 32236 6932 32276
rect 1228 32152 1268 32192
rect 2476 32152 2516 32192
rect 3436 32147 3476 32187
rect 3916 32152 3956 32192
rect 4876 32152 4916 32192
rect 4972 32152 5012 32192
rect 5260 32152 5300 32192
rect 6508 32152 6548 32192
rect 7084 32147 7124 32187
rect 7564 32152 7604 32192
rect 8044 32152 8084 32192
rect 8524 32152 8564 32192
rect 8620 32152 8660 32192
rect 9100 32152 9140 32192
rect 10348 32152 10388 32192
rect 10828 32152 10868 32192
rect 11116 32152 11156 32192
rect 11212 32152 11252 32192
rect 11692 32152 11732 32192
rect 11884 32152 11924 32192
rect 11980 32152 12020 32192
rect 12172 32152 12212 32192
rect 12364 32152 12404 32192
rect 12460 32152 12500 32192
rect 12652 32152 12692 32192
rect 12748 32152 12788 32192
rect 12940 32152 12980 32192
rect 13324 32152 13364 32192
rect 13708 32152 13748 32192
rect 13996 32152 14036 32192
rect 14380 32152 14420 32192
rect 14572 32152 14612 32192
rect 14668 32152 14708 32192
rect 15052 32152 15092 32192
rect 15148 32152 15188 32192
rect 15244 32152 15284 32192
rect 15340 32152 15380 32192
rect 15532 32152 15572 32192
rect 15724 32152 15764 32192
rect 15820 32152 15860 32192
rect 16204 32152 16244 32192
rect 17452 32131 17492 32171
rect 17836 32152 17876 32192
rect 18028 32152 18068 32192
rect 18220 32152 18260 32192
rect 18412 32152 18452 32192
rect 3052 32068 3092 32108
rect 4396 32068 4436 32108
rect 4492 32068 4532 32108
rect 8140 32068 8180 32108
rect 18604 32068 18644 32108
rect 18988 32068 19028 32108
rect 19372 32068 19412 32108
rect 19756 32068 19796 32108
rect 11500 31984 11540 32024
rect 13324 31984 13364 32024
rect 13996 31984 14036 32024
rect 18028 31984 18068 32024
rect 18220 31984 18260 32024
rect 2668 31900 2708 31940
rect 11692 31900 11732 31940
rect 12940 31900 12980 31940
rect 15532 31900 15572 31940
rect 17644 31900 17684 31940
rect 18796 31900 18836 31940
rect 19564 31900 19604 31940
rect 19948 31900 19988 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 4588 31564 4628 31604
rect 4780 31564 4820 31604
rect 17068 31564 17108 31604
rect 8044 31480 8084 31520
rect 8428 31480 8468 31520
rect 8812 31480 8852 31520
rect 10540 31480 10580 31520
rect 16300 31480 16340 31520
rect 8332 31396 8372 31436
rect 8524 31396 8564 31436
rect 13132 31396 13172 31436
rect 18028 31396 18068 31436
rect 1228 31312 1268 31352
rect 2476 31312 2516 31352
rect 3148 31312 3188 31352
rect 4396 31312 4436 31352
rect 4972 31312 5012 31352
rect 6220 31312 6260 31352
rect 6604 31312 6644 31352
rect 7852 31312 7892 31352
rect 8236 31312 8276 31352
rect 8620 31312 8660 31352
rect 9100 31312 9140 31352
rect 10348 31312 10388 31352
rect 10924 31312 10964 31352
rect 12172 31312 12212 31352
rect 12652 31312 12692 31352
rect 12748 31312 12788 31352
rect 13228 31312 13268 31352
rect 13708 31312 13748 31352
rect 14188 31317 14228 31357
rect 14860 31312 14900 31352
rect 16108 31312 16148 31352
rect 16492 31312 16532 31352
rect 16684 31354 16724 31394
rect 18124 31396 18164 31436
rect 19468 31396 19508 31436
rect 19852 31396 19892 31436
rect 16588 31312 16628 31352
rect 16972 31312 17012 31352
rect 17164 31299 17204 31339
rect 17548 31312 17588 31352
rect 17644 31312 17684 31352
rect 18604 31312 18644 31352
rect 19132 31321 19172 31361
rect 12364 31228 12404 31268
rect 14380 31228 14420 31268
rect 19276 31228 19316 31268
rect 2668 31144 2708 31184
rect 2956 31144 2996 31184
rect 4588 31144 4628 31184
rect 16780 31144 16820 31184
rect 19660 31144 19700 31184
rect 20044 31144 20084 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 1420 30808 1460 30848
rect 4876 30808 4916 30848
rect 7948 30808 7988 30848
rect 12364 30808 12404 30848
rect 13996 30808 14036 30848
rect 16108 30808 16148 30848
rect 19660 30808 19700 30848
rect 1612 30640 1652 30680
rect 2860 30640 2900 30680
rect 3436 30640 3476 30680
rect 4684 30640 4724 30680
rect 5356 30640 5396 30680
rect 5644 30640 5684 30680
rect 5740 30640 5780 30680
rect 6220 30640 6260 30680
rect 6508 30640 6548 30680
rect 7756 30640 7796 30680
rect 9100 30640 9140 30680
rect 9388 30640 9428 30680
rect 9772 30640 9812 30680
rect 9964 30640 10004 30680
rect 11212 30640 11252 30680
rect 11596 30640 11636 30680
rect 11980 30640 12020 30680
rect 12556 30640 12596 30680
rect 13804 30640 13844 30680
rect 14380 30640 14420 30680
rect 14476 30640 14516 30680
rect 14860 30640 14900 30680
rect 15436 30640 15476 30680
rect 15916 30635 15956 30675
rect 16300 30640 16340 30680
rect 17548 30640 17588 30680
rect 18220 30640 18260 30680
rect 19468 30640 19508 30680
rect 1228 30556 1268 30596
rect 5068 30556 5108 30596
rect 9484 30556 9524 30596
rect 9676 30556 9716 30596
rect 11692 30556 11732 30596
rect 11884 30556 11924 30596
rect 12172 30556 12212 30596
rect 14956 30556 14996 30596
rect 19852 30556 19892 30596
rect 9580 30472 9620 30512
rect 11788 30472 11828 30512
rect 3052 30388 3092 30428
rect 3244 30388 3284 30428
rect 6028 30388 6068 30428
rect 6316 30388 6356 30428
rect 8620 30388 8660 30428
rect 11404 30388 11444 30428
rect 17740 30388 17780 30428
rect 20044 30388 20084 30428
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 9868 30052 9908 30092
rect 12940 30052 12980 30092
rect 16204 30052 16244 30092
rect 16396 30052 16436 30092
rect 17068 30052 17108 30092
rect 8140 29968 8180 30008
rect 9196 29968 9236 30008
rect 11788 29968 11828 30008
rect 12748 29884 12788 29924
rect 17836 29884 17876 29924
rect 19372 29884 19412 29924
rect 19756 29884 19796 29924
rect 1324 29800 1364 29840
rect 1516 29800 1556 29840
rect 2764 29800 2804 29840
rect 3340 29800 3380 29840
rect 4588 29800 4628 29840
rect 5068 29800 5108 29840
rect 6316 29800 6356 29840
rect 6700 29800 6740 29840
rect 7948 29800 7988 29840
rect 8524 29800 8564 29840
rect 8812 29800 8852 29840
rect 9484 29800 9524 29840
rect 9580 29800 9620 29840
rect 10156 29800 10196 29840
rect 11404 29800 11444 29840
rect 12172 29800 12212 29840
rect 12460 29800 12500 29840
rect 13132 29800 13172 29840
rect 14380 29800 14420 29840
rect 14764 29800 14804 29840
rect 16012 29800 16052 29840
rect 16396 29800 16436 29840
rect 16588 29800 16628 29840
rect 16684 29800 16724 29840
rect 16876 29800 16916 29840
rect 17068 29800 17108 29840
rect 17356 29800 17396 29840
rect 17452 29800 17492 29840
rect 17932 29800 17972 29840
rect 18412 29800 18452 29840
rect 18940 29809 18980 29849
rect 8908 29716 8948 29756
rect 12076 29716 12116 29756
rect 14572 29716 14612 29756
rect 19084 29716 19124 29756
rect 1228 29632 1268 29672
rect 2956 29632 2996 29672
rect 3148 29632 3188 29672
rect 4876 29632 4916 29672
rect 9388 29628 9428 29668
rect 11596 29632 11636 29672
rect 19564 29632 19604 29672
rect 19948 29632 19988 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 15532 29296 15572 29336
rect 18988 29296 19028 29336
rect 12460 29212 12500 29252
rect 1228 29128 1268 29168
rect 2476 29128 2516 29168
rect 3244 29128 3284 29168
rect 4492 29128 4532 29168
rect 4876 29128 4916 29168
rect 6124 29128 6164 29168
rect 6508 29128 6548 29168
rect 7756 29128 7796 29168
rect 8140 29128 8180 29168
rect 8236 29128 8276 29168
rect 8428 29128 8468 29168
rect 8620 29128 8660 29168
rect 9868 29128 9908 29168
rect 10348 29128 10388 29168
rect 11596 29128 11636 29168
rect 12076 29128 12116 29168
rect 12364 29128 12404 29168
rect 12940 29128 12980 29168
rect 13324 29128 13364 29168
rect 13708 29128 13748 29168
rect 14956 29128 14996 29168
rect 15340 29128 15380 29168
rect 15628 29128 15668 29168
rect 15820 29128 15860 29168
rect 17068 29128 17108 29168
rect 17548 29128 17588 29168
rect 18796 29128 18836 29168
rect 2860 29044 2900 29084
rect 13036 29044 13076 29084
rect 13228 29044 13268 29084
rect 19372 29044 19412 29084
rect 19756 29044 19796 29084
rect 3052 28960 3092 29000
rect 11788 28960 11828 29000
rect 13132 28960 13172 29000
rect 19948 28960 19988 29000
rect 2668 28876 2708 28916
rect 4684 28876 4724 28916
rect 6316 28876 6356 28916
rect 7948 28876 7988 28916
rect 8428 28876 8468 28916
rect 10060 28876 10100 28916
rect 12748 28876 12788 28916
rect 15148 28876 15188 28916
rect 17260 28876 17300 28916
rect 19564 28876 19604 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 4204 28540 4244 28580
rect 7084 28540 7124 28580
rect 11308 28540 11348 28580
rect 12940 28540 12980 28580
rect 3820 28456 3860 28496
rect 12748 28456 12788 28496
rect 3628 28372 3668 28412
rect 4012 28372 4052 28412
rect 4588 28372 4628 28412
rect 6892 28372 6932 28412
rect 19372 28372 19412 28412
rect 19756 28372 19796 28412
rect 1228 28288 1268 28328
rect 2476 28288 2516 28328
rect 2857 28284 2897 28324
rect 2956 28288 2996 28328
rect 3148 28288 3188 28328
rect 3244 28288 3284 28328
rect 3345 28288 3385 28328
rect 5260 28288 5300 28328
rect 6508 28288 6548 28328
rect 7276 28288 7316 28328
rect 8524 28288 8564 28328
rect 9004 28288 9044 28328
rect 9196 28288 9236 28328
rect 10444 28288 10484 28328
rect 11020 28288 11060 28328
rect 11116 28288 11156 28328
rect 11308 28288 11348 28328
rect 11500 28288 11540 28328
rect 11596 28288 11636 28328
rect 11692 28288 11732 28328
rect 12076 28288 12116 28328
rect 12364 28288 12404 28328
rect 12940 28288 12980 28328
rect 13132 28288 13172 28328
rect 13228 28288 13268 28328
rect 13516 28288 13556 28328
rect 14764 28288 14804 28328
rect 15244 28288 15284 28328
rect 15340 28288 15380 28328
rect 15724 28288 15764 28328
rect 15820 28288 15860 28328
rect 16300 28288 16340 28328
rect 16780 28293 16820 28333
rect 17260 28288 17300 28328
rect 17356 28288 17396 28328
rect 17740 28288 17780 28328
rect 17836 28288 17876 28328
rect 18316 28288 18356 28328
rect 18796 28293 18836 28333
rect 12460 28204 12500 28244
rect 16972 28204 17012 28244
rect 18988 28204 19028 28244
rect 2668 28120 2708 28160
rect 3244 28120 3284 28160
rect 4876 28120 4916 28160
rect 6700 28120 6740 28160
rect 8716 28120 8756 28160
rect 8908 28120 8948 28160
rect 10636 28120 10676 28160
rect 11788 28120 11828 28160
rect 14956 28120 14996 28160
rect 19564 28120 19604 28160
rect 19948 28120 19988 28160
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 11884 27784 11924 27824
rect 12748 27784 12788 27824
rect 16780 27784 16820 27824
rect 5548 27700 5588 27740
rect 6796 27700 6836 27740
rect 8812 27700 8852 27740
rect 9100 27700 9140 27740
rect 9772 27700 9812 27740
rect 15148 27700 15188 27740
rect 19276 27700 19316 27740
rect 1324 27616 1364 27656
rect 1420 27616 1460 27656
rect 1612 27616 1652 27656
rect 1804 27616 1844 27656
rect 3052 27616 3092 27656
rect 3820 27616 3860 27656
rect 3916 27616 3956 27656
rect 4876 27616 4916 27656
rect 5356 27611 5396 27651
rect 6028 27616 6068 27656
rect 6124 27616 6164 27656
rect 6412 27616 6452 27656
rect 6700 27616 6740 27656
rect 7084 27616 7124 27656
rect 7180 27616 7220 27656
rect 8140 27616 8180 27656
rect 8668 27606 8708 27646
rect 9004 27616 9044 27656
rect 9196 27616 9236 27656
rect 9292 27616 9332 27656
rect 9484 27616 9524 27656
rect 9580 27616 9620 27656
rect 9676 27616 9716 27656
rect 10156 27616 10196 27656
rect 11404 27616 11444 27656
rect 11788 27616 11828 27656
rect 11980 27616 12020 27656
rect 12076 27616 12116 27656
rect 12460 27616 12500 27656
rect 12556 27616 12596 27656
rect 13420 27597 13460 27637
rect 13516 27616 13556 27656
rect 14476 27616 14516 27656
rect 14956 27611 14996 27651
rect 15340 27616 15380 27656
rect 16588 27616 16628 27656
rect 17836 27616 17876 27656
rect 19084 27616 19124 27656
rect 4300 27532 4340 27572
rect 4396 27532 4436 27572
rect 7564 27532 7604 27572
rect 7660 27532 7700 27572
rect 12940 27532 12980 27572
rect 13900 27532 13940 27572
rect 13996 27532 14036 27572
rect 17068 27532 17108 27572
rect 17452 27532 17492 27572
rect 19468 27532 19508 27572
rect 19852 27532 19892 27572
rect 3436 27448 3476 27488
rect 5740 27448 5780 27488
rect 13132 27448 13172 27488
rect 17260 27448 17300 27488
rect 17644 27448 17684 27488
rect 1612 27364 1652 27404
rect 3244 27364 3284 27404
rect 11596 27364 11636 27404
rect 19660 27364 19700 27404
rect 20044 27364 20084 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 8716 27028 8756 27068
rect 9196 27028 9236 27068
rect 13420 27028 13460 27068
rect 15532 27028 15572 27068
rect 6412 26944 6452 26984
rect 9772 26944 9812 26984
rect 17164 26944 17204 26984
rect 10540 26860 10580 26900
rect 10636 26860 10676 26900
rect 15340 26860 15380 26900
rect 19372 26860 19412 26900
rect 19756 26860 19796 26900
rect 1228 26776 1268 26816
rect 1324 26776 1364 26816
rect 1804 26776 1844 26816
rect 1900 26776 1940 26816
rect 2284 26776 2324 26816
rect 2380 26776 2420 26816
rect 2860 26776 2900 26816
rect 3388 26785 3428 26825
rect 4012 26776 4052 26816
rect 4108 26776 4148 26816
rect 4204 26776 4244 26816
rect 4300 26776 4340 26816
rect 4684 26776 4724 26816
rect 5932 26776 5972 26816
rect 6700 26776 6740 26816
rect 6796 26776 6836 26816
rect 7180 26776 7220 26816
rect 7276 26776 7316 26816
rect 7756 26776 7796 26816
rect 8236 26790 8276 26830
rect 8716 26776 8756 26816
rect 9004 26776 9044 26816
rect 9196 26776 9236 26816
rect 9388 26776 9428 26816
rect 9484 26776 9524 26816
rect 9676 26776 9716 26816
rect 10060 26776 10100 26816
rect 10156 26776 10196 26816
rect 11116 26776 11156 26816
rect 11596 26790 11636 26830
rect 11980 26776 12020 26816
rect 13228 26776 13268 26816
rect 13612 26776 13652 26816
rect 14860 26776 14900 26816
rect 15724 26776 15764 26816
rect 16972 26776 17012 26816
rect 17452 26776 17492 26816
rect 17548 26776 17588 26816
rect 17932 26776 17972 26816
rect 18028 26776 18068 26816
rect 18508 26776 18548 26816
rect 19036 26785 19076 26825
rect 3532 26692 3572 26732
rect 11788 26692 11828 26732
rect 1516 26608 1556 26648
rect 3820 26608 3860 26648
rect 6124 26608 6164 26648
rect 8428 26608 8468 26648
rect 15052 26608 15092 26648
rect 19180 26608 19220 26648
rect 19564 26608 19604 26648
rect 19948 26608 19988 26648
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 1420 26272 1460 26312
rect 4492 26272 4532 26312
rect 10924 26272 10964 26312
rect 14572 26272 14612 26312
rect 19564 26272 19604 26312
rect 3532 26188 3572 26228
rect 5356 26188 5396 26228
rect 7276 26188 7316 26228
rect 12556 26188 12596 26228
rect 1228 26104 1268 26144
rect 1324 26104 1364 26144
rect 1516 26104 1556 26144
rect 1804 26104 1844 26144
rect 1900 26104 1940 26144
rect 2284 26104 2324 26144
rect 2860 26104 2900 26144
rect 3340 26099 3380 26139
rect 4972 26104 5012 26144
rect 5260 26104 5300 26144
rect 5836 26104 5876 26144
rect 7084 26104 7124 26144
rect 7468 26104 7508 26144
rect 8716 26104 8756 26144
rect 9196 26104 9236 26144
rect 9292 26104 9332 26144
rect 9676 26104 9716 26144
rect 10252 26104 10292 26144
rect 10732 26099 10772 26139
rect 11116 26104 11156 26144
rect 12364 26104 12404 26144
rect 12844 26104 12884 26144
rect 12940 26104 12980 26144
rect 13324 26104 13364 26144
rect 13420 26104 13460 26144
rect 13900 26104 13940 26144
rect 14380 26090 14420 26130
rect 14956 26104 14996 26144
rect 16204 26104 16244 26144
rect 16396 26104 16436 26144
rect 17644 26104 17684 26144
rect 18124 26104 18164 26144
rect 19372 26104 19412 26144
rect 2380 26020 2420 26060
rect 4204 26020 4244 26060
rect 4684 26020 4724 26060
rect 9772 26020 9812 26060
rect 19756 26020 19796 26060
rect 3820 25936 3860 25976
rect 5644 25936 5684 25976
rect 4012 25852 4052 25892
rect 8908 25852 8948 25892
rect 14764 25852 14804 25892
rect 17836 25852 17876 25892
rect 19948 25852 19988 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 2860 25516 2900 25556
rect 6220 25516 6260 25556
rect 10540 25516 10580 25556
rect 12556 25516 12596 25556
rect 14668 25516 14708 25556
rect 3052 25348 3092 25388
rect 4684 25348 4724 25388
rect 6028 25348 6068 25388
rect 10348 25348 10388 25388
rect 12364 25348 12404 25388
rect 14476 25348 14516 25388
rect 15532 25348 15572 25388
rect 19372 25348 19412 25388
rect 19756 25348 19796 25388
rect 1228 25264 1268 25304
rect 2476 25264 2516 25304
rect 3628 25269 3668 25309
rect 4108 25264 4148 25304
rect 4588 25264 4628 25304
rect 5068 25264 5108 25304
rect 5164 25264 5204 25304
rect 5548 25264 5588 25304
rect 5644 25264 5684 25304
rect 6412 25264 6452 25304
rect 7660 25264 7700 25304
rect 8044 25264 8084 25304
rect 9292 25264 9332 25304
rect 10732 25264 10772 25304
rect 11980 25264 12020 25304
rect 12748 25264 12788 25304
rect 13996 25264 14036 25304
rect 14956 25264 14996 25304
rect 15052 25264 15092 25304
rect 15436 25264 15476 25304
rect 16012 25264 16052 25304
rect 16540 25273 16580 25313
rect 17260 25264 17300 25304
rect 17356 25264 17396 25304
rect 17740 25264 17780 25304
rect 17836 25264 17876 25304
rect 18316 25264 18356 25304
rect 18796 25269 18836 25309
rect 3436 25180 3476 25220
rect 16684 25180 16724 25220
rect 18988 25180 19028 25220
rect 2668 25096 2708 25136
rect 5836 25096 5876 25136
rect 7852 25096 7892 25136
rect 9484 25096 9524 25136
rect 12172 25096 12212 25136
rect 14188 25096 14228 25136
rect 19564 25096 19604 25136
rect 19948 25096 19988 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 12172 24760 12212 24800
rect 14476 24760 14516 24800
rect 14956 24760 14996 24800
rect 16588 24760 16628 24800
rect 17260 24760 17300 24800
rect 19276 24760 19316 24800
rect 8140 24676 8180 24716
rect 1228 24592 1268 24632
rect 2476 24592 2516 24632
rect 3052 24592 3092 24632
rect 4300 24592 4340 24632
rect 4684 24592 4724 24632
rect 5932 24592 5972 24632
rect 6412 24592 6452 24632
rect 6508 24592 6548 24632
rect 6892 24592 6932 24632
rect 7468 24592 7508 24632
rect 7948 24587 7988 24627
rect 8716 24592 8756 24632
rect 9964 24592 10004 24632
rect 10444 24592 10484 24632
rect 10540 24592 10580 24632
rect 11500 24592 11540 24632
rect 12460 24592 12500 24632
rect 12748 24592 12788 24632
rect 6988 24508 7028 24548
rect 10924 24508 10964 24548
rect 11020 24508 11060 24548
rect 12028 24550 12068 24590
rect 12844 24592 12884 24632
rect 13804 24592 13844 24632
rect 14284 24587 14324 24627
rect 15148 24592 15188 24632
rect 16396 24592 16436 24632
rect 17836 24592 17876 24632
rect 19084 24592 19124 24632
rect 19852 24592 19892 24632
rect 20044 24592 20084 24632
rect 12364 24508 12404 24548
rect 13228 24508 13268 24548
rect 13324 24508 13364 24548
rect 14764 24508 14804 24548
rect 17068 24508 17108 24548
rect 17452 24508 17492 24548
rect 19468 24508 19508 24548
rect 17644 24424 17684 24464
rect 2668 24340 2708 24380
rect 4492 24340 4532 24380
rect 6124 24340 6164 24380
rect 10156 24340 10196 24380
rect 19660 24340 19700 24380
rect 19852 24340 19892 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 12748 24004 12788 24044
rect 13228 24004 13268 24044
rect 13612 24004 13652 24044
rect 19756 24004 19796 24044
rect 13996 23920 14036 23960
rect 14380 23920 14420 23960
rect 14764 23920 14804 23960
rect 19372 23920 19412 23960
rect 6700 23836 6740 23876
rect 9772 23836 9812 23876
rect 13036 23836 13076 23876
rect 13420 23836 13460 23876
rect 13804 23836 13844 23876
rect 14188 23836 14228 23876
rect 14572 23836 14612 23876
rect 15532 23836 15572 23876
rect 19948 23836 19988 23876
rect 1420 23752 1460 23792
rect 1516 23752 1556 23792
rect 1612 23752 1652 23792
rect 1900 23752 1940 23792
rect 1996 23752 2036 23792
rect 2092 23752 2132 23792
rect 2284 23752 2324 23792
rect 3532 23752 3572 23792
rect 4300 23752 4340 23792
rect 5548 23752 5588 23792
rect 6124 23752 6164 23792
rect 6220 23752 6260 23792
rect 6604 23752 6644 23792
rect 7180 23752 7220 23792
rect 7660 23766 7700 23806
rect 9292 23752 9332 23792
rect 9388 23752 9428 23792
rect 9868 23752 9908 23792
rect 10348 23752 10388 23792
rect 10828 23766 10868 23806
rect 11308 23752 11348 23792
rect 12556 23752 12596 23792
rect 15052 23752 15092 23792
rect 15148 23752 15188 23792
rect 15628 23752 15668 23792
rect 16108 23752 16148 23792
rect 16636 23761 16676 23801
rect 17260 23757 17300 23797
rect 17740 23752 17780 23792
rect 18220 23752 18260 23792
rect 18316 23752 18356 23792
rect 18700 23752 18740 23792
rect 18796 23752 18836 23792
rect 19084 23752 19124 23792
rect 19180 23752 19220 23792
rect 19372 23752 19412 23792
rect 19564 23752 19604 23792
rect 19756 23752 19796 23792
rect 11020 23668 11060 23708
rect 16780 23668 16820 23708
rect 1324 23584 1364 23624
rect 1804 23584 1844 23624
rect 3724 23584 3764 23624
rect 4012 23584 4052 23624
rect 5740 23584 5780 23624
rect 7852 23584 7892 23624
rect 17068 23584 17108 23624
rect 20140 23584 20180 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 1516 23248 1556 23288
rect 3628 23248 3668 23288
rect 6604 23248 6644 23288
rect 13324 23248 13364 23288
rect 14956 23248 14996 23288
rect 16684 23248 16724 23288
rect 17068 23248 17108 23288
rect 19468 23248 19508 23288
rect 5836 23164 5876 23204
rect 1708 23080 1748 23120
rect 2956 23080 2996 23120
rect 3340 23080 3380 23120
rect 3436 23080 3476 23120
rect 4108 23080 4148 23120
rect 4204 23080 4244 23120
rect 4684 23080 4724 23120
rect 5164 23080 5204 23120
rect 5692 23070 5732 23110
rect 7084 23080 7124 23120
rect 8332 23080 8372 23120
rect 9484 23080 9524 23120
rect 10732 23080 10772 23120
rect 11404 23080 11444 23120
rect 12652 23080 12692 23120
rect 13516 23080 13556 23120
rect 14764 23080 14804 23120
rect 15244 23080 15284 23120
rect 16492 23080 16532 23120
rect 16972 23080 17012 23120
rect 17164 23080 17204 23120
rect 17356 23080 17396 23120
rect 18604 23080 18644 23120
rect 18988 23080 19028 23120
rect 19180 23080 19220 23120
rect 19276 23080 19316 23120
rect 19564 23080 19604 23120
rect 19660 23080 19700 23120
rect 19756 23080 19796 23120
rect 19948 23069 19988 23109
rect 20140 23080 20180 23120
rect 20236 23080 20276 23120
rect 1324 22996 1364 23036
rect 4588 22996 4628 23036
rect 6028 22996 6068 23036
rect 6412 22996 6452 23036
rect 13132 22996 13172 23036
rect 3148 22828 3188 22868
rect 6220 22828 6260 22868
rect 8524 22828 8564 22868
rect 10924 22828 10964 22868
rect 12844 22828 12884 22868
rect 18796 22828 18836 22868
rect 19948 22828 19988 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 1516 22492 1556 22532
rect 1708 22492 1748 22532
rect 4492 22492 4532 22532
rect 13516 22492 13556 22532
rect 19276 22492 19316 22532
rect 4108 22408 4148 22448
rect 4684 22408 4724 22448
rect 1324 22324 1364 22364
rect 1900 22324 1940 22364
rect 4300 22324 4340 22364
rect 7276 22324 7316 22364
rect 2380 22282 2420 22322
rect 3628 22240 3668 22280
rect 4972 22240 5012 22280
rect 6220 22240 6260 22280
rect 6700 22240 6740 22280
rect 6796 22240 6836 22280
rect 8284 22282 8324 22322
rect 9676 22324 9716 22364
rect 13324 22324 13364 22364
rect 19948 22324 19988 22364
rect 7180 22240 7220 22280
rect 7756 22240 7796 22280
rect 9196 22240 9236 22280
rect 9292 22240 9332 22280
rect 9772 22240 9812 22280
rect 10252 22240 10292 22280
rect 10780 22249 10820 22289
rect 11212 22240 11252 22280
rect 11308 22240 11348 22280
rect 11692 22240 11732 22280
rect 11788 22240 11828 22280
rect 12268 22240 12308 22280
rect 12748 22254 12788 22294
rect 13804 22240 13844 22280
rect 13900 22240 13940 22280
rect 14284 22240 14324 22280
rect 14380 22240 14420 22280
rect 14860 22240 14900 22280
rect 15340 22245 15380 22285
rect 15916 22240 15956 22280
rect 17164 22240 17204 22280
rect 17548 22240 17588 22280
rect 17836 22240 17876 22280
rect 19084 22240 19124 22280
rect 19468 22240 19508 22280
rect 19564 22240 19604 22280
rect 19660 22240 19700 22280
rect 19756 22240 19796 22280
rect 2188 22156 2228 22196
rect 15532 22156 15572 22196
rect 17356 22156 17396 22196
rect 3820 22072 3860 22112
rect 6412 22072 6452 22112
rect 8428 22072 8468 22112
rect 10924 22072 10964 22112
rect 12940 22072 12980 22112
rect 17644 22072 17684 22112
rect 20140 22072 20180 22112
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 1516 21736 1556 21776
rect 1900 21736 1940 21776
rect 2284 21736 2324 21776
rect 4300 21736 4340 21776
rect 9484 21736 9524 21776
rect 11116 21736 11156 21776
rect 13708 21736 13748 21776
rect 15340 21736 15380 21776
rect 7852 21652 7892 21692
rect 18604 21652 18644 21692
rect 2572 21568 2612 21608
rect 2668 21568 2708 21608
rect 3052 21568 3092 21608
rect 3148 21568 3188 21608
rect 3628 21568 3668 21608
rect 4108 21563 4148 21603
rect 4588 21568 4628 21608
rect 4876 21568 4916 21608
rect 4972 21568 5012 21608
rect 6124 21568 6164 21608
rect 6220 21568 6260 21608
rect 6604 21568 6644 21608
rect 7180 21568 7220 21608
rect 7660 21563 7700 21603
rect 8044 21568 8084 21608
rect 9292 21568 9332 21608
rect 9676 21568 9716 21608
rect 10924 21568 10964 21608
rect 12268 21568 12308 21608
rect 13516 21568 13556 21608
rect 13900 21568 13940 21608
rect 15148 21568 15188 21608
rect 15532 21568 15572 21608
rect 16780 21568 16820 21608
rect 17164 21568 17204 21608
rect 18412 21568 18452 21608
rect 18796 21568 18836 21608
rect 19084 21575 19124 21615
rect 19276 21568 19316 21608
rect 19372 21568 19412 21608
rect 19468 21568 19508 21608
rect 19564 21568 19604 21608
rect 19756 21568 19796 21608
rect 19948 21568 19988 21608
rect 20044 21568 20084 21608
rect 1324 21484 1364 21524
rect 1708 21484 1748 21524
rect 2092 21484 2132 21524
rect 6700 21484 6740 21524
rect 5260 21400 5300 21440
rect 19756 21400 19796 21440
rect 16972 21316 17012 21356
rect 19084 21316 19124 21356
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 1516 20980 1556 21020
rect 6796 20980 6836 21020
rect 15340 20980 15380 21020
rect 4492 20896 4532 20936
rect 5164 20896 5204 20936
rect 15724 20896 15764 20936
rect 19276 20896 19316 20936
rect 20044 20896 20084 20936
rect 1324 20812 1364 20852
rect 2860 20812 2900 20852
rect 2956 20812 2996 20852
rect 4300 20812 4340 20852
rect 13516 20812 13556 20852
rect 2380 20728 2420 20768
rect 3964 20770 4004 20810
rect 15148 20812 15188 20852
rect 16972 20812 17012 20852
rect 17068 20812 17108 20852
rect 19180 20812 19220 20852
rect 19372 20812 19412 20852
rect 2476 20728 2516 20768
rect 3436 20728 3476 20768
rect 5356 20728 5396 20768
rect 6604 20728 6644 20768
rect 8044 20728 8084 20768
rect 9292 20728 9332 20768
rect 9676 20728 9716 20768
rect 10924 20728 10964 20768
rect 11308 20728 11348 20768
rect 12556 20728 12596 20768
rect 13036 20728 13076 20768
rect 13132 20728 13172 20768
rect 13612 20728 13652 20768
rect 14092 20728 14132 20768
rect 14620 20737 14660 20777
rect 15532 20728 15572 20768
rect 15724 20728 15764 20768
rect 15916 20728 15956 20768
rect 16012 20728 16052 20768
rect 16204 20728 16244 20768
rect 16492 20728 16532 20768
rect 16588 20728 16628 20768
rect 17548 20728 17588 20768
rect 18028 20742 18068 20782
rect 18508 20728 18548 20768
rect 18604 20728 18644 20768
rect 18700 20728 18740 20768
rect 19084 20728 19124 20768
rect 19468 20728 19508 20768
rect 19660 20728 19700 20768
rect 19852 20728 19892 20768
rect 20044 20728 20084 20768
rect 20236 20728 20276 20768
rect 4108 20644 4148 20684
rect 12748 20644 12788 20684
rect 18220 20644 18260 20684
rect 1708 20560 1748 20600
rect 9484 20560 9524 20600
rect 11116 20560 11156 20600
rect 14764 20560 14804 20600
rect 16204 20560 16244 20600
rect 18412 20560 18452 20600
rect 19756 20560 19796 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 12652 20224 12692 20264
rect 18028 20224 18068 20264
rect 2956 20140 2996 20180
rect 6892 20140 6932 20180
rect 7084 20140 7124 20180
rect 11692 20140 11732 20180
rect 14764 20140 14804 20180
rect 17452 20140 17492 20180
rect 1516 20056 1556 20096
rect 2764 20056 2804 20096
rect 3148 20056 3188 20096
rect 4396 20056 4436 20096
rect 5164 20056 5204 20096
rect 5260 20056 5300 20096
rect 6220 20056 6260 20096
rect 6700 20042 6740 20082
rect 7276 20042 7316 20082
rect 7756 20056 7796 20096
rect 8716 20056 8756 20096
rect 8812 20056 8852 20096
rect 9964 20056 10004 20096
rect 10060 20056 10100 20096
rect 11020 20056 11060 20096
rect 11500 20051 11540 20091
rect 12172 20056 12212 20096
rect 12268 20056 12308 20096
rect 12460 20056 12500 20096
rect 12556 20056 12596 20096
rect 12713 20041 12753 20081
rect 13036 20056 13076 20096
rect 13132 20056 13172 20096
rect 14092 20056 14132 20096
rect 4876 19972 4916 20012
rect 5644 19972 5684 20012
rect 5740 19972 5780 20012
rect 8236 19972 8276 20012
rect 8332 19972 8372 20012
rect 10444 19972 10484 20012
rect 10540 19972 10580 20012
rect 13516 19972 13556 20012
rect 13612 19972 13652 20012
rect 14620 20014 14660 20054
rect 14956 20056 14996 20096
rect 15148 20056 15188 20096
rect 15436 20056 15476 20096
rect 15820 20056 15860 20096
rect 16012 20056 16052 20096
rect 17260 20056 17300 20096
rect 17836 20056 17876 20096
rect 17932 20056 17972 20096
rect 18124 20056 18164 20096
rect 18700 20056 18740 20096
rect 15532 19972 15572 20012
rect 18316 20014 18356 20054
rect 19180 20056 19220 20096
rect 19276 20056 19316 20096
rect 19564 20056 19604 20096
rect 19852 20056 19892 20096
rect 19948 20056 19988 20096
rect 15724 19972 15764 20012
rect 18412 19972 18452 20012
rect 20140 20014 20180 20054
rect 18604 19972 18644 20012
rect 1324 19888 1364 19928
rect 4588 19888 4628 19928
rect 15628 19888 15668 19928
rect 18892 19888 18932 19928
rect 15148 19804 15188 19844
rect 18508 19846 18548 19886
rect 19948 19804 19988 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 1708 19468 1748 19508
rect 7372 19468 7412 19508
rect 13036 19468 13076 19508
rect 14764 19468 14804 19508
rect 16396 19468 16436 19508
rect 17548 19468 17588 19508
rect 5164 19384 5204 19424
rect 1324 19300 1364 19340
rect 1516 19300 1556 19340
rect 3244 19300 3284 19340
rect 2764 19216 2804 19256
rect 2860 19216 2900 19256
rect 3340 19216 3380 19256
rect 3820 19216 3860 19256
rect 4300 19221 4340 19261
rect 5740 19216 5780 19256
rect 6988 19216 7028 19256
rect 7564 19216 7604 19256
rect 8812 19216 8852 19256
rect 9676 19216 9716 19256
rect 9772 19216 9812 19256
rect 10156 19216 10196 19256
rect 10252 19216 10292 19256
rect 10732 19216 10772 19256
rect 11212 19221 11252 19261
rect 11596 19216 11636 19256
rect 12844 19216 12884 19256
rect 13324 19216 13364 19256
rect 14572 19216 14612 19256
rect 14956 19216 14996 19256
rect 16204 19216 16244 19256
rect 16588 19216 16628 19256
rect 16684 19216 16724 19256
rect 16876 19216 16916 19256
rect 16972 19216 17012 19256
rect 17127 19216 17167 19256
rect 17356 19216 17396 19256
rect 17548 19216 17588 19256
rect 17740 19216 17780 19256
rect 18988 19216 19028 19256
rect 19468 19216 19508 19256
rect 19756 19216 19796 19256
rect 11404 19132 11444 19172
rect 19180 19132 19220 19172
rect 19852 19132 19892 19172
rect 4492 19048 4532 19088
rect 7180 19048 7220 19088
rect 16396 19048 16436 19088
rect 16972 19048 17012 19088
rect 20140 19006 20180 19046
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 6988 18712 7028 18752
rect 9484 18712 9524 18752
rect 11116 18712 11156 18752
rect 13228 18712 13268 18752
rect 14860 18712 14900 18752
rect 19180 18712 19220 18752
rect 19564 18712 19604 18752
rect 4396 18628 4436 18668
rect 5068 18628 5108 18668
rect 2092 18544 2132 18584
rect 2668 18544 2708 18584
rect 2764 18544 2804 18584
rect 3724 18544 3764 18584
rect 4204 18530 4244 18570
rect 4684 18544 4724 18584
rect 4972 18544 5012 18584
rect 5548 18544 5588 18584
rect 6796 18544 6836 18584
rect 8044 18544 8084 18584
rect 9292 18544 9332 18584
rect 9676 18544 9716 18584
rect 10924 18544 10964 18584
rect 11308 18544 11348 18584
rect 15052 18586 15092 18626
rect 11404 18544 11444 18584
rect 11596 18544 11636 18584
rect 11788 18544 11828 18584
rect 13036 18544 13076 18584
rect 13420 18544 13460 18584
rect 14668 18544 14708 18584
rect 16300 18544 16340 18584
rect 16780 18544 16820 18584
rect 17068 18544 17108 18584
rect 17164 18544 17204 18584
rect 17740 18544 17780 18584
rect 18988 18544 19028 18584
rect 19372 18544 19412 18584
rect 19468 18544 19508 18584
rect 19660 18544 19700 18584
rect 19756 18544 19796 18584
rect 19911 18544 19951 18584
rect 20140 18544 20180 18584
rect 3148 18460 3188 18500
rect 3244 18460 3284 18500
rect 1516 18376 1556 18416
rect 1804 18376 1844 18416
rect 16492 18376 16532 18416
rect 17452 18376 17492 18416
rect 1996 18292 2036 18332
rect 5356 18292 5396 18332
rect 11596 18292 11636 18332
rect 20236 18292 20276 18332
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 2668 17956 2708 17996
rect 4300 17956 4340 17996
rect 13132 17956 13172 17996
rect 13324 17956 13364 17996
rect 14476 17914 14516 17954
rect 16300 17956 16340 17996
rect 16492 17956 16532 17996
rect 17548 17956 17588 17996
rect 19180 17956 19220 17996
rect 19948 17956 19988 17996
rect 8908 17872 8948 17912
rect 6700 17788 6740 17828
rect 6796 17788 6836 17828
rect 14380 17830 14420 17870
rect 1228 17704 1268 17744
rect 2476 17704 2516 17744
rect 2860 17704 2900 17744
rect 4108 17704 4148 17744
rect 4492 17704 4532 17744
rect 5740 17704 5780 17744
rect 6220 17704 6260 17744
rect 6316 17704 6356 17744
rect 7276 17704 7316 17744
rect 7756 17709 7796 17749
rect 8236 17704 8276 17744
rect 8524 17704 8564 17744
rect 9196 17704 9236 17744
rect 9580 17704 9620 17744
rect 10828 17704 10868 17744
rect 11404 17704 11444 17744
rect 12652 17704 12692 17744
rect 13036 17704 13076 17744
rect 14284 17746 14324 17786
rect 14572 17788 14612 17828
rect 19372 17788 19412 17828
rect 19756 17788 19796 17828
rect 13708 17704 13748 17744
rect 13996 17704 14036 17744
rect 14668 17746 14708 17786
rect 14860 17704 14900 17744
rect 16108 17704 16148 17744
rect 16876 17704 16916 17744
rect 17164 17704 17204 17744
rect 17452 17704 17492 17744
rect 17740 17704 17780 17744
rect 18988 17704 19028 17744
rect 5932 17620 5972 17660
rect 7948 17620 7988 17660
rect 8620 17620 8660 17660
rect 12844 17620 12884 17660
rect 13612 17620 13652 17660
rect 16780 17620 16820 17660
rect 9100 17536 9140 17576
rect 11020 17536 11060 17576
rect 19564 17536 19604 17576
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 5932 17200 5972 17240
rect 7948 17200 7988 17240
rect 12844 17200 12884 17240
rect 1420 17116 1460 17156
rect 4108 17116 4148 17156
rect 9580 17116 9620 17156
rect 18796 17116 18836 17156
rect 1324 17032 1364 17072
rect 1516 17032 1556 17072
rect 1612 17032 1652 17072
rect 1804 17032 1844 17072
rect 1900 17032 1940 17072
rect 1996 17032 2036 17072
rect 2092 17032 2132 17072
rect 2380 17032 2420 17072
rect 2476 17032 2516 17072
rect 2956 17032 2996 17072
rect 3436 17032 3476 17072
rect 3916 17027 3956 17067
rect 4492 17032 4532 17072
rect 5740 17032 5780 17072
rect 6220 17032 6260 17072
rect 6316 17032 6356 17072
rect 7276 17032 7316 17072
rect 7756 17027 7796 17067
rect 8236 17032 8276 17072
rect 8716 17032 8756 17072
rect 9004 17032 9044 17072
rect 9100 17032 9140 17072
rect 9772 17032 9812 17072
rect 11020 17032 11060 17072
rect 11404 17032 11444 17072
rect 12652 17032 12692 17072
rect 13420 17032 13460 17072
rect 13708 17032 13748 17072
rect 13804 17032 13844 17072
rect 14476 17032 14516 17072
rect 15724 17032 15764 17072
rect 16108 17032 16148 17072
rect 16492 17032 16532 17072
rect 16684 17032 16724 17072
rect 17068 17032 17108 17072
rect 17356 17032 17396 17072
rect 18604 17032 18644 17072
rect 18988 17032 19028 17072
rect 19372 17032 19412 17072
rect 19564 17032 19604 17072
rect 19948 17032 19988 17072
rect 20127 17043 20167 17083
rect 2860 16948 2900 16988
rect 6700 16948 6740 16988
rect 6796 16948 6836 16988
rect 16204 16948 16244 16988
rect 16396 16948 16436 16988
rect 16780 16948 16820 16988
rect 16972 16948 17012 16988
rect 19084 16948 19124 16988
rect 19276 16948 19316 16988
rect 19660 16948 19700 16988
rect 19852 16948 19892 16988
rect 20236 16948 20276 16988
rect 14092 16864 14132 16904
rect 16300 16864 16340 16904
rect 16876 16864 16916 16904
rect 19180 16864 19220 16904
rect 19756 16864 19796 16904
rect 8140 16780 8180 16820
rect 9388 16780 9428 16820
rect 15916 16780 15956 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 19948 16444 19988 16484
rect 8524 16360 8564 16400
rect 18892 16360 18932 16400
rect 2860 16276 2900 16316
rect 9676 16276 9716 16316
rect 15724 16276 15764 16316
rect 15820 16276 15860 16316
rect 1228 16192 1268 16232
rect 1324 16192 1364 16232
rect 1516 16192 1556 16232
rect 1708 16192 1748 16232
rect 1900 16192 1940 16232
rect 1996 16192 2036 16232
rect 2284 16192 2324 16232
rect 2380 16192 2420 16232
rect 2764 16192 2804 16232
rect 3340 16192 3380 16232
rect 3820 16197 3860 16237
rect 4204 16192 4244 16232
rect 4300 16192 4340 16232
rect 4588 16192 4628 16232
rect 5836 16192 5876 16232
rect 6311 16192 6351 16232
rect 6412 16192 6452 16232
rect 6508 16192 6548 16232
rect 6700 16192 6740 16232
rect 6796 16192 6836 16232
rect 7084 16192 7124 16232
rect 8332 16192 8372 16232
rect 8716 16192 8756 16232
rect 8908 16192 8948 16232
rect 9196 16192 9236 16232
rect 9292 16192 9332 16232
rect 9772 16192 9812 16232
rect 10252 16192 10292 16232
rect 10732 16206 10772 16246
rect 11596 16192 11636 16232
rect 12844 16192 12884 16232
rect 13516 16192 13556 16232
rect 14764 16192 14804 16232
rect 15244 16192 15284 16232
rect 15340 16192 15380 16232
rect 16300 16192 16340 16232
rect 16780 16197 16820 16237
rect 17260 16192 17300 16232
rect 17452 16192 17492 16232
rect 18700 16192 18740 16232
rect 19180 16192 19220 16232
rect 19276 16192 19316 16232
rect 19468 16192 19508 16232
rect 19564 16192 19604 16232
rect 19721 16199 19761 16239
rect 20140 16234 20180 16274
rect 19948 16192 19988 16232
rect 20236 16192 20276 16232
rect 10924 16108 10964 16148
rect 1420 16024 1460 16064
rect 1804 16024 1844 16064
rect 4012 16024 4052 16064
rect 6028 16024 6068 16064
rect 6316 16024 6356 16064
rect 8812 16024 8852 16064
rect 13036 16024 13076 16064
rect 14956 16024 14996 16064
rect 16972 16024 17012 16064
rect 17164 16024 17204 16064
rect 19372 16024 19412 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 2668 15688 2708 15728
rect 10924 15688 10964 15728
rect 14956 15688 14996 15728
rect 3340 15604 3380 15644
rect 6892 15604 6932 15644
rect 8908 15604 8948 15644
rect 13420 15604 13460 15644
rect 17452 15604 17492 15644
rect 1228 15520 1268 15560
rect 2476 15520 2516 15560
rect 2956 15520 2996 15560
rect 3244 15520 3284 15560
rect 3820 15520 3860 15560
rect 5068 15520 5108 15560
rect 5452 15520 5492 15560
rect 6700 15520 6740 15560
rect 7180 15520 7220 15560
rect 7276 15520 7316 15560
rect 8236 15520 8276 15560
rect 8716 15506 8756 15546
rect 9196 15520 9236 15560
rect 9292 15520 9332 15560
rect 9676 15520 9716 15560
rect 9772 15520 9812 15560
rect 10252 15520 10292 15560
rect 10732 15515 10772 15555
rect 11116 15507 11156 15547
rect 11404 15520 11444 15560
rect 11788 15520 11828 15560
rect 11980 15520 12020 15560
rect 13228 15520 13268 15560
rect 13900 15520 13940 15560
rect 13996 15520 14036 15560
rect 14284 15520 14324 15560
rect 14606 15505 14646 15545
rect 14764 15520 14804 15560
rect 14860 15520 14900 15560
rect 15052 15520 15092 15560
rect 15148 15520 15188 15560
rect 15724 15520 15764 15560
rect 15820 15520 15860 15560
rect 16204 15520 16244 15560
rect 16780 15520 16820 15560
rect 17260 15515 17300 15555
rect 17644 15520 17684 15560
rect 18892 15520 18932 15560
rect 19372 15520 19412 15560
rect 19660 15520 19700 15560
rect 19756 15520 19796 15560
rect 7660 15436 7700 15476
rect 7756 15436 7796 15476
rect 11500 15436 11540 15476
rect 11692 15436 11732 15476
rect 16300 15436 16340 15476
rect 5260 15352 5300 15392
rect 11596 15352 11636 15392
rect 13612 15352 13652 15392
rect 20044 15352 20084 15392
rect 3628 15268 3668 15308
rect 11212 15268 11252 15308
rect 19084 15268 19124 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 3340 14932 3380 14972
rect 3532 14932 3572 14972
rect 9004 14932 9044 14972
rect 13324 14932 13364 14972
rect 14284 14932 14324 14972
rect 16972 14932 17012 14972
rect 18316 14932 18356 14972
rect 19852 14932 19892 14972
rect 20236 14932 20276 14972
rect 1516 14848 1556 14888
rect 5164 14848 5204 14888
rect 6316 14848 6356 14888
rect 6892 14848 6932 14888
rect 10828 14848 10868 14888
rect 14668 14848 14708 14888
rect 1420 14764 1460 14804
rect 1612 14764 1652 14804
rect 6220 14764 6260 14804
rect 6412 14764 6452 14804
rect 10732 14764 10772 14804
rect 10924 14764 10964 14804
rect 14572 14764 14612 14804
rect 14764 14764 14804 14804
rect 18124 14764 18164 14804
rect 1324 14680 1364 14720
rect 1708 14680 1748 14720
rect 1900 14680 1940 14720
rect 3148 14680 3188 14720
rect 3724 14680 3764 14720
rect 4972 14680 5012 14720
rect 5452 14680 5492 14720
rect 5548 14680 5588 14720
rect 5836 14680 5876 14720
rect 6124 14680 6164 14720
rect 6508 14680 6548 14720
rect 6796 14680 6836 14720
rect 6988 14680 7028 14720
rect 7084 14680 7124 14720
rect 7564 14680 7604 14720
rect 8812 14680 8852 14720
rect 9196 14680 9236 14720
rect 9292 14680 9332 14720
rect 9676 14680 9716 14720
rect 9772 14680 9812 14720
rect 9868 14680 9908 14720
rect 9964 14680 10004 14720
rect 10156 14680 10196 14720
rect 10348 14680 10388 14720
rect 10444 14680 10484 14720
rect 10636 14680 10676 14720
rect 11020 14680 11060 14720
rect 11212 14680 11252 14720
rect 11404 14680 11444 14720
rect 11596 14680 11636 14720
rect 12844 14680 12884 14720
rect 13228 14680 13268 14720
rect 13612 14680 13652 14720
rect 13900 14680 13940 14720
rect 14476 14680 14516 14720
rect 17260 14722 17300 14762
rect 14860 14680 14900 14720
rect 15340 14680 15380 14720
rect 16588 14680 16628 14720
rect 17356 14680 17396 14720
rect 17644 14680 17684 14720
rect 18508 14680 18548 14720
rect 18604 14680 18644 14720
rect 18796 14680 18836 14720
rect 19180 14680 19220 14720
rect 19468 14680 19508 14720
rect 20044 14680 20084 14720
rect 20236 14680 20276 14720
rect 11308 14596 11348 14636
rect 13996 14596 14036 14636
rect 16780 14596 16820 14636
rect 19564 14596 19604 14636
rect 3532 14512 3572 14552
rect 9484 14512 9524 14552
rect 10252 14512 10292 14552
rect 13036 14512 13076 14552
rect 18796 14512 18836 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 2668 14176 2708 14216
rect 4300 14176 4340 14216
rect 12268 14176 12308 14216
rect 12844 14176 12884 14216
rect 16204 14176 16244 14216
rect 16588 14176 16628 14216
rect 17068 14176 17108 14216
rect 20236 14176 20276 14216
rect 4780 14092 4820 14132
rect 8908 14092 8948 14132
rect 11788 14092 11828 14132
rect 14476 14092 14516 14132
rect 14956 14092 14996 14132
rect 1228 14008 1268 14048
rect 2476 14008 2516 14048
rect 2860 14008 2900 14048
rect 4108 14008 4148 14048
rect 4876 14008 4916 14048
rect 5164 14008 5204 14048
rect 5548 14008 5588 14048
rect 5932 14008 5972 14048
rect 7180 14008 7220 14048
rect 7468 14008 7508 14048
rect 8716 14008 8756 14048
rect 10348 14008 10388 14048
rect 10828 14008 10868 14048
rect 11116 14008 11156 14048
rect 9100 13966 9140 14006
rect 11212 14008 11252 14048
rect 11692 14008 11732 14048
rect 11884 14008 11924 14048
rect 11980 14008 12020 14048
rect 12172 14008 12212 14048
rect 12364 14008 12404 14048
rect 12556 14008 12596 14048
rect 12652 14008 12692 14048
rect 12844 14008 12884 14048
rect 13036 14008 13076 14048
rect 14284 14008 14324 14048
rect 14668 14008 14708 14048
rect 14764 14008 14804 14048
rect 14860 14008 14900 14048
rect 15148 14008 15188 14048
rect 15340 14008 15380 14048
rect 15436 14008 15476 14048
rect 15628 14008 15668 14048
rect 15724 14008 15764 14048
rect 15820 14008 15860 14048
rect 15916 14008 15956 14048
rect 16108 14008 16148 14048
rect 16300 14008 16340 14048
rect 16492 14008 16532 14048
rect 16684 14008 16724 14048
rect 17260 14008 17300 14048
rect 18508 14008 18548 14048
rect 18892 14008 18932 14048
rect 19276 14008 19316 14048
rect 19468 14008 19508 14048
rect 19852 14008 19892 14048
rect 16876 13924 16916 13964
rect 18988 13924 19028 13964
rect 19180 13924 19220 13964
rect 19564 13924 19604 13964
rect 19756 13924 19796 13964
rect 20044 13924 20084 13964
rect 4492 13840 4532 13880
rect 10540 13840 10580 13880
rect 11500 13840 11540 13880
rect 18700 13840 18740 13880
rect 19084 13840 19124 13880
rect 19660 13840 19700 13880
rect 4300 13756 4340 13796
rect 5452 13756 5492 13796
rect 5740 13756 5780 13796
rect 15148 13756 15188 13796
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 2668 13420 2708 13460
rect 9964 13420 10004 13460
rect 10828 13420 10868 13460
rect 16876 13420 16916 13460
rect 18508 13420 18548 13460
rect 19468 13420 19508 13460
rect 19660 13420 19700 13460
rect 7180 13252 7220 13292
rect 10444 13252 10484 13292
rect 1228 13168 1268 13208
rect 2476 13168 2516 13208
rect 3052 13168 3092 13208
rect 4300 13168 4340 13208
rect 4876 13168 4916 13208
rect 6124 13168 6164 13208
rect 6604 13168 6644 13208
rect 6700 13168 6740 13208
rect 7084 13168 7124 13208
rect 7660 13168 7700 13208
rect 8188 13177 8228 13217
rect 9772 13210 9812 13250
rect 13612 13252 13652 13292
rect 13708 13252 13748 13292
rect 8524 13168 8564 13208
rect 10348 13168 10388 13208
rect 10636 13168 10676 13208
rect 11116 13168 11156 13208
rect 11212 13168 11252 13208
rect 11500 13168 11540 13208
rect 11692 13168 11732 13208
rect 11788 13168 11828 13208
rect 12076 13168 12116 13208
rect 12172 13168 12212 13208
rect 12268 13168 12308 13208
rect 12556 13168 12596 13208
rect 12844 13168 12884 13208
rect 13132 13168 13172 13208
rect 13228 13168 13268 13208
rect 14188 13168 14228 13208
rect 14716 13177 14756 13217
rect 15052 13168 15092 13208
rect 15244 13168 15284 13208
rect 15436 13168 15476 13208
rect 16684 13168 16724 13208
rect 17068 13168 17108 13208
rect 18316 13168 18356 13208
rect 18796 13168 18836 13208
rect 19084 13168 19124 13208
rect 19180 13168 19220 13208
rect 19660 13168 19700 13208
rect 19756 13168 19796 13208
rect 19948 13168 19988 13208
rect 20044 13168 20084 13208
rect 20145 13168 20185 13208
rect 8332 13084 8372 13124
rect 12748 13084 12788 13124
rect 2860 13000 2900 13040
rect 4492 13000 4532 13040
rect 6316 13000 6356 13040
rect 9964 13000 10004 13040
rect 11596 13000 11636 13040
rect 12364 13000 12404 13040
rect 14860 13000 14900 13040
rect 15148 13000 15188 13040
rect 11308 12942 11348 12982
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 2668 12664 2708 12704
rect 5836 12664 5876 12704
rect 9772 12664 9812 12704
rect 10636 12664 10676 12704
rect 18700 12664 18740 12704
rect 5644 12580 5684 12620
rect 13612 12580 13652 12620
rect 13900 12580 13940 12620
rect 15724 12580 15764 12620
rect 1228 12496 1268 12536
rect 2476 12496 2516 12536
rect 2956 12496 2996 12536
rect 3532 12496 3572 12536
rect 3628 12496 3668 12536
rect 3916 12496 3956 12536
rect 4204 12496 4244 12536
rect 5452 12496 5492 12536
rect 5980 12486 6020 12526
rect 6508 12496 6548 12536
rect 6988 12496 7028 12536
rect 7468 12496 7508 12536
rect 7564 12496 7604 12536
rect 7852 12496 7892 12536
rect 8044 12496 8084 12536
rect 8140 12496 8180 12536
rect 8332 12496 8372 12536
rect 9580 12496 9620 12536
rect 9964 12496 10004 12536
rect 10156 12496 10196 12536
rect 10252 12496 10292 12536
rect 10732 12496 10772 12536
rect 10828 12496 10868 12536
rect 10924 12496 10964 12536
rect 7084 12412 7124 12452
rect 11212 12451 11252 12491
rect 11308 12496 11348 12536
rect 11404 12496 11444 12536
rect 11500 12496 11540 12536
rect 11692 12496 11732 12536
rect 11884 12496 11924 12536
rect 11980 12496 12020 12536
rect 12172 12496 12212 12536
rect 13420 12496 13460 12536
rect 13804 12496 13844 12536
rect 13996 12496 14036 12536
rect 14092 12496 14132 12536
rect 14284 12496 14324 12536
rect 15532 12496 15572 12536
rect 15916 12496 15956 12536
rect 16108 12496 16148 12536
rect 16300 12496 16340 12536
rect 16684 12496 16724 12536
rect 17260 12496 17300 12536
rect 18508 12496 18548 12536
rect 19180 12496 19220 12536
rect 19468 12496 19508 12536
rect 19564 12496 19604 12536
rect 16396 12412 16436 12452
rect 16588 12412 16628 12452
rect 16876 12412 16916 12452
rect 20044 12412 20084 12452
rect 3244 12328 3284 12368
rect 9964 12328 10004 12368
rect 16108 12328 16148 12368
rect 16492 12328 16532 12368
rect 17068 12328 17108 12368
rect 19852 12328 19892 12368
rect 20236 12328 20276 12368
rect 3052 12244 3092 12284
rect 7852 12244 7892 12284
rect 11692 12244 11732 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 1516 11908 1556 11948
rect 8332 11908 8372 11948
rect 11404 11908 11444 11948
rect 13036 11908 13076 11948
rect 16588 11908 16628 11948
rect 17644 11908 17684 11948
rect 17836 11908 17876 11948
rect 20044 11908 20084 11948
rect 8140 11824 8180 11864
rect 9580 11824 9620 11864
rect 9484 11740 9524 11780
rect 2956 11698 2996 11738
rect 9676 11740 9716 11780
rect 17452 11740 17492 11780
rect 19852 11740 19892 11780
rect 1324 11656 1364 11696
rect 1708 11656 1748 11696
rect 3148 11656 3188 11696
rect 4396 11656 4436 11696
rect 4876 11656 4916 11696
rect 5260 11656 5300 11696
rect 6508 11656 6548 11696
rect 6700 11656 6740 11696
rect 7948 11656 7988 11696
rect 8620 11656 8660 11696
rect 8716 11656 8756 11696
rect 9004 11656 9044 11696
rect 9388 11656 9428 11696
rect 9772 11656 9812 11696
rect 9964 11656 10004 11696
rect 11212 11656 11252 11696
rect 11596 11656 11636 11696
rect 12844 11656 12884 11696
rect 13420 11656 13460 11696
rect 14668 11656 14708 11696
rect 15052 11656 15092 11696
rect 16300 11656 16340 11696
rect 16588 11656 16628 11696
rect 16684 11656 16724 11696
rect 16876 11656 16916 11696
rect 16972 11656 17012 11696
rect 17127 11656 17167 11696
rect 17836 11656 17876 11696
rect 18028 11656 18068 11696
rect 18220 11656 18260 11696
rect 19468 11656 19508 11696
rect 4780 11572 4820 11612
rect 1228 11488 1268 11528
rect 1516 11488 1556 11528
rect 4588 11488 4628 11528
rect 5068 11488 5108 11528
rect 11404 11488 11444 11528
rect 13036 11488 13076 11528
rect 13228 11488 13268 11528
rect 14860 11488 14900 11528
rect 19660 11488 19700 11528
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 1324 11152 1364 11192
rect 2956 11152 2996 11192
rect 18124 11152 18164 11192
rect 20236 11152 20276 11192
rect 6604 11068 6644 11108
rect 6796 11068 6836 11108
rect 9292 11068 9332 11108
rect 12748 11068 12788 11108
rect 1516 10984 1556 11024
rect 2764 10984 2804 11024
rect 3148 10984 3188 11024
rect 3249 10974 3289 11014
rect 3724 10984 3764 11024
rect 4972 10984 5012 11024
rect 5164 10984 5204 11024
rect 6412 10984 6452 11024
rect 6988 10979 7028 11019
rect 7468 10984 7508 11024
rect 7948 10984 7988 11024
rect 8428 10984 8468 11024
rect 8524 10984 8564 11024
rect 8812 10984 8852 11024
rect 9100 10984 9140 11024
rect 9484 10984 9524 11024
rect 10732 10984 10772 11024
rect 11020 10984 11060 11024
rect 11116 10984 11156 11024
rect 12076 10984 12116 11024
rect 12556 10979 12596 11019
rect 13036 10984 13076 11024
rect 14284 10984 14324 11024
rect 14860 10984 14900 11024
rect 15052 10984 15092 11024
rect 16300 10984 16340 11024
rect 16780 10984 16820 11024
rect 17068 10984 17108 11024
rect 17164 10984 17204 11024
rect 17644 10984 17684 11024
rect 17836 10984 17876 11024
rect 18028 10984 18068 11024
rect 18220 10984 18260 11024
rect 18412 10984 18452 11024
rect 19660 10984 19700 11024
rect 8044 10900 8084 10940
rect 11500 10900 11540 10940
rect 11596 10900 11636 10940
rect 20044 10900 20084 10940
rect 17452 10816 17492 10856
rect 3532 10732 3572 10772
rect 9100 10732 9140 10772
rect 14476 10732 14516 10772
rect 14764 10732 14804 10772
rect 16492 10732 16532 10772
rect 17644 10732 17684 10772
rect 19852 10732 19892 10772
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 2668 10396 2708 10436
rect 2860 10396 2900 10436
rect 9868 10396 9908 10436
rect 15820 10396 15860 10436
rect 11404 10312 11444 10352
rect 11980 10312 12020 10352
rect 16204 10312 16244 10352
rect 16588 10312 16628 10352
rect 17740 10312 17780 10352
rect 5068 10228 5108 10268
rect 10924 10228 10964 10268
rect 11308 10228 11348 10268
rect 11500 10228 11540 10268
rect 11884 10228 11924 10268
rect 12076 10228 12116 10268
rect 13708 10228 13748 10268
rect 1228 10144 1268 10184
rect 2476 10144 2516 10184
rect 3244 10144 3284 10184
rect 3532 10144 3572 10184
rect 4012 10158 4052 10198
rect 4492 10144 4532 10184
rect 4972 10144 5012 10184
rect 5452 10144 5492 10184
rect 5548 10144 5588 10184
rect 5932 10144 5972 10184
rect 7180 10144 7220 10184
rect 7756 10144 7796 10184
rect 7852 10144 7892 10184
rect 7948 10144 7988 10184
rect 8044 10144 8084 10184
rect 8236 10144 8276 10184
rect 9484 10144 9524 10184
rect 10156 10144 10196 10184
rect 10252 10144 10292 10184
rect 10540 10144 10580 10184
rect 10828 10144 10868 10184
rect 11020 10144 11060 10184
rect 11212 10144 11252 10184
rect 11596 10144 11636 10184
rect 11788 10144 11828 10184
rect 12364 10186 12404 10226
rect 13804 10228 13844 10268
rect 16108 10228 16148 10268
rect 16300 10228 16340 10268
rect 12172 10144 12212 10184
rect 12556 10144 12596 10184
rect 12652 10144 12692 10184
rect 12844 10144 12884 10184
rect 13228 10144 13268 10184
rect 13324 10144 13364 10184
rect 14284 10144 14324 10184
rect 14764 10158 14804 10198
rect 15244 10144 15284 10184
rect 15532 10144 15572 10184
rect 15628 10144 15668 10184
rect 15820 10144 15860 10184
rect 16012 10144 16052 10184
rect 16396 10144 16436 10184
rect 16876 10144 16916 10184
rect 16972 10144 17012 10184
rect 17260 10144 17300 10184
rect 17740 10144 17780 10184
rect 18124 10144 18164 10184
rect 19372 10144 19412 10184
rect 19852 10186 19892 10226
rect 19756 10144 19796 10184
rect 19948 10144 19988 10184
rect 3148 10060 3188 10100
rect 3820 10060 3860 10100
rect 7372 10060 7412 10100
rect 9676 9976 9716 10016
rect 12364 9976 12404 10016
rect 12940 9976 12980 10016
rect 14956 9976 14996 10016
rect 15340 9976 15380 10016
rect 17932 9976 17972 10016
rect 19564 9976 19604 10016
rect 20044 9976 20084 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 3244 9640 3284 9680
rect 4492 9640 4532 9680
rect 9964 9640 10004 9680
rect 12076 9640 12116 9680
rect 12652 9640 12692 9680
rect 17932 9640 17972 9680
rect 3724 9556 3764 9596
rect 13516 9556 13556 9596
rect 17068 9556 17108 9596
rect 1324 9472 1364 9512
rect 1516 9472 1556 9512
rect 1612 9472 1652 9512
rect 1804 9472 1844 9512
rect 3052 9472 3092 9512
rect 3820 9472 3860 9512
rect 4108 9472 4148 9512
rect 4396 9472 4436 9512
rect 4588 9472 4628 9512
rect 4684 9472 4724 9512
rect 4876 9472 4916 9512
rect 6124 9472 6164 9512
rect 6508 9472 6548 9512
rect 7756 9472 7796 9512
rect 8332 9472 8372 9512
rect 9580 9472 9620 9512
rect 9772 9472 9812 9512
rect 9868 9472 9908 9512
rect 10060 9472 10100 9512
rect 10156 9472 10196 9512
rect 10257 9472 10297 9512
rect 10636 9472 10676 9512
rect 11884 9472 11924 9512
rect 12268 9472 12308 9512
rect 12412 9449 12452 9489
rect 12556 9472 12596 9512
rect 12652 9443 12692 9483
rect 12809 9457 12849 9497
rect 13036 9472 13076 9512
rect 13228 9472 13268 9512
rect 13708 9467 13748 9507
rect 14188 9472 14228 9512
rect 14764 9472 14804 9512
rect 15148 9472 15188 9512
rect 15244 9472 15284 9512
rect 15628 9472 15668 9512
rect 16012 9472 16052 9512
rect 16204 9472 16244 9512
rect 16588 9472 16628 9512
rect 17164 9472 17204 9512
rect 17452 9472 17492 9512
rect 17740 9472 17780 9512
rect 17836 9472 17876 9512
rect 18028 9472 18068 9512
rect 18124 9472 18164 9512
rect 18225 9472 18265 9512
rect 18796 9472 18836 9512
rect 19084 9472 19124 9512
rect 19180 9472 19220 9512
rect 19660 9472 19700 9512
rect 19756 9472 19796 9512
rect 19948 9472 19988 9512
rect 20127 9483 20167 9523
rect 14668 9388 14708 9428
rect 15724 9388 15764 9428
rect 15916 9388 15956 9428
rect 16300 9388 16340 9428
rect 16492 9388 16532 9428
rect 20236 9388 20276 9428
rect 8140 9304 8180 9344
rect 13036 9304 13076 9344
rect 15820 9304 15860 9344
rect 16396 9304 16436 9344
rect 19468 9304 19508 9344
rect 19948 9304 19988 9344
rect 1324 9220 1364 9260
rect 3436 9220 3476 9260
rect 6316 9220 6356 9260
rect 7948 9220 7988 9260
rect 16780 9220 16820 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 3244 8884 3284 8924
rect 10156 8884 10196 8924
rect 11404 8884 11444 8924
rect 13132 8884 13172 8924
rect 16780 8884 16820 8924
rect 17836 8884 17876 8924
rect 6220 8800 6260 8840
rect 2860 8716 2900 8756
rect 18124 8716 18164 8756
rect 1228 8632 1268 8672
rect 2476 8632 2516 8672
rect 3532 8632 3572 8672
rect 3628 8632 3668 8672
rect 3916 8632 3956 8672
rect 4300 8632 4340 8672
rect 4396 8632 4436 8672
rect 4780 8632 4820 8672
rect 4876 8632 4916 8672
rect 5356 8632 5396 8672
rect 5836 8637 5876 8677
rect 6604 8632 6644 8672
rect 6700 8632 6740 8672
rect 7084 8632 7124 8672
rect 7180 8632 7220 8672
rect 7660 8632 7700 8672
rect 8140 8646 8180 8686
rect 8524 8632 8564 8672
rect 9772 8632 9812 8672
rect 10444 8632 10484 8672
rect 10540 8632 10580 8672
rect 10828 8632 10868 8672
rect 11116 8632 11156 8672
rect 11212 8632 11252 8672
rect 11788 8632 11828 8672
rect 12076 8632 12116 8672
rect 12460 8632 12500 8672
rect 14668 8674 14708 8714
rect 12748 8632 12788 8672
rect 13420 8632 13460 8672
rect 15052 8632 15092 8672
rect 15340 8632 15380 8672
rect 16588 8632 16628 8672
rect 17164 8632 17204 8672
rect 17452 8632 17492 8672
rect 18028 8632 18068 8672
rect 18412 8651 18452 8691
rect 18508 8651 18548 8691
rect 18892 8632 18932 8672
rect 18988 8632 19028 8672
rect 19468 8632 19508 8672
rect 19948 8646 19988 8686
rect 6028 8548 6068 8588
rect 9964 8548 10004 8588
rect 11692 8548 11732 8588
rect 12844 8548 12884 8588
rect 17548 8548 17588 8588
rect 2668 8464 2708 8504
rect 3052 8464 3092 8504
rect 8332 8464 8372 8504
rect 14860 8464 14900 8504
rect 15148 8464 15188 8504
rect 20140 8464 20180 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 2956 8128 2996 8168
rect 5164 8128 5204 8168
rect 2668 8044 2708 8084
rect 5836 8086 5876 8126
rect 12748 8128 12788 8168
rect 14092 8128 14132 8168
rect 17644 8128 17684 8168
rect 18412 8128 18452 8168
rect 11884 8044 11924 8084
rect 1228 7960 1268 8000
rect 2476 7960 2516 8000
rect 3100 7950 3140 7990
rect 3628 7960 3668 8000
rect 4588 7960 4628 8000
rect 4684 7960 4724 8000
rect 4972 7960 5012 8000
rect 5068 7960 5108 8000
rect 5260 7960 5300 8000
rect 5356 7960 5396 8000
rect 5457 7960 5497 8000
rect 5980 7950 6020 7990
rect 6508 7960 6548 8000
rect 6988 7960 7028 8000
rect 7084 7960 7124 8000
rect 7468 7960 7508 8000
rect 9676 8002 9716 8042
rect 14956 8044 14996 8084
rect 16876 8044 16916 8084
rect 7564 7960 7604 8000
rect 8044 7960 8084 8000
rect 9292 7960 9332 8000
rect 10060 7960 10100 8000
rect 10444 7960 10484 8000
rect 11692 7960 11732 8000
rect 12076 7960 12116 8000
rect 12268 7960 12308 8000
rect 12364 7960 12404 8000
rect 12652 7960 12692 8000
rect 12844 7960 12884 8000
rect 13036 7960 13076 8000
rect 13324 7960 13364 8000
rect 13516 7960 13556 8000
rect 13612 7960 13652 8000
rect 13708 7960 13748 8000
rect 13804 7960 13844 8000
rect 13996 7960 14036 8000
rect 14188 7960 14228 8000
rect 14572 7960 14612 8000
rect 14860 7960 14900 8000
rect 15436 7960 15476 8000
rect 16684 7960 16724 8000
rect 17068 7960 17108 8000
rect 17164 7960 17204 8000
rect 17356 7960 17396 8000
rect 17548 7960 17588 8000
rect 17740 7960 17780 8000
rect 18508 7960 18548 8000
rect 18604 7960 18644 8000
rect 18700 7960 18740 8000
rect 18892 7960 18932 8000
rect 19276 7960 19316 8000
rect 19468 7960 19508 8000
rect 19852 7960 19892 8000
rect 20044 7960 20084 8000
rect 20236 7960 20276 8000
rect 4108 7876 4148 7916
rect 4204 7876 4244 7916
rect 9772 7876 9812 7916
rect 9964 7876 10004 7916
rect 18028 7876 18068 7916
rect 18988 7876 19028 7916
rect 19180 7876 19220 7916
rect 19564 7876 19604 7916
rect 19756 7876 19796 7916
rect 9484 7792 9524 7832
rect 9868 7792 9908 7832
rect 12268 7792 12308 7832
rect 17164 7792 17204 7832
rect 19084 7792 19124 7832
rect 19660 7792 19700 7832
rect 20236 7792 20276 7832
rect 13324 7708 13364 7748
rect 15244 7708 15284 7748
rect 18220 7708 18260 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 3628 7372 3668 7412
rect 5644 7372 5684 7412
rect 5836 7372 5876 7412
rect 13996 7372 14036 7412
rect 14668 7372 14708 7412
rect 17452 7372 17492 7412
rect 19276 7372 19316 7412
rect 8140 7288 8180 7328
rect 8332 7262 8372 7302
rect 15052 7288 15092 7328
rect 15628 7288 15668 7328
rect 9484 7204 9524 7244
rect 9580 7204 9620 7244
rect 11116 7204 11156 7244
rect 11500 7204 11540 7244
rect 15532 7204 15572 7244
rect 15724 7204 15764 7244
rect 1228 7120 1268 7160
rect 1420 7120 1460 7160
rect 1516 7120 1556 7160
rect 1708 7120 1748 7160
rect 1804 7120 1844 7160
rect 1900 7120 1940 7160
rect 1996 7120 2036 7160
rect 2188 7120 2228 7160
rect 3436 7120 3476 7160
rect 3820 7120 3860 7160
rect 4012 7120 4052 7160
rect 4204 7120 4244 7160
rect 5452 7120 5492 7160
rect 6028 7120 6068 7160
rect 7276 7120 7316 7160
rect 7660 7120 7700 7160
rect 7756 7120 7796 7160
rect 7852 7120 7892 7160
rect 7948 7120 7988 7160
rect 8332 7112 8372 7152
rect 8716 7120 8756 7160
rect 9004 7120 9044 7160
rect 9100 7120 9140 7160
rect 10060 7120 10100 7160
rect 10540 7125 10580 7165
rect 11788 7120 11828 7160
rect 12076 7120 12116 7160
rect 12172 7120 12212 7160
rect 12556 7120 12596 7160
rect 12652 7120 12692 7160
rect 13132 7120 13172 7160
rect 13612 7125 13652 7165
rect 13996 7120 14036 7160
rect 14188 7120 14228 7160
rect 14284 7120 14324 7160
rect 14476 7120 14516 7160
rect 14668 7120 14708 7160
rect 14956 7120 14996 7160
rect 15052 7120 15092 7160
rect 15244 7120 15284 7160
rect 15436 7120 15476 7160
rect 15820 7120 15860 7160
rect 16012 7120 16052 7160
rect 17260 7120 17300 7160
rect 17836 7120 17876 7160
rect 19084 7120 19124 7160
rect 19468 7120 19508 7160
rect 19564 7120 19604 7160
rect 19756 7120 19796 7160
rect 19852 7120 19892 7160
rect 19953 7120 19993 7160
rect 1324 7036 1364 7076
rect 8620 7036 8660 7076
rect 3916 6952 3956 6992
rect 10732 6952 10772 6992
rect 10924 6952 10964 6992
rect 11308 6952 11348 6992
rect 11692 6952 11732 6992
rect 13804 6952 13844 6992
rect 19660 6952 19700 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 1612 6616 1652 6656
rect 2380 6616 2420 6656
rect 2572 6616 2612 6656
rect 6028 6616 6068 6656
rect 10252 6616 10292 6656
rect 11884 6616 11924 6656
rect 13516 6616 13556 6656
rect 14380 6616 14420 6656
rect 16108 6616 16148 6656
rect 6412 6532 6452 6572
rect 17260 6574 17300 6614
rect 1228 6448 1268 6488
rect 1420 6448 1460 6488
rect 1804 6448 1844 6488
rect 1905 6457 1945 6497
rect 2092 6448 2132 6488
rect 2188 6448 2228 6488
rect 2764 6443 2804 6483
rect 3244 6448 3284 6488
rect 3724 6448 3764 6488
rect 3820 6448 3860 6488
rect 4204 6448 4244 6488
rect 4300 6448 4340 6488
rect 4588 6448 4628 6488
rect 5836 6448 5876 6488
rect 6604 6434 6644 6474
rect 7084 6448 7124 6488
rect 7564 6448 7604 6488
rect 8044 6448 8084 6488
rect 8140 6448 8180 6488
rect 8428 6448 8468 6488
rect 8620 6448 8660 6488
rect 8812 6448 8852 6488
rect 10060 6448 10100 6488
rect 10444 6448 10484 6488
rect 11692 6448 11732 6488
rect 13324 6448 13364 6488
rect 13708 6448 13748 6488
rect 12076 6406 12116 6446
rect 13900 6448 13940 6488
rect 13996 6448 14036 6488
rect 14284 6448 14324 6488
rect 14476 6448 14516 6488
rect 14668 6448 14708 6488
rect 15916 6448 15956 6488
rect 16300 6448 16340 6488
rect 16396 6448 16436 6488
rect 16588 6448 16628 6488
rect 16684 6448 16724 6488
rect 16828 6447 16868 6487
rect 17068 6448 17108 6488
rect 17452 6448 17492 6488
rect 17740 6448 17780 6488
rect 18988 6448 19028 6488
rect 19660 6448 19700 6488
rect 19756 6448 19796 6488
rect 20044 6448 20084 6488
rect 7660 6364 7700 6404
rect 17164 6364 17204 6404
rect 17356 6364 17396 6404
rect 8620 6280 8660 6320
rect 19372 6280 19412 6320
rect 1420 6196 1460 6236
rect 13708 6196 13748 6236
rect 16300 6196 16340 6236
rect 19180 6196 19220 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 2764 5860 2804 5900
rect 5932 5860 5972 5900
rect 7564 5860 7604 5900
rect 11884 5860 11924 5900
rect 15532 5860 15572 5900
rect 16876 5860 16916 5900
rect 19852 5860 19892 5900
rect 20236 5860 20276 5900
rect 1804 5776 1844 5816
rect 2380 5776 2420 5816
rect 9868 5776 9908 5816
rect 2284 5692 2324 5732
rect 2476 5692 2516 5732
rect 8908 5692 8948 5732
rect 9004 5692 9044 5732
rect 10060 5692 10100 5732
rect 13516 5692 13556 5732
rect 17164 5692 17204 5732
rect 1228 5608 1268 5648
rect 1324 5608 1364 5648
rect 1516 5608 1556 5648
rect 1708 5608 1748 5648
rect 1900 5608 1940 5648
rect 1996 5608 2036 5648
rect 2188 5608 2228 5648
rect 2572 5608 2612 5648
rect 2956 5608 2996 5648
rect 4204 5608 4244 5648
rect 4492 5608 4532 5648
rect 5740 5608 5780 5648
rect 6124 5608 6164 5648
rect 7372 5608 7412 5648
rect 7948 5613 7988 5653
rect 8428 5608 8468 5648
rect 9388 5608 9428 5648
rect 9484 5608 9524 5648
rect 10444 5608 10484 5648
rect 11692 5608 11732 5648
rect 12364 5608 12404 5648
rect 12460 5608 12500 5648
rect 12556 5608 12596 5648
rect 12940 5608 12980 5648
rect 13036 5608 13076 5648
rect 13132 5608 13172 5648
rect 13228 5608 13268 5648
rect 13420 5608 13460 5648
rect 13612 5608 13652 5648
rect 13900 5608 13940 5648
rect 14092 5608 14132 5648
rect 15340 5608 15380 5648
rect 15724 5608 15764 5648
rect 15916 5608 15956 5648
rect 16204 5608 16244 5648
rect 16492 5608 16532 5648
rect 16588 5608 16628 5648
rect 17068 5608 17108 5648
rect 17260 5608 17300 5648
rect 17452 5608 17492 5648
rect 18700 5608 18740 5648
rect 19180 5608 19220 5648
rect 19468 5608 19508 5648
rect 19564 5608 19604 5648
rect 20044 5608 20084 5648
rect 20236 5608 20276 5648
rect 1420 5440 1460 5480
rect 7756 5440 7796 5480
rect 9772 5440 9812 5480
rect 10252 5440 10292 5480
rect 12172 5440 12212 5480
rect 12652 5440 12692 5480
rect 13804 5440 13844 5480
rect 15532 5440 15572 5480
rect 15820 5440 15860 5480
rect 18892 5440 18932 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 15628 5104 15668 5144
rect 15916 5104 15956 5144
rect 17356 5104 17396 5144
rect 17740 5104 17780 5144
rect 6316 5020 6356 5060
rect 7372 5020 7412 5060
rect 8332 5020 8372 5060
rect 10348 5020 10388 5060
rect 11116 5020 11156 5060
rect 16588 5020 16628 5060
rect 19180 5020 19220 5060
rect 1228 4936 1268 4976
rect 1420 4936 1460 4976
rect 1612 4936 1652 4976
rect 2860 4936 2900 4976
rect 3244 4936 3284 4976
rect 4492 4936 4532 4976
rect 4876 4936 4916 4976
rect 6124 4936 6164 4976
rect 7660 4936 7700 4976
rect 7756 4936 7796 4976
rect 7948 4936 7988 4976
rect 8524 4922 8564 4962
rect 9004 4936 9044 4976
rect 9580 4936 9620 4976
rect 9964 4936 10004 4976
rect 10060 4936 10100 4976
rect 10636 4936 10676 4976
rect 10924 4936 10964 4976
rect 11308 4922 11348 4962
rect 11788 4936 11828 4976
rect 12268 4936 12308 4976
rect 12364 4936 12404 4976
rect 12748 4936 12788 4976
rect 12844 4936 12884 4976
rect 13132 4936 13172 4976
rect 13324 4936 13364 4976
rect 13420 4936 13460 4976
rect 13708 4936 13748 4976
rect 13804 4936 13844 4976
rect 13900 4936 13940 4976
rect 13996 4936 14036 4976
rect 14188 4936 14228 4976
rect 15436 4936 15476 4976
rect 15820 4936 15860 4976
rect 16204 4936 16244 4976
rect 16492 4936 16532 4976
rect 17068 4936 17108 4976
rect 17164 4936 17204 4976
rect 17836 4936 17876 4976
rect 18412 4936 18452 4976
rect 18508 4936 18548 4976
rect 18700 4936 18740 4976
rect 19276 4936 19316 4976
rect 19564 4936 19604 4976
rect 6508 4852 6548 4892
rect 6988 4852 7028 4892
rect 9484 4852 9524 4892
rect 19852 4852 19892 4892
rect 7756 4768 7796 4808
rect 10924 4768 10964 4808
rect 16876 4768 16916 4808
rect 18508 4768 18548 4808
rect 20044 4768 20084 4808
rect 1324 4684 1364 4724
rect 3052 4684 3092 4724
rect 4684 4684 4724 4724
rect 7180 4684 7220 4724
rect 13132 4684 13172 4724
rect 18028 4684 18068 4724
rect 18892 4684 18932 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 3436 4348 3476 4388
rect 6988 4348 7028 4388
rect 10924 4348 10964 4388
rect 13516 4348 13556 4388
rect 18220 4348 18260 4388
rect 5644 4264 5684 4304
rect 5932 4264 5972 4304
rect 6220 4264 6260 4304
rect 9100 4264 9140 4304
rect 9292 4264 9332 4304
rect 18604 4264 18644 4304
rect 19756 4264 19796 4304
rect 1228 4180 1268 4220
rect 4780 4180 4820 4220
rect 4876 4180 4916 4220
rect 9580 4191 9620 4231
rect 9964 4180 10004 4220
rect 10444 4180 10484 4220
rect 11596 4180 11636 4220
rect 16588 4180 16628 4220
rect 18508 4180 18548 4220
rect 18700 4180 18740 4220
rect 1516 4096 1556 4136
rect 1612 4096 1652 4136
rect 1708 4096 1748 4136
rect 1804 4096 1844 4136
rect 1996 4096 2036 4136
rect 3244 4096 3284 4136
rect 3820 4101 3860 4141
rect 4300 4096 4340 4136
rect 5260 4096 5300 4136
rect 5356 4096 5396 4136
rect 6508 4096 6548 4136
rect 6604 4096 6644 4136
rect 6700 4075 6740 4115
rect 6796 4096 6836 4136
rect 7084 4096 7124 4136
rect 7276 4096 7316 4136
rect 7468 4096 7508 4136
rect 7660 4096 7700 4136
rect 8908 4096 8948 4136
rect 10348 4096 10388 4136
rect 10540 4096 10580 4136
rect 10732 4096 10772 4136
rect 10924 4096 10964 4136
rect 11116 4096 11156 4136
rect 11308 4096 11348 4136
rect 11404 4096 11444 4136
rect 12076 4096 12116 4136
rect 13324 4096 13364 4136
rect 13708 4096 13748 4136
rect 13804 4096 13844 4136
rect 13900 4096 13940 4136
rect 14284 4096 14324 4136
rect 15532 4096 15572 4136
rect 16012 4096 16052 4136
rect 16108 4096 16148 4136
rect 16492 4096 16532 4136
rect 17068 4096 17108 4136
rect 17548 4101 17588 4141
rect 17932 4096 17972 4136
rect 18028 4096 18068 4136
rect 18220 4096 18260 4136
rect 18412 4096 18452 4136
rect 18796 4096 18836 4136
rect 19084 4096 19124 4136
rect 19372 4096 19412 4136
rect 19468 4096 19508 4136
rect 19948 4096 19988 4136
rect 20122 4101 20162 4141
rect 3628 4012 3668 4052
rect 15724 4012 15764 4052
rect 7372 3928 7412 3968
rect 9772 3928 9812 3968
rect 10156 3928 10196 3968
rect 11212 3928 11252 3968
rect 11788 3928 11828 3968
rect 13996 3928 14036 3968
rect 17740 3928 17780 3968
rect 20044 3928 20084 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 1420 3592 1460 3632
rect 3628 3592 3668 3632
rect 6508 3592 6548 3632
rect 8236 3592 8276 3632
rect 12076 3592 12116 3632
rect 17068 3592 17108 3632
rect 3436 3508 3476 3548
rect 6316 3508 6356 3548
rect 8524 3508 8564 3548
rect 15820 3508 15860 3548
rect 20044 3508 20084 3548
rect 1996 3424 2036 3464
rect 3244 3424 3284 3464
rect 3724 3424 3764 3464
rect 3820 3424 3860 3464
rect 3916 3424 3956 3464
rect 4588 3424 4628 3464
rect 4684 3405 4724 3445
rect 5644 3424 5684 3464
rect 6124 3410 6164 3450
rect 6796 3424 6836 3464
rect 8044 3424 8084 3464
rect 9196 3424 9236 3464
rect 9676 3424 9716 3464
rect 5068 3340 5108 3380
rect 5164 3340 5204 3380
rect 8668 3382 8708 3422
rect 10156 3424 10196 3464
rect 10252 3424 10292 3464
rect 11500 3424 11540 3464
rect 11596 3424 11636 3464
rect 11692 3424 11732 3464
rect 11788 3424 11828 3464
rect 12268 3424 12308 3464
rect 13516 3424 13556 3464
rect 13900 3424 13940 3464
rect 15148 3424 15188 3464
rect 15436 3424 15476 3464
rect 15724 3424 15764 3464
rect 16684 3424 16724 3464
rect 16780 3424 16820 3464
rect 16876 3424 16916 3464
rect 17260 3424 17300 3464
rect 17356 3424 17396 3464
rect 17548 3424 17588 3464
rect 17740 3424 17780 3464
rect 17932 3424 17972 3464
rect 18028 3424 18068 3464
rect 18220 3424 18260 3464
rect 18412 3424 18452 3464
rect 18604 3424 18644 3464
rect 18988 3424 19028 3464
rect 19180 3424 19220 3464
rect 19276 3424 19316 3464
rect 19468 3424 19508 3464
rect 19564 3424 19604 3464
rect 19708 3424 19748 3464
rect 19948 3424 19988 3464
rect 20129 3411 20169 3451
rect 9772 3340 9812 3380
rect 10732 3340 10772 3380
rect 11116 3340 11156 3380
rect 18700 3340 18740 3380
rect 18892 3340 18932 3380
rect 1708 3256 1748 3296
rect 4300 3256 4340 3296
rect 16300 3256 16340 3296
rect 17740 3256 17780 3296
rect 18796 3256 18836 3296
rect 10924 3172 10964 3212
rect 11308 3172 11348 3212
rect 13708 3172 13748 3212
rect 16108 3172 16148 3212
rect 17548 3172 17588 3212
rect 18220 3172 18260 3212
rect 19180 3172 19220 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 3628 2836 3668 2876
rect 5740 2836 5780 2876
rect 14092 2836 14132 2876
rect 17356 2836 17396 2876
rect 19468 2836 19508 2876
rect 1612 2752 1652 2792
rect 1900 2752 1940 2792
rect 4876 2752 4916 2792
rect 6124 2752 6164 2792
rect 6508 2752 6548 2792
rect 9292 2752 9332 2792
rect 17548 2752 17588 2792
rect 5068 2668 5108 2708
rect 6028 2668 6068 2708
rect 6220 2668 6260 2708
rect 7372 2668 7412 2708
rect 7468 2668 7508 2708
rect 11212 2679 11252 2719
rect 11884 2668 11924 2708
rect 12172 2668 12212 2708
rect 1420 2584 1460 2624
rect 2188 2584 2228 2624
rect 3436 2584 3476 2624
rect 4396 2584 4436 2624
rect 4492 2584 4532 2624
rect 5452 2584 5492 2624
rect 5548 2584 5588 2624
rect 5740 2584 5780 2624
rect 5932 2584 5972 2624
rect 6316 2584 6356 2624
rect 6892 2584 6932 2624
rect 6988 2584 7028 2624
rect 7948 2584 7988 2624
rect 8428 2598 8468 2638
rect 9004 2584 9044 2624
rect 9100 2584 9140 2624
rect 9772 2584 9812 2624
rect 11020 2584 11060 2624
rect 12076 2597 12116 2637
rect 12268 2584 12308 2624
rect 12652 2584 12692 2624
rect 13900 2584 13940 2624
rect 14284 2584 14324 2624
rect 15532 2584 15572 2624
rect 15724 2584 15764 2624
rect 16972 2584 17012 2624
rect 17548 2584 17588 2624
rect 18028 2584 18068 2624
rect 19276 2584 19316 2624
rect 19660 2584 19700 2624
rect 19756 2584 19796 2624
rect 19948 2584 19988 2624
rect 4012 2500 4052 2540
rect 4780 2500 4820 2540
rect 8620 2500 8660 2540
rect 17164 2500 17204 2540
rect 19852 2500 19892 2540
rect 20140 2500 20180 2540
rect 4204 2416 4244 2456
rect 5260 2416 5300 2456
rect 8812 2416 8852 2456
rect 9580 2416 9620 2456
rect 11404 2416 11444 2456
rect 11692 2416 11732 2456
rect 12460 2416 12500 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 1612 2080 1652 2120
rect 1900 2080 1940 2120
rect 5740 2080 5780 2120
rect 8332 2080 8372 2120
rect 9964 2080 10004 2120
rect 11980 2080 12020 2120
rect 17356 2080 17396 2120
rect 19372 2080 19412 2120
rect 19660 2080 19700 2120
rect 20236 2080 20276 2120
rect 8140 1996 8180 2036
rect 15532 1996 15572 2036
rect 2188 1912 2228 1952
rect 3436 1912 3476 1952
rect 4012 1912 4052 1952
rect 4108 1912 4148 1952
rect 4492 1912 4532 1952
rect 5068 1912 5108 1952
rect 5548 1907 5588 1947
rect 6412 1912 6452 1952
rect 6508 1912 6548 1952
rect 6988 1912 7028 1952
rect 7468 1912 7508 1952
rect 7948 1898 7988 1938
rect 8524 1912 8564 1952
rect 9772 1912 9812 1952
rect 10156 1912 10196 1952
rect 11404 1912 11444 1952
rect 12172 1912 12212 1952
rect 13420 1912 13460 1952
rect 13612 1912 13652 1952
rect 14860 1912 14900 1952
rect 15244 1912 15284 1952
rect 15340 1912 15380 1952
rect 15436 1912 15476 1952
rect 15916 1912 15956 1952
rect 17164 1912 17204 1952
rect 17932 1912 17972 1952
rect 19180 1912 19220 1952
rect 19660 1912 19700 1952
rect 19852 1912 19892 1952
rect 19948 1912 19988 1952
rect 20127 1912 20167 1952
rect 1228 1828 1268 1868
rect 4588 1828 4628 1868
rect 5932 1828 5972 1868
rect 6892 1828 6932 1868
rect 11596 1828 11636 1868
rect 17740 1828 17780 1868
rect 1708 1744 1748 1784
rect 3628 1744 3668 1784
rect 1420 1660 1460 1700
rect 6124 1660 6164 1700
rect 11788 1660 11828 1700
rect 15052 1660 15092 1700
rect 17548 1660 17588 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 9100 1324 9140 1364
rect 11116 1324 11156 1364
rect 12748 1324 12788 1364
rect 19468 1324 19508 1364
rect 1324 1240 1364 1280
rect 3916 1240 3956 1280
rect 4204 1240 4244 1280
rect 4684 1240 4724 1280
rect 7468 1240 7508 1280
rect 12940 1240 12980 1280
rect 1516 1156 1556 1196
rect 2476 1156 2516 1196
rect 2572 1156 2612 1196
rect 4876 1156 4916 1196
rect 5260 1156 5300 1196
rect 5644 1156 5684 1196
rect 9292 1156 9332 1196
rect 13900 1156 13940 1196
rect 19852 1156 19892 1196
rect 20236 1156 20276 1196
rect 1996 1072 2036 1112
rect 2092 1072 2132 1112
rect 3052 1072 3092 1112
rect 3532 1077 3572 1117
rect 6028 1072 6068 1112
rect 7276 1072 7316 1112
rect 7660 1072 7700 1112
rect 8908 1072 8948 1112
rect 9676 1072 9716 1112
rect 10924 1072 10964 1112
rect 11308 1072 11348 1112
rect 12556 1072 12596 1112
rect 12940 1072 12980 1112
rect 13132 1072 13172 1112
rect 13228 1072 13268 1112
rect 13420 1072 13460 1112
rect 13516 1072 13556 1112
rect 13612 1072 13652 1112
rect 13708 1072 13748 1112
rect 14380 1072 14420 1112
rect 15628 1072 15668 1112
rect 16012 1072 16052 1112
rect 17260 1072 17300 1112
rect 17452 1072 17492 1112
rect 17644 1072 17684 1112
rect 17740 1072 17780 1112
rect 18028 1072 18068 1112
rect 19276 1072 19316 1112
rect 3724 988 3764 1028
rect 17548 988 17588 1028
rect 1708 904 1748 944
rect 5068 904 5108 944
rect 5452 904 5492 944
rect 5836 904 5876 944
rect 9484 904 9524 944
rect 14188 904 14228 944
rect 15820 904 15860 944
rect 19660 904 19700 944
rect 20044 904 20084 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1227 42944 1269 42953
rect 1227 42904 1228 42944
rect 1268 42904 1269 42944
rect 1784 42928 1864 43008
rect 1976 42928 2056 43008
rect 2168 42928 2248 43008
rect 2360 42928 2440 43008
rect 2552 42928 2632 43008
rect 2744 42928 2824 43008
rect 2936 42928 3016 43008
rect 3128 42928 3208 43008
rect 3320 42928 3400 43008
rect 3512 42928 3592 43008
rect 3704 42928 3784 43008
rect 3896 42928 3976 43008
rect 4088 42928 4168 43008
rect 4280 42928 4360 43008
rect 4472 42928 4552 43008
rect 4664 42928 4744 43008
rect 4856 42928 4936 43008
rect 5048 42928 5128 43008
rect 5240 42928 5320 43008
rect 5432 42928 5512 43008
rect 5624 42928 5704 43008
rect 5816 42928 5896 43008
rect 6008 42928 6088 43008
rect 6200 42928 6280 43008
rect 6392 42928 6472 43008
rect 6584 42928 6664 43008
rect 6776 42928 6856 43008
rect 6968 42928 7048 43008
rect 7160 42928 7240 43008
rect 7352 42928 7432 43008
rect 7544 42928 7624 43008
rect 7736 42928 7816 43008
rect 7928 42928 8008 43008
rect 8120 42928 8200 43008
rect 8312 42928 8392 43008
rect 8504 42928 8584 43008
rect 8696 42928 8776 43008
rect 8888 42928 8968 43008
rect 9080 42928 9160 43008
rect 9272 42928 9352 43008
rect 9464 42928 9544 43008
rect 9656 42928 9736 43008
rect 9848 42928 9928 43008
rect 10040 42928 10120 43008
rect 10232 42928 10312 43008
rect 10424 42928 10504 43008
rect 10616 42928 10696 43008
rect 10808 42928 10888 43008
rect 11000 42928 11080 43008
rect 11192 42928 11272 43008
rect 11384 42928 11464 43008
rect 11576 42928 11656 43008
rect 11768 42928 11848 43008
rect 11960 42928 12040 43008
rect 12152 42928 12232 43008
rect 12344 42928 12424 43008
rect 12536 42928 12616 43008
rect 12728 42928 12808 43008
rect 12920 42928 13000 43008
rect 13112 42928 13192 43008
rect 13304 42928 13384 43008
rect 13496 42928 13576 43008
rect 13688 42928 13768 43008
rect 13880 42928 13960 43008
rect 14072 42928 14152 43008
rect 14264 42928 14344 43008
rect 14456 42928 14536 43008
rect 14648 42944 14728 43008
rect 14648 42928 14668 42944
rect 1227 42895 1269 42904
rect 1131 41600 1173 41609
rect 1131 41560 1132 41600
rect 1172 41560 1173 41600
rect 1131 41551 1173 41560
rect 1035 40340 1077 40349
rect 1035 40300 1036 40340
rect 1076 40300 1077 40340
rect 1035 40291 1077 40300
rect 75 39416 117 39425
rect 75 39376 76 39416
rect 116 39376 117 39416
rect 75 39367 117 39376
rect 76 39089 116 39367
rect 75 39080 117 39089
rect 75 39040 76 39080
rect 116 39040 117 39080
rect 75 39031 117 39040
rect 939 37232 981 37241
rect 939 37192 940 37232
rect 980 37192 981 37232
rect 939 37183 981 37192
rect 171 35384 213 35393
rect 171 35344 172 35384
rect 212 35344 213 35384
rect 171 35335 213 35344
rect 75 33284 117 33293
rect 75 33244 76 33284
rect 116 33244 117 33284
rect 75 33235 117 33244
rect 76 33041 116 33235
rect 75 33032 117 33041
rect 75 32992 76 33032
rect 116 32992 117 33032
rect 75 32983 117 32992
rect 75 32528 117 32537
rect 75 32488 76 32528
rect 116 32488 117 32528
rect 75 32479 117 32488
rect 76 32369 116 32479
rect 75 32360 117 32369
rect 75 32320 76 32360
rect 116 32320 117 32360
rect 75 32311 117 32320
rect 172 25229 212 35335
rect 555 34040 597 34049
rect 555 34000 556 34040
rect 596 34000 597 34040
rect 555 33991 597 34000
rect 363 31520 405 31529
rect 363 31480 364 31520
rect 404 31480 405 31520
rect 363 31471 405 31480
rect 364 31361 404 31471
rect 363 31352 405 31361
rect 363 31312 364 31352
rect 404 31312 405 31352
rect 363 31303 405 31312
rect 364 29000 404 31303
rect 556 30437 596 33991
rect 747 33704 789 33713
rect 747 33664 748 33704
rect 788 33664 789 33704
rect 747 33655 789 33664
rect 651 31520 693 31529
rect 651 31480 652 31520
rect 692 31480 693 31520
rect 651 31471 693 31480
rect 555 30428 597 30437
rect 555 30388 556 30428
rect 596 30388 597 30428
rect 555 30379 597 30388
rect 364 28960 500 29000
rect 171 25220 213 25229
rect 171 25180 172 25220
rect 212 25180 213 25220
rect 171 25171 213 25180
rect 267 21860 309 21869
rect 267 21820 268 21860
rect 308 21820 309 21860
rect 267 21811 309 21820
rect 75 20936 117 20945
rect 75 20896 76 20936
rect 116 20896 117 20936
rect 75 20887 117 20896
rect 76 20273 116 20887
rect 75 20264 117 20273
rect 75 20224 76 20264
rect 116 20224 117 20264
rect 75 20215 117 20224
rect 75 17408 117 17417
rect 75 17368 76 17408
rect 116 17368 117 17408
rect 75 17359 117 17368
rect 76 16661 116 17359
rect 171 17324 213 17333
rect 171 17284 172 17324
rect 212 17284 213 17324
rect 171 17275 213 17284
rect 75 16652 117 16661
rect 75 16612 76 16652
rect 116 16612 117 16652
rect 75 16603 117 16612
rect 75 10184 117 10193
rect 75 10144 76 10184
rect 116 10144 117 10184
rect 75 10135 117 10144
rect 76 8849 116 10135
rect 75 8840 117 8849
rect 75 8800 76 8840
rect 116 8800 117 8840
rect 75 8791 117 8800
rect 172 3305 212 17275
rect 268 4313 308 21811
rect 460 19265 500 28960
rect 555 23960 597 23969
rect 555 23920 556 23960
rect 596 23920 597 23960
rect 555 23911 597 23920
rect 556 19517 596 23911
rect 555 19508 597 19517
rect 555 19468 556 19508
rect 596 19468 597 19508
rect 555 19459 597 19468
rect 459 19256 501 19265
rect 459 19216 460 19256
rect 500 19216 501 19256
rect 459 19207 501 19216
rect 459 18584 501 18593
rect 459 18544 460 18584
rect 500 18544 501 18584
rect 459 18535 501 18544
rect 363 12116 405 12125
rect 363 12076 364 12116
rect 404 12076 405 12116
rect 363 12067 405 12076
rect 364 6329 404 12067
rect 460 11873 500 18535
rect 652 15821 692 31471
rect 748 26069 788 33655
rect 940 30605 980 37183
rect 939 30596 981 30605
rect 939 30556 940 30596
rect 980 30556 981 30596
rect 939 30547 981 30556
rect 939 30428 981 30437
rect 939 30388 940 30428
rect 980 30388 981 30428
rect 939 30379 981 30388
rect 843 30176 885 30185
rect 843 30136 844 30176
rect 884 30136 885 30176
rect 843 30127 885 30136
rect 747 26060 789 26069
rect 747 26020 748 26060
rect 788 26020 789 26060
rect 747 26011 789 26020
rect 747 25892 789 25901
rect 747 25852 748 25892
rect 788 25852 789 25892
rect 747 25843 789 25852
rect 748 20180 788 25843
rect 844 25565 884 30127
rect 843 25556 885 25565
rect 843 25516 844 25556
rect 884 25516 885 25556
rect 843 25507 885 25516
rect 748 20140 884 20180
rect 747 16988 789 16997
rect 747 16948 748 16988
rect 788 16948 789 16988
rect 747 16939 789 16948
rect 651 15812 693 15821
rect 651 15772 652 15812
rect 692 15772 693 15812
rect 651 15763 693 15772
rect 459 11864 501 11873
rect 459 11824 460 11864
rect 500 11824 501 11864
rect 459 11815 501 11824
rect 555 9008 597 9017
rect 555 8968 556 9008
rect 596 8968 597 9008
rect 555 8959 597 8968
rect 556 7337 596 8959
rect 555 7328 597 7337
rect 555 7288 556 7328
rect 596 7288 597 7328
rect 555 7279 597 7288
rect 363 6320 405 6329
rect 363 6280 364 6320
rect 404 6280 405 6320
rect 363 6271 405 6280
rect 748 4817 788 16939
rect 844 4901 884 20140
rect 940 17585 980 30379
rect 1036 23297 1076 40291
rect 1132 30185 1172 41551
rect 1228 41180 1268 42895
rect 1228 41131 1268 41140
rect 1612 41264 1652 41273
rect 1420 41012 1460 41021
rect 1420 40769 1460 40972
rect 1612 40937 1652 41224
rect 1611 40928 1653 40937
rect 1611 40888 1612 40928
rect 1652 40888 1653 40928
rect 1611 40879 1653 40888
rect 1419 40760 1461 40769
rect 1419 40720 1420 40760
rect 1460 40720 1461 40760
rect 1419 40711 1461 40720
rect 1323 40424 1365 40433
rect 1323 40384 1324 40424
rect 1364 40384 1365 40424
rect 1323 40375 1365 40384
rect 1324 40290 1364 40375
rect 1228 39752 1268 39761
rect 1323 39752 1365 39761
rect 1268 39712 1324 39752
rect 1364 39712 1365 39752
rect 1228 39703 1268 39712
rect 1323 39703 1365 39712
rect 1419 39416 1461 39425
rect 1419 39376 1420 39416
rect 1460 39376 1461 39416
rect 1419 39367 1461 39376
rect 1323 38996 1365 39005
rect 1323 38956 1324 38996
rect 1364 38956 1365 38996
rect 1323 38947 1365 38956
rect 1324 38862 1364 38947
rect 1323 38156 1365 38165
rect 1323 38116 1324 38156
rect 1364 38116 1365 38156
rect 1323 38107 1365 38116
rect 1324 38022 1364 38107
rect 1420 37820 1460 39367
rect 1515 38744 1557 38753
rect 1515 38704 1516 38744
rect 1556 38704 1557 38744
rect 1515 38695 1557 38704
rect 1516 38610 1556 38695
rect 1515 38408 1557 38417
rect 1515 38368 1516 38408
rect 1556 38368 1557 38408
rect 1515 38359 1557 38368
rect 1516 38274 1556 38359
rect 1324 37780 1460 37820
rect 1228 37484 1268 37493
rect 1228 35813 1268 37444
rect 1324 37400 1364 37780
rect 1419 37652 1461 37661
rect 1419 37612 1420 37652
rect 1460 37612 1461 37652
rect 1612 37652 1652 40879
rect 1804 40517 1844 42928
rect 1899 42104 1941 42113
rect 1899 42064 1900 42104
rect 1940 42064 1941 42104
rect 1899 42055 1941 42064
rect 1803 40508 1845 40517
rect 1803 40468 1804 40508
rect 1844 40468 1845 40508
rect 1803 40459 1845 40468
rect 1707 39080 1749 39089
rect 1707 39040 1708 39080
rect 1748 39040 1749 39080
rect 1707 39031 1749 39040
rect 1708 38954 1748 39031
rect 1708 38905 1748 38914
rect 1900 38408 1940 42055
rect 1996 40349 2036 42928
rect 2188 40424 2228 42928
rect 2283 42188 2325 42197
rect 2283 42148 2284 42188
rect 2324 42148 2325 42188
rect 2283 42139 2325 42148
rect 2092 40384 2228 40424
rect 1995 40340 2037 40349
rect 1995 40300 1996 40340
rect 2036 40300 2037 40340
rect 1995 40291 2037 40300
rect 1995 40172 2037 40181
rect 1995 40132 1996 40172
rect 2036 40132 2037 40172
rect 1995 40123 2037 40132
rect 1900 38359 1940 38368
rect 1899 38240 1941 38249
rect 1899 38200 1900 38240
rect 1940 38200 1941 38240
rect 1899 38191 1941 38200
rect 1707 38156 1749 38165
rect 1707 38116 1708 38156
rect 1748 38116 1749 38156
rect 1707 38107 1749 38116
rect 1708 38022 1748 38107
rect 1803 37988 1845 37997
rect 1803 37948 1804 37988
rect 1844 37948 1845 37988
rect 1803 37939 1845 37948
rect 1612 37612 1748 37652
rect 1419 37603 1461 37612
rect 1420 37518 1460 37603
rect 1324 37360 1460 37400
rect 1420 36728 1460 37360
rect 1708 37316 1748 37612
rect 1804 37414 1844 37939
rect 1804 37365 1844 37374
rect 1708 37276 1844 37316
rect 1611 37232 1653 37241
rect 1611 37192 1612 37232
rect 1652 37192 1653 37232
rect 1611 37183 1653 37192
rect 1612 37098 1652 37183
rect 1515 36980 1557 36989
rect 1515 36940 1516 36980
rect 1556 36940 1557 36980
rect 1515 36931 1557 36940
rect 1516 36896 1556 36931
rect 1516 36845 1556 36856
rect 1708 36728 1748 36737
rect 1420 36688 1708 36728
rect 1708 36679 1748 36688
rect 1324 36644 1364 36653
rect 1227 35804 1269 35813
rect 1227 35764 1228 35804
rect 1268 35764 1269 35804
rect 1227 35755 1269 35764
rect 1324 35225 1364 36604
rect 1804 36560 1844 37276
rect 1516 36520 1844 36560
rect 1419 35972 1461 35981
rect 1419 35932 1420 35972
rect 1460 35932 1461 35972
rect 1419 35923 1461 35932
rect 1420 35838 1460 35923
rect 1516 35300 1556 36520
rect 1612 36140 1652 36149
rect 1900 36140 1940 38191
rect 1652 36100 1940 36140
rect 1612 36091 1652 36100
rect 1611 35972 1653 35981
rect 1611 35932 1612 35972
rect 1652 35932 1653 35972
rect 1611 35923 1653 35932
rect 1803 35972 1845 35981
rect 1803 35932 1804 35972
rect 1844 35932 1845 35972
rect 1803 35923 1845 35932
rect 1420 35260 1556 35300
rect 1323 35216 1365 35225
rect 1323 35176 1324 35216
rect 1364 35176 1365 35216
rect 1323 35167 1365 35176
rect 1324 35048 1364 35059
rect 1420 35057 1460 35260
rect 1515 35132 1557 35141
rect 1515 35092 1516 35132
rect 1556 35092 1557 35132
rect 1515 35083 1557 35092
rect 1324 34973 1364 35008
rect 1419 35048 1461 35057
rect 1419 35008 1420 35048
rect 1460 35008 1461 35048
rect 1419 34999 1461 35008
rect 1516 34998 1556 35083
rect 1323 34964 1365 34973
rect 1323 34924 1324 34964
rect 1364 34924 1365 34964
rect 1323 34915 1365 34924
rect 1612 34796 1652 35923
rect 1804 35838 1844 35923
rect 1996 35888 2036 40123
rect 2092 36140 2132 40384
rect 2284 38249 2324 42139
rect 2380 41609 2420 42928
rect 2572 41945 2612 42928
rect 2571 41936 2613 41945
rect 2571 41896 2572 41936
rect 2612 41896 2613 41936
rect 2571 41887 2613 41896
rect 2379 41600 2421 41609
rect 2379 41560 2380 41600
rect 2420 41560 2421 41600
rect 2379 41551 2421 41560
rect 2379 41096 2421 41105
rect 2379 41056 2380 41096
rect 2420 41056 2421 41096
rect 2379 41047 2421 41056
rect 2380 38417 2420 41047
rect 2572 40424 2612 40433
rect 2764 40424 2804 42928
rect 2859 41264 2901 41273
rect 2859 41224 2860 41264
rect 2900 41224 2901 41264
rect 2859 41215 2901 41224
rect 2860 41130 2900 41215
rect 2956 40601 2996 42928
rect 3148 41609 3188 42928
rect 3340 42197 3380 42928
rect 3339 42188 3381 42197
rect 3339 42148 3340 42188
rect 3380 42148 3381 42188
rect 3339 42139 3381 42148
rect 3532 41768 3572 42928
rect 3244 41728 3572 41768
rect 3147 41600 3189 41609
rect 3147 41560 3148 41600
rect 3188 41560 3189 41600
rect 3147 41551 3189 41560
rect 3244 41432 3284 41728
rect 3339 41600 3381 41609
rect 3339 41560 3340 41600
rect 3380 41560 3381 41600
rect 3339 41551 3381 41560
rect 3148 41392 3284 41432
rect 3051 41096 3093 41105
rect 3051 41056 3052 41096
rect 3092 41056 3093 41096
rect 3051 41047 3093 41056
rect 3052 40962 3092 41047
rect 3148 40844 3188 41392
rect 3052 40804 3188 40844
rect 3244 41264 3284 41273
rect 2955 40592 2997 40601
rect 2955 40552 2956 40592
rect 2996 40552 2997 40592
rect 2955 40543 2997 40552
rect 2476 39752 2516 39761
rect 2572 39752 2612 40384
rect 2668 40384 2804 40424
rect 2955 40424 2997 40433
rect 2955 40384 2956 40424
rect 2996 40384 2997 40424
rect 2668 40088 2708 40384
rect 2955 40375 2997 40384
rect 2859 40340 2901 40349
rect 2764 40300 2860 40340
rect 2900 40300 2901 40340
rect 2764 40256 2804 40300
rect 2859 40291 2901 40300
rect 2956 40290 2996 40375
rect 2764 40207 2804 40216
rect 2668 40048 2804 40088
rect 2516 39712 2612 39752
rect 2476 39089 2516 39712
rect 2668 39500 2708 39509
rect 2475 39080 2517 39089
rect 2475 39040 2476 39080
rect 2516 39040 2517 39080
rect 2475 39031 2517 39040
rect 2571 38912 2613 38921
rect 2571 38872 2572 38912
rect 2612 38872 2613 38912
rect 2571 38863 2613 38872
rect 2379 38408 2421 38417
rect 2379 38368 2380 38408
rect 2420 38368 2421 38408
rect 2379 38359 2421 38368
rect 2283 38240 2325 38249
rect 2572 38240 2612 38863
rect 2283 38200 2284 38240
rect 2324 38200 2325 38240
rect 2283 38191 2325 38200
rect 2476 38200 2572 38240
rect 2187 38156 2229 38165
rect 2187 38116 2188 38156
rect 2228 38116 2229 38156
rect 2187 38107 2229 38116
rect 2188 38022 2228 38107
rect 2380 37988 2420 37997
rect 2284 37948 2380 37988
rect 2284 37568 2324 37948
rect 2380 37939 2420 37948
rect 2188 37528 2324 37568
rect 2188 36317 2228 37528
rect 2284 37400 2324 37409
rect 2187 36308 2229 36317
rect 2187 36268 2188 36308
rect 2228 36268 2229 36308
rect 2187 36259 2229 36268
rect 2092 36100 2228 36140
rect 2091 35972 2133 35981
rect 2091 35932 2092 35972
rect 2132 35932 2133 35972
rect 2091 35923 2133 35932
rect 1900 35848 2036 35888
rect 1900 35384 1940 35848
rect 1995 35720 2037 35729
rect 1995 35680 1996 35720
rect 2036 35680 2037 35720
rect 1995 35671 2037 35680
rect 1996 35586 2036 35671
rect 1708 35344 1940 35384
rect 1708 35048 1748 35344
rect 2092 35225 2132 35923
rect 1803 35216 1845 35225
rect 1803 35176 1804 35216
rect 1844 35176 1845 35216
rect 1803 35167 1845 35176
rect 1900 35216 1940 35225
rect 1708 34999 1748 35008
rect 1420 34756 1652 34796
rect 1323 34712 1365 34721
rect 1323 34672 1324 34712
rect 1364 34672 1365 34712
rect 1323 34663 1365 34672
rect 1324 34376 1364 34663
rect 1324 34327 1364 34336
rect 1228 34208 1268 34217
rect 1228 32873 1268 34168
rect 1324 33704 1364 33713
rect 1324 33545 1364 33664
rect 1420 33704 1460 34756
rect 1515 34628 1557 34637
rect 1515 34588 1516 34628
rect 1556 34588 1557 34628
rect 1515 34579 1557 34588
rect 1516 34376 1556 34579
rect 1516 34327 1556 34336
rect 1707 33872 1749 33881
rect 1707 33832 1708 33872
rect 1748 33832 1749 33872
rect 1707 33823 1749 33832
rect 1612 33713 1652 33798
rect 1611 33704 1653 33713
rect 1460 33664 1556 33704
rect 1420 33655 1460 33664
rect 1323 33536 1365 33545
rect 1323 33496 1324 33536
rect 1364 33496 1365 33536
rect 1323 33487 1365 33496
rect 1420 33536 1460 33545
rect 1227 32864 1269 32873
rect 1227 32824 1228 32864
rect 1268 32824 1269 32864
rect 1227 32815 1269 32824
rect 1420 32864 1460 33496
rect 1420 32815 1460 32824
rect 1516 32864 1556 33664
rect 1611 33664 1612 33704
rect 1652 33664 1653 33704
rect 1611 33655 1653 33664
rect 1611 33452 1653 33461
rect 1611 33412 1612 33452
rect 1652 33412 1653 33452
rect 1611 33403 1653 33412
rect 1516 32815 1556 32824
rect 1612 32453 1652 33403
rect 1708 32864 1748 33823
rect 1804 33041 1844 35167
rect 1900 35048 1940 35176
rect 2091 35216 2133 35225
rect 2091 35176 2092 35216
rect 2132 35176 2133 35216
rect 2091 35167 2133 35176
rect 1900 35008 2132 35048
rect 1899 34880 1941 34889
rect 1899 34840 1900 34880
rect 1940 34840 1941 34880
rect 1899 34831 1941 34840
rect 1900 33704 1940 34831
rect 1900 33629 1940 33664
rect 1899 33620 1941 33629
rect 1899 33580 1900 33620
rect 1940 33580 1941 33620
rect 1899 33571 1941 33580
rect 1995 33536 2037 33545
rect 1995 33496 1996 33536
rect 2036 33496 2037 33536
rect 1995 33487 2037 33496
rect 1996 33200 2036 33487
rect 2092 33461 2132 35008
rect 2091 33452 2133 33461
rect 2091 33412 2092 33452
rect 2132 33412 2133 33452
rect 2091 33403 2133 33412
rect 1961 33160 2036 33200
rect 1803 33032 1845 33041
rect 1803 32992 1804 33032
rect 1844 32992 1845 33032
rect 1803 32983 1845 32992
rect 1961 32879 2001 33160
rect 2188 33116 2228 36100
rect 1708 32815 1748 32824
rect 1803 32864 1845 32873
rect 1803 32824 1804 32864
rect 1844 32824 1845 32864
rect 1961 32830 2001 32839
rect 2092 33076 2228 33116
rect 1803 32815 1845 32824
rect 1804 32730 1844 32815
rect 1900 32696 1940 32705
rect 1900 32453 1940 32656
rect 1611 32444 1653 32453
rect 1611 32404 1612 32444
rect 1652 32404 1653 32444
rect 1611 32395 1653 32404
rect 1899 32444 1941 32453
rect 1899 32404 1900 32444
rect 1940 32404 1941 32444
rect 1899 32395 1941 32404
rect 1323 32276 1365 32285
rect 2092 32276 2132 33076
rect 2187 32948 2229 32957
rect 2187 32908 2188 32948
rect 2228 32908 2229 32948
rect 2187 32899 2229 32908
rect 2188 32814 2228 32899
rect 2284 32883 2324 37360
rect 2476 36737 2516 38200
rect 2572 38191 2612 38200
rect 2668 37652 2708 39460
rect 2764 38072 2804 40048
rect 2859 39584 2901 39593
rect 2859 39544 2860 39584
rect 2900 39544 2901 39584
rect 2859 39535 2901 39544
rect 2860 39450 2900 39535
rect 2955 38912 2997 38921
rect 2955 38872 2956 38912
rect 2996 38872 2997 38912
rect 2955 38863 2997 38872
rect 2956 38778 2996 38863
rect 2764 38032 2996 38072
rect 2572 37612 2708 37652
rect 2572 37400 2612 37612
rect 2764 37400 2804 37409
rect 2572 37360 2708 37400
rect 2475 36728 2517 36737
rect 2475 36688 2476 36728
rect 2516 36688 2517 36728
rect 2475 36679 2517 36688
rect 2571 36476 2613 36485
rect 2571 36436 2572 36476
rect 2612 36436 2613 36476
rect 2571 36427 2613 36436
rect 2572 36140 2612 36427
rect 2572 36091 2612 36100
rect 2380 35972 2420 35981
rect 2380 35393 2420 35932
rect 2571 35804 2613 35813
rect 2571 35764 2572 35804
rect 2612 35764 2613 35804
rect 2571 35755 2613 35764
rect 2379 35384 2421 35393
rect 2379 35344 2380 35384
rect 2420 35344 2421 35384
rect 2379 35335 2421 35344
rect 2475 35216 2517 35225
rect 2475 35176 2476 35216
rect 2516 35176 2517 35216
rect 2475 35167 2517 35176
rect 2379 33116 2421 33125
rect 2379 33076 2380 33116
rect 2420 33076 2421 33116
rect 2379 33067 2421 33076
rect 2380 32982 2420 33067
rect 2284 32843 2420 32883
rect 2187 32696 2229 32705
rect 2187 32656 2188 32696
rect 2228 32656 2229 32696
rect 2187 32647 2229 32656
rect 1228 32236 1324 32276
rect 1364 32236 1365 32276
rect 1228 32192 1268 32236
rect 1323 32227 1365 32236
rect 1420 32236 2132 32276
rect 1228 32143 1268 32152
rect 1323 32108 1365 32117
rect 1323 32068 1324 32108
rect 1364 32068 1365 32108
rect 1323 32059 1365 32068
rect 1227 31352 1269 31361
rect 1227 31312 1228 31352
rect 1268 31312 1269 31352
rect 1227 31303 1269 31312
rect 1228 31218 1268 31303
rect 1324 30680 1364 32059
rect 1420 30848 1460 32236
rect 1707 32108 1749 32117
rect 1707 32068 1708 32108
rect 1748 32068 1749 32108
rect 1707 32059 1749 32068
rect 2091 32108 2133 32117
rect 2091 32068 2092 32108
rect 2132 32068 2133 32108
rect 2091 32059 2133 32068
rect 1611 32024 1653 32033
rect 1611 31984 1612 32024
rect 1652 31984 1653 32024
rect 1611 31975 1653 31984
rect 1420 30799 1460 30808
rect 1612 30680 1652 31975
rect 1324 30640 1460 30680
rect 1227 30596 1269 30605
rect 1227 30556 1228 30596
rect 1268 30556 1269 30596
rect 1227 30547 1269 30556
rect 1228 30462 1268 30547
rect 1131 30176 1173 30185
rect 1131 30136 1132 30176
rect 1172 30136 1173 30176
rect 1131 30127 1173 30136
rect 1420 30017 1460 30640
rect 1612 30017 1652 30640
rect 1419 30008 1461 30017
rect 1419 29968 1420 30008
rect 1460 29968 1461 30008
rect 1419 29959 1461 29968
rect 1611 30008 1653 30017
rect 1611 29968 1612 30008
rect 1652 29968 1653 30008
rect 1611 29959 1653 29968
rect 1323 29840 1365 29849
rect 1323 29800 1324 29840
rect 1364 29800 1365 29840
rect 1323 29791 1365 29800
rect 1324 29706 1364 29791
rect 1228 29672 1268 29681
rect 1132 29632 1228 29672
rect 1132 29093 1172 29632
rect 1228 29623 1268 29632
rect 1228 29168 1268 29177
rect 1268 29128 1364 29168
rect 1228 29119 1268 29128
rect 1131 29084 1173 29093
rect 1131 29044 1132 29084
rect 1172 29044 1173 29084
rect 1131 29035 1173 29044
rect 1324 28925 1364 29128
rect 1323 28916 1365 28925
rect 1323 28876 1324 28916
rect 1364 28876 1365 28916
rect 1323 28867 1365 28876
rect 1420 28421 1460 29959
rect 1516 29840 1556 29849
rect 1516 29681 1556 29800
rect 1515 29672 1557 29681
rect 1515 29632 1516 29672
rect 1556 29632 1557 29672
rect 1515 29623 1557 29632
rect 1516 29009 1556 29623
rect 1708 29597 1748 32059
rect 1899 31352 1941 31361
rect 1899 31312 1900 31352
rect 1940 31312 1941 31352
rect 1899 31303 1941 31312
rect 1803 30680 1845 30689
rect 1803 30640 1804 30680
rect 1844 30640 1845 30680
rect 1803 30631 1845 30640
rect 1707 29588 1749 29597
rect 1707 29548 1708 29588
rect 1748 29548 1749 29588
rect 1707 29539 1749 29548
rect 1707 29252 1749 29261
rect 1707 29212 1708 29252
rect 1748 29212 1749 29252
rect 1707 29203 1749 29212
rect 1515 29000 1557 29009
rect 1515 28960 1516 29000
rect 1556 28960 1557 29000
rect 1515 28951 1557 28960
rect 1419 28412 1461 28421
rect 1419 28372 1420 28412
rect 1460 28372 1461 28412
rect 1419 28363 1461 28372
rect 1228 28328 1268 28337
rect 1132 28288 1228 28328
rect 1132 26237 1172 28288
rect 1228 28279 1268 28288
rect 1515 28244 1557 28253
rect 1515 28204 1516 28244
rect 1556 28204 1557 28244
rect 1515 28195 1557 28204
rect 1324 27656 1364 27665
rect 1324 27497 1364 27616
rect 1420 27656 1460 27665
rect 1323 27488 1365 27497
rect 1323 27448 1324 27488
rect 1364 27448 1365 27488
rect 1323 27439 1365 27448
rect 1227 27068 1269 27077
rect 1227 27028 1228 27068
rect 1268 27028 1269 27068
rect 1227 27019 1269 27028
rect 1228 26816 1268 27019
rect 1420 26909 1460 27616
rect 1419 26900 1461 26909
rect 1419 26860 1420 26900
rect 1460 26860 1461 26900
rect 1419 26851 1461 26860
rect 1131 26228 1173 26237
rect 1131 26188 1132 26228
rect 1172 26188 1173 26228
rect 1131 26179 1173 26188
rect 1228 26144 1268 26776
rect 1324 26816 1364 26825
rect 1324 26489 1364 26776
rect 1516 26648 1556 28195
rect 1611 27656 1653 27665
rect 1611 27616 1612 27656
rect 1652 27616 1653 27656
rect 1611 27607 1653 27616
rect 1612 27522 1652 27607
rect 1612 27404 1652 27413
rect 1612 26825 1652 27364
rect 1611 26816 1653 26825
rect 1611 26776 1612 26816
rect 1652 26776 1653 26816
rect 1611 26767 1653 26776
rect 1516 26599 1556 26608
rect 1323 26480 1365 26489
rect 1323 26440 1324 26480
rect 1364 26440 1365 26480
rect 1323 26431 1365 26440
rect 1419 26312 1461 26321
rect 1419 26272 1420 26312
rect 1460 26272 1461 26312
rect 1419 26263 1461 26272
rect 1420 26178 1460 26263
rect 1228 26095 1268 26104
rect 1323 26144 1365 26153
rect 1323 26104 1324 26144
rect 1364 26104 1365 26144
rect 1323 26095 1365 26104
rect 1515 26144 1557 26153
rect 1515 26104 1516 26144
rect 1556 26104 1557 26144
rect 1708 26144 1748 29203
rect 1804 28505 1844 30631
rect 1803 28496 1845 28505
rect 1803 28456 1804 28496
rect 1844 28456 1845 28496
rect 1803 28447 1845 28456
rect 1804 27749 1844 28447
rect 1803 27740 1845 27749
rect 1803 27700 1804 27740
rect 1844 27700 1845 27740
rect 1803 27691 1845 27700
rect 1804 27656 1844 27691
rect 1804 27605 1844 27616
rect 1900 27488 1940 31303
rect 2092 29000 2132 32059
rect 2188 30857 2228 32647
rect 2283 32360 2325 32369
rect 2283 32320 2284 32360
rect 2324 32320 2325 32360
rect 2283 32311 2325 32320
rect 2187 30848 2229 30857
rect 2187 30808 2188 30848
rect 2228 30808 2229 30848
rect 2187 30799 2229 30808
rect 2092 28960 2228 29000
rect 1995 28160 2037 28169
rect 1995 28120 1996 28160
rect 2036 28120 2037 28160
rect 1995 28111 2037 28120
rect 1804 27448 1940 27488
rect 1804 26816 1844 27448
rect 1904 26984 1946 26993
rect 1804 26767 1844 26776
rect 1900 26944 1905 26984
rect 1945 26944 1946 26984
rect 1900 26935 1946 26944
rect 1900 26816 1940 26935
rect 1804 26144 1844 26153
rect 1708 26104 1804 26144
rect 1515 26095 1557 26104
rect 1804 26095 1844 26104
rect 1900 26144 1940 26776
rect 1996 26237 2036 28111
rect 2091 27740 2133 27749
rect 2091 27700 2092 27740
rect 2132 27700 2133 27740
rect 2091 27691 2133 27700
rect 1995 26228 2037 26237
rect 1995 26188 1996 26228
rect 2036 26188 2037 26228
rect 1995 26179 2037 26188
rect 1324 26010 1364 26095
rect 1516 26010 1556 26095
rect 1227 25976 1269 25985
rect 1227 25936 1228 25976
rect 1268 25936 1269 25976
rect 1227 25927 1269 25936
rect 1228 25472 1268 25927
rect 1323 25640 1365 25649
rect 1323 25600 1324 25640
rect 1364 25600 1365 25640
rect 1323 25591 1365 25600
rect 1324 25481 1364 25591
rect 1132 25432 1268 25472
rect 1323 25472 1365 25481
rect 1323 25432 1324 25472
rect 1364 25432 1365 25472
rect 1035 23288 1077 23297
rect 1035 23248 1036 23288
rect 1076 23248 1077 23288
rect 1035 23239 1077 23248
rect 1132 23120 1172 25432
rect 1323 25423 1365 25432
rect 1228 25304 1268 25313
rect 1324 25304 1364 25423
rect 1268 25264 1364 25304
rect 1228 25255 1268 25264
rect 1900 25061 1940 26104
rect 2092 25892 2132 27691
rect 1996 25852 2132 25892
rect 1899 25052 1941 25061
rect 1899 25012 1900 25052
rect 1940 25012 1941 25052
rect 1899 25003 1941 25012
rect 1323 24968 1365 24977
rect 1323 24928 1324 24968
rect 1364 24928 1365 24968
rect 1323 24919 1365 24928
rect 1228 24632 1268 24641
rect 1324 24632 1364 24919
rect 1268 24592 1364 24632
rect 1228 24583 1268 24592
rect 1324 24473 1364 24592
rect 1323 24464 1365 24473
rect 1323 24424 1324 24464
rect 1364 24424 1365 24464
rect 1323 24415 1365 24424
rect 1996 24221 2036 25852
rect 2091 25472 2133 25481
rect 2091 25432 2092 25472
rect 2132 25432 2133 25472
rect 2091 25423 2133 25432
rect 1995 24212 2037 24221
rect 1995 24172 1996 24212
rect 2036 24172 2037 24212
rect 1995 24163 2037 24172
rect 2092 23969 2132 25423
rect 1515 23960 1557 23969
rect 1515 23920 1516 23960
rect 1556 23920 1557 23960
rect 1515 23911 1557 23920
rect 2091 23960 2133 23969
rect 2091 23920 2092 23960
rect 2132 23920 2133 23960
rect 2091 23911 2133 23920
rect 1420 23801 1460 23886
rect 1419 23792 1461 23801
rect 1419 23752 1420 23792
rect 1460 23752 1461 23792
rect 1419 23743 1461 23752
rect 1516 23792 1556 23911
rect 1708 23836 1940 23876
rect 1516 23743 1556 23752
rect 1612 23792 1652 23801
rect 1324 23633 1364 23718
rect 1323 23624 1365 23633
rect 1323 23584 1324 23624
rect 1364 23584 1365 23624
rect 1323 23575 1365 23584
rect 1323 23372 1365 23381
rect 1323 23332 1324 23372
rect 1364 23332 1365 23372
rect 1323 23323 1365 23332
rect 1036 23080 1172 23120
rect 1036 21617 1076 23080
rect 1324 23036 1364 23323
rect 1515 23288 1557 23297
rect 1515 23248 1516 23288
rect 1556 23248 1557 23288
rect 1515 23239 1557 23248
rect 1516 23154 1556 23239
rect 1324 22987 1364 22996
rect 1612 22793 1652 23752
rect 1708 23633 1748 23836
rect 1900 23792 1940 23836
rect 1900 23743 1940 23752
rect 1996 23792 2036 23801
rect 1707 23624 1749 23633
rect 1707 23584 1708 23624
rect 1748 23584 1749 23624
rect 1707 23575 1749 23584
rect 1804 23624 1844 23633
rect 1707 23120 1749 23129
rect 1707 23080 1708 23120
rect 1748 23080 1749 23120
rect 1707 23071 1749 23080
rect 1708 22986 1748 23071
rect 1804 22961 1844 23584
rect 1899 23624 1941 23633
rect 1899 23584 1900 23624
rect 1940 23584 1941 23624
rect 1899 23575 1941 23584
rect 1900 23120 1940 23575
rect 1996 23297 2036 23752
rect 2092 23792 2132 23911
rect 2188 23792 2228 28960
rect 2284 28925 2324 32311
rect 2283 28916 2325 28925
rect 2283 28876 2284 28916
rect 2324 28876 2325 28916
rect 2283 28867 2325 28876
rect 2284 28160 2324 28867
rect 2380 28589 2420 32843
rect 2476 32369 2516 35167
rect 2572 35141 2612 35755
rect 2571 35132 2613 35141
rect 2571 35092 2572 35132
rect 2612 35092 2613 35132
rect 2571 35083 2613 35092
rect 2668 32864 2708 37360
rect 2764 35981 2804 37360
rect 2860 37400 2900 37409
rect 2860 37157 2900 37360
rect 2859 37148 2901 37157
rect 2859 37108 2860 37148
rect 2900 37108 2901 37148
rect 2859 37099 2901 37108
rect 2956 36812 2996 38032
rect 3052 36905 3092 40804
rect 3147 40424 3189 40433
rect 3147 40384 3148 40424
rect 3188 40384 3189 40424
rect 3147 40375 3189 40384
rect 3148 39761 3188 40375
rect 3147 39752 3189 39761
rect 3147 39712 3148 39752
rect 3188 39712 3189 39752
rect 3147 39703 3189 39712
rect 3148 39618 3188 39703
rect 3244 39005 3284 41224
rect 3340 40676 3380 41551
rect 3724 41012 3764 42928
rect 3916 42449 3956 42928
rect 3915 42440 3957 42449
rect 3915 42400 3916 42440
rect 3956 42400 3957 42440
rect 3915 42391 3957 42400
rect 3532 40972 3764 41012
rect 3340 40636 3476 40676
rect 3339 39920 3381 39929
rect 3339 39880 3340 39920
rect 3380 39880 3381 39920
rect 3339 39871 3381 39880
rect 3340 39425 3380 39871
rect 3339 39416 3381 39425
rect 3339 39376 3340 39416
rect 3380 39376 3381 39416
rect 3339 39367 3381 39376
rect 3243 38996 3285 39005
rect 3243 38956 3244 38996
rect 3284 38956 3285 38996
rect 3243 38947 3285 38956
rect 3340 38996 3380 39005
rect 3148 38744 3188 38753
rect 3148 37829 3188 38704
rect 3340 38333 3380 38956
rect 3339 38324 3381 38333
rect 3339 38284 3340 38324
rect 3380 38284 3381 38324
rect 3339 38275 3381 38284
rect 3147 37820 3189 37829
rect 3147 37780 3148 37820
rect 3188 37780 3189 37820
rect 3147 37771 3189 37780
rect 3436 37568 3476 40636
rect 3532 39089 3572 40972
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 3627 39164 3669 39173
rect 3627 39124 3628 39164
rect 3668 39124 3669 39164
rect 3627 39115 3669 39124
rect 3531 39080 3573 39089
rect 3531 39040 3532 39080
rect 3572 39040 3573 39080
rect 3531 39031 3573 39040
rect 3531 38744 3573 38753
rect 3531 38704 3532 38744
rect 3572 38704 3573 38744
rect 3531 38695 3573 38704
rect 3532 38610 3572 38695
rect 3628 38492 3668 39115
rect 3915 38912 3957 38921
rect 3915 38872 3916 38912
rect 3956 38872 3957 38912
rect 3915 38863 3957 38872
rect 3819 38744 3861 38753
rect 3819 38704 3820 38744
rect 3860 38704 3861 38744
rect 3819 38695 3861 38704
rect 3820 38610 3860 38695
rect 3148 37528 3476 37568
rect 3532 38452 3668 38492
rect 3051 36896 3093 36905
rect 3051 36856 3052 36896
rect 3092 36856 3093 36896
rect 3051 36847 3093 36856
rect 2860 36772 2996 36812
rect 2763 35972 2805 35981
rect 2763 35932 2764 35972
rect 2804 35932 2805 35972
rect 2763 35923 2805 35932
rect 2764 35804 2804 35923
rect 2764 35755 2804 35764
rect 2763 34796 2805 34805
rect 2763 34756 2764 34796
rect 2804 34756 2805 34796
rect 2763 34747 2805 34756
rect 2764 34376 2804 34747
rect 2764 33041 2804 34336
rect 2763 33032 2805 33041
rect 2763 32992 2764 33032
rect 2804 32992 2805 33032
rect 2763 32983 2805 32992
rect 2668 32815 2708 32824
rect 2763 32864 2805 32873
rect 2763 32824 2764 32864
rect 2804 32824 2805 32864
rect 2763 32815 2805 32824
rect 2764 32730 2804 32815
rect 2763 32612 2805 32621
rect 2763 32572 2764 32612
rect 2804 32572 2805 32612
rect 2763 32563 2805 32572
rect 2475 32360 2517 32369
rect 2475 32320 2476 32360
rect 2516 32320 2517 32360
rect 2475 32311 2517 32320
rect 2476 32192 2516 32201
rect 2476 31529 2516 32152
rect 2764 32033 2804 32563
rect 2860 32360 2900 36772
rect 3051 36728 3093 36737
rect 2956 36707 3052 36728
rect 2996 36688 3052 36707
rect 3092 36688 3093 36728
rect 3051 36679 3093 36688
rect 2956 36658 2996 36667
rect 3148 36644 3188 37528
rect 3340 37400 3380 37409
rect 3244 37380 3284 37389
rect 3244 37241 3284 37340
rect 3243 37232 3285 37241
rect 3243 37192 3244 37232
rect 3284 37192 3285 37232
rect 3243 37183 3285 37192
rect 3340 37064 3380 37360
rect 3532 37148 3572 38452
rect 3819 38240 3861 38249
rect 3916 38240 3956 38863
rect 3819 38200 3820 38240
rect 3860 38200 3956 38240
rect 4012 38744 4052 38753
rect 3819 38191 3861 38200
rect 3820 38106 3860 38191
rect 4012 38156 4052 38704
rect 4108 38240 4148 42928
rect 4204 40424 4244 40433
rect 4204 39425 4244 40384
rect 4203 39416 4245 39425
rect 4203 39376 4204 39416
rect 4244 39376 4245 39416
rect 4203 39367 4245 39376
rect 4203 39080 4245 39089
rect 4203 39040 4204 39080
rect 4244 39040 4245 39080
rect 4203 39031 4245 39040
rect 4204 38585 4244 39031
rect 4203 38576 4245 38585
rect 4203 38536 4204 38576
rect 4244 38536 4245 38576
rect 4203 38527 4245 38536
rect 4204 38408 4244 38417
rect 4300 38408 4340 42928
rect 4492 41609 4532 42928
rect 4684 42113 4724 42928
rect 4683 42104 4725 42113
rect 4683 42064 4684 42104
rect 4724 42064 4725 42104
rect 4683 42055 4725 42064
rect 4876 41768 4916 42928
rect 5068 41777 5108 42928
rect 5260 42533 5300 42928
rect 5259 42524 5301 42533
rect 5259 42484 5260 42524
rect 5300 42484 5301 42524
rect 5259 42475 5301 42484
rect 4780 41728 4916 41768
rect 5067 41768 5109 41777
rect 5067 41728 5068 41768
rect 5108 41728 5109 41768
rect 4491 41600 4533 41609
rect 4491 41560 4492 41600
rect 4532 41560 4533 41600
rect 4491 41551 4533 41560
rect 4491 41264 4533 41273
rect 4491 41224 4492 41264
rect 4532 41224 4533 41264
rect 4491 41215 4533 41224
rect 4492 40853 4532 41215
rect 4683 41012 4725 41021
rect 4683 40972 4684 41012
rect 4724 40972 4725 41012
rect 4683 40963 4725 40972
rect 4684 40878 4724 40963
rect 4491 40844 4533 40853
rect 4491 40804 4492 40844
rect 4532 40804 4533 40844
rect 4491 40795 4533 40804
rect 4780 40517 4820 41728
rect 5067 41719 5109 41728
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 5067 41432 5109 41441
rect 5067 41392 5068 41432
rect 5108 41392 5109 41432
rect 5067 41383 5109 41392
rect 4971 41264 5013 41273
rect 4971 41224 4972 41264
rect 5012 41224 5013 41264
rect 4971 41215 5013 41224
rect 5068 41264 5108 41383
rect 5260 41273 5300 41358
rect 5068 41215 5108 41224
rect 5259 41264 5301 41273
rect 5259 41224 5260 41264
rect 5300 41224 5301 41264
rect 5259 41215 5301 41224
rect 4972 41130 5012 41215
rect 5452 41180 5492 42928
rect 5644 41525 5684 42928
rect 5739 42524 5781 42533
rect 5739 42484 5740 42524
rect 5780 42484 5781 42524
rect 5739 42475 5781 42484
rect 5643 41516 5685 41525
rect 5643 41476 5644 41516
rect 5684 41476 5685 41516
rect 5643 41467 5685 41476
rect 5644 41264 5684 41273
rect 5452 41140 5588 41180
rect 5260 41012 5300 41021
rect 5260 40601 5300 40972
rect 5355 41012 5397 41021
rect 5355 40972 5356 41012
rect 5396 40972 5397 41012
rect 5355 40963 5397 40972
rect 5452 41012 5492 41021
rect 5259 40592 5301 40601
rect 5259 40552 5260 40592
rect 5300 40552 5301 40592
rect 5259 40543 5301 40552
rect 4779 40508 4821 40517
rect 4779 40468 4780 40508
rect 4820 40468 4821 40508
rect 4779 40459 4821 40468
rect 4875 40424 4917 40433
rect 4875 40384 4876 40424
rect 4916 40384 4917 40424
rect 4875 40375 4917 40384
rect 4876 40290 4916 40375
rect 4396 40256 4436 40265
rect 4684 40256 4724 40265
rect 4436 40216 4532 40256
rect 4396 40207 4436 40216
rect 4396 39752 4436 39761
rect 4396 39425 4436 39712
rect 4395 39416 4437 39425
rect 4395 39376 4396 39416
rect 4436 39376 4437 39416
rect 4395 39367 4437 39376
rect 4395 39164 4437 39173
rect 4395 39124 4396 39164
rect 4436 39124 4437 39164
rect 4395 39115 4437 39124
rect 4396 38996 4436 39115
rect 4396 38947 4436 38956
rect 4395 38576 4437 38585
rect 4395 38536 4396 38576
rect 4436 38536 4437 38576
rect 4395 38527 4437 38536
rect 4244 38368 4340 38408
rect 4396 38408 4436 38527
rect 4204 38359 4244 38368
rect 4396 38359 4436 38368
rect 4395 38240 4437 38249
rect 4108 38200 4244 38240
rect 4052 38116 4148 38156
rect 4012 38107 4052 38116
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3723 37652 3765 37661
rect 3723 37612 3724 37652
rect 3764 37612 3765 37652
rect 3723 37603 3765 37612
rect 3627 37484 3669 37493
rect 3627 37444 3628 37484
rect 3668 37444 3669 37484
rect 3627 37435 3669 37444
rect 3628 37350 3668 37435
rect 3627 37232 3669 37241
rect 3627 37192 3628 37232
rect 3668 37192 3669 37232
rect 3627 37183 3669 37192
rect 3244 37024 3380 37064
rect 3436 37108 3572 37148
rect 3244 36905 3284 37024
rect 3243 36896 3285 36905
rect 3243 36856 3244 36896
rect 3284 36856 3285 36896
rect 3243 36847 3285 36856
rect 3339 36728 3381 36737
rect 3339 36688 3340 36728
rect 3380 36688 3381 36728
rect 3339 36679 3381 36688
rect 3436 36728 3476 37108
rect 3532 36821 3572 36843
rect 3531 36812 3573 36821
rect 3628 36812 3668 37183
rect 3531 36772 3532 36812
rect 3572 36772 3668 36812
rect 3531 36763 3573 36772
rect 3532 36748 3572 36763
rect 3532 36699 3572 36708
rect 3436 36679 3476 36688
rect 3148 36604 3284 36644
rect 2955 36476 2997 36485
rect 3148 36476 3188 36485
rect 2955 36436 2956 36476
rect 2996 36436 2997 36476
rect 2955 36427 2997 36436
rect 3052 36436 3148 36476
rect 2956 35902 2996 36427
rect 2956 35853 2996 35862
rect 3052 34628 3092 36436
rect 3148 36427 3188 36436
rect 2956 34588 3092 34628
rect 3148 35216 3188 35225
rect 2956 34385 2996 34588
rect 3148 34544 3188 35176
rect 3244 34712 3284 36604
rect 3340 35477 3380 36679
rect 3435 36560 3477 36569
rect 3435 36520 3436 36560
rect 3476 36520 3477 36560
rect 3435 36511 3477 36520
rect 3436 35888 3476 36511
rect 3724 36476 3764 37603
rect 3819 37232 3861 37241
rect 3819 37192 3820 37232
rect 3860 37192 3861 37232
rect 3819 37183 3861 37192
rect 4108 37232 4148 38116
rect 3820 37098 3860 37183
rect 3915 36812 3957 36821
rect 3915 36772 3916 36812
rect 3956 36772 3957 36812
rect 3915 36763 3957 36772
rect 3916 36728 3956 36763
rect 3916 36677 3956 36688
rect 4011 36644 4053 36653
rect 4011 36604 4012 36644
rect 4052 36604 4053 36644
rect 4011 36595 4053 36604
rect 4012 36510 4052 36595
rect 3436 35839 3476 35848
rect 3532 36436 3764 36476
rect 3532 35720 3572 36436
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3915 36140 3957 36149
rect 3915 36100 3916 36140
rect 3956 36100 3957 36140
rect 3915 36091 3957 36100
rect 3916 35972 3956 36091
rect 3916 35923 3956 35932
rect 4012 35888 4052 35899
rect 4012 35813 4052 35848
rect 4011 35804 4053 35813
rect 4011 35764 4012 35804
rect 4052 35764 4053 35804
rect 4011 35755 4053 35764
rect 3436 35680 3572 35720
rect 3339 35468 3381 35477
rect 3339 35428 3340 35468
rect 3380 35428 3381 35468
rect 3339 35419 3381 35428
rect 3339 34964 3381 34973
rect 3339 34924 3340 34964
rect 3380 34924 3381 34964
rect 3339 34915 3381 34924
rect 3340 34830 3380 34915
rect 3244 34672 3380 34712
rect 3340 34628 3380 34672
rect 3340 34579 3380 34588
rect 3052 34504 3188 34544
rect 2955 34376 2997 34385
rect 2955 34336 2956 34376
rect 2996 34336 2997 34376
rect 2955 34327 2997 34336
rect 2956 34208 2996 34217
rect 2956 33629 2996 34168
rect 3052 33704 3092 34504
rect 3436 34460 3476 35680
rect 4011 35384 4053 35393
rect 4011 35344 4012 35384
rect 4052 35344 4053 35384
rect 4011 35335 4053 35344
rect 3819 35132 3861 35141
rect 3819 35092 3820 35132
rect 3860 35092 3861 35132
rect 3819 35083 3861 35092
rect 3531 35048 3573 35057
rect 3531 35008 3532 35048
rect 3572 35008 3573 35048
rect 3531 34999 3573 35008
rect 3532 34914 3572 34999
rect 3820 34998 3860 35083
rect 4012 35048 4052 35335
rect 4108 35057 4148 37192
rect 4204 36989 4244 38200
rect 4395 38200 4396 38240
rect 4436 38200 4437 38240
rect 4395 38191 4437 38200
rect 4300 37484 4340 37493
rect 4203 36980 4245 36989
rect 4203 36940 4204 36980
rect 4244 36940 4245 36980
rect 4203 36931 4245 36940
rect 4203 36644 4245 36653
rect 4203 36604 4204 36644
rect 4244 36604 4245 36644
rect 4203 36595 4245 36604
rect 4204 36149 4244 36595
rect 4203 36140 4245 36149
rect 4203 36100 4204 36140
rect 4244 36100 4245 36140
rect 4203 36091 4245 36100
rect 4203 35216 4245 35225
rect 4203 35176 4204 35216
rect 4244 35176 4245 35216
rect 4203 35167 4245 35176
rect 4204 35082 4244 35167
rect 4012 34999 4052 35008
rect 4107 35048 4149 35057
rect 4107 35008 4108 35048
rect 4148 35008 4149 35048
rect 4107 34999 4149 35008
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 4203 34796 4245 34805
rect 4203 34756 4204 34796
rect 4244 34756 4245 34796
rect 4203 34747 4245 34756
rect 3148 34447 3188 34456
rect 3436 34420 3716 34460
rect 3148 34217 3188 34407
rect 3676 34418 3716 34420
rect 3243 34376 3285 34385
rect 3243 34336 3244 34376
rect 3284 34336 3285 34376
rect 3676 34369 3716 34378
rect 4204 34376 4244 34747
rect 3243 34327 3285 34336
rect 4204 34327 4244 34336
rect 3147 34208 3189 34217
rect 3147 34168 3148 34208
rect 3188 34168 3189 34208
rect 3147 34159 3189 34168
rect 3148 33704 3188 33713
rect 3052 33664 3148 33704
rect 2955 33620 2997 33629
rect 2955 33580 2956 33620
rect 2996 33580 2997 33620
rect 2955 33571 2997 33580
rect 3148 33461 3188 33664
rect 3147 33452 3189 33461
rect 3147 33412 3148 33452
rect 3188 33412 3189 33452
rect 3147 33403 3189 33412
rect 2955 33368 2997 33377
rect 2955 33328 2956 33368
rect 2996 33328 2997 33368
rect 2955 33319 2997 33328
rect 2860 32311 2900 32320
rect 2763 32024 2805 32033
rect 2763 31984 2764 32024
rect 2804 31984 2805 32024
rect 2763 31975 2805 31984
rect 2668 31940 2708 31949
rect 2475 31520 2517 31529
rect 2475 31480 2476 31520
rect 2516 31480 2517 31520
rect 2475 31471 2517 31480
rect 2668 31361 2708 31900
rect 2476 31352 2516 31361
rect 2476 30605 2516 31312
rect 2667 31352 2709 31361
rect 2667 31312 2668 31352
rect 2708 31312 2709 31352
rect 2667 31303 2709 31312
rect 2668 31184 2708 31193
rect 2475 30596 2517 30605
rect 2475 30556 2476 30596
rect 2516 30556 2517 30596
rect 2475 30547 2517 30556
rect 2476 29168 2516 30547
rect 2668 29261 2708 31144
rect 2764 29840 2804 31975
rect 2956 31352 2996 33319
rect 3148 32957 3188 33042
rect 3244 33041 3284 34327
rect 3531 34292 3573 34301
rect 3531 34252 3532 34292
rect 3572 34252 3573 34292
rect 3531 34243 3573 34252
rect 3532 34158 3572 34243
rect 4203 34208 4245 34217
rect 4203 34168 4204 34208
rect 4244 34168 4245 34208
rect 4203 34159 4245 34168
rect 3531 34040 3573 34049
rect 3531 34000 3532 34040
rect 3572 34000 3573 34040
rect 3531 33991 3573 34000
rect 3532 33872 3572 33991
rect 3532 33823 3572 33832
rect 3819 33872 3861 33881
rect 3819 33832 3820 33872
rect 3860 33832 3861 33872
rect 3819 33823 3861 33832
rect 3820 33738 3860 33823
rect 4012 33704 4052 33713
rect 3435 33620 3477 33629
rect 3435 33580 3436 33620
rect 3476 33580 3477 33620
rect 3435 33571 3477 33580
rect 3340 33452 3380 33461
rect 3243 33032 3285 33041
rect 3243 32992 3244 33032
rect 3284 32992 3285 33032
rect 3243 32983 3285 32992
rect 3147 32948 3189 32957
rect 3147 32908 3148 32948
rect 3188 32908 3189 32948
rect 3147 32899 3189 32908
rect 3243 32864 3285 32873
rect 3243 32824 3244 32864
rect 3284 32824 3285 32864
rect 3243 32815 3285 32824
rect 3244 32730 3284 32815
rect 3051 32696 3093 32705
rect 3051 32656 3052 32696
rect 3092 32656 3093 32696
rect 3051 32647 3093 32656
rect 3052 32108 3092 32647
rect 3340 32621 3380 33412
rect 3339 32612 3381 32621
rect 3339 32572 3340 32612
rect 3380 32572 3381 32612
rect 3339 32563 3381 32572
rect 3243 32360 3285 32369
rect 3243 32320 3244 32360
rect 3284 32320 3285 32360
rect 3243 32311 3285 32320
rect 3244 32226 3284 32311
rect 3436 32187 3476 33571
rect 4012 33452 4052 33664
rect 4107 33704 4149 33713
rect 4107 33664 4108 33704
rect 4148 33664 4149 33704
rect 4107 33655 4149 33664
rect 4108 33570 4148 33655
rect 4012 33412 4148 33452
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 3531 33032 3573 33041
rect 3531 32992 3532 33032
rect 3572 32992 3573 33032
rect 3531 32983 3573 32992
rect 3436 32138 3476 32147
rect 3052 32059 3092 32068
rect 3148 31352 3188 31361
rect 2956 31312 3148 31352
rect 2955 31184 2997 31193
rect 2955 31144 2956 31184
rect 2996 31144 2997 31184
rect 2955 31135 2997 31144
rect 2956 31050 2996 31135
rect 2860 30680 2900 30691
rect 2860 30605 2900 30640
rect 2859 30596 2901 30605
rect 2859 30556 2860 30596
rect 2900 30556 2901 30596
rect 2859 30547 2901 30556
rect 2667 29252 2709 29261
rect 2667 29212 2668 29252
rect 2708 29212 2709 29252
rect 2667 29203 2709 29212
rect 2379 28580 2421 28589
rect 2379 28540 2380 28580
rect 2420 28540 2421 28580
rect 2379 28531 2421 28540
rect 2476 28328 2516 29128
rect 2668 28916 2708 28925
rect 2476 28279 2516 28288
rect 2572 28876 2668 28916
rect 2284 28120 2516 28160
rect 2284 26816 2324 26825
rect 2284 26741 2324 26776
rect 2380 26816 2420 26825
rect 2283 26732 2325 26741
rect 2283 26692 2284 26732
rect 2324 26692 2325 26732
rect 2283 26683 2325 26692
rect 2284 26144 2324 26683
rect 2380 26657 2420 26776
rect 2379 26648 2421 26657
rect 2379 26608 2380 26648
rect 2420 26608 2421 26648
rect 2379 26599 2421 26608
rect 2284 26095 2324 26104
rect 2380 26060 2420 26599
rect 2284 23792 2324 23801
rect 2188 23752 2284 23792
rect 2092 23743 2132 23752
rect 2091 23624 2133 23633
rect 2091 23584 2092 23624
rect 2132 23584 2133 23624
rect 2091 23575 2133 23584
rect 1995 23288 2037 23297
rect 1995 23248 1996 23288
rect 2036 23248 2037 23288
rect 1995 23239 2037 23248
rect 1900 23080 2036 23120
rect 1803 22952 1845 22961
rect 1803 22912 1804 22952
rect 1844 22912 1845 22952
rect 1803 22903 1845 22912
rect 1611 22784 1653 22793
rect 1611 22744 1612 22784
rect 1652 22744 1653 22784
rect 1611 22735 1653 22744
rect 1516 22541 1556 22626
rect 1707 22616 1749 22625
rect 1707 22576 1708 22616
rect 1748 22576 1749 22616
rect 1707 22567 1749 22576
rect 1515 22532 1557 22541
rect 1515 22492 1516 22532
rect 1556 22492 1557 22532
rect 1515 22483 1557 22492
rect 1708 22532 1748 22567
rect 1708 22481 1748 22492
rect 1324 22364 1364 22373
rect 1900 22364 1940 22373
rect 1364 22324 1652 22364
rect 1324 22315 1364 22324
rect 1515 21776 1557 21785
rect 1515 21736 1516 21776
rect 1556 21736 1557 21776
rect 1515 21727 1557 21736
rect 1323 21692 1365 21701
rect 1323 21652 1324 21692
rect 1364 21652 1365 21692
rect 1323 21643 1365 21652
rect 1035 21608 1077 21617
rect 1035 21568 1036 21608
rect 1076 21568 1077 21608
rect 1035 21559 1077 21568
rect 939 17576 981 17585
rect 939 17536 940 17576
rect 980 17536 981 17576
rect 939 17527 981 17536
rect 939 15728 981 15737
rect 939 15688 940 15728
rect 980 15688 981 15728
rect 939 15679 981 15688
rect 940 11033 980 15679
rect 939 11024 981 11033
rect 939 10984 940 11024
rect 980 10984 981 11024
rect 939 10975 981 10984
rect 939 6320 981 6329
rect 939 6280 940 6320
rect 980 6280 981 6320
rect 939 6271 981 6280
rect 843 4892 885 4901
rect 843 4852 844 4892
rect 884 4852 885 4892
rect 843 4843 885 4852
rect 747 4808 789 4817
rect 747 4768 748 4808
rect 788 4768 789 4808
rect 747 4759 789 4768
rect 267 4304 309 4313
rect 267 4264 268 4304
rect 308 4264 309 4304
rect 267 4255 309 4264
rect 940 3977 980 6271
rect 939 3968 981 3977
rect 939 3928 940 3968
rect 980 3928 981 3968
rect 939 3919 981 3928
rect 171 3296 213 3305
rect 171 3256 172 3296
rect 212 3256 213 3296
rect 171 3247 213 3256
rect 1036 2540 1076 21559
rect 1324 21524 1364 21643
rect 1516 21642 1556 21727
rect 1324 21475 1364 21484
rect 1419 21524 1461 21533
rect 1419 21484 1420 21524
rect 1460 21484 1461 21524
rect 1419 21475 1461 21484
rect 1131 21440 1173 21449
rect 1131 21400 1132 21440
rect 1172 21400 1173 21440
rect 1131 21391 1173 21400
rect 1132 18257 1172 21391
rect 1323 20852 1365 20861
rect 1323 20812 1324 20852
rect 1364 20812 1365 20852
rect 1323 20803 1365 20812
rect 1324 20718 1364 20803
rect 1420 20096 1460 21475
rect 1515 21020 1557 21029
rect 1515 20980 1516 21020
rect 1556 20980 1557 21020
rect 1515 20971 1557 20980
rect 1516 20886 1556 20971
rect 1228 20056 1460 20096
rect 1516 20096 1556 20105
rect 1228 19760 1268 20056
rect 1324 19928 1364 19937
rect 1324 19844 1364 19888
rect 1419 19844 1461 19853
rect 1324 19804 1420 19844
rect 1460 19804 1461 19844
rect 1419 19795 1461 19804
rect 1516 19769 1556 20056
rect 1515 19760 1557 19769
rect 1228 19720 1364 19760
rect 1324 19676 1364 19720
rect 1515 19720 1516 19760
rect 1556 19720 1557 19760
rect 1515 19711 1557 19720
rect 1324 19636 1460 19676
rect 1323 19340 1365 19349
rect 1323 19300 1324 19340
rect 1364 19300 1365 19340
rect 1323 19291 1365 19300
rect 1324 19206 1364 19291
rect 1131 18248 1173 18257
rect 1131 18208 1132 18248
rect 1172 18208 1173 18248
rect 1131 18199 1173 18208
rect 1228 17744 1268 17753
rect 1420 17744 1460 19636
rect 1516 19340 1556 19349
rect 1516 19265 1556 19300
rect 1515 19256 1557 19265
rect 1515 19216 1516 19256
rect 1556 19216 1557 19256
rect 1515 19207 1557 19216
rect 1516 18668 1556 19207
rect 1612 18845 1652 22324
rect 1804 22324 1900 22364
rect 1708 21524 1748 21533
rect 1708 20609 1748 21484
rect 1707 20600 1749 20609
rect 1707 20560 1708 20600
rect 1748 20560 1749 20600
rect 1707 20551 1749 20560
rect 1708 20466 1748 20551
rect 1707 19508 1749 19517
rect 1707 19468 1708 19508
rect 1748 19468 1749 19508
rect 1707 19459 1749 19468
rect 1708 19374 1748 19459
rect 1804 19013 1844 22324
rect 1900 22315 1940 22324
rect 1899 21776 1941 21785
rect 1899 21736 1900 21776
rect 1940 21736 1941 21776
rect 1899 21727 1941 21736
rect 1900 21642 1940 21727
rect 1803 19004 1845 19013
rect 1803 18964 1804 19004
rect 1844 18964 1845 19004
rect 1803 18955 1845 18964
rect 1611 18836 1653 18845
rect 1611 18796 1612 18836
rect 1652 18796 1653 18836
rect 1611 18787 1653 18796
rect 1996 18668 2036 23080
rect 2092 21944 2132 23575
rect 2284 22364 2324 23752
rect 2380 23633 2420 26020
rect 2476 25649 2516 28120
rect 2475 25640 2517 25649
rect 2475 25600 2476 25640
rect 2516 25600 2517 25640
rect 2475 25591 2517 25600
rect 2475 25304 2517 25313
rect 2475 25264 2476 25304
rect 2516 25264 2517 25304
rect 2572 25304 2612 28876
rect 2668 28867 2708 28876
rect 2764 28841 2804 29800
rect 3052 30428 3092 30437
rect 2956 29672 2996 29681
rect 2859 29168 2901 29177
rect 2859 29128 2860 29168
rect 2900 29128 2901 29168
rect 2859 29119 2901 29128
rect 2860 29084 2900 29119
rect 2860 29033 2900 29044
rect 2763 28832 2805 28841
rect 2763 28792 2764 28832
rect 2804 28792 2805 28832
rect 2763 28783 2805 28792
rect 2956 28664 2996 29632
rect 3052 29504 3092 30388
rect 3148 30101 3188 31312
rect 3435 31352 3477 31361
rect 3435 31312 3436 31352
rect 3476 31312 3477 31352
rect 3435 31303 3477 31312
rect 3436 30680 3476 31303
rect 3340 30640 3436 30680
rect 3244 30428 3284 30437
rect 3147 30092 3189 30101
rect 3147 30052 3148 30092
rect 3188 30052 3189 30092
rect 3147 30043 3189 30052
rect 3244 29849 3284 30388
rect 3243 29840 3285 29849
rect 3243 29800 3244 29840
rect 3284 29800 3285 29840
rect 3243 29791 3285 29800
rect 3340 29840 3380 30640
rect 3436 30631 3476 30640
rect 3148 29672 3188 29681
rect 3188 29632 3284 29672
rect 3148 29623 3188 29632
rect 3052 29464 3188 29504
rect 3051 29000 3093 29009
rect 3051 28960 3052 29000
rect 3092 28960 3093 29000
rect 3051 28951 3093 28960
rect 3052 28866 3092 28951
rect 2956 28624 3092 28664
rect 2763 28496 2805 28505
rect 2763 28456 2764 28496
rect 2804 28456 2805 28496
rect 2763 28447 2805 28456
rect 2668 28160 2708 28169
rect 2668 25481 2708 28120
rect 2764 26657 2804 28447
rect 2857 28324 2897 28333
rect 2855 28284 2857 28324
rect 2855 28275 2897 28284
rect 2956 28328 2996 28339
rect 2855 28160 2895 28275
rect 2956 28253 2996 28288
rect 2955 28244 2997 28253
rect 2955 28204 2956 28244
rect 2996 28204 2997 28244
rect 2955 28195 2997 28204
rect 2855 28120 2900 28160
rect 2860 27404 2900 28120
rect 3052 28076 3092 28624
rect 3148 28505 3188 29464
rect 3244 29429 3284 29632
rect 3340 29513 3380 29800
rect 3532 29756 3572 32983
rect 3723 32864 3765 32873
rect 3723 32824 3724 32864
rect 3764 32824 3765 32864
rect 3723 32815 3765 32824
rect 3724 32730 3764 32815
rect 3915 32360 3957 32369
rect 3915 32320 3916 32360
rect 3956 32320 3957 32360
rect 3915 32311 3957 32320
rect 3916 32192 3956 32311
rect 3916 32143 3956 32152
rect 4108 32117 4148 33412
rect 4204 32878 4244 34159
rect 4204 32829 4244 32838
rect 4203 32696 4245 32705
rect 4203 32656 4204 32696
rect 4244 32656 4245 32696
rect 4203 32647 4245 32656
rect 4107 32108 4149 32117
rect 4107 32068 4108 32108
rect 4148 32068 4149 32108
rect 4107 32059 4149 32068
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 4204 31352 4244 32647
rect 4108 31312 4244 31352
rect 4108 30437 4148 31312
rect 4203 31184 4245 31193
rect 4203 31144 4204 31184
rect 4244 31144 4245 31184
rect 4203 31135 4245 31144
rect 4107 30428 4149 30437
rect 4107 30388 4108 30428
rect 4148 30388 4149 30428
rect 4107 30379 4149 30388
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3627 30092 3669 30101
rect 3627 30052 3628 30092
rect 3668 30052 3669 30092
rect 3627 30043 3669 30052
rect 3436 29716 3572 29756
rect 3339 29504 3381 29513
rect 3339 29464 3340 29504
rect 3380 29464 3381 29504
rect 3339 29455 3381 29464
rect 3243 29420 3285 29429
rect 3243 29380 3244 29420
rect 3284 29380 3285 29420
rect 3243 29371 3285 29380
rect 3243 29252 3285 29261
rect 3243 29212 3244 29252
rect 3284 29212 3285 29252
rect 3243 29203 3285 29212
rect 3244 29168 3284 29203
rect 3244 29117 3284 29128
rect 3243 29000 3285 29009
rect 3243 28960 3244 29000
rect 3284 28960 3285 29000
rect 3243 28951 3285 28960
rect 3147 28496 3189 28505
rect 3147 28456 3148 28496
rect 3188 28456 3189 28496
rect 3147 28447 3189 28456
rect 3147 28328 3189 28337
rect 3147 28288 3148 28328
rect 3188 28288 3189 28328
rect 3147 28279 3189 28288
rect 3244 28328 3284 28951
rect 3345 28328 3385 28337
rect 3436 28328 3476 29716
rect 3531 29420 3573 29429
rect 3531 29380 3532 29420
rect 3572 29380 3573 29420
rect 3531 29371 3573 29380
rect 3244 28279 3284 28288
rect 3340 28288 3345 28328
rect 3385 28288 3476 28328
rect 3340 28279 3385 28288
rect 3148 28194 3188 28279
rect 3244 28160 3284 28171
rect 3244 28085 3284 28120
rect 3243 28076 3285 28085
rect 3052 28036 3188 28076
rect 3051 27908 3093 27917
rect 3051 27868 3052 27908
rect 3092 27868 3093 27908
rect 3051 27859 3093 27868
rect 3052 27656 3092 27859
rect 2860 27364 2996 27404
rect 2860 26816 2900 26856
rect 2860 26741 2900 26776
rect 2859 26732 2901 26741
rect 2859 26692 2860 26732
rect 2900 26692 2901 26732
rect 2859 26683 2901 26692
rect 2763 26648 2805 26657
rect 2763 26608 2764 26648
rect 2804 26608 2805 26648
rect 2763 26599 2805 26608
rect 2860 26144 2900 26683
rect 2956 26321 2996 27364
rect 2955 26312 2997 26321
rect 2955 26272 2956 26312
rect 2996 26272 2997 26312
rect 2955 26263 2997 26272
rect 2860 26095 2900 26104
rect 3052 25817 3092 27616
rect 3148 26321 3188 28036
rect 3243 28036 3244 28076
rect 3284 28036 3285 28076
rect 3243 28027 3285 28036
rect 3244 27404 3284 27413
rect 3147 26312 3189 26321
rect 3147 26272 3148 26312
rect 3188 26272 3189 26312
rect 3147 26263 3189 26272
rect 3051 25808 3093 25817
rect 3051 25768 3052 25808
rect 3092 25768 3093 25808
rect 3051 25759 3093 25768
rect 2859 25556 2901 25565
rect 2859 25516 2860 25556
rect 2900 25516 2901 25556
rect 2859 25507 2901 25516
rect 2667 25472 2709 25481
rect 2667 25432 2668 25472
rect 2708 25432 2709 25472
rect 2667 25423 2709 25432
rect 2860 25422 2900 25507
rect 3052 25388 3092 25397
rect 2572 25264 2900 25304
rect 2475 25255 2517 25264
rect 2476 24632 2516 25255
rect 2668 25136 2708 25145
rect 2708 25096 2804 25136
rect 2668 25087 2708 25096
rect 2379 23624 2421 23633
rect 2379 23584 2380 23624
rect 2420 23584 2421 23624
rect 2379 23575 2421 23584
rect 2476 23213 2516 24592
rect 2668 24380 2708 24389
rect 2572 24340 2668 24380
rect 2475 23204 2517 23213
rect 2475 23164 2476 23204
rect 2516 23164 2517 23204
rect 2475 23155 2517 23164
rect 2380 22373 2420 22417
rect 2379 22364 2421 22373
rect 2284 22324 2380 22364
rect 2420 22324 2421 22364
rect 2379 22322 2421 22324
rect 2379 22315 2380 22322
rect 2420 22315 2421 22322
rect 2380 22273 2420 22282
rect 2187 22196 2229 22205
rect 2187 22156 2188 22196
rect 2228 22156 2229 22196
rect 2187 22147 2229 22156
rect 2188 22062 2228 22147
rect 2283 22028 2325 22037
rect 2283 21988 2284 22028
rect 2324 21988 2325 22028
rect 2283 21979 2325 21988
rect 2092 21904 2228 21944
rect 2091 21524 2133 21533
rect 2091 21484 2092 21524
rect 2132 21484 2133 21524
rect 2091 21475 2133 21484
rect 2092 21390 2132 21475
rect 1516 18628 1652 18668
rect 1515 18416 1557 18425
rect 1515 18376 1516 18416
rect 1556 18376 1557 18416
rect 1515 18367 1557 18376
rect 1516 18282 1556 18367
rect 1268 17704 1460 17744
rect 1228 16904 1268 17704
rect 1612 17669 1652 18628
rect 1708 18628 2036 18668
rect 1611 17660 1653 17669
rect 1611 17620 1612 17660
rect 1652 17620 1653 17660
rect 1611 17611 1653 17620
rect 1324 17081 1364 17166
rect 1419 17156 1461 17165
rect 1419 17116 1420 17156
rect 1460 17116 1461 17156
rect 1419 17107 1461 17116
rect 1323 17072 1365 17081
rect 1323 17032 1324 17072
rect 1364 17032 1365 17072
rect 1323 17023 1365 17032
rect 1420 17022 1460 17107
rect 1516 17072 1556 17081
rect 1228 16864 1364 16904
rect 1324 16493 1364 16864
rect 1323 16484 1365 16493
rect 1323 16444 1324 16484
rect 1364 16444 1365 16484
rect 1323 16435 1365 16444
rect 1516 16409 1556 17032
rect 1611 17072 1653 17081
rect 1611 17032 1612 17072
rect 1652 17032 1653 17072
rect 1611 17023 1653 17032
rect 1612 16938 1652 17023
rect 1708 16577 1748 18628
rect 2092 18584 2132 18593
rect 1804 18509 1844 18540
rect 1803 18500 1845 18509
rect 1803 18460 1804 18500
rect 1844 18460 1845 18500
rect 1803 18451 1845 18460
rect 1804 18416 1844 18451
rect 1804 17753 1844 18376
rect 1996 18332 2036 18341
rect 1803 17744 1845 17753
rect 1803 17704 1804 17744
rect 1844 17704 1845 17744
rect 1803 17695 1845 17704
rect 1996 17249 2036 18292
rect 2092 17333 2132 18544
rect 2188 17417 2228 21904
rect 2284 21776 2324 21979
rect 2284 21727 2324 21736
rect 2572 21608 2612 24340
rect 2668 24331 2708 24340
rect 2764 21701 2804 25096
rect 2860 23801 2900 25264
rect 3052 24809 3092 25348
rect 3244 25313 3284 27364
rect 3340 27077 3380 28279
rect 3435 27488 3477 27497
rect 3435 27448 3436 27488
rect 3476 27448 3477 27488
rect 3435 27439 3477 27448
rect 3436 27354 3476 27439
rect 3339 27068 3381 27077
rect 3339 27028 3340 27068
rect 3380 27028 3381 27068
rect 3339 27019 3381 27028
rect 3388 26830 3428 26834
rect 3532 26830 3572 29371
rect 3628 28925 3668 30043
rect 3915 29840 3957 29849
rect 3915 29800 3916 29840
rect 3956 29800 3957 29840
rect 3915 29791 3957 29800
rect 3916 29000 3956 29791
rect 4204 29000 4244 31135
rect 4300 29681 4340 37444
rect 4396 36728 4436 38191
rect 4492 37820 4532 40216
rect 4724 40216 4820 40256
rect 4684 40207 4724 40216
rect 4588 39500 4628 39509
rect 4628 39460 4724 39500
rect 4588 39451 4628 39460
rect 4587 38744 4629 38753
rect 4587 38704 4588 38744
rect 4628 38704 4629 38744
rect 4587 38695 4629 38704
rect 4588 38610 4628 38695
rect 4587 38156 4629 38165
rect 4587 38116 4588 38156
rect 4628 38116 4629 38156
rect 4587 38107 4629 38116
rect 4588 38022 4628 38107
rect 4684 37988 4724 39460
rect 4780 38996 4820 40216
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 4875 39836 4917 39845
rect 5356 39836 5396 40963
rect 5452 39845 5492 40972
rect 4875 39796 4876 39836
rect 4916 39796 4917 39836
rect 4875 39787 4917 39796
rect 5164 39796 5396 39836
rect 5451 39836 5493 39845
rect 5451 39796 5452 39836
rect 5492 39796 5493 39836
rect 4876 39752 4916 39787
rect 4876 39701 4916 39712
rect 4972 39752 5012 39761
rect 4972 39509 5012 39712
rect 5067 39668 5109 39677
rect 5067 39628 5068 39668
rect 5108 39628 5109 39668
rect 5067 39619 5109 39628
rect 4971 39500 5013 39509
rect 4971 39460 4972 39500
rect 5012 39460 5013 39500
rect 4971 39451 5013 39460
rect 5068 39173 5108 39619
rect 5067 39164 5109 39173
rect 5067 39124 5068 39164
rect 5108 39124 5109 39164
rect 5067 39115 5109 39124
rect 4971 39080 5013 39089
rect 4971 39040 4972 39080
rect 5012 39040 5013 39080
rect 4971 39031 5013 39040
rect 4780 38249 4820 38956
rect 4972 38946 5012 39031
rect 5164 38744 5204 39796
rect 5451 39787 5493 39796
rect 5355 39668 5397 39677
rect 5355 39628 5356 39668
rect 5396 39628 5397 39668
rect 5355 39619 5397 39628
rect 5452 39668 5492 39679
rect 5356 39534 5396 39619
rect 5452 39593 5492 39628
rect 5451 39584 5493 39593
rect 5451 39544 5452 39584
rect 5492 39544 5493 39584
rect 5451 39535 5493 39544
rect 5548 39089 5588 41140
rect 5644 40853 5684 41224
rect 5643 40844 5685 40853
rect 5643 40804 5644 40844
rect 5684 40804 5685 40844
rect 5643 40795 5685 40804
rect 5644 40097 5684 40795
rect 5643 40088 5685 40097
rect 5643 40048 5644 40088
rect 5684 40048 5685 40088
rect 5643 40039 5685 40048
rect 5547 39080 5589 39089
rect 5547 39040 5548 39080
rect 5588 39040 5589 39080
rect 5547 39031 5589 39040
rect 5260 38921 5300 39006
rect 5259 38912 5301 38921
rect 5259 38872 5260 38912
rect 5300 38872 5301 38912
rect 5259 38863 5301 38872
rect 5643 38912 5685 38921
rect 5643 38872 5644 38912
rect 5684 38872 5685 38912
rect 5643 38863 5685 38872
rect 5164 38704 5396 38744
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5356 38408 5396 38704
rect 5547 38660 5589 38669
rect 5547 38620 5548 38660
rect 5588 38620 5589 38660
rect 5547 38611 5589 38620
rect 5260 38368 5396 38408
rect 5067 38324 5109 38333
rect 5067 38284 5068 38324
rect 5108 38284 5109 38324
rect 5067 38275 5109 38284
rect 4779 38240 4821 38249
rect 4779 38200 4780 38240
rect 4820 38200 4821 38240
rect 4779 38191 4821 38200
rect 4780 38106 4820 38191
rect 5068 38190 5108 38275
rect 5260 38235 5300 38368
rect 5260 38186 5300 38195
rect 4684 37948 4916 37988
rect 4492 37780 4724 37820
rect 4684 37400 4724 37780
rect 4780 37577 4820 37662
rect 4876 37661 4916 37948
rect 4875 37652 4917 37661
rect 4875 37612 4876 37652
rect 4916 37612 4917 37652
rect 4875 37603 4917 37612
rect 4779 37568 4821 37577
rect 4779 37528 4780 37568
rect 4820 37528 4821 37568
rect 4779 37519 4821 37528
rect 4971 37484 5013 37493
rect 4971 37444 4972 37484
rect 5012 37444 5013 37484
rect 4971 37435 5013 37444
rect 4684 37360 4820 37400
rect 4491 37232 4533 37241
rect 4491 37192 4492 37232
rect 4532 37192 4533 37232
rect 4491 37183 4533 37192
rect 4492 37098 4532 37183
rect 4683 37064 4725 37073
rect 4683 37024 4684 37064
rect 4724 37024 4725 37064
rect 4683 37015 4725 37024
rect 4587 36812 4629 36821
rect 4587 36772 4588 36812
rect 4628 36772 4629 36812
rect 4587 36763 4629 36772
rect 4492 36728 4532 36737
rect 4396 36688 4492 36728
rect 4492 36569 4532 36688
rect 4491 36560 4533 36569
rect 4491 36520 4492 36560
rect 4532 36520 4533 36560
rect 4491 36511 4533 36520
rect 4395 35888 4437 35897
rect 4395 35848 4396 35888
rect 4436 35848 4437 35888
rect 4395 35839 4437 35848
rect 4492 35888 4532 35897
rect 4396 35754 4436 35839
rect 4492 35729 4532 35848
rect 4588 35813 4628 36763
rect 4587 35804 4629 35813
rect 4587 35764 4588 35804
rect 4628 35764 4629 35804
rect 4587 35755 4629 35764
rect 4491 35720 4533 35729
rect 4491 35680 4492 35720
rect 4532 35680 4533 35720
rect 4491 35671 4533 35680
rect 4587 35552 4629 35561
rect 4587 35512 4588 35552
rect 4628 35512 4629 35552
rect 4587 35503 4629 35512
rect 4491 35216 4533 35225
rect 4491 35176 4492 35216
rect 4532 35176 4533 35216
rect 4491 35167 4533 35176
rect 4395 34628 4437 34637
rect 4395 34588 4396 34628
rect 4436 34588 4437 34628
rect 4395 34579 4437 34588
rect 4396 33872 4436 34579
rect 4396 33823 4436 33832
rect 4395 32780 4437 32789
rect 4395 32740 4396 32780
rect 4436 32740 4437 32780
rect 4395 32731 4437 32740
rect 4396 32646 4436 32731
rect 4492 32621 4532 35167
rect 4491 32612 4533 32621
rect 4491 32572 4492 32612
rect 4532 32572 4533 32612
rect 4491 32563 4533 32572
rect 4396 32108 4436 32117
rect 4396 31865 4436 32068
rect 4491 32108 4533 32117
rect 4491 32068 4492 32108
rect 4532 32068 4533 32108
rect 4491 32059 4533 32068
rect 4492 31974 4532 32059
rect 4395 31856 4437 31865
rect 4395 31816 4396 31856
rect 4436 31816 4437 31856
rect 4395 31807 4437 31816
rect 4588 31772 4628 35503
rect 4684 34796 4724 37015
rect 4780 36896 4820 37360
rect 4972 37350 5012 37435
rect 5356 37400 5396 37409
rect 5548 37400 5588 38611
rect 5644 37409 5684 38863
rect 5740 38240 5780 42475
rect 5836 41693 5876 42928
rect 5835 41684 5877 41693
rect 5835 41644 5836 41684
rect 5876 41644 5877 41684
rect 5835 41635 5877 41644
rect 6028 40517 6068 42928
rect 6027 40508 6069 40517
rect 6027 40468 6028 40508
rect 6068 40468 6069 40508
rect 6027 40459 6069 40468
rect 6124 40424 6164 40433
rect 6124 40340 6164 40384
rect 6028 40300 6164 40340
rect 5931 40172 5973 40181
rect 5931 40132 5932 40172
rect 5972 40132 5973 40172
rect 5931 40123 5973 40132
rect 5932 39752 5972 40123
rect 6028 40097 6068 40300
rect 6220 40256 6260 42928
rect 6412 41357 6452 42928
rect 6604 41609 6644 42928
rect 6796 42029 6836 42928
rect 6795 42020 6837 42029
rect 6795 41980 6796 42020
rect 6836 41980 6837 42020
rect 6795 41971 6837 41980
rect 6603 41600 6645 41609
rect 6603 41560 6604 41600
rect 6644 41560 6645 41600
rect 6603 41551 6645 41560
rect 6795 41600 6837 41609
rect 6795 41560 6796 41600
rect 6836 41560 6837 41600
rect 6795 41551 6837 41560
rect 6411 41348 6453 41357
rect 6411 41308 6412 41348
rect 6452 41308 6453 41348
rect 6411 41299 6453 41308
rect 6411 41096 6453 41105
rect 6411 41056 6412 41096
rect 6452 41056 6453 41096
rect 6411 41047 6453 41056
rect 6124 40216 6260 40256
rect 6316 40256 6356 40265
rect 6027 40088 6069 40097
rect 6027 40048 6028 40088
rect 6068 40048 6069 40088
rect 6027 40039 6069 40048
rect 5932 39703 5972 39712
rect 5835 39164 5877 39173
rect 5835 39124 5836 39164
rect 5876 39124 5877 39164
rect 5835 39115 5877 39124
rect 5740 38191 5780 38200
rect 5739 37736 5781 37745
rect 5739 37696 5740 37736
rect 5780 37696 5781 37736
rect 5739 37687 5781 37696
rect 5396 37360 5588 37400
rect 5643 37400 5685 37409
rect 5643 37360 5644 37400
rect 5684 37360 5685 37400
rect 5164 37241 5204 37326
rect 5163 37232 5205 37241
rect 5163 37192 5164 37232
rect 5204 37192 5205 37232
rect 5163 37183 5205 37192
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4780 36856 5012 36896
rect 4972 36723 5012 36856
rect 5163 36812 5205 36821
rect 5163 36772 5164 36812
rect 5204 36772 5205 36812
rect 5163 36763 5205 36772
rect 4972 36674 5012 36683
rect 5164 36678 5204 36763
rect 5356 36233 5396 37360
rect 5643 37351 5685 37360
rect 5740 36896 5780 37687
rect 5740 36847 5780 36856
rect 5643 36812 5685 36821
rect 5643 36772 5644 36812
rect 5684 36772 5685 36812
rect 5643 36763 5685 36772
rect 5548 36653 5588 36738
rect 5547 36644 5589 36653
rect 5547 36604 5548 36644
rect 5588 36604 5589 36644
rect 5547 36595 5589 36604
rect 5547 36392 5589 36401
rect 5547 36352 5548 36392
rect 5588 36352 5589 36392
rect 5547 36343 5589 36352
rect 5355 36224 5397 36233
rect 5355 36184 5356 36224
rect 5396 36184 5397 36224
rect 5355 36175 5397 36184
rect 5164 36016 5492 36056
rect 5067 35888 5109 35897
rect 5067 35848 5068 35888
rect 5108 35848 5109 35888
rect 5067 35839 5109 35848
rect 5068 35754 5108 35839
rect 5164 35804 5204 36016
rect 5259 35888 5301 35897
rect 5259 35848 5260 35888
rect 5300 35848 5301 35888
rect 5259 35839 5301 35848
rect 5356 35888 5396 35897
rect 5164 35755 5204 35764
rect 5260 35754 5300 35839
rect 4780 35720 4820 35729
rect 4780 35309 4820 35680
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4779 35300 4821 35309
rect 4779 35260 4780 35300
rect 4820 35260 4821 35300
rect 4779 35251 4821 35260
rect 5163 35132 5205 35141
rect 5163 35092 5164 35132
rect 5204 35092 5205 35132
rect 5163 35083 5205 35092
rect 4684 34756 4916 34796
rect 4683 34628 4725 34637
rect 4683 34588 4684 34628
rect 4724 34588 4725 34628
rect 4683 34579 4725 34588
rect 4684 34460 4724 34579
rect 4684 34411 4724 34420
rect 4780 34385 4820 34470
rect 4779 34376 4821 34385
rect 4779 34336 4780 34376
rect 4820 34336 4821 34376
rect 4779 34327 4821 34336
rect 4876 34208 4916 34756
rect 5164 34376 5204 35083
rect 5259 34544 5301 34553
rect 5259 34504 5260 34544
rect 5300 34504 5301 34544
rect 5259 34495 5301 34504
rect 5164 34327 5204 34336
rect 5260 34376 5300 34495
rect 5260 34327 5300 34336
rect 4780 34168 4916 34208
rect 4683 33872 4725 33881
rect 4683 33832 4684 33872
rect 4724 33832 4725 33872
rect 4780 33872 4820 34168
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4780 33832 5012 33872
rect 4683 33823 4725 33832
rect 4684 33738 4724 33823
rect 4779 33704 4821 33713
rect 4779 33664 4780 33704
rect 4820 33664 4821 33704
rect 4779 33655 4821 33664
rect 4876 33704 4916 33715
rect 4683 33032 4725 33041
rect 4683 32992 4684 33032
rect 4724 32992 4725 33032
rect 4683 32983 4725 32992
rect 4684 32898 4724 32983
rect 4492 31732 4628 31772
rect 4396 31352 4436 31361
rect 4396 30941 4436 31312
rect 4395 30932 4437 30941
rect 4395 30892 4396 30932
rect 4436 30892 4437 30932
rect 4395 30883 4437 30892
rect 4492 30269 4532 31732
rect 4587 31604 4629 31613
rect 4587 31564 4588 31604
rect 4628 31564 4629 31604
rect 4587 31555 4629 31564
rect 4780 31604 4820 33655
rect 4876 33629 4916 33664
rect 4875 33620 4917 33629
rect 4875 33580 4876 33620
rect 4916 33580 4917 33620
rect 4875 33571 4917 33580
rect 4876 32864 4916 32873
rect 4972 32864 5012 33832
rect 4916 32824 5012 32864
rect 4876 32705 4916 32824
rect 4875 32696 4917 32705
rect 4875 32656 4876 32696
rect 4916 32656 4917 32696
rect 4875 32647 4917 32656
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 5356 32444 5396 35848
rect 5452 35384 5492 36016
rect 5548 35888 5588 36343
rect 5548 35645 5588 35848
rect 5547 35636 5589 35645
rect 5547 35596 5548 35636
rect 5588 35596 5589 35636
rect 5547 35587 5589 35596
rect 5452 35344 5588 35384
rect 5451 35216 5493 35225
rect 5451 35176 5452 35216
rect 5492 35176 5493 35216
rect 5451 35167 5493 35176
rect 5452 34889 5492 35167
rect 5451 34880 5493 34889
rect 5451 34840 5452 34880
rect 5492 34840 5493 34880
rect 5451 34831 5493 34840
rect 5451 34628 5493 34637
rect 5451 34588 5452 34628
rect 5492 34588 5493 34628
rect 5451 34579 5493 34588
rect 5452 34133 5492 34579
rect 5451 34124 5493 34133
rect 5451 34084 5452 34124
rect 5492 34084 5493 34124
rect 5451 34075 5493 34084
rect 5548 33209 5588 35344
rect 5644 35309 5684 36763
rect 5836 36728 5876 39115
rect 6027 38324 6069 38333
rect 6027 38284 6028 38324
rect 6068 38284 6069 38324
rect 6027 38275 6069 38284
rect 5932 36728 5972 36737
rect 5836 36688 5932 36728
rect 5932 36679 5972 36688
rect 6028 36485 6068 38275
rect 6027 36476 6069 36485
rect 6027 36436 6028 36476
rect 6068 36436 6069 36476
rect 6027 36427 6069 36436
rect 6027 35636 6069 35645
rect 6027 35596 6028 35636
rect 6068 35596 6069 35636
rect 6027 35587 6069 35596
rect 5835 35468 5877 35477
rect 5835 35428 5836 35468
rect 5876 35428 5877 35468
rect 5835 35419 5877 35428
rect 5836 35309 5876 35419
rect 6028 35309 6068 35587
rect 6124 35393 6164 40216
rect 6316 39089 6356 40216
rect 6412 39747 6452 41047
rect 6699 40676 6741 40685
rect 6699 40636 6700 40676
rect 6740 40636 6741 40676
rect 6699 40627 6741 40636
rect 6700 40542 6740 40627
rect 6507 40508 6549 40517
rect 6507 40468 6508 40508
rect 6548 40468 6549 40508
rect 6507 40459 6549 40468
rect 6508 40374 6548 40459
rect 6412 39698 6452 39707
rect 6604 39836 6644 39845
rect 6604 39584 6644 39796
rect 6412 39544 6644 39584
rect 6315 39080 6357 39089
rect 6315 39040 6316 39080
rect 6356 39040 6357 39080
rect 6315 39031 6357 39040
rect 6220 38156 6260 38167
rect 6220 38081 6260 38116
rect 6315 38156 6357 38165
rect 6315 38116 6316 38156
rect 6356 38116 6357 38156
rect 6315 38107 6357 38116
rect 6219 38072 6261 38081
rect 6219 38032 6220 38072
rect 6260 38032 6261 38072
rect 6219 38023 6261 38032
rect 6316 38022 6356 38107
rect 6219 35888 6261 35897
rect 6219 35848 6220 35888
rect 6260 35848 6261 35888
rect 6219 35839 6261 35848
rect 6123 35384 6165 35393
rect 6123 35344 6124 35384
rect 6164 35344 6165 35384
rect 6123 35335 6165 35344
rect 5643 35300 5685 35309
rect 5643 35260 5644 35300
rect 5684 35260 5685 35300
rect 5643 35251 5685 35260
rect 5835 35300 5877 35309
rect 5835 35260 5836 35300
rect 5876 35260 5877 35300
rect 5835 35251 5877 35260
rect 6027 35300 6069 35309
rect 6027 35260 6028 35300
rect 6068 35260 6069 35300
rect 6027 35251 6069 35260
rect 5931 35216 5973 35225
rect 5931 35176 5932 35216
rect 5972 35176 5973 35216
rect 5931 35167 5973 35176
rect 6028 35216 6068 35251
rect 6028 35167 6068 35176
rect 5739 35132 5781 35141
rect 5644 35092 5740 35132
rect 5780 35092 5781 35132
rect 5644 35048 5684 35092
rect 5739 35083 5781 35092
rect 5932 35082 5972 35167
rect 5644 34999 5684 35008
rect 5835 35048 5877 35057
rect 5835 35008 5836 35048
rect 5876 35008 5877 35048
rect 5835 34999 5877 35008
rect 6123 35048 6165 35057
rect 6123 35008 6124 35048
rect 6164 35008 6165 35048
rect 6123 34999 6165 35008
rect 5740 34376 5780 34385
rect 5740 34133 5780 34336
rect 5739 34124 5781 34133
rect 5739 34084 5740 34124
rect 5780 34084 5781 34124
rect 5739 34075 5781 34084
rect 5643 34040 5685 34049
rect 5643 34000 5644 34040
rect 5684 34000 5685 34040
rect 5643 33991 5685 34000
rect 5547 33200 5589 33209
rect 5547 33160 5548 33200
rect 5588 33160 5589 33200
rect 5547 33151 5589 33160
rect 5356 32404 5588 32444
rect 5451 32276 5493 32285
rect 5451 32236 5452 32276
rect 5492 32236 5493 32276
rect 5451 32227 5493 32236
rect 4876 32192 4916 32201
rect 4876 31781 4916 32152
rect 4971 32192 5013 32201
rect 4971 32152 4972 32192
rect 5012 32152 5013 32192
rect 4971 32143 5013 32152
rect 5259 32192 5301 32201
rect 5259 32152 5260 32192
rect 5300 32152 5301 32192
rect 5259 32143 5301 32152
rect 4972 32058 5012 32143
rect 5260 32058 5300 32143
rect 5355 31940 5397 31949
rect 5355 31900 5356 31940
rect 5396 31900 5397 31940
rect 5355 31891 5397 31900
rect 4875 31772 4917 31781
rect 4875 31732 4876 31772
rect 4916 31732 4917 31772
rect 4875 31723 4917 31732
rect 4780 31555 4820 31564
rect 4588 31470 4628 31555
rect 4683 31520 4725 31529
rect 4683 31480 4684 31520
rect 4724 31480 4725 31520
rect 4683 31471 4725 31480
rect 4588 31184 4628 31193
rect 4588 30428 4628 31144
rect 4684 30848 4724 31471
rect 4971 31352 5013 31361
rect 4971 31312 4972 31352
rect 5012 31312 5013 31352
rect 4971 31303 5013 31312
rect 4972 31218 5012 31303
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4876 30848 4916 30857
rect 4684 30808 4876 30848
rect 4876 30799 4916 30808
rect 4683 30680 4725 30689
rect 4683 30640 4684 30680
rect 4724 30640 4725 30680
rect 4683 30631 4725 30640
rect 5356 30680 5396 31891
rect 5356 30631 5396 30640
rect 4684 30546 4724 30631
rect 5068 30596 5108 30605
rect 4588 30388 4724 30428
rect 4491 30260 4533 30269
rect 4491 30220 4492 30260
rect 4532 30220 4533 30260
rect 4491 30211 4533 30220
rect 4587 29840 4629 29849
rect 4587 29800 4588 29840
rect 4628 29800 4629 29840
rect 4587 29791 4629 29800
rect 4588 29706 4628 29791
rect 4299 29672 4341 29681
rect 4299 29632 4300 29672
rect 4340 29632 4341 29672
rect 4299 29623 4341 29632
rect 4491 29672 4533 29681
rect 4491 29632 4492 29672
rect 4532 29632 4533 29672
rect 4491 29623 4533 29632
rect 4492 29513 4532 29623
rect 4684 29588 4724 30388
rect 5068 30353 5108 30556
rect 5067 30344 5109 30353
rect 5067 30304 5068 30344
rect 5108 30304 5109 30344
rect 5067 30295 5109 30304
rect 5068 29840 5108 29849
rect 5068 29681 5108 29800
rect 4876 29672 4916 29681
rect 4588 29548 4724 29588
rect 4780 29632 4876 29672
rect 4491 29504 4533 29513
rect 4491 29464 4492 29504
rect 4532 29464 4533 29504
rect 4491 29455 4533 29464
rect 4492 29177 4532 29455
rect 4491 29168 4533 29177
rect 4491 29128 4492 29168
rect 4532 29128 4533 29168
rect 4491 29119 4533 29128
rect 4492 29034 4532 29119
rect 3916 28960 4148 29000
rect 4204 28960 4340 29000
rect 3627 28916 3669 28925
rect 3627 28876 3628 28916
rect 3668 28876 3669 28916
rect 3627 28867 3669 28876
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3723 28580 3765 28589
rect 3723 28540 3724 28580
rect 3764 28540 3765 28580
rect 3723 28531 3765 28540
rect 3627 28412 3669 28421
rect 3627 28372 3628 28412
rect 3668 28372 3669 28412
rect 3627 28363 3669 28372
rect 3628 28278 3668 28363
rect 3724 28085 3764 28531
rect 3819 28496 3861 28505
rect 3819 28456 3820 28496
rect 3860 28456 3861 28496
rect 3819 28447 3861 28456
rect 3820 28362 3860 28447
rect 4011 28412 4053 28421
rect 4011 28372 4012 28412
rect 4052 28372 4053 28412
rect 4011 28363 4053 28372
rect 4012 28278 4052 28363
rect 3723 28076 3765 28085
rect 3723 28036 3724 28076
rect 3764 28036 3765 28076
rect 3723 28027 3765 28036
rect 4108 27992 4148 28960
rect 4203 28580 4245 28589
rect 4203 28540 4204 28580
rect 4244 28540 4245 28580
rect 4203 28531 4245 28540
rect 4204 28446 4244 28531
rect 4300 28496 4340 28960
rect 4491 28748 4533 28757
rect 4491 28708 4492 28748
rect 4532 28708 4533 28748
rect 4491 28699 4533 28708
rect 4300 28456 4436 28496
rect 3820 27952 4148 27992
rect 3820 27656 3860 27952
rect 3820 27607 3860 27616
rect 3916 27656 3956 27665
rect 3916 27497 3956 27616
rect 4300 27581 4340 27666
rect 4299 27572 4341 27581
rect 4299 27532 4300 27572
rect 4340 27532 4341 27572
rect 4299 27523 4341 27532
rect 4396 27572 4436 28456
rect 4492 27908 4532 28699
rect 4588 28664 4628 29548
rect 4683 28916 4725 28925
rect 4683 28876 4684 28916
rect 4724 28876 4725 28916
rect 4683 28867 4725 28876
rect 4684 28782 4724 28867
rect 4588 28624 4724 28664
rect 4588 28412 4628 28423
rect 4588 28337 4628 28372
rect 4587 28328 4629 28337
rect 4587 28288 4588 28328
rect 4628 28288 4629 28328
rect 4587 28279 4629 28288
rect 4492 27868 4628 27908
rect 4491 27740 4533 27749
rect 4491 27700 4492 27740
rect 4532 27700 4533 27740
rect 4491 27691 4533 27700
rect 3915 27488 3957 27497
rect 3915 27448 3916 27488
rect 3956 27448 3957 27488
rect 3915 27439 3957 27448
rect 4107 27404 4149 27413
rect 4107 27364 4108 27404
rect 4148 27364 4149 27404
rect 4107 27355 4149 27364
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 4011 27068 4053 27077
rect 4011 27028 4012 27068
rect 4052 27028 4053 27068
rect 4011 27019 4053 27028
rect 3627 26984 3669 26993
rect 3627 26944 3628 26984
rect 3668 26944 3669 26984
rect 3627 26935 3669 26944
rect 3388 26825 3572 26830
rect 3428 26790 3572 26825
rect 3388 26776 3428 26785
rect 3531 26732 3573 26741
rect 3531 26692 3532 26732
rect 3572 26692 3573 26732
rect 3531 26683 3573 26692
rect 3339 26648 3381 26657
rect 3339 26608 3340 26648
rect 3380 26608 3381 26648
rect 3339 26599 3381 26608
rect 3340 26139 3380 26599
rect 3532 26598 3572 26683
rect 3628 26657 3668 26935
rect 4012 26816 4052 27019
rect 4012 26767 4052 26776
rect 4108 26816 4148 27355
rect 4299 27320 4341 27329
rect 4299 27280 4300 27320
rect 4340 27280 4341 27320
rect 4299 27271 4341 27280
rect 3627 26648 3669 26657
rect 3627 26608 3628 26648
rect 3668 26608 3669 26648
rect 3627 26599 3669 26608
rect 3820 26648 3860 26657
rect 3820 26489 3860 26608
rect 4108 26573 4148 26776
rect 4203 26816 4245 26825
rect 4203 26776 4204 26816
rect 4244 26776 4245 26816
rect 4203 26767 4245 26776
rect 4300 26816 4340 27271
rect 4300 26767 4340 26776
rect 4204 26682 4244 26767
rect 4107 26564 4149 26573
rect 4107 26524 4108 26564
rect 4148 26524 4149 26564
rect 4107 26515 4149 26524
rect 4396 26489 4436 27532
rect 3819 26480 3861 26489
rect 3819 26440 3820 26480
rect 3860 26440 3861 26480
rect 3819 26431 3861 26440
rect 4395 26480 4437 26489
rect 4395 26440 4396 26480
rect 4436 26440 4437 26480
rect 4395 26431 4437 26440
rect 3340 26090 3380 26099
rect 3532 26228 3572 26237
rect 3532 25472 3572 26188
rect 3820 25976 3860 26431
rect 4492 26312 4532 27691
rect 4492 26263 4532 26272
rect 4204 26069 4244 26154
rect 4203 26060 4245 26069
rect 4203 26020 4204 26060
rect 4244 26020 4245 26060
rect 4203 26011 4245 26020
rect 3820 25901 3860 25936
rect 3819 25892 3861 25901
rect 3819 25852 3820 25892
rect 3860 25852 3861 25892
rect 3819 25843 3861 25852
rect 4012 25892 4052 25901
rect 4052 25852 4244 25892
rect 4012 25843 4052 25852
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 4107 25556 4149 25565
rect 4107 25516 4108 25556
rect 4148 25516 4149 25556
rect 4107 25507 4149 25516
rect 3532 25432 3764 25472
rect 3628 25313 3668 25318
rect 3243 25304 3285 25313
rect 3243 25264 3244 25304
rect 3284 25264 3285 25304
rect 3243 25255 3285 25264
rect 3627 25309 3669 25313
rect 3627 25264 3628 25309
rect 3668 25264 3669 25309
rect 3627 25255 3669 25264
rect 3435 25220 3477 25229
rect 3435 25180 3436 25220
rect 3476 25180 3477 25220
rect 3435 25171 3477 25180
rect 3628 25174 3668 25255
rect 3436 25086 3476 25171
rect 3147 25052 3189 25061
rect 3147 25012 3148 25052
rect 3188 25012 3189 25052
rect 3147 25003 3189 25012
rect 3051 24800 3093 24809
rect 3051 24760 3052 24800
rect 3092 24760 3093 24800
rect 3051 24751 3093 24760
rect 3052 24632 3092 24643
rect 3052 24557 3092 24592
rect 3051 24548 3093 24557
rect 3051 24508 3052 24548
rect 3092 24508 3093 24548
rect 3051 24499 3093 24508
rect 2859 23792 2901 23801
rect 2859 23752 2860 23792
rect 2900 23752 2901 23792
rect 2859 23743 2901 23752
rect 3051 23540 3093 23549
rect 3051 23500 3052 23540
rect 3092 23500 3093 23540
rect 3051 23491 3093 23500
rect 2955 23204 2997 23213
rect 2955 23164 2956 23204
rect 2996 23164 2997 23204
rect 2955 23155 2997 23164
rect 2859 23120 2901 23129
rect 2859 23080 2860 23120
rect 2900 23080 2901 23120
rect 2859 23071 2901 23080
rect 2956 23120 2996 23155
rect 2763 21692 2805 21701
rect 2763 21652 2764 21692
rect 2804 21652 2805 21692
rect 2763 21643 2805 21652
rect 2572 21440 2612 21568
rect 2667 21608 2709 21617
rect 2667 21568 2668 21608
rect 2708 21568 2709 21608
rect 2667 21559 2709 21568
rect 2668 21474 2708 21559
rect 2380 21400 2612 21440
rect 2283 21020 2325 21029
rect 2283 20980 2284 21020
rect 2324 20980 2325 21020
rect 2283 20971 2325 20980
rect 2284 18509 2324 20971
rect 2380 20768 2420 21400
rect 2860 20852 2900 23071
rect 2956 23069 2996 23080
rect 3052 22616 3092 23491
rect 3148 23129 3188 25003
rect 3531 24632 3573 24641
rect 3531 24592 3532 24632
rect 3572 24592 3573 24632
rect 3531 24583 3573 24592
rect 3339 23792 3381 23801
rect 3339 23752 3340 23792
rect 3380 23752 3381 23792
rect 3339 23743 3381 23752
rect 3532 23792 3572 24583
rect 3724 24389 3764 25432
rect 4108 25304 4148 25507
rect 4108 25255 4148 25264
rect 3723 24380 3765 24389
rect 3723 24340 3724 24380
rect 3764 24340 3765 24380
rect 3723 24331 3765 24340
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 3147 23120 3189 23129
rect 3147 23080 3148 23120
rect 3188 23080 3189 23120
rect 3147 23071 3189 23080
rect 3340 23120 3380 23743
rect 3340 23071 3380 23080
rect 3436 23120 3476 23129
rect 3147 22868 3189 22877
rect 3147 22828 3148 22868
rect 3188 22828 3189 22868
rect 3147 22819 3189 22828
rect 3148 22734 3188 22819
rect 3052 22576 3284 22616
rect 3147 22028 3189 22037
rect 3147 21988 3148 22028
rect 3188 21988 3189 22028
rect 3147 21979 3189 21988
rect 3148 21869 3188 21979
rect 3147 21860 3189 21869
rect 3147 21820 3148 21860
rect 3188 21820 3189 21860
rect 3147 21811 3189 21820
rect 3051 21608 3093 21617
rect 3051 21568 3052 21608
rect 3092 21568 3093 21608
rect 3051 21559 3093 21568
rect 3148 21608 3188 21811
rect 3148 21559 3188 21568
rect 3052 21474 3092 21559
rect 3244 21440 3284 22576
rect 3436 21533 3476 23080
rect 3435 21524 3477 21533
rect 3435 21484 3436 21524
rect 3476 21484 3477 21524
rect 3435 21475 3477 21484
rect 3148 21400 3284 21440
rect 2955 21104 2997 21113
rect 2955 21064 2956 21104
rect 2996 21064 2997 21104
rect 2955 21055 2997 21064
rect 2956 20861 2996 21055
rect 2380 20719 2420 20728
rect 2475 20768 2517 20777
rect 2475 20728 2476 20768
rect 2516 20728 2517 20768
rect 2475 20719 2517 20728
rect 2476 20634 2516 20719
rect 2379 20516 2421 20525
rect 2379 20476 2380 20516
rect 2420 20476 2421 20516
rect 2379 20467 2421 20476
rect 2283 18500 2325 18509
rect 2283 18460 2284 18500
rect 2324 18460 2325 18500
rect 2283 18451 2325 18460
rect 2283 17660 2325 17669
rect 2283 17620 2284 17660
rect 2324 17620 2325 17660
rect 2283 17611 2325 17620
rect 2187 17408 2229 17417
rect 2187 17368 2188 17408
rect 2228 17368 2229 17408
rect 2187 17359 2229 17368
rect 2284 17333 2324 17611
rect 2091 17324 2133 17333
rect 2091 17284 2092 17324
rect 2132 17284 2133 17324
rect 2091 17275 2133 17284
rect 2283 17324 2325 17333
rect 2283 17284 2284 17324
rect 2324 17284 2325 17324
rect 2380 17324 2420 20467
rect 2764 20096 2804 20105
rect 2764 19769 2804 20056
rect 2571 19760 2613 19769
rect 2571 19720 2572 19760
rect 2612 19720 2613 19760
rect 2571 19711 2613 19720
rect 2763 19760 2805 19769
rect 2763 19720 2764 19760
rect 2804 19720 2805 19760
rect 2763 19711 2805 19720
rect 2572 19181 2612 19711
rect 2860 19424 2900 20812
rect 2955 20852 2997 20861
rect 2955 20812 2956 20852
rect 2996 20812 2997 20852
rect 2955 20803 2997 20812
rect 2956 20718 2996 20803
rect 3148 20357 3188 21400
rect 3339 20852 3381 20861
rect 3339 20812 3340 20852
rect 3380 20812 3381 20852
rect 3339 20803 3381 20812
rect 3243 20432 3285 20441
rect 3243 20392 3244 20432
rect 3284 20392 3285 20432
rect 3243 20383 3285 20392
rect 3147 20348 3189 20357
rect 3147 20308 3148 20348
rect 3188 20308 3189 20348
rect 3147 20299 3189 20308
rect 2956 20189 2996 20274
rect 2955 20180 2997 20189
rect 2955 20140 2956 20180
rect 2996 20140 2997 20180
rect 2955 20131 2997 20140
rect 3148 20096 3188 20105
rect 2956 20056 3148 20082
rect 2956 20042 3188 20056
rect 2956 19937 2996 20042
rect 2955 19928 2997 19937
rect 2955 19888 2956 19928
rect 2996 19888 2997 19928
rect 2955 19879 2997 19888
rect 3147 19928 3189 19937
rect 3147 19888 3148 19928
rect 3188 19888 3189 19928
rect 3147 19879 3189 19888
rect 2860 19384 3092 19424
rect 2764 19256 2804 19265
rect 2668 19216 2764 19256
rect 2571 19172 2613 19181
rect 2571 19132 2572 19172
rect 2612 19132 2613 19172
rect 2571 19123 2613 19132
rect 2668 18584 2708 19216
rect 2764 19207 2804 19216
rect 2859 19256 2901 19265
rect 2859 19216 2860 19256
rect 2900 19216 2901 19256
rect 2859 19207 2901 19216
rect 2860 19122 2900 19207
rect 2955 18752 2997 18761
rect 2955 18712 2956 18752
rect 2996 18712 2997 18752
rect 2955 18703 2997 18712
rect 2572 18544 2668 18584
rect 2475 17828 2517 17837
rect 2475 17788 2476 17828
rect 2516 17788 2517 17828
rect 2475 17779 2517 17788
rect 2476 17744 2516 17779
rect 2476 17693 2516 17704
rect 2380 17284 2516 17324
rect 2283 17275 2325 17284
rect 1995 17240 2037 17249
rect 1995 17200 1996 17240
rect 2036 17200 2037 17240
rect 1995 17191 2037 17200
rect 1804 17072 1844 17081
rect 1707 16568 1749 16577
rect 1707 16528 1708 16568
rect 1748 16528 1749 16568
rect 1707 16519 1749 16528
rect 1515 16400 1557 16409
rect 1804 16400 1844 17032
rect 1900 17072 1940 17081
rect 1900 16745 1940 17032
rect 1996 17072 2036 17081
rect 1899 16736 1941 16745
rect 1899 16696 1900 16736
rect 1940 16696 1941 16736
rect 1899 16687 1941 16696
rect 1996 16577 2036 17032
rect 2092 17072 2132 17083
rect 2092 16997 2132 17032
rect 2187 17072 2229 17081
rect 2380 17072 2420 17081
rect 2187 17032 2188 17072
rect 2228 17032 2229 17072
rect 2187 17023 2229 17032
rect 2284 17032 2380 17072
rect 2091 16988 2133 16997
rect 2091 16948 2092 16988
rect 2132 16948 2133 16988
rect 2091 16939 2133 16948
rect 1995 16568 2037 16577
rect 1995 16528 1996 16568
rect 2036 16528 2037 16568
rect 1995 16519 2037 16528
rect 1515 16360 1516 16400
rect 1556 16360 1557 16400
rect 1515 16351 1557 16360
rect 1612 16360 1844 16400
rect 2091 16400 2133 16409
rect 2091 16360 2092 16400
rect 2132 16360 2133 16400
rect 1228 16232 1268 16241
rect 1131 15980 1173 15989
rect 1131 15940 1132 15980
rect 1172 15940 1173 15980
rect 1131 15931 1173 15940
rect 1132 14393 1172 15931
rect 1228 15737 1268 16192
rect 1323 16232 1365 16241
rect 1323 16192 1324 16232
rect 1364 16192 1365 16232
rect 1323 16183 1365 16192
rect 1516 16232 1556 16241
rect 1324 16098 1364 16183
rect 1516 16073 1556 16192
rect 1420 16064 1460 16073
rect 1227 15728 1269 15737
rect 1227 15688 1228 15728
rect 1268 15688 1269 15728
rect 1227 15679 1269 15688
rect 1228 15560 1268 15571
rect 1228 15485 1268 15520
rect 1227 15476 1269 15485
rect 1227 15436 1228 15476
rect 1268 15436 1269 15476
rect 1227 15427 1269 15436
rect 1420 14804 1460 16024
rect 1515 16064 1557 16073
rect 1515 16024 1516 16064
rect 1556 16024 1557 16064
rect 1515 16015 1557 16024
rect 1515 14888 1557 14897
rect 1515 14848 1516 14888
rect 1556 14848 1557 14888
rect 1515 14839 1557 14848
rect 1420 14755 1460 14764
rect 1516 14754 1556 14839
rect 1612 14804 1652 16360
rect 2091 16351 2133 16360
rect 1707 16232 1749 16241
rect 1707 16192 1708 16232
rect 1748 16192 1749 16232
rect 1707 16183 1749 16192
rect 1900 16232 1940 16243
rect 1708 16098 1748 16183
rect 1900 16157 1940 16192
rect 1996 16232 2036 16241
rect 1899 16148 1941 16157
rect 1899 16108 1900 16148
rect 1940 16108 1941 16148
rect 1899 16099 1941 16108
rect 1612 14755 1652 14764
rect 1804 16064 1844 16073
rect 1324 14720 1364 14729
rect 1324 14636 1364 14680
rect 1708 14720 1748 14729
rect 1515 14636 1557 14645
rect 1324 14596 1516 14636
rect 1556 14596 1557 14636
rect 1515 14587 1557 14596
rect 1131 14384 1173 14393
rect 1131 14344 1132 14384
rect 1172 14344 1173 14384
rect 1131 14335 1173 14344
rect 1323 14300 1365 14309
rect 1323 14260 1324 14300
rect 1364 14260 1365 14300
rect 1323 14251 1365 14260
rect 1228 14048 1268 14057
rect 1324 14048 1364 14251
rect 1268 14008 1364 14048
rect 1228 13999 1268 14008
rect 1323 13796 1365 13805
rect 1323 13756 1324 13796
rect 1364 13756 1365 13796
rect 1323 13747 1365 13756
rect 1324 13217 1364 13747
rect 1228 13208 1268 13217
rect 1323 13208 1365 13217
rect 1268 13168 1324 13208
rect 1364 13168 1365 13208
rect 1228 13159 1268 13168
rect 1323 13159 1365 13168
rect 1324 13074 1364 13159
rect 1515 12788 1557 12797
rect 1515 12748 1516 12788
rect 1556 12748 1557 12788
rect 1515 12739 1557 12748
rect 1228 12536 1268 12545
rect 1323 12536 1365 12545
rect 1268 12496 1324 12536
rect 1364 12496 1365 12536
rect 1228 12487 1268 12496
rect 1323 12487 1365 12496
rect 1516 11948 1556 12739
rect 1516 11899 1556 11908
rect 1708 11873 1748 14680
rect 1804 14645 1844 16024
rect 1996 15317 2036 16192
rect 1995 15308 2037 15317
rect 1995 15268 1996 15308
rect 2036 15268 2037 15308
rect 1995 15259 2037 15268
rect 1995 15056 2037 15065
rect 1995 15016 1996 15056
rect 2036 15016 2037 15056
rect 1995 15007 2037 15016
rect 1899 14720 1941 14729
rect 1899 14680 1900 14720
rect 1940 14680 1941 14720
rect 1899 14671 1941 14680
rect 1803 14636 1845 14645
rect 1803 14596 1804 14636
rect 1844 14596 1845 14636
rect 1803 14587 1845 14596
rect 1900 14586 1940 14671
rect 1996 14393 2036 15007
rect 1803 14384 1845 14393
rect 1803 14344 1804 14384
rect 1844 14344 1845 14384
rect 1803 14335 1845 14344
rect 1995 14384 2037 14393
rect 1995 14344 1996 14384
rect 2036 14344 2037 14384
rect 1995 14335 2037 14344
rect 1707 11864 1749 11873
rect 1707 11824 1708 11864
rect 1748 11824 1749 11864
rect 1707 11815 1749 11824
rect 1323 11696 1365 11705
rect 1707 11696 1749 11705
rect 1323 11656 1324 11696
rect 1364 11656 1365 11696
rect 1323 11647 1365 11656
rect 1612 11656 1708 11696
rect 1748 11656 1749 11696
rect 1228 11528 1268 11537
rect 1228 11360 1268 11488
rect 1132 11320 1268 11360
rect 1132 7160 1172 11320
rect 1324 11192 1364 11647
rect 1516 11528 1556 11537
rect 1516 11360 1556 11488
rect 1324 11143 1364 11152
rect 1420 11320 1556 11360
rect 1420 10352 1460 11320
rect 1516 11024 1556 11033
rect 1612 11024 1652 11656
rect 1707 11647 1749 11656
rect 1708 11562 1748 11647
rect 1556 10984 1652 11024
rect 1516 10975 1556 10984
rect 1611 10688 1653 10697
rect 1611 10648 1612 10688
rect 1652 10648 1653 10688
rect 1611 10639 1653 10648
rect 1324 10312 1460 10352
rect 1228 10184 1268 10193
rect 1228 10025 1268 10144
rect 1227 10016 1269 10025
rect 1227 9976 1228 10016
rect 1268 9976 1269 10016
rect 1227 9967 1269 9976
rect 1324 9512 1364 10312
rect 1419 10016 1461 10025
rect 1419 9976 1420 10016
rect 1460 9976 1461 10016
rect 1419 9967 1461 9976
rect 1324 9428 1364 9472
rect 1420 9437 1460 9967
rect 1515 9512 1557 9521
rect 1515 9472 1516 9512
rect 1556 9472 1557 9512
rect 1515 9463 1557 9472
rect 1612 9512 1652 10639
rect 1804 9773 1844 14335
rect 1899 14300 1941 14309
rect 1899 14260 1900 14300
rect 1940 14260 1941 14300
rect 1899 14251 1941 14260
rect 1803 9764 1845 9773
rect 1803 9724 1804 9764
rect 1844 9724 1845 9764
rect 1803 9715 1845 9724
rect 1803 9596 1845 9605
rect 1803 9556 1804 9596
rect 1844 9556 1845 9596
rect 1803 9547 1845 9556
rect 1228 9388 1364 9428
rect 1419 9428 1461 9437
rect 1419 9388 1420 9428
rect 1460 9388 1461 9428
rect 1228 9092 1268 9388
rect 1419 9379 1461 9388
rect 1516 9378 1556 9463
rect 1324 9260 1364 9269
rect 1364 9220 1556 9260
rect 1324 9211 1364 9220
rect 1228 9052 1460 9092
rect 1227 8672 1269 8681
rect 1227 8632 1228 8672
rect 1268 8632 1269 8672
rect 1227 8623 1269 8632
rect 1228 8538 1268 8623
rect 1228 8000 1268 8009
rect 1323 8000 1365 8009
rect 1268 7960 1324 8000
rect 1364 7960 1365 8000
rect 1228 7951 1268 7960
rect 1323 7951 1365 7960
rect 1228 7160 1268 7169
rect 1132 7120 1228 7160
rect 1228 7111 1268 7120
rect 1420 7160 1460 9052
rect 1516 7589 1556 9220
rect 1612 7673 1652 9472
rect 1804 9512 1844 9547
rect 1804 9461 1844 9472
rect 1900 7757 1940 14251
rect 1995 14216 2037 14225
rect 1995 14176 1996 14216
rect 2036 14176 2037 14216
rect 1995 14167 2037 14176
rect 1996 12209 2036 14167
rect 2092 12797 2132 16351
rect 2188 14225 2228 17023
rect 2284 16232 2324 17032
rect 2380 17023 2420 17032
rect 2476 17072 2516 17284
rect 2379 16316 2421 16325
rect 2379 16276 2380 16316
rect 2420 16276 2421 16316
rect 2379 16267 2421 16276
rect 2187 14216 2229 14225
rect 2187 14176 2188 14216
rect 2228 14176 2229 14216
rect 2187 14167 2229 14176
rect 2284 13889 2324 16192
rect 2380 16232 2420 16267
rect 2380 16181 2420 16192
rect 2476 16064 2516 17032
rect 2380 16024 2516 16064
rect 2283 13880 2325 13889
rect 2283 13840 2284 13880
rect 2324 13840 2325 13880
rect 2283 13831 2325 13840
rect 2283 13712 2325 13721
rect 2283 13672 2284 13712
rect 2324 13672 2325 13712
rect 2283 13663 2325 13672
rect 2187 13460 2229 13469
rect 2187 13420 2188 13460
rect 2228 13420 2229 13460
rect 2187 13411 2229 13420
rect 2091 12788 2133 12797
rect 2091 12748 2092 12788
rect 2132 12748 2133 12788
rect 2091 12739 2133 12748
rect 2188 12368 2228 13411
rect 2092 12328 2228 12368
rect 1995 12200 2037 12209
rect 1995 12160 1996 12200
rect 2036 12160 2037 12200
rect 1995 12151 2037 12160
rect 1995 9512 2037 9521
rect 1995 9472 1996 9512
rect 2036 9472 2037 9512
rect 1995 9463 2037 9472
rect 1996 9185 2036 9463
rect 1995 9176 2037 9185
rect 1995 9136 1996 9176
rect 2036 9136 2037 9176
rect 1995 9127 2037 9136
rect 1899 7748 1941 7757
rect 1899 7708 1900 7748
rect 1940 7708 1941 7748
rect 1899 7699 1941 7708
rect 1611 7664 1653 7673
rect 1611 7624 1612 7664
rect 1652 7624 1653 7664
rect 1611 7615 1653 7624
rect 1803 7664 1845 7673
rect 1803 7624 1804 7664
rect 1844 7624 1845 7664
rect 1803 7615 1845 7624
rect 1515 7580 1557 7589
rect 1515 7540 1516 7580
rect 1556 7540 1557 7580
rect 1515 7531 1557 7540
rect 1611 7496 1653 7505
rect 1611 7456 1612 7496
rect 1652 7456 1653 7496
rect 1611 7447 1653 7456
rect 1515 7328 1557 7337
rect 1515 7288 1516 7328
rect 1556 7288 1557 7328
rect 1515 7279 1557 7288
rect 1323 7076 1365 7085
rect 1323 7036 1324 7076
rect 1364 7036 1365 7076
rect 1323 7027 1365 7036
rect 1324 6942 1364 7027
rect 1420 6749 1460 7120
rect 1516 7160 1556 7279
rect 1516 7111 1556 7120
rect 1419 6740 1461 6749
rect 1419 6700 1420 6740
rect 1460 6700 1461 6740
rect 1419 6691 1461 6700
rect 1612 6656 1652 7447
rect 1708 7160 1748 7169
rect 1708 7001 1748 7120
rect 1804 7160 1844 7615
rect 1899 7580 1941 7589
rect 1899 7540 1900 7580
rect 1940 7540 1941 7580
rect 1899 7531 1941 7540
rect 1804 7111 1844 7120
rect 1900 7160 1940 7531
rect 1995 7412 2037 7421
rect 1995 7372 1996 7412
rect 2036 7372 2037 7412
rect 1995 7363 2037 7372
rect 1900 7111 1940 7120
rect 1996 7160 2036 7363
rect 1996 7111 2036 7120
rect 2092 7085 2132 12328
rect 2187 12200 2229 12209
rect 2187 12160 2188 12200
rect 2228 12160 2229 12200
rect 2187 12151 2229 12160
rect 2188 8933 2228 12151
rect 2187 8924 2229 8933
rect 2187 8884 2188 8924
rect 2228 8884 2229 8924
rect 2187 8875 2229 8884
rect 2187 8672 2229 8681
rect 2187 8632 2188 8672
rect 2228 8632 2229 8672
rect 2187 8623 2229 8632
rect 2188 8009 2228 8623
rect 2187 8000 2229 8009
rect 2187 7960 2188 8000
rect 2228 7960 2229 8000
rect 2187 7951 2229 7960
rect 2188 7160 2228 7951
rect 2188 7111 2228 7120
rect 2091 7076 2133 7085
rect 2091 7036 2092 7076
rect 2132 7036 2133 7076
rect 2091 7027 2133 7036
rect 1707 6992 1749 7001
rect 1707 6952 1708 6992
rect 1748 6952 1749 6992
rect 1707 6943 1749 6952
rect 1707 6824 1749 6833
rect 1707 6784 1708 6824
rect 1748 6784 1749 6824
rect 1707 6775 1749 6784
rect 1612 6607 1652 6616
rect 1228 6488 1268 6497
rect 1132 6448 1228 6488
rect 1132 4061 1172 6448
rect 1228 6439 1268 6448
rect 1420 6488 1460 6497
rect 1460 6448 1556 6488
rect 1420 6439 1460 6448
rect 1419 6236 1461 6245
rect 1419 6196 1420 6236
rect 1460 6196 1461 6236
rect 1419 6187 1461 6196
rect 1420 6102 1460 6187
rect 1516 5825 1556 6448
rect 1611 6068 1653 6077
rect 1611 6028 1612 6068
rect 1652 6028 1653 6068
rect 1611 6019 1653 6028
rect 1515 5816 1557 5825
rect 1515 5776 1516 5816
rect 1556 5776 1557 5816
rect 1515 5767 1557 5776
rect 1612 5732 1652 6019
rect 1708 5816 1748 6775
rect 2091 6740 2133 6749
rect 2091 6700 2092 6740
rect 2132 6700 2133 6740
rect 2091 6691 2133 6700
rect 1899 6572 1941 6581
rect 1899 6532 1900 6572
rect 1940 6532 1945 6572
rect 1899 6523 1945 6532
rect 1905 6497 1945 6523
rect 1803 6488 1845 6497
rect 1803 6448 1804 6488
rect 1844 6448 1845 6488
rect 1803 6439 1845 6448
rect 2092 6488 2132 6691
rect 1945 6457 2036 6483
rect 1905 6443 2036 6457
rect 1905 6442 1945 6443
rect 1804 6354 1844 6439
rect 1899 6152 1941 6161
rect 1899 6112 1900 6152
rect 1940 6112 1941 6152
rect 1899 6103 1941 6112
rect 1804 5816 1844 5825
rect 1708 5776 1804 5816
rect 1804 5767 1844 5776
rect 1612 5692 1748 5732
rect 1228 5648 1268 5657
rect 1228 5405 1268 5608
rect 1323 5648 1365 5657
rect 1323 5608 1324 5648
rect 1364 5608 1365 5648
rect 1323 5599 1365 5608
rect 1516 5648 1556 5657
rect 1708 5648 1748 5692
rect 1556 5608 1652 5648
rect 1516 5599 1556 5608
rect 1324 5514 1364 5599
rect 1420 5480 1460 5489
rect 1460 5440 1556 5480
rect 1420 5431 1460 5440
rect 1227 5396 1269 5405
rect 1227 5356 1228 5396
rect 1268 5356 1269 5396
rect 1227 5347 1269 5356
rect 1419 5144 1461 5153
rect 1419 5104 1420 5144
rect 1460 5104 1461 5144
rect 1419 5095 1461 5104
rect 1228 4976 1268 4985
rect 1228 4817 1268 4936
rect 1420 4976 1460 5095
rect 1420 4927 1460 4936
rect 1227 4808 1269 4817
rect 1227 4768 1228 4808
rect 1268 4768 1269 4808
rect 1227 4759 1269 4768
rect 1324 4724 1364 4733
rect 1227 4220 1269 4229
rect 1227 4180 1228 4220
rect 1268 4180 1269 4220
rect 1227 4171 1269 4180
rect 1228 4086 1268 4171
rect 1131 4052 1173 4061
rect 1131 4012 1132 4052
rect 1172 4012 1173 4052
rect 1131 4003 1173 4012
rect 1227 3968 1269 3977
rect 1227 3928 1228 3968
rect 1268 3928 1269 3968
rect 1324 3968 1364 4684
rect 1516 4136 1556 5440
rect 1612 5144 1652 5608
rect 1708 5599 1748 5608
rect 1900 5648 1940 6103
rect 1900 5599 1940 5608
rect 1996 5648 2036 6443
rect 2092 6439 2132 6448
rect 2188 6488 2228 6497
rect 2284 6488 2324 13663
rect 2380 8429 2420 16024
rect 2572 15728 2612 18544
rect 2668 18535 2708 18544
rect 2763 18584 2805 18593
rect 2763 18544 2764 18584
rect 2804 18544 2805 18584
rect 2763 18535 2805 18544
rect 2764 18450 2804 18535
rect 2859 18500 2901 18509
rect 2859 18460 2860 18500
rect 2900 18460 2901 18500
rect 2859 18451 2901 18460
rect 2667 17996 2709 18005
rect 2667 17956 2668 17996
rect 2708 17956 2709 17996
rect 2667 17947 2709 17956
rect 2668 17862 2708 17947
rect 2860 17912 2900 18451
rect 2956 18425 2996 18703
rect 2955 18416 2997 18425
rect 2955 18376 2956 18416
rect 2996 18376 2997 18416
rect 2955 18367 2997 18376
rect 2764 17872 2900 17912
rect 2764 16232 2804 17872
rect 2859 17744 2901 17753
rect 2859 17704 2860 17744
rect 2900 17704 2901 17744
rect 2859 17695 2901 17704
rect 2860 17610 2900 17695
rect 2955 17492 2997 17501
rect 2955 17452 2956 17492
rect 2996 17452 2997 17492
rect 2955 17443 2997 17452
rect 2859 17408 2901 17417
rect 2859 17368 2860 17408
rect 2900 17368 2901 17408
rect 2859 17359 2901 17368
rect 2860 16988 2900 17359
rect 2956 17072 2996 17443
rect 2956 17023 2996 17032
rect 2860 16913 2900 16948
rect 2859 16904 2901 16913
rect 2859 16864 2860 16904
rect 2900 16864 2901 16904
rect 2859 16855 2901 16864
rect 2859 16484 2901 16493
rect 2859 16444 2860 16484
rect 2900 16444 2901 16484
rect 2859 16435 2901 16444
rect 2860 16316 2900 16435
rect 3052 16325 3092 19384
rect 3148 18668 3188 19879
rect 3244 19340 3284 20383
rect 3340 20180 3380 20803
rect 3436 20768 3476 20777
rect 3436 20357 3476 20728
rect 3435 20348 3477 20357
rect 3435 20308 3436 20348
rect 3476 20308 3477 20348
rect 3435 20299 3477 20308
rect 3340 20140 3476 20180
rect 3244 19291 3284 19300
rect 3340 19256 3380 19265
rect 3340 18929 3380 19216
rect 3339 18920 3381 18929
rect 3339 18880 3340 18920
rect 3380 18880 3381 18920
rect 3339 18871 3381 18880
rect 3148 18628 3380 18668
rect 3147 18500 3189 18509
rect 3147 18460 3148 18500
rect 3188 18460 3189 18500
rect 3147 18451 3189 18460
rect 3244 18500 3284 18511
rect 3148 18366 3188 18451
rect 3244 18425 3284 18460
rect 3243 18416 3285 18425
rect 3243 18376 3244 18416
rect 3284 18376 3285 18416
rect 3243 18367 3285 18376
rect 3147 16568 3189 16577
rect 3147 16528 3148 16568
rect 3188 16528 3189 16568
rect 3147 16519 3189 16528
rect 2860 16267 2900 16276
rect 3051 16316 3093 16325
rect 3051 16276 3052 16316
rect 3092 16276 3093 16316
rect 3051 16267 3093 16276
rect 2668 15728 2708 15737
rect 2572 15688 2668 15728
rect 2668 15679 2708 15688
rect 2476 15560 2516 15569
rect 2476 14897 2516 15520
rect 2475 14888 2517 14897
rect 2475 14848 2476 14888
rect 2516 14848 2517 14888
rect 2475 14839 2517 14848
rect 2476 14048 2516 14839
rect 2764 14393 2804 16192
rect 3051 16064 3093 16073
rect 3051 16024 3052 16064
rect 3092 16024 3093 16064
rect 3051 16015 3093 16024
rect 2956 15560 2996 15569
rect 2860 15520 2956 15560
rect 2763 14384 2805 14393
rect 2763 14344 2764 14384
rect 2804 14344 2805 14384
rect 2763 14335 2805 14344
rect 2668 14216 2708 14225
rect 2860 14216 2900 15520
rect 2956 15511 2996 15520
rect 3052 15392 3092 16015
rect 2708 14176 2900 14216
rect 2956 15352 3092 15392
rect 2668 14167 2708 14176
rect 2476 13208 2516 14008
rect 2860 14048 2900 14059
rect 2860 13973 2900 14008
rect 2859 13964 2901 13973
rect 2859 13924 2860 13964
rect 2900 13924 2901 13964
rect 2859 13915 2901 13924
rect 2571 13880 2613 13889
rect 2571 13840 2572 13880
rect 2612 13840 2613 13880
rect 2571 13831 2613 13840
rect 2572 13460 2612 13831
rect 2668 13460 2708 13469
rect 2572 13420 2668 13460
rect 2668 13411 2708 13420
rect 2956 13292 2996 15352
rect 3148 15233 3188 16519
rect 3244 16493 3284 18367
rect 3340 16829 3380 18628
rect 3436 18341 3476 20140
rect 3532 19769 3572 23752
rect 3724 23624 3764 23633
rect 3627 23288 3669 23297
rect 3627 23248 3628 23288
rect 3668 23248 3669 23288
rect 3627 23239 3669 23248
rect 3628 23154 3668 23239
rect 3724 23129 3764 23584
rect 4012 23624 4052 23633
rect 4012 23381 4052 23584
rect 4204 23465 4244 25852
rect 4588 25472 4628 27868
rect 4684 27665 4724 28624
rect 4780 28253 4820 29632
rect 4876 29623 4916 29632
rect 5067 29672 5109 29681
rect 5067 29632 5068 29672
rect 5108 29632 5109 29672
rect 5067 29623 5109 29632
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 4875 29168 4917 29177
rect 4875 29128 4876 29168
rect 4916 29128 4917 29168
rect 4875 29119 4917 29128
rect 4876 29034 4916 29119
rect 5355 28916 5397 28925
rect 5355 28876 5356 28916
rect 5396 28876 5397 28916
rect 5355 28867 5397 28876
rect 5260 28328 5300 28339
rect 4779 28244 4821 28253
rect 4779 28204 4780 28244
rect 4820 28204 4821 28244
rect 4779 28195 4821 28204
rect 4876 28169 4916 28254
rect 5260 28253 5300 28288
rect 5259 28244 5301 28253
rect 5259 28204 5260 28244
rect 5300 28204 5301 28244
rect 5259 28195 5301 28204
rect 4875 28160 4917 28169
rect 4875 28120 4876 28160
rect 4916 28120 4917 28160
rect 4875 28111 4917 28120
rect 4779 27992 4821 28001
rect 4779 27952 4780 27992
rect 4820 27952 4821 27992
rect 4779 27943 4821 27952
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4683 27656 4725 27665
rect 4683 27616 4684 27656
rect 4724 27616 4725 27656
rect 4683 27607 4725 27616
rect 4684 27077 4724 27607
rect 4683 27068 4725 27077
rect 4683 27028 4684 27068
rect 4724 27028 4725 27068
rect 4683 27019 4725 27028
rect 4684 26816 4724 26825
rect 4780 26816 4820 27943
rect 4875 27656 4917 27665
rect 4875 27616 4876 27656
rect 4916 27616 4917 27656
rect 4875 27607 4917 27616
rect 5356 27651 5396 28867
rect 4876 27522 4916 27607
rect 5356 27602 5396 27611
rect 4724 26776 4820 26816
rect 5355 26816 5397 26825
rect 5355 26776 5356 26816
rect 5396 26776 5397 26816
rect 4684 26237 4724 26776
rect 5355 26767 5397 26776
rect 4779 26564 4821 26573
rect 4779 26524 4780 26564
rect 4820 26524 4821 26564
rect 4779 26515 4821 26524
rect 4780 26312 4820 26515
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 5163 26312 5205 26321
rect 4780 26272 5012 26312
rect 4683 26228 4725 26237
rect 4683 26188 4684 26228
rect 4724 26188 4725 26228
rect 4683 26179 4725 26188
rect 4972 26144 5012 26272
rect 5163 26272 5164 26312
rect 5204 26272 5205 26312
rect 5163 26263 5205 26272
rect 4972 26095 5012 26104
rect 4684 26060 4724 26069
rect 4684 25733 4724 26020
rect 4683 25724 4725 25733
rect 4683 25684 4684 25724
rect 4724 25684 4725 25724
rect 4683 25675 4725 25684
rect 4396 25432 4628 25472
rect 4299 24632 4341 24641
rect 4299 24592 4300 24632
rect 4340 24592 4341 24632
rect 4299 24583 4341 24592
rect 4300 24498 4340 24583
rect 4300 23792 4340 23801
rect 4396 23792 4436 25432
rect 4683 25388 4725 25397
rect 4683 25348 4684 25388
rect 4724 25348 4725 25388
rect 4683 25339 4725 25348
rect 4588 25304 4628 25313
rect 4491 25220 4533 25229
rect 4588 25220 4628 25264
rect 4684 25254 4724 25339
rect 5067 25304 5109 25313
rect 5067 25264 5068 25304
rect 5108 25264 5109 25304
rect 5067 25255 5109 25264
rect 5164 25304 5204 26263
rect 5356 26228 5396 26767
rect 5356 26179 5396 26188
rect 5260 26144 5300 26153
rect 5260 25649 5300 26104
rect 5259 25640 5301 25649
rect 5259 25600 5260 25640
rect 5300 25600 5301 25640
rect 5259 25591 5301 25600
rect 5164 25255 5204 25264
rect 4491 25180 4492 25220
rect 4532 25180 4628 25220
rect 4491 25171 4533 25180
rect 5068 25170 5108 25255
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 4684 24632 4724 24641
rect 4684 24473 4724 24592
rect 4683 24464 4725 24473
rect 4683 24424 4684 24464
rect 4724 24424 4725 24464
rect 4683 24415 4725 24424
rect 4491 24380 4533 24389
rect 4491 24340 4492 24380
rect 4532 24340 4533 24380
rect 4491 24331 4533 24340
rect 4492 24246 4532 24331
rect 4340 23752 4436 23792
rect 4300 23743 4340 23752
rect 4203 23456 4245 23465
rect 4203 23416 4204 23456
rect 4244 23416 4245 23456
rect 4203 23407 4245 23416
rect 4011 23372 4053 23381
rect 4011 23332 4012 23372
rect 4052 23332 4053 23372
rect 4011 23323 4053 23332
rect 3723 23120 3765 23129
rect 3723 23080 3724 23120
rect 3764 23080 3765 23120
rect 3723 23071 3765 23080
rect 4012 22868 4052 23323
rect 4107 23120 4149 23129
rect 4107 23080 4108 23120
rect 4148 23080 4149 23120
rect 4107 23071 4149 23080
rect 4204 23120 4244 23129
rect 4108 22986 4148 23071
rect 4204 23036 4244 23080
rect 4299 23036 4341 23045
rect 4204 22996 4300 23036
rect 4340 22996 4341 23036
rect 4299 22987 4341 22996
rect 4396 22877 4436 23752
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4683 23372 4725 23381
rect 4683 23332 4684 23372
rect 4724 23332 4725 23372
rect 4683 23323 4725 23332
rect 4684 23120 4724 23323
rect 4684 23071 4724 23080
rect 5163 23120 5205 23129
rect 5163 23080 5164 23120
rect 5204 23080 5205 23120
rect 5163 23071 5205 23080
rect 4587 23036 4629 23045
rect 4587 22996 4588 23036
rect 4628 22996 4629 23036
rect 4587 22987 4629 22996
rect 4588 22902 4628 22987
rect 5164 22986 5204 23071
rect 4203 22868 4245 22877
rect 4012 22828 4148 22868
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3723 22532 3765 22541
rect 3723 22492 3724 22532
rect 3764 22492 3765 22532
rect 3723 22483 3765 22492
rect 3627 22280 3669 22289
rect 3627 22240 3628 22280
rect 3668 22240 3669 22280
rect 3627 22231 3669 22240
rect 3628 22146 3668 22231
rect 3628 21608 3668 21617
rect 3724 21608 3764 22483
rect 4108 22448 4148 22828
rect 4203 22828 4204 22868
rect 4244 22828 4245 22868
rect 4203 22819 4245 22828
rect 4395 22868 4437 22877
rect 4395 22828 4396 22868
rect 4436 22828 4437 22868
rect 4395 22819 4437 22828
rect 4971 22868 5013 22877
rect 4971 22828 4972 22868
rect 5012 22828 5013 22868
rect 4971 22819 5013 22828
rect 4108 22399 4148 22408
rect 3820 22112 3860 22121
rect 3820 21617 3860 22072
rect 4107 21692 4149 21701
rect 4107 21652 4108 21692
rect 4148 21652 4149 21692
rect 4107 21643 4149 21652
rect 3668 21568 3764 21608
rect 3819 21608 3861 21617
rect 3819 21568 3820 21608
rect 3860 21568 3861 21608
rect 3628 21449 3668 21568
rect 3819 21559 3861 21568
rect 4108 21603 4148 21643
rect 4204 21608 4244 22819
rect 4491 22532 4533 22541
rect 4491 22492 4492 22532
rect 4532 22492 4533 22532
rect 4491 22483 4533 22492
rect 4492 22398 4532 22483
rect 4683 22448 4725 22457
rect 4683 22408 4684 22448
rect 4724 22408 4725 22448
rect 4683 22399 4725 22408
rect 4299 22364 4341 22373
rect 4299 22324 4300 22364
rect 4340 22324 4341 22364
rect 4299 22315 4341 22324
rect 4300 22230 4340 22315
rect 4684 22314 4724 22399
rect 4972 22280 5012 22819
rect 4780 22240 4972 22280
rect 4300 21785 4340 21870
rect 4299 21776 4341 21785
rect 4299 21736 4300 21776
rect 4340 21736 4341 21776
rect 4299 21727 4341 21736
rect 4588 21608 4628 21617
rect 4204 21568 4588 21608
rect 3627 21440 3669 21449
rect 3627 21400 3628 21440
rect 3668 21400 3669 21440
rect 3627 21391 3669 21400
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 4108 20936 4148 21563
rect 4588 21559 4628 21568
rect 4203 21104 4245 21113
rect 4203 21064 4204 21104
rect 4244 21064 4245 21104
rect 4203 21055 4245 21064
rect 4012 20896 4148 20936
rect 4012 20852 4052 20896
rect 3964 20812 4052 20852
rect 3964 20810 4004 20812
rect 3964 20761 4004 20770
rect 4108 20693 4148 20778
rect 4107 20684 4149 20693
rect 4107 20644 4108 20684
rect 4148 20644 4149 20684
rect 4107 20635 4149 20644
rect 3819 20600 3861 20609
rect 3819 20560 3820 20600
rect 3860 20560 3861 20600
rect 3819 20551 3861 20560
rect 3820 19853 3860 20551
rect 3819 19844 3861 19853
rect 3819 19804 3820 19844
rect 3860 19804 3861 19844
rect 3819 19795 3861 19804
rect 3531 19760 3573 19769
rect 3531 19720 3532 19760
rect 3572 19720 3573 19760
rect 3531 19711 3573 19720
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 3531 19256 3573 19265
rect 3531 19216 3532 19256
rect 3572 19216 3573 19256
rect 3531 19207 3573 19216
rect 3820 19256 3860 19265
rect 3532 18509 3572 19207
rect 3627 19172 3669 19181
rect 3627 19132 3628 19172
rect 3668 19132 3669 19172
rect 3627 19123 3669 19132
rect 3531 18500 3573 18509
rect 3531 18460 3532 18500
rect 3572 18460 3573 18500
rect 3531 18451 3573 18460
rect 3435 18332 3477 18341
rect 3628 18332 3668 19123
rect 3820 19097 3860 19216
rect 4204 19097 4244 21055
rect 4491 20936 4533 20945
rect 4491 20896 4492 20936
rect 4532 20896 4533 20936
rect 4491 20887 4533 20896
rect 4299 20852 4341 20861
rect 4299 20812 4300 20852
rect 4340 20812 4341 20852
rect 4299 20803 4341 20812
rect 4300 20718 4340 20803
rect 4492 20802 4532 20887
rect 4396 20096 4436 20105
rect 4396 19769 4436 20056
rect 4587 19928 4629 19937
rect 4587 19888 4588 19928
rect 4628 19888 4629 19928
rect 4587 19879 4629 19888
rect 4588 19794 4628 19879
rect 4395 19760 4437 19769
rect 4395 19720 4396 19760
rect 4436 19720 4437 19760
rect 4395 19711 4437 19720
rect 4300 19261 4340 19270
rect 3819 19088 3861 19097
rect 3819 19048 3820 19088
rect 3860 19048 3861 19088
rect 3819 19039 3861 19048
rect 4203 19088 4245 19097
rect 4203 19048 4204 19088
rect 4244 19048 4245 19088
rect 4203 19039 4245 19048
rect 3724 18584 3764 18593
rect 4300 18584 4340 19221
rect 4396 18929 4436 19711
rect 4780 19349 4820 22240
rect 4972 22231 5012 22240
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4875 21692 4917 21701
rect 4875 21652 4876 21692
rect 4916 21652 4917 21692
rect 4875 21643 4917 21652
rect 4876 21608 4916 21643
rect 4876 21557 4916 21568
rect 4972 21608 5012 21617
rect 4972 20693 5012 21568
rect 5259 21440 5301 21449
rect 5259 21400 5260 21440
rect 5300 21400 5301 21440
rect 5259 21391 5301 21400
rect 5163 21356 5205 21365
rect 5163 21316 5164 21356
rect 5204 21316 5205 21356
rect 5163 21307 5205 21316
rect 5164 20936 5204 21307
rect 5260 21306 5300 21391
rect 5355 21272 5397 21281
rect 5355 21232 5356 21272
rect 5396 21232 5397 21272
rect 5355 21223 5397 21232
rect 5204 20896 5300 20936
rect 5164 20887 5204 20896
rect 4971 20684 5013 20693
rect 4971 20644 4972 20684
rect 5012 20644 5013 20684
rect 4971 20635 5013 20644
rect 5260 20600 5300 20896
rect 5356 20861 5396 21223
rect 5355 20852 5397 20861
rect 5355 20812 5356 20852
rect 5396 20812 5397 20852
rect 5355 20803 5397 20812
rect 5356 20768 5396 20803
rect 5356 20718 5396 20728
rect 5260 20560 5396 20600
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 5356 20264 5396 20560
rect 5260 20224 5396 20264
rect 5163 20096 5205 20105
rect 5163 20056 5164 20096
rect 5204 20056 5205 20096
rect 5163 20047 5205 20056
rect 5260 20096 5300 20224
rect 4875 20012 4917 20021
rect 4875 19972 4876 20012
rect 4916 19972 4917 20012
rect 4875 19963 4917 19972
rect 4876 19878 4916 19963
rect 5164 19962 5204 20047
rect 5164 19424 5204 19433
rect 5260 19424 5300 20056
rect 5204 19384 5300 19424
rect 5164 19375 5204 19384
rect 4779 19340 4821 19349
rect 4779 19300 4780 19340
rect 4820 19300 4821 19340
rect 4779 19291 4821 19300
rect 5260 19181 5300 19384
rect 5259 19172 5301 19181
rect 5259 19132 5260 19172
rect 5300 19132 5301 19172
rect 5259 19123 5301 19132
rect 4492 19088 4532 19097
rect 4532 19048 4820 19088
rect 4492 19039 4532 19048
rect 4395 18920 4437 18929
rect 4395 18880 4396 18920
rect 4436 18880 4437 18920
rect 4395 18871 4437 18880
rect 4395 18668 4437 18677
rect 4395 18628 4396 18668
rect 4436 18628 4437 18668
rect 4395 18619 4437 18628
rect 3724 18341 3764 18544
rect 4204 18570 4340 18584
rect 4244 18544 4340 18570
rect 4396 18534 4436 18619
rect 4684 18584 4724 18593
rect 4492 18544 4684 18584
rect 4780 18584 4820 19048
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 5067 18668 5109 18677
rect 5067 18628 5068 18668
rect 5108 18628 5109 18668
rect 5067 18619 5109 18628
rect 4972 18584 5012 18593
rect 4780 18544 4972 18584
rect 3435 18292 3436 18332
rect 3476 18292 3477 18332
rect 3435 18283 3477 18292
rect 3532 18292 3668 18332
rect 3723 18332 3765 18341
rect 3723 18292 3724 18332
rect 3764 18292 3765 18332
rect 3436 17072 3476 17083
rect 3436 16997 3476 17032
rect 3435 16988 3477 16997
rect 3435 16948 3436 16988
rect 3476 16948 3477 16988
rect 3435 16939 3477 16948
rect 3339 16820 3381 16829
rect 3339 16780 3340 16820
rect 3380 16780 3381 16820
rect 3339 16771 3381 16780
rect 3243 16484 3285 16493
rect 3243 16444 3244 16484
rect 3284 16444 3476 16484
rect 3243 16435 3285 16444
rect 3340 16232 3380 16241
rect 3340 15989 3380 16192
rect 3339 15980 3381 15989
rect 3339 15940 3340 15980
rect 3380 15940 3381 15980
rect 3339 15931 3381 15940
rect 3339 15644 3381 15653
rect 3339 15604 3340 15644
rect 3380 15604 3381 15644
rect 3339 15595 3381 15604
rect 3243 15560 3285 15569
rect 3243 15520 3244 15560
rect 3284 15520 3285 15560
rect 3243 15511 3285 15520
rect 3244 15426 3284 15511
rect 3340 15510 3380 15595
rect 3243 15308 3285 15317
rect 3243 15268 3244 15308
rect 3284 15268 3285 15308
rect 3243 15259 3285 15268
rect 3147 15224 3189 15233
rect 3147 15184 3148 15224
rect 3188 15184 3189 15224
rect 3147 15175 3189 15184
rect 3147 14888 3189 14897
rect 3147 14848 3148 14888
rect 3188 14848 3189 14888
rect 3147 14839 3189 14848
rect 3148 14720 3188 14839
rect 3148 14671 3188 14680
rect 2476 12536 2516 13168
rect 2668 13252 2996 13292
rect 3051 13292 3093 13301
rect 3051 13252 3052 13292
rect 3092 13252 3093 13292
rect 2571 12872 2613 12881
rect 2571 12832 2572 12872
rect 2612 12832 2613 12872
rect 2571 12823 2613 12832
rect 2476 11705 2516 12496
rect 2475 11696 2517 11705
rect 2475 11656 2476 11696
rect 2516 11656 2517 11696
rect 2475 11647 2517 11656
rect 2476 10184 2516 11647
rect 2476 10135 2516 10144
rect 2475 8756 2517 8765
rect 2475 8716 2476 8756
rect 2516 8716 2517 8756
rect 2475 8707 2517 8716
rect 2476 8672 2516 8707
rect 2572 8681 2612 12823
rect 2668 12704 2708 13252
rect 3051 13243 3093 13252
rect 3052 13208 3092 13243
rect 3052 13157 3092 13168
rect 2668 12655 2708 12664
rect 2860 13040 2900 13049
rect 2860 11192 2900 13000
rect 2956 12536 2996 12545
rect 2956 12377 2996 12496
rect 2955 12368 2997 12377
rect 2955 12328 2956 12368
rect 2996 12328 2997 12368
rect 2955 12319 2997 12328
rect 3244 12368 3284 15259
rect 3339 14972 3381 14981
rect 3339 14932 3340 14972
rect 3380 14932 3381 14972
rect 3339 14923 3381 14932
rect 3340 14838 3380 14923
rect 3436 14636 3476 16444
rect 3532 16325 3572 18292
rect 3723 18283 3765 18292
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 4204 18089 4244 18530
rect 4203 18080 4245 18089
rect 4203 18040 4204 18080
rect 4244 18040 4245 18080
rect 4203 18031 4245 18040
rect 4300 17996 4340 18005
rect 4492 17996 4532 18544
rect 4684 18535 4724 18544
rect 4972 18535 5012 18544
rect 5068 18534 5108 18619
rect 4779 18332 4821 18341
rect 4779 18292 4780 18332
rect 4820 18292 4821 18332
rect 4779 18283 4821 18292
rect 5356 18332 5396 18341
rect 4683 18080 4725 18089
rect 4683 18040 4684 18080
rect 4724 18040 4725 18080
rect 4683 18031 4725 18040
rect 4340 17956 4532 17996
rect 4300 17947 4340 17956
rect 4108 17753 4148 17838
rect 4395 17828 4437 17837
rect 4395 17788 4396 17828
rect 4436 17788 4437 17828
rect 4395 17779 4437 17788
rect 4587 17828 4629 17837
rect 4587 17788 4588 17828
rect 4628 17788 4629 17828
rect 4587 17779 4629 17788
rect 4107 17744 4149 17753
rect 4107 17704 4108 17744
rect 4148 17704 4149 17744
rect 4107 17695 4149 17704
rect 4299 17744 4341 17753
rect 4299 17704 4300 17744
rect 4340 17704 4341 17744
rect 4299 17695 4341 17704
rect 3915 17156 3957 17165
rect 3915 17116 3916 17156
rect 3956 17116 3957 17156
rect 3915 17107 3957 17116
rect 4108 17156 4148 17165
rect 3916 17067 3956 17107
rect 3916 17018 3956 17027
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 4108 16484 4148 17116
rect 4300 16577 4340 17695
rect 4299 16568 4341 16577
rect 4299 16528 4300 16568
rect 4340 16528 4341 16568
rect 4299 16519 4341 16528
rect 4100 16444 4148 16484
rect 3819 16400 3861 16409
rect 3819 16360 3820 16400
rect 3860 16360 3861 16400
rect 3819 16351 3861 16360
rect 3531 16316 3573 16325
rect 3531 16276 3532 16316
rect 3572 16276 3573 16316
rect 3531 16267 3573 16276
rect 3820 16237 3860 16351
rect 4100 16316 4140 16444
rect 4100 16276 4148 16316
rect 3531 16148 3573 16157
rect 3531 16108 3532 16148
rect 3572 16108 3573 16148
rect 3531 16099 3573 16108
rect 3532 14972 3572 16099
rect 3820 15980 3860 16197
rect 4012 16064 4052 16073
rect 3820 15940 3956 15980
rect 3819 15728 3861 15737
rect 3819 15688 3820 15728
rect 3860 15688 3861 15728
rect 3819 15679 3861 15688
rect 3820 15560 3860 15679
rect 3820 15511 3860 15520
rect 3628 15317 3668 15402
rect 3916 15392 3956 15940
rect 4012 15653 4052 16024
rect 4011 15644 4053 15653
rect 4011 15604 4012 15644
rect 4052 15604 4053 15644
rect 4011 15595 4053 15604
rect 4108 15569 4148 16276
rect 4204 16232 4244 16243
rect 4204 16157 4244 16192
rect 4299 16232 4341 16241
rect 4299 16192 4300 16232
rect 4340 16192 4341 16232
rect 4299 16183 4341 16192
rect 4203 16148 4245 16157
rect 4203 16108 4204 16148
rect 4244 16108 4245 16148
rect 4203 16099 4245 16108
rect 4300 16098 4340 16183
rect 4396 15737 4436 17779
rect 4491 17744 4533 17753
rect 4491 17704 4492 17744
rect 4532 17704 4533 17744
rect 4491 17695 4533 17704
rect 4492 17610 4532 17695
rect 4492 17072 4532 17081
rect 4588 17072 4628 17779
rect 4532 17032 4628 17072
rect 4492 17023 4532 17032
rect 4587 16232 4629 16241
rect 4587 16192 4588 16232
rect 4628 16192 4629 16232
rect 4587 16183 4629 16192
rect 4588 16098 4628 16183
rect 4395 15728 4437 15737
rect 4395 15688 4396 15728
rect 4436 15688 4437 15728
rect 4395 15679 4437 15688
rect 4107 15560 4149 15569
rect 4107 15520 4108 15560
rect 4148 15520 4149 15560
rect 4107 15511 4149 15520
rect 4587 15560 4629 15569
rect 4684 15560 4724 18031
rect 4587 15520 4588 15560
rect 4628 15520 4724 15560
rect 4587 15511 4629 15520
rect 4203 15476 4245 15485
rect 4203 15436 4204 15476
rect 4244 15436 4245 15476
rect 4203 15427 4245 15436
rect 3916 15352 4148 15392
rect 3627 15308 3669 15317
rect 3627 15268 3628 15308
rect 3668 15268 3669 15308
rect 3627 15259 3669 15268
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 4108 14981 4148 15352
rect 4204 15317 4244 15427
rect 4203 15308 4245 15317
rect 4203 15268 4204 15308
rect 4244 15268 4245 15308
rect 4203 15259 4245 15268
rect 4299 15224 4341 15233
rect 4299 15184 4300 15224
rect 4340 15184 4341 15224
rect 4299 15175 4341 15184
rect 3532 14923 3572 14932
rect 4107 14972 4149 14981
rect 4107 14932 4108 14972
rect 4148 14932 4149 14972
rect 4107 14923 4149 14932
rect 3723 14888 3765 14897
rect 3723 14848 3724 14888
rect 3764 14848 3765 14888
rect 3723 14839 3765 14848
rect 3724 14720 3764 14839
rect 4107 14804 4149 14813
rect 4107 14764 4108 14804
rect 4148 14764 4149 14804
rect 4107 14755 4149 14764
rect 3724 14671 3764 14680
rect 3340 14596 3476 14636
rect 3340 12881 3380 14596
rect 3532 14552 3572 14561
rect 3436 14512 3532 14552
rect 3339 12872 3381 12881
rect 3339 12832 3340 12872
rect 3380 12832 3381 12872
rect 3339 12823 3381 12832
rect 3436 12704 3476 14512
rect 3532 14503 3572 14512
rect 4108 14048 4148 14755
rect 4300 14729 4340 15175
rect 4299 14720 4341 14729
rect 4299 14680 4300 14720
rect 4340 14680 4341 14720
rect 4299 14671 4341 14680
rect 4300 14216 4340 14671
rect 4300 14167 4340 14176
rect 4108 13999 4148 14008
rect 3531 13964 3573 13973
rect 3531 13924 3532 13964
rect 3572 13924 3573 13964
rect 3531 13915 3573 13924
rect 3532 12881 3572 13915
rect 4491 13880 4533 13889
rect 4491 13840 4492 13880
rect 4532 13840 4533 13880
rect 4491 13831 4533 13840
rect 4300 13796 4340 13805
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 4300 13385 4340 13756
rect 4492 13746 4532 13831
rect 3915 13376 3957 13385
rect 3915 13336 3916 13376
rect 3956 13336 3957 13376
rect 3915 13327 3957 13336
rect 4299 13376 4341 13385
rect 4299 13336 4300 13376
rect 4340 13336 4341 13376
rect 4299 13327 4341 13336
rect 3627 13208 3669 13217
rect 3627 13168 3628 13208
rect 3668 13168 3669 13208
rect 3627 13159 3669 13168
rect 3531 12872 3573 12881
rect 3531 12832 3532 12872
rect 3572 12832 3573 12872
rect 3531 12823 3573 12832
rect 3244 12319 3284 12328
rect 3340 12664 3476 12704
rect 2956 12125 2996 12319
rect 3052 12284 3092 12293
rect 2955 12116 2997 12125
rect 2955 12076 2956 12116
rect 2996 12076 2997 12116
rect 2955 12067 2997 12076
rect 2955 11948 2997 11957
rect 2955 11908 2956 11948
rect 2996 11908 2997 11948
rect 2955 11899 2997 11908
rect 2956 11738 2996 11899
rect 2956 11689 2996 11698
rect 2955 11612 2997 11621
rect 2955 11572 2956 11612
rect 2996 11572 2997 11612
rect 2955 11563 2997 11572
rect 2668 11152 2900 11192
rect 2956 11192 2996 11563
rect 3052 11444 3092 12244
rect 3147 12032 3189 12041
rect 3147 11992 3148 12032
rect 3188 11992 3189 12032
rect 3147 11983 3189 11992
rect 3148 11696 3188 11983
rect 3148 11647 3188 11656
rect 3147 11444 3189 11453
rect 3052 11404 3148 11444
rect 3188 11404 3189 11444
rect 3147 11395 3189 11404
rect 2668 10856 2708 11152
rect 2956 11143 2996 11152
rect 3051 11192 3093 11201
rect 3051 11152 3052 11192
rect 3092 11152 3093 11192
rect 3051 11143 3093 11152
rect 2764 11024 2804 11033
rect 2804 10984 2996 11024
rect 2764 10975 2804 10984
rect 2859 10856 2901 10865
rect 2668 10816 2804 10856
rect 2667 10688 2709 10697
rect 2667 10648 2668 10688
rect 2708 10648 2709 10688
rect 2667 10639 2709 10648
rect 2668 10436 2708 10639
rect 2668 10387 2708 10396
rect 2379 8420 2421 8429
rect 2379 8380 2380 8420
rect 2420 8380 2421 8420
rect 2379 8371 2421 8380
rect 2379 8168 2421 8177
rect 2379 8128 2380 8168
rect 2420 8128 2421 8168
rect 2379 8119 2421 8128
rect 2380 6833 2420 8119
rect 2476 8000 2516 8632
rect 2571 8672 2613 8681
rect 2571 8632 2572 8672
rect 2612 8632 2613 8672
rect 2571 8623 2613 8632
rect 2668 8504 2708 8513
rect 2668 8261 2708 8464
rect 2667 8252 2709 8261
rect 2476 7951 2516 7960
rect 2572 8212 2668 8252
rect 2708 8212 2709 8252
rect 2379 6824 2421 6833
rect 2572 6824 2612 8212
rect 2667 8203 2709 8212
rect 2668 8084 2708 8095
rect 2668 8009 2708 8044
rect 2667 8000 2709 8009
rect 2667 7960 2668 8000
rect 2708 7960 2709 8000
rect 2667 7951 2709 7960
rect 2667 6908 2709 6917
rect 2667 6868 2668 6908
rect 2708 6868 2709 6908
rect 2667 6859 2709 6868
rect 2379 6784 2380 6824
rect 2420 6784 2421 6824
rect 2379 6775 2421 6784
rect 2500 6784 2612 6824
rect 2500 6740 2540 6784
rect 2476 6700 2540 6740
rect 2379 6656 2421 6665
rect 2379 6616 2380 6656
rect 2420 6616 2421 6656
rect 2379 6607 2421 6616
rect 2380 6522 2420 6607
rect 2476 6581 2516 6700
rect 2572 6656 2612 6665
rect 2668 6656 2708 6859
rect 2612 6616 2708 6656
rect 2572 6607 2612 6616
rect 2475 6572 2517 6581
rect 2475 6532 2476 6572
rect 2516 6532 2517 6572
rect 2475 6523 2517 6532
rect 2228 6448 2324 6488
rect 2764 6483 2804 10816
rect 2859 10816 2860 10856
rect 2900 10816 2901 10856
rect 2859 10807 2901 10816
rect 2860 10436 2900 10807
rect 2860 10387 2900 10396
rect 2859 9932 2901 9941
rect 2859 9892 2860 9932
rect 2900 9892 2901 9932
rect 2859 9883 2901 9892
rect 2860 8756 2900 9883
rect 2956 9773 2996 10984
rect 3052 10025 3092 11143
rect 3340 11108 3380 12664
rect 3532 12536 3572 12545
rect 3435 11444 3477 11453
rect 3435 11404 3436 11444
rect 3476 11404 3477 11444
rect 3435 11395 3477 11404
rect 3436 11201 3476 11395
rect 3435 11192 3477 11201
rect 3435 11152 3436 11192
rect 3476 11152 3477 11192
rect 3435 11143 3477 11152
rect 3532 11117 3572 12496
rect 3628 12536 3668 13159
rect 3628 12293 3668 12496
rect 3916 12536 3956 13327
rect 4300 13208 4340 13217
rect 4300 13049 4340 13168
rect 4299 13040 4341 13049
rect 4299 13000 4300 13040
rect 4340 13000 4341 13040
rect 4299 12991 4341 13000
rect 4491 13040 4533 13049
rect 4491 13000 4492 13040
rect 4532 13000 4533 13040
rect 4491 12991 4533 13000
rect 4492 12906 4532 12991
rect 4203 12872 4245 12881
rect 4203 12832 4204 12872
rect 4244 12832 4245 12872
rect 4203 12823 4245 12832
rect 3916 12293 3956 12496
rect 4204 12536 4244 12823
rect 4204 12487 4244 12496
rect 3627 12284 3669 12293
rect 3627 12244 3628 12284
rect 3668 12244 3669 12284
rect 3627 12235 3669 12244
rect 3915 12284 3957 12293
rect 3915 12244 3916 12284
rect 3956 12244 3957 12284
rect 3915 12235 3957 12244
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 4588 11705 4628 15511
rect 4683 14972 4725 14981
rect 4683 14932 4684 14972
rect 4724 14932 4725 14972
rect 4683 14923 4725 14932
rect 4684 14132 4724 14923
rect 4780 14720 4820 18283
rect 5356 18089 5396 18292
rect 5355 18080 5397 18089
rect 5355 18040 5356 18080
rect 5396 18040 5397 18080
rect 5355 18031 5397 18040
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 5452 15737 5492 32227
rect 5548 29000 5588 32404
rect 5644 30680 5684 33991
rect 5836 33956 5876 34999
rect 5931 34880 5973 34889
rect 5931 34840 5932 34880
rect 5972 34840 5973 34880
rect 5931 34831 5973 34840
rect 5740 33916 5876 33956
rect 5740 33797 5780 33916
rect 5739 33788 5781 33797
rect 5739 33748 5740 33788
rect 5780 33748 5781 33788
rect 5739 33739 5781 33748
rect 5835 33704 5877 33713
rect 5835 33664 5836 33704
rect 5876 33664 5877 33704
rect 5835 33655 5877 33664
rect 5644 30631 5684 30640
rect 5740 30680 5780 30689
rect 5740 30512 5780 30640
rect 5644 30472 5780 30512
rect 5644 29177 5684 30472
rect 5643 29168 5685 29177
rect 5643 29128 5644 29168
rect 5684 29128 5685 29168
rect 5643 29119 5685 29128
rect 5836 29084 5876 33655
rect 5932 32033 5972 34831
rect 6124 33704 6164 34999
rect 6124 32864 6164 33664
rect 6220 33629 6260 35839
rect 6412 35309 6452 39544
rect 6796 39425 6836 41551
rect 6892 41264 6932 41273
rect 6892 40424 6932 41224
rect 6892 40349 6932 40384
rect 6891 40340 6933 40349
rect 6891 40300 6892 40340
rect 6932 40300 6933 40340
rect 6891 40291 6933 40300
rect 6891 39668 6933 39677
rect 6891 39628 6892 39668
rect 6932 39628 6933 39668
rect 6891 39619 6933 39628
rect 6892 39534 6932 39619
rect 6507 39416 6549 39425
rect 6507 39376 6508 39416
rect 6548 39376 6549 39416
rect 6507 39367 6549 39376
rect 6795 39416 6837 39425
rect 6795 39376 6796 39416
rect 6836 39376 6837 39416
rect 6795 39367 6837 39376
rect 6508 38921 6548 39367
rect 6603 39080 6645 39089
rect 6603 39040 6604 39080
rect 6644 39040 6645 39080
rect 6603 39031 6645 39040
rect 6700 39080 6740 39089
rect 6891 39080 6933 39089
rect 6740 39040 6892 39080
rect 6932 39040 6933 39080
rect 6700 39031 6740 39040
rect 6891 39031 6933 39040
rect 6507 38912 6549 38921
rect 6507 38872 6508 38912
rect 6548 38872 6549 38912
rect 6507 38863 6549 38872
rect 6508 38576 6548 38863
rect 6604 38660 6644 39031
rect 6892 38912 6932 38923
rect 6892 38837 6932 38872
rect 6891 38828 6933 38837
rect 6891 38788 6892 38828
rect 6932 38788 6933 38828
rect 6891 38779 6933 38788
rect 6604 38620 6836 38660
rect 6508 38536 6559 38576
rect 6519 38492 6559 38536
rect 6508 38452 6559 38492
rect 6508 38408 6548 38452
rect 6508 38368 6644 38408
rect 6507 38072 6549 38081
rect 6507 38032 6508 38072
rect 6548 38032 6549 38072
rect 6507 38023 6549 38032
rect 6411 35300 6453 35309
rect 6411 35260 6412 35300
rect 6452 35260 6453 35300
rect 6508 35300 6548 38023
rect 6604 37400 6644 38368
rect 6699 38240 6741 38249
rect 6699 38200 6700 38240
rect 6740 38200 6741 38240
rect 6699 38191 6741 38200
rect 6796 38240 6836 38620
rect 6796 38191 6836 38200
rect 6700 38106 6740 38191
rect 6892 38081 6932 38779
rect 6891 38072 6933 38081
rect 6891 38032 6892 38072
rect 6932 38032 6933 38072
rect 6891 38023 6933 38032
rect 6988 37913 7028 42928
rect 7180 41609 7220 42928
rect 7275 42440 7317 42449
rect 7275 42400 7276 42440
rect 7316 42400 7317 42440
rect 7275 42391 7317 42400
rect 7179 41600 7221 41609
rect 7179 41560 7180 41600
rect 7220 41560 7221 41600
rect 7179 41551 7221 41560
rect 7084 41264 7124 41273
rect 7084 40265 7124 41224
rect 7083 40256 7125 40265
rect 7083 40216 7084 40256
rect 7124 40216 7125 40256
rect 7083 40207 7125 40216
rect 7276 39752 7316 42391
rect 7372 41609 7412 42928
rect 7564 41861 7604 42928
rect 7563 41852 7605 41861
rect 7563 41812 7564 41852
rect 7604 41812 7605 41852
rect 7563 41803 7605 41812
rect 7659 41768 7701 41777
rect 7659 41728 7660 41768
rect 7700 41728 7701 41768
rect 7659 41719 7701 41728
rect 7371 41600 7413 41609
rect 7371 41560 7372 41600
rect 7412 41560 7413 41600
rect 7371 41551 7413 41560
rect 7467 41516 7509 41525
rect 7467 41476 7468 41516
rect 7508 41476 7509 41516
rect 7467 41467 7509 41476
rect 7468 39920 7508 41467
rect 7660 41180 7700 41719
rect 7756 41264 7796 42928
rect 7948 41609 7988 42928
rect 8140 42785 8180 42928
rect 8139 42776 8181 42785
rect 8139 42736 8140 42776
rect 8180 42736 8181 42776
rect 8139 42727 8181 42736
rect 8332 41693 8372 42928
rect 8524 41861 8564 42928
rect 8523 41852 8565 41861
rect 8523 41812 8524 41852
rect 8564 41812 8565 41852
rect 8523 41803 8565 41812
rect 8331 41684 8373 41693
rect 8331 41644 8332 41684
rect 8372 41644 8373 41684
rect 8331 41635 8373 41644
rect 7947 41600 7989 41609
rect 7947 41560 7948 41600
rect 7988 41560 7989 41600
rect 7947 41551 7989 41560
rect 8332 41264 8372 41273
rect 7756 41224 8276 41264
rect 7660 41140 7988 41180
rect 7468 39871 7508 39880
rect 7276 39712 7412 39752
rect 7083 39668 7125 39677
rect 7083 39628 7084 39668
rect 7124 39628 7125 39668
rect 7083 39619 7125 39628
rect 7084 39534 7124 39619
rect 7275 39584 7317 39593
rect 7275 39544 7276 39584
rect 7316 39544 7317 39584
rect 7275 39535 7317 39544
rect 7276 39450 7316 39535
rect 7083 39416 7125 39425
rect 7083 39376 7084 39416
rect 7124 39376 7125 39416
rect 7083 39367 7125 39376
rect 6987 37904 7029 37913
rect 6987 37864 6988 37904
rect 7028 37864 7029 37904
rect 6987 37855 7029 37864
rect 6699 37820 6741 37829
rect 7084 37820 7124 39367
rect 7275 39164 7317 39173
rect 7275 39124 7276 39164
rect 7316 39124 7317 39164
rect 7275 39115 7317 39124
rect 7276 38156 7316 39115
rect 6699 37780 6700 37820
rect 6740 37780 6932 37820
rect 7084 37780 7220 37820
rect 6699 37771 6741 37780
rect 6892 37484 6932 37780
rect 7180 37652 7220 37780
rect 7276 37745 7316 38116
rect 7372 37988 7412 39712
rect 7660 39668 7700 39677
rect 7851 39668 7893 39677
rect 7700 39628 7796 39668
rect 7660 39619 7700 39628
rect 7467 39080 7509 39089
rect 7467 39040 7468 39080
rect 7508 39040 7509 39080
rect 7467 39031 7509 39040
rect 7468 38156 7508 39031
rect 7659 38408 7701 38417
rect 7659 38368 7660 38408
rect 7700 38368 7701 38408
rect 7659 38359 7701 38368
rect 7660 38240 7700 38359
rect 7660 38191 7700 38200
rect 7468 38116 7604 38156
rect 7468 37988 7508 37997
rect 7372 37948 7468 37988
rect 7468 37939 7508 37948
rect 7564 37820 7604 38116
rect 7756 37820 7796 39628
rect 7851 39628 7852 39668
rect 7892 39628 7893 39668
rect 7851 39619 7893 39628
rect 7852 39534 7892 39619
rect 7948 37820 7988 41140
rect 8139 41012 8181 41021
rect 8139 40972 8140 41012
rect 8180 40972 8181 41012
rect 8139 40963 8181 40972
rect 8140 40424 8180 40963
rect 8044 39500 8084 39509
rect 8044 39257 8084 39460
rect 8043 39248 8085 39257
rect 8043 39208 8044 39248
rect 8084 39208 8085 39248
rect 8043 39199 8085 39208
rect 8140 38921 8180 40384
rect 8236 39920 8276 41224
rect 8332 41021 8372 41224
rect 8716 41180 8756 42928
rect 8908 41777 8948 42928
rect 8907 41768 8949 41777
rect 8907 41728 8908 41768
rect 8948 41728 8949 41768
rect 8907 41719 8949 41728
rect 8428 41140 8756 41180
rect 8908 41264 8948 41273
rect 8331 41012 8373 41021
rect 8331 40972 8332 41012
rect 8372 40972 8373 41012
rect 8331 40963 8373 40972
rect 8332 40265 8372 40350
rect 8331 40256 8373 40265
rect 8331 40216 8332 40256
rect 8372 40216 8373 40256
rect 8331 40207 8373 40216
rect 8428 40088 8468 41140
rect 8524 41012 8564 41021
rect 8564 40972 8660 41012
rect 8524 40963 8564 40972
rect 8523 40256 8565 40265
rect 8523 40216 8524 40256
rect 8564 40216 8565 40256
rect 8523 40207 8565 40216
rect 8236 39871 8276 39880
rect 8332 40048 8468 40088
rect 8332 39416 8372 40048
rect 8427 39668 8469 39677
rect 8427 39628 8428 39668
rect 8468 39628 8469 39668
rect 8427 39619 8469 39628
rect 8428 39534 8468 39619
rect 8332 39376 8468 39416
rect 8139 38912 8181 38921
rect 8139 38872 8140 38912
rect 8180 38872 8181 38912
rect 8139 38863 8181 38872
rect 8140 38778 8180 38863
rect 8332 38744 8372 38753
rect 7564 37780 7700 37820
rect 7756 37780 7892 37820
rect 7948 37780 8084 37820
rect 7275 37736 7317 37745
rect 7275 37696 7276 37736
rect 7316 37696 7317 37736
rect 7275 37687 7317 37696
rect 7180 37603 7220 37612
rect 7467 37652 7509 37661
rect 7467 37612 7468 37652
rect 7508 37612 7509 37652
rect 7467 37603 7509 37612
rect 6988 37484 7028 37493
rect 6892 37444 6988 37484
rect 6644 37360 6740 37400
rect 6604 37351 6644 37360
rect 6700 35888 6740 37360
rect 6796 37232 6836 37241
rect 6796 36065 6836 37192
rect 6795 36056 6837 36065
rect 6795 36016 6796 36056
rect 6836 36016 6837 36056
rect 6795 36007 6837 36016
rect 6796 35888 6836 35897
rect 6700 35848 6796 35888
rect 6508 35260 6644 35300
rect 6411 35251 6453 35260
rect 6411 35132 6453 35141
rect 6411 35092 6412 35132
rect 6452 35092 6453 35132
rect 6411 35083 6453 35092
rect 6508 35132 6548 35141
rect 6412 34998 6452 35083
rect 6508 35057 6548 35092
rect 6507 35048 6549 35057
rect 6507 35008 6508 35048
rect 6548 35008 6549 35048
rect 6507 34999 6549 35008
rect 6508 34721 6548 34999
rect 6507 34712 6549 34721
rect 6507 34672 6508 34712
rect 6548 34672 6549 34712
rect 6507 34663 6549 34672
rect 6604 34637 6644 35260
rect 6603 34628 6645 34637
rect 6603 34588 6604 34628
rect 6644 34588 6645 34628
rect 6603 34579 6645 34588
rect 6507 33704 6549 33713
rect 6507 33664 6508 33704
rect 6548 33664 6549 33704
rect 6507 33655 6549 33664
rect 6604 33704 6644 33715
rect 6219 33620 6261 33629
rect 6219 33580 6220 33620
rect 6260 33580 6261 33620
rect 6219 33571 6261 33580
rect 6028 32824 6124 32864
rect 6028 32285 6068 32824
rect 6124 32815 6164 32824
rect 6123 32444 6165 32453
rect 6123 32404 6124 32444
rect 6164 32404 6165 32444
rect 6123 32395 6165 32404
rect 6027 32276 6069 32285
rect 6027 32236 6028 32276
rect 6068 32236 6069 32276
rect 6027 32227 6069 32236
rect 5931 32024 5973 32033
rect 5931 31984 5932 32024
rect 5972 31984 5973 32024
rect 5931 31975 5973 31984
rect 6124 30680 6164 32395
rect 6220 31613 6260 33571
rect 6508 33570 6548 33655
rect 6604 33629 6644 33664
rect 6603 33620 6645 33629
rect 6603 33580 6604 33620
rect 6644 33580 6645 33620
rect 6603 33571 6645 33580
rect 6315 33452 6357 33461
rect 6315 33412 6316 33452
rect 6356 33412 6357 33452
rect 6315 33403 6357 33412
rect 6316 33318 6356 33403
rect 6700 33125 6740 35848
rect 6796 35839 6836 35848
rect 6892 34208 6932 37444
rect 6988 37435 7028 37444
rect 7468 37400 7508 37603
rect 7468 37351 7508 37360
rect 7564 37400 7604 37409
rect 7180 36728 7220 36737
rect 7084 36688 7180 36728
rect 6987 35804 7029 35813
rect 6987 35764 6988 35804
rect 7028 35764 7029 35804
rect 6987 35755 7029 35764
rect 6988 35670 7028 35755
rect 6987 35552 7029 35561
rect 6987 35512 6988 35552
rect 7028 35512 7029 35552
rect 6987 35503 7029 35512
rect 6988 35216 7028 35503
rect 6988 35167 7028 35176
rect 7084 34889 7124 36688
rect 7180 36679 7220 36688
rect 7371 36476 7413 36485
rect 7371 36436 7372 36476
rect 7412 36436 7413 36476
rect 7371 36427 7413 36436
rect 7372 36342 7412 36427
rect 7564 36233 7604 37360
rect 7660 36728 7700 37780
rect 7660 36679 7700 36688
rect 7756 36728 7796 36737
rect 7371 36224 7413 36233
rect 7371 36184 7372 36224
rect 7412 36184 7413 36224
rect 7371 36175 7413 36184
rect 7563 36224 7605 36233
rect 7756 36224 7796 36688
rect 7563 36184 7564 36224
rect 7604 36184 7796 36224
rect 7563 36175 7605 36184
rect 7275 36056 7317 36065
rect 7275 36016 7276 36056
rect 7316 36016 7317 36056
rect 7275 36007 7317 36016
rect 7276 35888 7316 36007
rect 7276 35839 7316 35848
rect 7372 35888 7412 36175
rect 7852 36140 7892 37780
rect 7948 37400 7988 37409
rect 7948 36728 7988 37360
rect 8044 37400 8084 37780
rect 8332 37661 8372 38704
rect 8331 37652 8373 37661
rect 8331 37612 8332 37652
rect 8372 37612 8373 37652
rect 8331 37603 8373 37612
rect 8084 37360 8276 37400
rect 8044 37351 8084 37360
rect 8140 36737 8180 36822
rect 8139 36728 8181 36737
rect 7948 36688 8140 36728
rect 8180 36688 8181 36728
rect 7947 36308 7989 36317
rect 7947 36268 7948 36308
rect 7988 36268 7989 36308
rect 7947 36259 7989 36268
rect 7660 36100 7892 36140
rect 7372 35645 7412 35848
rect 7563 35888 7605 35897
rect 7563 35848 7564 35888
rect 7604 35848 7605 35888
rect 7563 35839 7605 35848
rect 7371 35636 7413 35645
rect 7371 35596 7372 35636
rect 7412 35596 7413 35636
rect 7371 35587 7413 35596
rect 7564 35384 7604 35839
rect 7660 35477 7700 36100
rect 7852 35897 7892 35982
rect 7756 35888 7796 35897
rect 7756 35720 7796 35848
rect 7851 35888 7893 35897
rect 7948 35888 7988 36259
rect 7851 35848 7852 35888
rect 7892 35848 7988 35888
rect 7851 35839 7893 35848
rect 8044 35720 8084 36688
rect 8139 36679 8181 36688
rect 8236 36644 8276 37360
rect 8139 36476 8181 36485
rect 8139 36436 8140 36476
rect 8180 36436 8181 36476
rect 8139 36427 8181 36436
rect 7756 35680 8084 35720
rect 7659 35468 7701 35477
rect 7659 35428 7660 35468
rect 7700 35428 7701 35468
rect 7659 35419 7701 35428
rect 7756 35393 7796 35680
rect 7468 35344 7604 35384
rect 7755 35384 7797 35393
rect 7755 35344 7756 35384
rect 7796 35344 7797 35384
rect 7468 35300 7508 35344
rect 7755 35335 7797 35344
rect 7372 35260 7508 35300
rect 7660 35300 7700 35309
rect 7372 35057 7412 35260
rect 7660 35225 7700 35260
rect 7659 35216 7701 35225
rect 7468 35202 7508 35211
rect 7659 35176 7660 35216
rect 7700 35176 7701 35216
rect 7659 35167 7701 35176
rect 7852 35216 7892 35227
rect 7660 35165 7700 35167
rect 7371 35048 7413 35057
rect 7371 35008 7372 35048
rect 7412 35008 7413 35048
rect 7371 34999 7413 35008
rect 7083 34880 7125 34889
rect 7083 34840 7084 34880
rect 7124 34840 7125 34880
rect 7083 34831 7125 34840
rect 6988 34385 7028 34470
rect 6987 34376 7029 34385
rect 6987 34336 6988 34376
rect 7028 34336 7029 34376
rect 6987 34327 7029 34336
rect 6892 34168 7028 34208
rect 6796 33704 6836 33713
rect 6836 33664 6932 33704
rect 6796 33655 6836 33664
rect 6796 33452 6836 33461
rect 6699 33116 6741 33125
rect 6699 33076 6700 33116
rect 6740 33076 6741 33116
rect 6699 33067 6741 33076
rect 6652 32906 6692 32915
rect 6604 32866 6652 32883
rect 6604 32843 6692 32866
rect 6316 32780 6356 32789
rect 6604 32780 6644 32843
rect 6796 32789 6836 33412
rect 6356 32740 6644 32780
rect 6795 32780 6837 32789
rect 6795 32740 6796 32780
rect 6836 32740 6837 32780
rect 6316 32731 6356 32740
rect 6795 32731 6837 32740
rect 6508 32654 6548 32663
rect 6508 32537 6548 32614
rect 6507 32528 6549 32537
rect 6507 32488 6508 32528
rect 6548 32488 6549 32528
rect 6507 32479 6549 32488
rect 6892 32444 6932 33664
rect 6796 32404 6932 32444
rect 6699 32276 6741 32285
rect 6699 32236 6700 32276
rect 6740 32236 6741 32276
rect 6699 32227 6741 32236
rect 6508 32192 6548 32201
rect 6508 32033 6548 32152
rect 6700 32142 6740 32227
rect 6507 32024 6549 32033
rect 6507 31984 6508 32024
rect 6548 31984 6549 32024
rect 6507 31975 6549 31984
rect 6219 31604 6261 31613
rect 6219 31564 6220 31604
rect 6260 31564 6261 31604
rect 6219 31555 6261 31564
rect 6219 31436 6261 31445
rect 6219 31396 6220 31436
rect 6260 31396 6261 31436
rect 6219 31387 6261 31396
rect 6220 31352 6260 31387
rect 6220 31301 6260 31312
rect 6604 31352 6644 31361
rect 6507 31268 6549 31277
rect 6507 31228 6508 31268
rect 6548 31228 6549 31268
rect 6507 31219 6549 31228
rect 6508 30857 6548 31219
rect 6604 31109 6644 31312
rect 6603 31100 6645 31109
rect 6603 31060 6604 31100
rect 6644 31060 6645 31100
rect 6603 31051 6645 31060
rect 6507 30848 6549 30857
rect 6507 30808 6508 30848
rect 6548 30808 6549 30848
rect 6507 30799 6549 30808
rect 6220 30680 6260 30689
rect 6124 30640 6220 30680
rect 6220 30631 6260 30640
rect 6508 30680 6548 30799
rect 6508 30631 6548 30640
rect 5740 29044 5876 29084
rect 6028 30428 6068 30437
rect 5548 28960 5684 29000
rect 5547 28832 5589 28841
rect 5547 28792 5548 28832
rect 5588 28792 5589 28832
rect 5547 28783 5589 28792
rect 5548 28160 5588 28783
rect 5644 28664 5684 28960
rect 5740 28841 5780 29044
rect 6028 29000 6068 30388
rect 6316 30428 6356 30437
rect 6316 30269 6356 30388
rect 6507 30428 6549 30437
rect 6507 30388 6508 30428
rect 6548 30388 6549 30428
rect 6507 30379 6549 30388
rect 6315 30260 6357 30269
rect 6315 30220 6316 30260
rect 6356 30220 6357 30260
rect 6315 30211 6357 30220
rect 6316 29840 6356 29851
rect 6316 29765 6356 29800
rect 6315 29756 6357 29765
rect 6315 29716 6316 29756
rect 6356 29716 6357 29756
rect 6315 29707 6357 29716
rect 6508 29504 6548 30379
rect 6699 30008 6741 30017
rect 6699 29968 6700 30008
rect 6740 29968 6741 30008
rect 6699 29959 6741 29968
rect 6700 29840 6740 29959
rect 6700 29681 6740 29800
rect 6699 29672 6741 29681
rect 6699 29632 6700 29672
rect 6740 29632 6741 29672
rect 6699 29623 6741 29632
rect 6508 29464 6740 29504
rect 6123 29420 6165 29429
rect 6123 29380 6124 29420
rect 6164 29380 6165 29420
rect 6123 29371 6165 29380
rect 5836 28960 6068 29000
rect 6124 29168 6164 29371
rect 6507 29336 6549 29345
rect 6507 29296 6508 29336
rect 6548 29296 6549 29336
rect 6507 29287 6549 29296
rect 5739 28832 5781 28841
rect 5739 28792 5740 28832
rect 5780 28792 5781 28832
rect 5739 28783 5781 28792
rect 5644 28624 5780 28664
rect 5548 28120 5684 28160
rect 5548 27740 5588 27749
rect 5548 27245 5588 27700
rect 5547 27236 5589 27245
rect 5547 27196 5548 27236
rect 5588 27196 5589 27236
rect 5547 27187 5589 27196
rect 5547 27068 5589 27077
rect 5547 27028 5548 27068
rect 5588 27028 5589 27068
rect 5547 27019 5589 27028
rect 5548 25304 5588 27019
rect 5644 25976 5684 28120
rect 5740 27488 5780 28624
rect 5740 27439 5780 27448
rect 5836 27152 5876 28960
rect 6124 28757 6164 29128
rect 6508 29168 6548 29287
rect 6508 29119 6548 29128
rect 6315 28916 6357 28925
rect 6315 28876 6316 28916
rect 6356 28876 6357 28916
rect 6315 28867 6357 28876
rect 6316 28782 6356 28867
rect 5931 28748 5973 28757
rect 5931 28708 5932 28748
rect 5972 28708 5973 28748
rect 5931 28699 5973 28708
rect 6123 28748 6165 28757
rect 6123 28708 6124 28748
rect 6164 28708 6165 28748
rect 6123 28699 6165 28708
rect 6507 28748 6549 28757
rect 6507 28708 6508 28748
rect 6548 28708 6549 28748
rect 6507 28699 6549 28708
rect 5644 25927 5684 25936
rect 5740 27112 5876 27152
rect 5548 25255 5588 25264
rect 5644 25304 5684 25313
rect 5740 25304 5780 27112
rect 5932 26816 5972 28699
rect 6219 28580 6261 28589
rect 6219 28540 6220 28580
rect 6260 28540 6261 28580
rect 6219 28531 6261 28540
rect 6123 28412 6165 28421
rect 6123 28372 6124 28412
rect 6164 28372 6165 28412
rect 6123 28363 6165 28372
rect 6124 28001 6164 28363
rect 6220 28085 6260 28531
rect 6315 28412 6357 28421
rect 6315 28372 6316 28412
rect 6356 28372 6357 28412
rect 6315 28363 6357 28372
rect 6219 28076 6261 28085
rect 6219 28036 6220 28076
rect 6260 28036 6261 28076
rect 6219 28027 6261 28036
rect 6123 27992 6165 28001
rect 6123 27952 6124 27992
rect 6164 27952 6165 27992
rect 6123 27943 6165 27952
rect 5932 26767 5972 26776
rect 6028 27656 6068 27665
rect 5836 26144 5876 26153
rect 5876 26104 5972 26144
rect 5836 26095 5876 26104
rect 5835 25892 5877 25901
rect 5835 25852 5836 25892
rect 5876 25852 5877 25892
rect 5835 25843 5877 25852
rect 5684 25264 5780 25304
rect 5644 25255 5684 25264
rect 5836 25136 5876 25843
rect 5836 25087 5876 25096
rect 5932 24968 5972 26104
rect 6028 25556 6068 27616
rect 6124 27656 6164 27665
rect 6124 27077 6164 27616
rect 6123 27068 6165 27077
rect 6123 27028 6124 27068
rect 6164 27028 6165 27068
rect 6123 27019 6165 27028
rect 6220 26825 6260 28027
rect 6219 26816 6261 26825
rect 6219 26776 6220 26816
rect 6260 26776 6261 26816
rect 6219 26767 6261 26776
rect 6124 26648 6164 26657
rect 6124 26480 6164 26608
rect 6316 26564 6356 28363
rect 6508 28328 6548 28699
rect 6700 28421 6740 29464
rect 6699 28412 6741 28421
rect 6699 28372 6700 28412
rect 6740 28372 6741 28412
rect 6699 28363 6741 28372
rect 6508 28279 6548 28288
rect 6699 28160 6741 28169
rect 6699 28120 6700 28160
rect 6740 28120 6741 28160
rect 6699 28111 6741 28120
rect 6700 28026 6740 28111
rect 6700 27665 6740 27750
rect 6796 27740 6836 32404
rect 6892 32276 6932 32285
rect 6892 31697 6932 32236
rect 6988 32201 7028 34168
rect 7084 33797 7124 34831
rect 7468 34712 7508 35162
rect 7852 35141 7892 35176
rect 8044 35216 8084 35225
rect 7851 35132 7893 35141
rect 7756 35092 7852 35132
rect 7892 35092 7893 35132
rect 7659 35048 7701 35057
rect 7659 35008 7660 35048
rect 7700 35008 7701 35048
rect 7659 34999 7701 35008
rect 7180 34672 7508 34712
rect 7180 34628 7220 34672
rect 7180 34579 7220 34588
rect 7660 34376 7700 34999
rect 7468 34355 7508 34364
rect 7371 34208 7413 34217
rect 7371 34168 7372 34208
rect 7412 34168 7413 34208
rect 7371 34159 7413 34168
rect 7372 34074 7412 34159
rect 7083 33788 7125 33797
rect 7083 33748 7084 33788
rect 7124 33748 7125 33788
rect 7083 33739 7125 33748
rect 7275 33788 7317 33797
rect 7275 33748 7276 33788
rect 7316 33748 7317 33788
rect 7275 33739 7317 33748
rect 7276 33704 7316 33739
rect 7276 33629 7316 33664
rect 7371 33704 7413 33713
rect 7371 33664 7372 33704
rect 7412 33664 7413 33704
rect 7371 33655 7413 33664
rect 7275 33620 7317 33629
rect 7275 33580 7276 33620
rect 7316 33580 7317 33620
rect 7275 33571 7317 33580
rect 7084 33452 7124 33461
rect 6987 32192 7029 32201
rect 6987 32152 6988 32192
rect 7028 32152 7029 32192
rect 6987 32143 7029 32152
rect 7084 32187 7124 33412
rect 7180 32864 7220 32873
rect 7180 32453 7220 32824
rect 7179 32444 7221 32453
rect 7179 32404 7180 32444
rect 7220 32404 7221 32444
rect 7179 32395 7221 32404
rect 7084 32138 7124 32147
rect 7083 32024 7125 32033
rect 7083 31984 7084 32024
rect 7124 31984 7125 32024
rect 7083 31975 7125 31984
rect 6987 31940 7029 31949
rect 6987 31900 6988 31940
rect 7028 31900 7029 31940
rect 6987 31891 7029 31900
rect 6891 31688 6933 31697
rect 6891 31648 6892 31688
rect 6932 31648 6933 31688
rect 6891 31639 6933 31648
rect 6891 31520 6933 31529
rect 6891 31480 6892 31520
rect 6932 31480 6933 31520
rect 6891 31471 6933 31480
rect 6892 28757 6932 31471
rect 6891 28748 6933 28757
rect 6891 28708 6892 28748
rect 6932 28708 6933 28748
rect 6891 28699 6933 28708
rect 6891 28412 6933 28421
rect 6891 28372 6892 28412
rect 6932 28372 6933 28412
rect 6891 28363 6933 28372
rect 6892 28278 6932 28363
rect 6891 27992 6933 28001
rect 6891 27952 6892 27992
rect 6932 27952 6933 27992
rect 6891 27943 6933 27952
rect 6796 27691 6836 27700
rect 6412 27656 6452 27665
rect 6412 27413 6452 27616
rect 6699 27656 6741 27665
rect 6699 27616 6700 27656
rect 6740 27616 6741 27656
rect 6699 27607 6741 27616
rect 6603 27488 6645 27497
rect 6603 27448 6604 27488
rect 6644 27448 6645 27488
rect 6603 27439 6645 27448
rect 6411 27404 6453 27413
rect 6411 27364 6412 27404
rect 6452 27364 6453 27404
rect 6411 27355 6453 27364
rect 6412 26984 6452 26993
rect 6604 26984 6644 27439
rect 6699 27404 6741 27413
rect 6699 27364 6700 27404
rect 6740 27364 6741 27404
rect 6699 27355 6741 27364
rect 6452 26944 6644 26984
rect 6412 26935 6452 26944
rect 6507 26816 6549 26825
rect 6507 26776 6508 26816
rect 6548 26776 6549 26816
rect 6507 26767 6549 26776
rect 6508 26573 6548 26767
rect 6507 26564 6549 26573
rect 6316 26524 6452 26564
rect 6124 26440 6356 26480
rect 6219 25556 6261 25565
rect 6028 25516 6164 25556
rect 6027 25388 6069 25397
rect 6027 25348 6028 25388
rect 6068 25348 6069 25388
rect 6027 25339 6069 25348
rect 6028 25254 6068 25339
rect 5836 24928 5972 24968
rect 5643 24884 5685 24893
rect 5643 24844 5644 24884
rect 5684 24844 5685 24884
rect 5643 24835 5685 24844
rect 5547 24632 5589 24641
rect 5547 24592 5548 24632
rect 5588 24592 5589 24632
rect 5547 24583 5589 24592
rect 5548 23792 5588 24583
rect 5548 23743 5588 23752
rect 5644 23204 5684 24835
rect 5836 24557 5876 24928
rect 6124 24893 6164 25516
rect 6219 25516 6220 25556
rect 6260 25516 6261 25556
rect 6219 25507 6261 25516
rect 6220 25422 6260 25507
rect 6123 24884 6165 24893
rect 6123 24844 6124 24884
rect 6164 24844 6165 24884
rect 6123 24835 6165 24844
rect 5931 24632 5973 24641
rect 5931 24592 5932 24632
rect 5972 24592 5973 24632
rect 6316 24632 6356 26440
rect 6412 25304 6452 26524
rect 6507 26524 6508 26564
rect 6548 26524 6549 26564
rect 6507 26515 6549 26524
rect 6604 26489 6644 26944
rect 6700 26816 6740 27355
rect 6795 27152 6837 27161
rect 6795 27112 6796 27152
rect 6836 27112 6837 27152
rect 6795 27103 6837 27112
rect 6700 26767 6740 26776
rect 6796 26816 6836 27103
rect 6796 26767 6836 26776
rect 6699 26564 6741 26573
rect 6699 26524 6700 26564
rect 6740 26524 6741 26564
rect 6699 26515 6741 26524
rect 6603 26480 6645 26489
rect 6603 26440 6604 26480
rect 6644 26440 6645 26480
rect 6603 26431 6645 26440
rect 6412 24809 6452 25264
rect 6700 24809 6740 26515
rect 6892 26153 6932 27943
rect 6891 26144 6933 26153
rect 6891 26104 6892 26144
rect 6932 26104 6933 26144
rect 6891 26095 6933 26104
rect 6988 24977 7028 31891
rect 7084 28580 7124 31975
rect 7372 31529 7412 33655
rect 7468 32780 7508 34315
rect 7564 34355 7604 34364
rect 7564 33797 7604 34315
rect 7563 33788 7605 33797
rect 7563 33748 7564 33788
rect 7604 33748 7605 33788
rect 7563 33739 7605 33748
rect 7563 33116 7605 33125
rect 7563 33076 7564 33116
rect 7604 33076 7605 33116
rect 7563 33067 7605 33076
rect 7564 32864 7604 33067
rect 7660 33041 7700 34336
rect 7756 34301 7796 35092
rect 7851 35083 7893 35092
rect 8044 35057 8084 35176
rect 8043 35048 8085 35057
rect 8043 35008 8044 35048
rect 8084 35008 8085 35048
rect 8043 34999 8085 35008
rect 7948 34964 7988 34973
rect 7852 34924 7948 34964
rect 7755 34292 7797 34301
rect 7755 34252 7756 34292
rect 7796 34252 7797 34292
rect 7755 34243 7797 34252
rect 7659 33032 7701 33041
rect 7659 32992 7660 33032
rect 7700 32992 7701 33032
rect 7659 32983 7701 32992
rect 7660 32864 7700 32873
rect 7564 32824 7660 32864
rect 7660 32815 7700 32824
rect 7755 32864 7797 32873
rect 7755 32824 7756 32864
rect 7796 32824 7797 32864
rect 7755 32815 7797 32824
rect 7468 32740 7604 32780
rect 7467 32612 7509 32621
rect 7467 32572 7468 32612
rect 7508 32572 7509 32612
rect 7564 32612 7604 32740
rect 7756 32730 7796 32815
rect 7564 32572 7796 32612
rect 7467 32563 7509 32572
rect 7468 32201 7508 32563
rect 7563 32444 7605 32453
rect 7563 32404 7564 32444
rect 7604 32404 7605 32444
rect 7563 32395 7605 32404
rect 7467 32192 7509 32201
rect 7467 32152 7468 32192
rect 7508 32152 7509 32192
rect 7467 32143 7509 32152
rect 7564 32192 7604 32395
rect 7564 32143 7604 32152
rect 7371 31520 7413 31529
rect 7371 31480 7372 31520
rect 7412 31480 7413 31520
rect 7371 31471 7413 31480
rect 7371 30764 7413 30773
rect 7371 30724 7372 30764
rect 7412 30724 7413 30764
rect 7371 30715 7413 30724
rect 7275 28748 7317 28757
rect 7275 28708 7276 28748
rect 7316 28708 7317 28748
rect 7275 28699 7317 28708
rect 7084 28531 7124 28540
rect 7276 28328 7316 28699
rect 7276 28279 7316 28288
rect 7083 28160 7125 28169
rect 7083 28120 7084 28160
rect 7124 28120 7125 28160
rect 7083 28111 7125 28120
rect 7084 27656 7124 28111
rect 7084 27607 7124 27616
rect 7180 27656 7220 27665
rect 7180 27161 7220 27616
rect 7275 27572 7317 27581
rect 7275 27532 7276 27572
rect 7316 27532 7317 27572
rect 7275 27523 7317 27532
rect 7179 27152 7221 27161
rect 7179 27112 7180 27152
rect 7220 27112 7221 27152
rect 7179 27103 7221 27112
rect 7276 26825 7316 27523
rect 7180 26816 7220 26825
rect 7180 26657 7220 26776
rect 7275 26816 7317 26825
rect 7275 26776 7276 26816
rect 7316 26776 7317 26816
rect 7275 26767 7317 26776
rect 7276 26682 7316 26767
rect 7179 26648 7221 26657
rect 7179 26608 7180 26648
rect 7220 26608 7221 26648
rect 7179 26599 7221 26608
rect 7179 26480 7221 26489
rect 7179 26440 7180 26480
rect 7220 26440 7221 26480
rect 7179 26431 7221 26440
rect 7083 26312 7125 26321
rect 7083 26272 7084 26312
rect 7124 26272 7125 26312
rect 7083 26263 7125 26272
rect 7084 26144 7124 26263
rect 7084 26095 7124 26104
rect 7180 25976 7220 26431
rect 7275 26228 7317 26237
rect 7275 26188 7276 26228
rect 7316 26188 7317 26228
rect 7275 26179 7317 26188
rect 7276 26094 7316 26179
rect 7180 25936 7316 25976
rect 7179 25220 7221 25229
rect 7179 25180 7180 25220
rect 7220 25180 7221 25220
rect 7179 25171 7221 25180
rect 7180 24977 7220 25171
rect 6987 24968 7029 24977
rect 6987 24928 6988 24968
rect 7028 24928 7029 24968
rect 6987 24919 7029 24928
rect 7179 24968 7221 24977
rect 7179 24928 7180 24968
rect 7220 24928 7221 24968
rect 7179 24919 7221 24928
rect 6411 24800 6453 24809
rect 6411 24760 6412 24800
rect 6452 24760 6453 24800
rect 6411 24751 6453 24760
rect 6699 24800 6741 24809
rect 6699 24760 6700 24800
rect 6740 24760 6741 24800
rect 6699 24751 6741 24760
rect 6987 24800 7029 24809
rect 6987 24760 6988 24800
rect 7028 24760 7029 24800
rect 6987 24751 7029 24760
rect 6412 24632 6452 24641
rect 6316 24592 6412 24632
rect 5931 24583 5973 24592
rect 6412 24583 6452 24592
rect 6508 24632 6548 24641
rect 5835 24548 5877 24557
rect 5835 24508 5836 24548
rect 5876 24508 5877 24548
rect 5835 24499 5877 24508
rect 5548 23164 5684 23204
rect 5740 23624 5780 23633
rect 5548 21197 5588 23164
rect 5740 23120 5780 23584
rect 5836 23456 5876 24499
rect 5932 24498 5972 24583
rect 6027 24380 6069 24389
rect 6027 24340 6028 24380
rect 6068 24340 6069 24380
rect 6027 24331 6069 24340
rect 6124 24380 6164 24389
rect 6028 23792 6068 24331
rect 6124 23969 6164 24340
rect 6123 23960 6165 23969
rect 6123 23920 6124 23960
rect 6164 23920 6165 23960
rect 6123 23911 6165 23920
rect 6124 23792 6164 23801
rect 6028 23752 6124 23792
rect 6124 23743 6164 23752
rect 6220 23792 6260 23801
rect 6508 23792 6548 24592
rect 6603 24632 6645 24641
rect 6603 24592 6604 24632
rect 6644 24592 6645 24632
rect 6603 24583 6645 24592
rect 6795 24632 6837 24641
rect 6892 24632 6932 24641
rect 6795 24592 6796 24632
rect 6836 24592 6892 24632
rect 6795 24583 6837 24592
rect 6892 24583 6932 24592
rect 6260 23752 6548 23792
rect 6604 23792 6644 24583
rect 6988 24548 7028 24751
rect 7179 24632 7221 24641
rect 7179 24592 7180 24632
rect 7220 24592 7221 24632
rect 7179 24583 7221 24592
rect 6988 24499 7028 24508
rect 6987 24380 7029 24389
rect 6987 24340 6988 24380
rect 7028 24340 7029 24380
rect 6987 24331 7029 24340
rect 6699 23876 6741 23885
rect 6699 23836 6700 23876
rect 6740 23836 6741 23876
rect 6699 23827 6741 23836
rect 6220 23743 6260 23752
rect 5836 23416 5972 23456
rect 5692 23110 5780 23120
rect 5732 23080 5780 23110
rect 5836 23204 5876 23213
rect 5692 23061 5732 23070
rect 5836 22961 5876 23164
rect 5835 22952 5877 22961
rect 5835 22912 5836 22952
rect 5876 22912 5877 22952
rect 5835 22903 5877 22912
rect 5547 21188 5589 21197
rect 5547 21148 5548 21188
rect 5588 21148 5589 21188
rect 5547 21139 5589 21148
rect 5644 20012 5684 20021
rect 5547 18752 5589 18761
rect 5547 18712 5548 18752
rect 5588 18712 5589 18752
rect 5547 18703 5589 18712
rect 5548 18584 5588 18703
rect 5548 17249 5588 18544
rect 5547 17240 5589 17249
rect 5547 17200 5548 17240
rect 5588 17200 5589 17240
rect 5547 17191 5589 17200
rect 5547 16232 5589 16241
rect 5547 16192 5548 16232
rect 5588 16192 5589 16232
rect 5547 16183 5589 16192
rect 5451 15728 5493 15737
rect 5451 15688 5452 15728
rect 5492 15688 5493 15728
rect 5451 15679 5493 15688
rect 5548 15569 5588 16183
rect 5067 15560 5109 15569
rect 5067 15520 5068 15560
rect 5108 15520 5109 15560
rect 5067 15511 5109 15520
rect 5452 15560 5492 15569
rect 5068 15426 5108 15511
rect 5259 15476 5301 15485
rect 5259 15436 5260 15476
rect 5300 15436 5301 15476
rect 5259 15427 5301 15436
rect 5260 15392 5300 15427
rect 5260 15341 5300 15352
rect 5452 15317 5492 15520
rect 5547 15560 5589 15569
rect 5547 15520 5548 15560
rect 5588 15520 5589 15560
rect 5547 15511 5589 15520
rect 5451 15308 5493 15317
rect 5451 15268 5452 15308
rect 5492 15268 5493 15308
rect 5451 15259 5493 15268
rect 5451 14972 5493 14981
rect 5451 14932 5452 14972
rect 5492 14932 5493 14972
rect 5451 14923 5493 14932
rect 5164 14888 5204 14897
rect 5204 14848 5396 14888
rect 5164 14839 5204 14848
rect 4972 14720 5012 14729
rect 4780 14680 4972 14720
rect 4780 14309 4820 14680
rect 4972 14671 5012 14680
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4779 14300 4821 14309
rect 4779 14260 4780 14300
rect 4820 14260 4821 14300
rect 4779 14251 4821 14260
rect 4875 14216 4917 14225
rect 4875 14176 4876 14216
rect 4916 14176 4917 14216
rect 4875 14167 4917 14176
rect 4780 14132 4820 14141
rect 4684 14092 4780 14132
rect 4780 11789 4820 14092
rect 4876 14048 4916 14167
rect 4876 13999 4916 14008
rect 5164 14048 5204 14057
rect 4875 13880 4917 13889
rect 4875 13840 4876 13880
rect 4916 13840 4917 13880
rect 4875 13831 4917 13840
rect 4876 13208 4916 13831
rect 4876 13159 4916 13168
rect 5164 13049 5204 14008
rect 5356 13964 5396 14848
rect 5452 14720 5492 14923
rect 5452 14671 5492 14680
rect 5548 14720 5588 14729
rect 5548 14393 5588 14680
rect 5547 14384 5589 14393
rect 5547 14344 5548 14384
rect 5588 14344 5589 14384
rect 5547 14335 5589 14344
rect 5644 14225 5684 19972
rect 5739 20012 5781 20021
rect 5739 19972 5740 20012
rect 5780 19972 5781 20012
rect 5739 19963 5781 19972
rect 5740 19878 5780 19963
rect 5739 19340 5781 19349
rect 5739 19300 5740 19340
rect 5780 19300 5781 19340
rect 5739 19291 5781 19300
rect 5740 19256 5780 19291
rect 5740 19205 5780 19216
rect 5739 19088 5781 19097
rect 5739 19048 5740 19088
rect 5780 19048 5781 19088
rect 5739 19039 5781 19048
rect 5740 17744 5780 19039
rect 5740 17501 5780 17704
rect 5739 17492 5781 17501
rect 5739 17452 5740 17492
rect 5780 17452 5781 17492
rect 5739 17443 5781 17452
rect 5740 17072 5780 17443
rect 5740 17023 5780 17032
rect 5739 16904 5781 16913
rect 5739 16864 5740 16904
rect 5780 16864 5781 16904
rect 5739 16855 5781 16864
rect 5643 14216 5685 14225
rect 5643 14176 5644 14216
rect 5684 14176 5685 14216
rect 5643 14167 5685 14176
rect 5548 14048 5588 14057
rect 5740 14048 5780 16855
rect 5836 16409 5876 22903
rect 5932 22784 5972 23416
rect 6027 23036 6069 23045
rect 6027 22996 6028 23036
rect 6068 22996 6069 23036
rect 6027 22987 6069 22996
rect 6028 22902 6068 22987
rect 6219 22868 6261 22877
rect 6219 22828 6220 22868
rect 6260 22828 6261 22868
rect 6219 22819 6261 22828
rect 5932 22744 6068 22784
rect 5931 22196 5973 22205
rect 5931 22156 5932 22196
rect 5972 22156 5973 22196
rect 5931 22147 5973 22156
rect 5932 20180 5972 22147
rect 6028 21701 6068 22744
rect 6220 22734 6260 22819
rect 6219 22280 6261 22289
rect 6219 22240 6220 22280
rect 6260 22240 6261 22280
rect 6219 22231 6261 22240
rect 6220 22146 6260 22231
rect 6027 21692 6069 21701
rect 6027 21652 6028 21692
rect 6068 21652 6069 21692
rect 6027 21643 6069 21652
rect 6123 21608 6165 21617
rect 6123 21568 6124 21608
rect 6164 21568 6165 21608
rect 6123 21559 6165 21568
rect 6220 21608 6260 21617
rect 6316 21608 6356 23752
rect 6604 23633 6644 23752
rect 6603 23624 6645 23633
rect 6603 23584 6604 23624
rect 6644 23584 6645 23624
rect 6603 23575 6645 23584
rect 6603 23288 6645 23297
rect 6603 23248 6604 23288
rect 6644 23248 6645 23288
rect 6603 23239 6645 23248
rect 6604 23154 6644 23239
rect 6411 23036 6453 23045
rect 6411 22996 6412 23036
rect 6452 22996 6453 23036
rect 6411 22987 6453 22996
rect 6412 22902 6452 22987
rect 6700 22457 6740 23827
rect 6988 22868 7028 24331
rect 7083 23792 7125 23801
rect 7083 23752 7084 23792
rect 7124 23752 7125 23792
rect 7083 23743 7125 23752
rect 7180 23792 7220 24583
rect 7276 24389 7316 25936
rect 7275 24380 7317 24389
rect 7275 24340 7276 24380
rect 7316 24340 7317 24380
rect 7275 24331 7317 24340
rect 7372 24053 7412 30715
rect 7468 29765 7508 32143
rect 7563 32024 7605 32033
rect 7563 31984 7564 32024
rect 7604 31984 7605 32024
rect 7563 31975 7605 31984
rect 7467 29756 7509 29765
rect 7467 29716 7468 29756
rect 7508 29716 7509 29756
rect 7467 29707 7509 29716
rect 7564 29093 7604 31975
rect 7659 31352 7701 31361
rect 7659 31312 7660 31352
rect 7700 31312 7701 31352
rect 7659 31303 7701 31312
rect 7563 29084 7605 29093
rect 7563 29044 7564 29084
rect 7604 29044 7605 29084
rect 7563 29035 7605 29044
rect 7467 27992 7509 28001
rect 7467 27952 7468 27992
rect 7508 27952 7509 27992
rect 7467 27943 7509 27952
rect 7468 26489 7508 27943
rect 7660 27824 7700 31303
rect 7756 31016 7796 32572
rect 7852 31529 7892 34924
rect 7948 34915 7988 34924
rect 8140 34796 8180 36427
rect 8236 36317 8276 36604
rect 8235 36308 8277 36317
rect 8235 36268 8236 36308
rect 8276 36268 8277 36308
rect 8235 36259 8277 36268
rect 8235 35888 8277 35897
rect 8235 35848 8236 35888
rect 8276 35848 8277 35888
rect 8235 35839 8277 35848
rect 8332 35888 8372 35897
rect 7948 34756 8180 34796
rect 8236 35216 8276 35839
rect 8332 35561 8372 35848
rect 8331 35552 8373 35561
rect 8331 35512 8332 35552
rect 8372 35512 8373 35552
rect 8331 35503 8373 35512
rect 7948 34376 7988 34756
rect 7948 34327 7988 34336
rect 8043 34376 8085 34385
rect 8043 34336 8044 34376
rect 8084 34336 8085 34376
rect 8043 34327 8085 34336
rect 8044 34242 8084 34327
rect 8139 34292 8181 34301
rect 8139 34252 8140 34292
rect 8180 34252 8181 34292
rect 8139 34243 8181 34252
rect 8043 33116 8085 33125
rect 8043 33076 8044 33116
rect 8084 33076 8085 33116
rect 8043 33067 8085 33076
rect 7947 32948 7989 32957
rect 7947 32908 7948 32948
rect 7988 32908 7989 32948
rect 7947 32899 7989 32908
rect 7948 31604 7988 32899
rect 8044 32192 8084 33067
rect 8140 32864 8180 34243
rect 8236 33713 8276 35176
rect 8428 34628 8468 39376
rect 8524 38912 8564 40207
rect 8620 39752 8660 40972
rect 8715 40928 8757 40937
rect 8715 40888 8716 40928
rect 8756 40888 8757 40928
rect 8715 40879 8757 40888
rect 8716 40433 8756 40879
rect 8715 40424 8757 40433
rect 8715 40384 8716 40424
rect 8756 40384 8757 40424
rect 8715 40375 8757 40384
rect 8716 40290 8756 40375
rect 8908 39929 8948 41224
rect 8907 39920 8949 39929
rect 8907 39880 8908 39920
rect 8948 39880 8949 39920
rect 8907 39871 8949 39880
rect 9100 39836 9140 42928
rect 9292 41609 9332 42928
rect 9387 41936 9429 41945
rect 9387 41896 9388 41936
rect 9428 41896 9429 41936
rect 9387 41887 9429 41896
rect 9291 41600 9333 41609
rect 9291 41560 9292 41600
rect 9332 41560 9333 41600
rect 9291 41551 9333 41560
rect 9100 39796 9332 39836
rect 8716 39752 8756 39761
rect 8620 39712 8716 39752
rect 8716 39703 8756 39712
rect 8812 39752 8852 39761
rect 8812 39164 8852 39712
rect 9292 39752 9332 39796
rect 9196 39668 9236 39677
rect 8716 39124 8852 39164
rect 9100 39628 9196 39668
rect 8620 38912 8660 38921
rect 8524 38872 8620 38912
rect 8620 38863 8660 38872
rect 8716 38912 8756 39124
rect 8716 38576 8756 38872
rect 8907 38912 8949 38921
rect 9100 38912 9140 39628
rect 9196 39619 9236 39628
rect 8907 38872 8908 38912
rect 8948 38872 8949 38912
rect 8907 38863 8949 38872
rect 9004 38872 9100 38912
rect 8620 38536 8756 38576
rect 8524 37400 8564 37409
rect 8524 36485 8564 37360
rect 8620 37325 8660 38536
rect 8715 38408 8757 38417
rect 8715 38368 8716 38408
rect 8756 38368 8757 38408
rect 8715 38359 8757 38368
rect 8716 38249 8756 38359
rect 8715 38240 8757 38249
rect 8715 38200 8716 38240
rect 8756 38200 8757 38240
rect 8715 38191 8757 38200
rect 8908 38240 8948 38863
rect 8908 38191 8948 38200
rect 8619 37316 8661 37325
rect 8619 37276 8620 37316
rect 8660 37276 8661 37316
rect 8619 37267 8661 37276
rect 8716 36896 8756 38191
rect 8907 38072 8949 38081
rect 8907 38032 8908 38072
rect 8948 38032 8949 38072
rect 8907 38023 8949 38032
rect 8811 37400 8853 37409
rect 8811 37360 8812 37400
rect 8852 37360 8853 37400
rect 8811 37351 8853 37360
rect 8812 36989 8852 37351
rect 8811 36980 8853 36989
rect 8811 36940 8812 36980
rect 8852 36940 8853 36980
rect 8811 36931 8853 36940
rect 8620 36856 8756 36896
rect 8523 36476 8565 36485
rect 8523 36436 8524 36476
rect 8564 36436 8565 36476
rect 8523 36427 8565 36436
rect 8523 36224 8565 36233
rect 8523 36184 8524 36224
rect 8564 36184 8565 36224
rect 8523 36175 8565 36184
rect 8524 35981 8564 36175
rect 8523 35972 8565 35981
rect 8523 35932 8524 35972
rect 8564 35932 8565 35972
rect 8523 35923 8565 35932
rect 8332 34588 8468 34628
rect 8235 33704 8277 33713
rect 8235 33664 8236 33704
rect 8276 33664 8277 33704
rect 8235 33655 8277 33664
rect 8235 33452 8277 33461
rect 8235 33412 8236 33452
rect 8276 33412 8277 33452
rect 8235 33403 8277 33412
rect 8140 32537 8180 32824
rect 8236 32864 8276 33403
rect 8236 32815 8276 32824
rect 8235 32696 8277 32705
rect 8235 32656 8236 32696
rect 8276 32656 8277 32696
rect 8235 32647 8277 32656
rect 8139 32528 8181 32537
rect 8139 32488 8140 32528
rect 8180 32488 8181 32528
rect 8139 32479 8181 32488
rect 8044 32143 8084 32152
rect 8140 32108 8180 32117
rect 8140 31949 8180 32068
rect 8139 31940 8181 31949
rect 8139 31900 8140 31940
rect 8180 31900 8181 31940
rect 8139 31891 8181 31900
rect 7948 31564 8084 31604
rect 7851 31520 7893 31529
rect 7851 31480 7852 31520
rect 7892 31480 7893 31520
rect 7851 31471 7893 31480
rect 8044 31520 8084 31564
rect 7852 31352 7892 31363
rect 7852 31277 7892 31312
rect 7851 31268 7893 31277
rect 7851 31228 7852 31268
rect 7892 31228 7893 31268
rect 7851 31219 7893 31228
rect 7756 30976 7988 31016
rect 7755 30680 7797 30689
rect 7755 30640 7756 30680
rect 7796 30640 7797 30680
rect 7755 30631 7797 30640
rect 7756 29933 7796 30631
rect 7755 29924 7797 29933
rect 7755 29884 7756 29924
rect 7796 29884 7797 29924
rect 7755 29875 7797 29884
rect 7852 29429 7892 30976
rect 7948 30848 7988 30976
rect 8044 30848 8084 31480
rect 8236 31352 8276 32647
rect 8332 32033 8372 34588
rect 8427 34460 8469 34469
rect 8427 34420 8428 34460
rect 8468 34420 8469 34460
rect 8427 34411 8469 34420
rect 8524 34460 8564 35923
rect 8428 34326 8468 34411
rect 8524 33965 8564 34420
rect 8523 33956 8565 33965
rect 8523 33916 8524 33956
rect 8564 33916 8565 33956
rect 8523 33907 8565 33916
rect 8523 33704 8565 33713
rect 8523 33664 8524 33704
rect 8564 33664 8565 33704
rect 8523 33655 8565 33664
rect 8524 33570 8564 33655
rect 8427 33200 8469 33209
rect 8427 33160 8428 33200
rect 8468 33160 8469 33200
rect 8427 33151 8469 33160
rect 8331 32024 8373 32033
rect 8331 31984 8332 32024
rect 8372 31984 8373 32024
rect 8331 31975 8373 31984
rect 8428 31856 8468 33151
rect 8620 32873 8660 36856
rect 8716 36728 8756 36737
rect 8716 36485 8756 36688
rect 8812 36653 8852 36931
rect 8811 36644 8853 36653
rect 8811 36604 8812 36644
rect 8852 36604 8853 36644
rect 8811 36595 8853 36604
rect 8908 36569 8948 38023
rect 9004 37820 9044 38872
rect 9100 38863 9140 38872
rect 9196 38996 9236 39005
rect 9292 38996 9332 39712
rect 9236 38956 9332 38996
rect 9196 38165 9236 38956
rect 9291 38744 9333 38753
rect 9291 38704 9292 38744
rect 9332 38704 9333 38744
rect 9291 38695 9333 38704
rect 9292 38240 9332 38695
rect 9292 38191 9332 38200
rect 9195 38156 9237 38165
rect 9195 38116 9196 38156
rect 9236 38116 9237 38156
rect 9195 38107 9237 38116
rect 9100 37988 9140 37997
rect 9140 37948 9332 37988
rect 9100 37939 9140 37948
rect 9004 37780 9140 37820
rect 9003 37652 9045 37661
rect 9003 37612 9004 37652
rect 9044 37612 9045 37652
rect 9003 37603 9045 37612
rect 9004 37414 9044 37603
rect 9100 37493 9140 37780
rect 9099 37484 9141 37493
rect 9099 37444 9100 37484
rect 9140 37444 9141 37484
rect 9099 37435 9141 37444
rect 9004 37365 9044 37374
rect 9100 37316 9140 37435
rect 9004 37276 9140 37316
rect 9004 36821 9044 37276
rect 9196 37232 9236 37241
rect 9100 37192 9196 37232
rect 9003 36812 9045 36821
rect 9003 36772 9004 36812
rect 9044 36772 9045 36812
rect 9003 36763 9045 36772
rect 8907 36560 8949 36569
rect 8907 36520 8908 36560
rect 8948 36520 8949 36560
rect 8907 36511 8949 36520
rect 8715 36476 8757 36485
rect 8715 36436 8716 36476
rect 8756 36436 8757 36476
rect 8715 36427 8757 36436
rect 8716 35561 8756 36427
rect 8812 35893 8852 35902
rect 8812 35813 8852 35853
rect 8811 35804 8853 35813
rect 8811 35764 8812 35804
rect 8852 35764 8853 35804
rect 8811 35755 8853 35764
rect 9004 35720 9044 35729
rect 8715 35552 8757 35561
rect 8715 35512 8716 35552
rect 8756 35512 8757 35552
rect 8715 35503 8757 35512
rect 9004 35225 9044 35680
rect 8811 35216 8853 35225
rect 8811 35176 8812 35216
rect 8852 35176 8853 35216
rect 8811 35167 8853 35176
rect 9003 35216 9045 35225
rect 9003 35176 9004 35216
rect 9044 35176 9045 35216
rect 9003 35167 9045 35176
rect 8812 35057 8852 35167
rect 8811 35048 8853 35057
rect 8811 35008 8812 35048
rect 8852 35008 8853 35048
rect 8811 34999 8853 35008
rect 9004 34628 9044 35167
rect 9100 34721 9140 37192
rect 9196 37183 9236 37192
rect 9292 37064 9332 37948
rect 9388 37661 9428 41887
rect 9387 37652 9429 37661
rect 9387 37612 9388 37652
rect 9428 37612 9429 37652
rect 9387 37603 9429 37612
rect 9387 37484 9429 37493
rect 9387 37444 9388 37484
rect 9428 37444 9429 37484
rect 9387 37435 9429 37444
rect 9388 37350 9428 37435
rect 9387 37148 9429 37157
rect 9387 37108 9388 37148
rect 9428 37108 9429 37148
rect 9387 37099 9429 37108
rect 9196 37024 9332 37064
rect 9196 36723 9236 37024
rect 9388 36896 9428 37099
rect 9388 36847 9428 36856
rect 9196 36674 9236 36683
rect 9291 36560 9333 36569
rect 9291 36520 9292 36560
rect 9332 36520 9333 36560
rect 9291 36511 9333 36520
rect 9195 36140 9237 36149
rect 9195 36100 9196 36140
rect 9236 36100 9237 36140
rect 9195 36091 9237 36100
rect 9196 35972 9236 36091
rect 9196 35923 9236 35932
rect 9099 34712 9141 34721
rect 9099 34672 9100 34712
rect 9140 34672 9141 34712
rect 9099 34663 9141 34672
rect 8716 34588 9044 34628
rect 8619 32864 8661 32873
rect 8619 32824 8620 32864
rect 8660 32824 8661 32864
rect 8619 32815 8661 32824
rect 8716 32864 8756 34588
rect 9004 34376 9044 34385
rect 9044 34336 9140 34376
rect 9004 34327 9044 34336
rect 8811 34208 8853 34217
rect 8811 34168 8812 34208
rect 8852 34168 8853 34208
rect 8811 34159 8853 34168
rect 8812 33032 8852 34159
rect 8908 33704 8948 33713
rect 8908 33377 8948 33664
rect 8907 33368 8949 33377
rect 8907 33328 8908 33368
rect 8948 33328 8949 33368
rect 8907 33319 8949 33328
rect 8812 32992 8948 33032
rect 8716 32815 8756 32824
rect 8811 32864 8853 32873
rect 8811 32824 8812 32864
rect 8852 32824 8853 32864
rect 8811 32815 8853 32824
rect 8812 32730 8852 32815
rect 8524 32696 8564 32705
rect 8564 32656 8756 32696
rect 8524 32647 8564 32656
rect 8523 32528 8565 32537
rect 8523 32488 8524 32528
rect 8564 32488 8565 32528
rect 8523 32479 8565 32488
rect 8524 32201 8564 32479
rect 8619 32276 8661 32285
rect 8619 32236 8620 32276
rect 8660 32236 8661 32276
rect 8619 32227 8661 32236
rect 8523 32192 8565 32201
rect 8523 32152 8524 32192
rect 8564 32152 8565 32192
rect 8523 32143 8565 32152
rect 8620 32192 8660 32227
rect 8524 32058 8564 32143
rect 8620 32141 8660 32152
rect 8332 31816 8468 31856
rect 8332 31436 8372 31816
rect 8427 31688 8469 31697
rect 8427 31648 8428 31688
rect 8468 31648 8469 31688
rect 8427 31639 8469 31648
rect 8428 31520 8468 31639
rect 8428 31471 8468 31480
rect 8332 31387 8372 31396
rect 8524 31436 8564 31445
rect 8236 31303 8276 31312
rect 8044 30808 8372 30848
rect 7948 30799 7988 30808
rect 8043 30428 8085 30437
rect 8043 30388 8044 30428
rect 8084 30388 8085 30428
rect 8043 30379 8085 30388
rect 7947 29924 7989 29933
rect 7947 29884 7948 29924
rect 7988 29884 7989 29924
rect 7947 29875 7989 29884
rect 7948 29840 7988 29875
rect 7948 29789 7988 29800
rect 7851 29420 7893 29429
rect 7851 29380 7852 29420
rect 7892 29380 7893 29420
rect 7851 29371 7893 29380
rect 7756 29168 7796 29177
rect 7756 28841 7796 29128
rect 7851 29084 7893 29093
rect 7851 29044 7852 29084
rect 7892 29044 7893 29084
rect 7851 29035 7893 29044
rect 7755 28832 7797 28841
rect 7755 28792 7756 28832
rect 7796 28792 7797 28832
rect 7755 28783 7797 28792
rect 7756 28337 7796 28783
rect 7755 28328 7797 28337
rect 7755 28288 7756 28328
rect 7796 28288 7797 28328
rect 7755 28279 7797 28288
rect 7660 27784 7796 27824
rect 7660 27581 7700 27666
rect 7564 27572 7604 27581
rect 7564 26657 7604 27532
rect 7659 27572 7701 27581
rect 7659 27532 7660 27572
rect 7700 27532 7701 27572
rect 7659 27523 7701 27532
rect 7756 27404 7796 27784
rect 7660 27364 7796 27404
rect 7563 26648 7605 26657
rect 7563 26608 7564 26648
rect 7604 26608 7605 26648
rect 7563 26599 7605 26608
rect 7467 26480 7509 26489
rect 7467 26440 7468 26480
rect 7508 26440 7509 26480
rect 7467 26431 7509 26440
rect 7467 26144 7509 26153
rect 7467 26104 7468 26144
rect 7508 26104 7509 26144
rect 7467 26095 7509 26104
rect 7468 24809 7508 26095
rect 7660 25901 7700 27364
rect 7755 26984 7797 26993
rect 7755 26944 7756 26984
rect 7796 26944 7797 26984
rect 7755 26935 7797 26944
rect 7756 26825 7796 26935
rect 7755 26816 7797 26825
rect 7755 26776 7756 26816
rect 7796 26776 7797 26816
rect 7755 26767 7797 26776
rect 7756 26682 7796 26767
rect 7852 26573 7892 29035
rect 7947 28916 7989 28925
rect 7947 28876 7948 28916
rect 7988 28876 7989 28916
rect 7947 28867 7989 28876
rect 7948 28782 7988 28867
rect 7947 28328 7989 28337
rect 7947 28288 7948 28328
rect 7988 28288 7989 28328
rect 7947 28279 7989 28288
rect 7851 26564 7893 26573
rect 7851 26524 7852 26564
rect 7892 26524 7893 26564
rect 7851 26515 7893 26524
rect 7659 25892 7701 25901
rect 7659 25852 7660 25892
rect 7700 25852 7701 25892
rect 7659 25843 7701 25852
rect 7563 25724 7605 25733
rect 7563 25684 7564 25724
rect 7604 25684 7605 25724
rect 7563 25675 7605 25684
rect 7467 24800 7509 24809
rect 7467 24760 7468 24800
rect 7508 24760 7509 24800
rect 7467 24751 7509 24760
rect 7467 24632 7509 24641
rect 7467 24592 7468 24632
rect 7508 24592 7509 24632
rect 7467 24583 7509 24592
rect 7468 24498 7508 24583
rect 7467 24212 7509 24221
rect 7467 24172 7468 24212
rect 7508 24172 7509 24212
rect 7467 24163 7509 24172
rect 7371 24044 7413 24053
rect 7371 24004 7372 24044
rect 7412 24004 7413 24044
rect 7371 23995 7413 24004
rect 7220 23752 7316 23792
rect 7180 23743 7220 23752
rect 7084 23120 7124 23743
rect 7179 23624 7221 23633
rect 7179 23584 7180 23624
rect 7220 23584 7221 23624
rect 7179 23575 7221 23584
rect 7084 23071 7124 23080
rect 6988 22828 7124 22868
rect 6699 22448 6741 22457
rect 6699 22408 6700 22448
rect 6740 22408 6741 22448
rect 6699 22399 6741 22408
rect 6987 22448 7029 22457
rect 6987 22408 6988 22448
rect 7028 22408 7029 22448
rect 6987 22399 7029 22408
rect 6700 22280 6740 22289
rect 6411 22112 6453 22121
rect 6411 22072 6412 22112
rect 6452 22072 6453 22112
rect 6411 22063 6453 22072
rect 6412 21978 6452 22063
rect 6507 21944 6549 21953
rect 6507 21904 6508 21944
rect 6548 21904 6549 21944
rect 6507 21895 6549 21904
rect 6411 21860 6453 21869
rect 6411 21820 6412 21860
rect 6452 21820 6453 21860
rect 6411 21811 6453 21820
rect 6412 21608 6452 21811
rect 6260 21568 6452 21608
rect 6220 21559 6260 21568
rect 6124 21474 6164 21559
rect 6315 21356 6357 21365
rect 6315 21316 6316 21356
rect 6356 21316 6357 21356
rect 6315 21307 6357 21316
rect 6027 20852 6069 20861
rect 6027 20812 6028 20852
rect 6068 20812 6069 20852
rect 6027 20803 6069 20812
rect 6219 20852 6261 20861
rect 6219 20812 6220 20852
rect 6260 20812 6261 20852
rect 6219 20803 6261 20812
rect 6028 20441 6068 20803
rect 6123 20684 6165 20693
rect 6123 20644 6124 20684
rect 6164 20644 6165 20684
rect 6123 20635 6165 20644
rect 6027 20432 6069 20441
rect 6027 20392 6028 20432
rect 6068 20392 6069 20432
rect 6027 20383 6069 20392
rect 5932 20140 6068 20180
rect 5931 17660 5973 17669
rect 5931 17620 5932 17660
rect 5972 17620 5973 17660
rect 5931 17611 5973 17620
rect 5932 17526 5972 17611
rect 6028 17417 6068 20140
rect 6124 19433 6164 20635
rect 6220 20096 6260 20803
rect 6220 20047 6260 20056
rect 6123 19424 6165 19433
rect 6123 19384 6124 19424
rect 6164 19384 6165 19424
rect 6123 19375 6165 19384
rect 6124 18929 6164 19375
rect 6123 18920 6165 18929
rect 6123 18880 6124 18920
rect 6164 18880 6165 18920
rect 6123 18871 6165 18880
rect 6316 18005 6356 21307
rect 6315 17996 6357 18005
rect 6315 17956 6316 17996
rect 6356 17956 6357 17996
rect 6315 17947 6357 17956
rect 6220 17744 6260 17753
rect 6027 17408 6069 17417
rect 6027 17368 6028 17408
rect 6068 17368 6069 17408
rect 6027 17359 6069 17368
rect 5932 17240 5972 17249
rect 6220 17240 6260 17704
rect 6316 17744 6356 17753
rect 6412 17744 6452 21568
rect 6356 17704 6452 17744
rect 6316 17695 6356 17704
rect 5972 17200 6260 17240
rect 5932 17191 5972 17200
rect 6123 17072 6165 17081
rect 6123 17032 6124 17072
rect 6164 17032 6165 17072
rect 6123 17023 6165 17032
rect 6220 17072 6260 17200
rect 6315 17156 6357 17165
rect 6315 17116 6316 17156
rect 6356 17116 6357 17156
rect 6315 17107 6357 17116
rect 6220 17023 6260 17032
rect 6316 17072 6356 17107
rect 5835 16400 5877 16409
rect 5835 16360 5836 16400
rect 5876 16360 5877 16400
rect 5835 16351 5877 16360
rect 5835 16232 5877 16241
rect 5835 16192 5836 16232
rect 5876 16192 5877 16232
rect 5835 16183 5877 16192
rect 6027 16232 6069 16241
rect 6027 16192 6028 16232
rect 6068 16192 6069 16232
rect 6027 16183 6069 16192
rect 5836 16098 5876 16183
rect 6028 16064 6068 16183
rect 5931 15728 5973 15737
rect 5931 15688 5932 15728
rect 5972 15688 5973 15728
rect 5931 15679 5973 15688
rect 5835 14720 5877 14729
rect 5835 14680 5836 14720
rect 5876 14680 5877 14720
rect 5835 14671 5877 14680
rect 5836 14586 5876 14671
rect 5588 14008 5780 14048
rect 5932 14048 5972 15679
rect 6028 14729 6068 16024
rect 6124 15812 6164 17023
rect 6316 17021 6356 17032
rect 6412 16409 6452 17704
rect 6508 16661 6548 21895
rect 6700 21692 6740 22240
rect 6796 22280 6836 22289
rect 6796 21869 6836 22240
rect 6891 22280 6933 22289
rect 6891 22240 6892 22280
rect 6932 22240 6933 22280
rect 6891 22231 6933 22240
rect 6795 21860 6837 21869
rect 6795 21820 6796 21860
rect 6836 21820 6837 21860
rect 6795 21811 6837 21820
rect 6700 21652 6836 21692
rect 6603 21608 6645 21617
rect 6603 21568 6604 21608
rect 6644 21568 6645 21608
rect 6603 21559 6645 21568
rect 6604 21474 6644 21559
rect 6699 21524 6741 21533
rect 6699 21484 6700 21524
rect 6740 21484 6741 21524
rect 6699 21475 6741 21484
rect 6603 21188 6645 21197
rect 6603 21148 6604 21188
rect 6644 21148 6645 21188
rect 6603 21139 6645 21148
rect 6604 20768 6644 21139
rect 6507 16652 6549 16661
rect 6507 16612 6508 16652
rect 6548 16612 6549 16652
rect 6507 16603 6549 16612
rect 6604 16577 6644 20728
rect 6700 20180 6740 21475
rect 6796 21020 6836 21652
rect 6892 21197 6932 22231
rect 6988 21533 7028 22399
rect 6987 21524 7029 21533
rect 6987 21484 6988 21524
rect 7028 21484 7029 21524
rect 6987 21475 7029 21484
rect 7084 21365 7124 22828
rect 7180 22280 7220 23575
rect 7276 22709 7316 23752
rect 7468 23129 7508 24163
rect 7564 23633 7604 25675
rect 7660 25304 7700 25313
rect 7948 25304 7988 28279
rect 8044 26069 8084 30379
rect 8332 30101 8372 30808
rect 8524 30353 8564 31396
rect 8619 31352 8661 31361
rect 8619 31312 8620 31352
rect 8660 31312 8661 31352
rect 8619 31303 8661 31312
rect 8620 31218 8660 31303
rect 8619 30428 8661 30437
rect 8619 30388 8620 30428
rect 8660 30388 8661 30428
rect 8619 30379 8661 30388
rect 8523 30344 8565 30353
rect 8523 30304 8524 30344
rect 8564 30304 8565 30344
rect 8523 30295 8565 30304
rect 8620 30294 8660 30379
rect 8331 30092 8373 30101
rect 8331 30052 8332 30092
rect 8372 30052 8373 30092
rect 8331 30043 8373 30052
rect 8140 30008 8180 30017
rect 8235 30008 8277 30017
rect 8180 29968 8236 30008
rect 8276 29968 8277 30008
rect 8140 29959 8180 29968
rect 8235 29959 8277 29968
rect 8332 29840 8372 30043
rect 8524 29840 8564 29849
rect 8332 29800 8524 29840
rect 8524 29791 8564 29800
rect 8716 29672 8756 32656
rect 8811 31520 8853 31529
rect 8811 31480 8812 31520
rect 8852 31480 8853 31520
rect 8811 31471 8853 31480
rect 8812 31386 8852 31471
rect 8811 30680 8853 30689
rect 8811 30640 8812 30680
rect 8852 30640 8853 30680
rect 8811 30631 8853 30640
rect 8812 30269 8852 30631
rect 8811 30260 8853 30269
rect 8811 30220 8812 30260
rect 8852 30220 8853 30260
rect 8811 30211 8853 30220
rect 8812 30017 8852 30211
rect 8811 30008 8853 30017
rect 8811 29968 8812 30008
rect 8852 29968 8853 30008
rect 8811 29959 8853 29968
rect 8908 29933 8948 32992
rect 9004 32864 9044 32873
rect 9004 32621 9044 32824
rect 9003 32612 9045 32621
rect 9003 32572 9004 32612
rect 9044 32572 9045 32612
rect 9003 32563 9045 32572
rect 9100 32360 9140 34336
rect 9292 33881 9332 36511
rect 9388 35720 9428 35729
rect 9388 35561 9428 35680
rect 9387 35552 9429 35561
rect 9387 35512 9388 35552
rect 9428 35512 9429 35552
rect 9387 35503 9429 35512
rect 9484 35384 9524 42928
rect 9676 42617 9716 42928
rect 9675 42608 9717 42617
rect 9675 42568 9676 42608
rect 9716 42568 9717 42608
rect 9675 42559 9717 42568
rect 9868 41609 9908 42928
rect 9867 41600 9909 41609
rect 9867 41560 9868 41600
rect 9908 41560 9909 41600
rect 9867 41551 9909 41560
rect 9963 40928 10005 40937
rect 9963 40888 9964 40928
rect 10004 40888 10005 40928
rect 9963 40879 10005 40888
rect 9964 40424 10004 40879
rect 9964 40375 10004 40384
rect 10060 40349 10100 42928
rect 10252 41609 10292 42928
rect 10444 41852 10484 42928
rect 10636 42029 10676 42928
rect 10635 42020 10677 42029
rect 10635 41980 10636 42020
rect 10676 41980 10677 42020
rect 10635 41971 10677 41980
rect 10444 41812 10676 41852
rect 10443 41684 10485 41693
rect 10443 41644 10444 41684
rect 10484 41644 10485 41684
rect 10443 41635 10485 41644
rect 10251 41600 10293 41609
rect 10251 41560 10252 41600
rect 10292 41560 10293 41600
rect 10251 41551 10293 41560
rect 10156 41264 10196 41273
rect 10156 40937 10196 41224
rect 10348 41012 10388 41021
rect 10252 40972 10348 41012
rect 10155 40928 10197 40937
rect 10155 40888 10156 40928
rect 10196 40888 10197 40928
rect 10155 40879 10197 40888
rect 10059 40340 10101 40349
rect 10059 40300 10060 40340
rect 10100 40300 10101 40340
rect 10059 40291 10101 40300
rect 10156 40256 10196 40265
rect 9772 39752 9812 39761
rect 9772 38921 9812 39712
rect 10156 38926 10196 40216
rect 10252 39747 10292 40972
rect 10348 40963 10388 40972
rect 10444 40844 10484 41635
rect 10348 40804 10484 40844
rect 10540 41012 10580 41021
rect 10348 40676 10388 40804
rect 10540 40760 10580 40972
rect 10348 40627 10388 40636
rect 10444 40720 10580 40760
rect 10444 40424 10484 40720
rect 10539 40592 10581 40601
rect 10539 40552 10540 40592
rect 10580 40552 10581 40592
rect 10539 40543 10581 40552
rect 10540 40508 10580 40543
rect 10540 40457 10580 40468
rect 10252 39698 10292 39707
rect 10348 40384 10484 40424
rect 10348 39341 10388 40384
rect 10443 40256 10485 40265
rect 10443 40216 10444 40256
rect 10484 40216 10485 40256
rect 10443 40207 10485 40216
rect 10444 39836 10484 40207
rect 10636 40004 10676 41812
rect 10732 41264 10772 41273
rect 10732 40937 10772 41224
rect 10731 40928 10773 40937
rect 10731 40888 10732 40928
rect 10772 40888 10773 40928
rect 10731 40879 10773 40888
rect 10731 40424 10773 40433
rect 10731 40384 10732 40424
rect 10772 40384 10773 40424
rect 10731 40375 10773 40384
rect 10732 40290 10772 40375
rect 10347 39332 10389 39341
rect 10347 39292 10348 39332
rect 10388 39292 10389 39332
rect 10347 39283 10389 39292
rect 9676 38912 9716 38921
rect 9771 38912 9813 38921
rect 9716 38872 9772 38912
rect 9812 38872 9813 38912
rect 10156 38877 10196 38886
rect 9676 38585 9716 38872
rect 9771 38863 9813 38872
rect 9772 38778 9812 38863
rect 10347 38828 10389 38837
rect 10347 38788 10348 38828
rect 10388 38788 10389 38828
rect 10347 38779 10389 38788
rect 10348 38694 10388 38779
rect 9675 38576 9717 38585
rect 9675 38536 9676 38576
rect 9716 38536 9717 38576
rect 9675 38527 9717 38536
rect 10347 38576 10389 38585
rect 10347 38536 10348 38576
rect 10388 38536 10389 38576
rect 10347 38527 10389 38536
rect 9963 37904 10005 37913
rect 9963 37864 9964 37904
rect 10004 37864 10005 37904
rect 9963 37855 10005 37864
rect 9579 37652 9621 37661
rect 9579 37612 9580 37652
rect 9620 37612 9621 37652
rect 9579 37603 9621 37612
rect 9964 37652 10004 37855
rect 10059 37736 10101 37745
rect 10059 37696 10060 37736
rect 10100 37696 10101 37736
rect 10059 37687 10101 37696
rect 9964 37603 10004 37612
rect 9580 37518 9620 37603
rect 9772 37484 9812 37493
rect 9675 37232 9717 37241
rect 9675 37192 9676 37232
rect 9716 37192 9717 37232
rect 9675 37183 9717 37192
rect 9579 36644 9621 36653
rect 9579 36604 9580 36644
rect 9620 36604 9621 36644
rect 9579 36595 9621 36604
rect 9580 36510 9620 36595
rect 9676 36149 9716 37183
rect 9772 36989 9812 37444
rect 9771 36980 9813 36989
rect 9771 36940 9772 36980
rect 9812 36940 9813 36980
rect 9771 36931 9813 36940
rect 10060 36728 10100 37687
rect 10348 37577 10388 38527
rect 10444 38072 10484 39796
rect 10540 39964 10676 40004
rect 10540 39089 10580 39964
rect 10635 39836 10677 39845
rect 10635 39796 10636 39836
rect 10676 39796 10677 39836
rect 10635 39787 10677 39796
rect 10636 39752 10676 39787
rect 10636 39701 10676 39712
rect 10635 39164 10677 39173
rect 10635 39124 10636 39164
rect 10676 39124 10677 39164
rect 10635 39115 10677 39124
rect 10539 39080 10581 39089
rect 10539 39040 10540 39080
rect 10580 39040 10581 39080
rect 10539 39031 10581 39040
rect 10540 38912 10580 38921
rect 10636 38912 10676 39115
rect 10580 38872 10676 38912
rect 10540 38863 10580 38872
rect 10540 38249 10580 38334
rect 10539 38240 10581 38249
rect 10539 38200 10540 38240
rect 10580 38200 10581 38240
rect 10539 38191 10581 38200
rect 10444 38032 10676 38072
rect 10539 37652 10581 37661
rect 10539 37612 10540 37652
rect 10580 37612 10581 37652
rect 10539 37603 10581 37612
rect 10347 37568 10389 37577
rect 10347 37528 10348 37568
rect 10388 37528 10389 37568
rect 10347 37519 10389 37528
rect 10251 37400 10293 37409
rect 10251 37360 10252 37400
rect 10292 37360 10293 37400
rect 10348 37400 10388 37519
rect 10444 37400 10484 37409
rect 10348 37360 10444 37400
rect 10251 37351 10293 37360
rect 10252 37266 10292 37351
rect 10156 37232 10196 37241
rect 10156 36896 10196 37192
rect 10156 36856 10388 36896
rect 10060 36679 10100 36688
rect 10155 36728 10197 36737
rect 10155 36688 10156 36728
rect 10196 36688 10197 36728
rect 10155 36679 10197 36688
rect 10156 36594 10196 36679
rect 9771 36560 9813 36569
rect 9771 36520 9772 36560
rect 9812 36520 9813 36560
rect 9771 36511 9813 36520
rect 9772 36426 9812 36511
rect 10251 36308 10293 36317
rect 10251 36268 10252 36308
rect 10292 36268 10293 36308
rect 10251 36259 10293 36268
rect 9675 36140 9717 36149
rect 9675 36100 9676 36140
rect 9716 36100 9717 36140
rect 9675 36091 9717 36100
rect 9675 35972 9717 35981
rect 9675 35932 9676 35972
rect 9716 35932 9717 35972
rect 9675 35923 9717 35932
rect 9676 35888 9716 35923
rect 9580 35720 9620 35729
rect 9580 35393 9620 35680
rect 9388 35344 9524 35384
rect 9579 35384 9621 35393
rect 9579 35344 9580 35384
rect 9620 35344 9621 35384
rect 9676 35384 9716 35848
rect 9771 35888 9813 35897
rect 9771 35848 9772 35888
rect 9812 35848 9813 35888
rect 9771 35839 9813 35848
rect 9868 35888 9908 35897
rect 10059 35888 10101 35897
rect 9908 35848 10004 35888
rect 9868 35839 9908 35848
rect 9772 35754 9812 35839
rect 9868 35384 9908 35393
rect 9676 35344 9868 35384
rect 9291 33872 9333 33881
rect 9291 33832 9292 33872
rect 9332 33832 9333 33872
rect 9291 33823 9333 33832
rect 9291 33704 9333 33713
rect 9291 33664 9292 33704
rect 9332 33664 9333 33704
rect 9291 33655 9333 33664
rect 9195 32864 9237 32873
rect 9195 32824 9196 32864
rect 9236 32824 9237 32864
rect 9195 32815 9237 32824
rect 9004 32320 9140 32360
rect 9004 30437 9044 32320
rect 9099 32192 9141 32201
rect 9099 32152 9100 32192
rect 9140 32152 9141 32192
rect 9099 32143 9141 32152
rect 9100 32058 9140 32143
rect 9099 31352 9141 31361
rect 9099 31312 9100 31352
rect 9140 31312 9141 31352
rect 9099 31303 9141 31312
rect 9100 31218 9140 31303
rect 9100 30680 9140 30689
rect 9196 30680 9236 32815
rect 9292 32201 9332 33655
rect 9291 32192 9333 32201
rect 9291 32152 9292 32192
rect 9332 32152 9333 32192
rect 9291 32143 9333 32152
rect 9388 31193 9428 35344
rect 9579 35335 9621 35344
rect 9868 35335 9908 35344
rect 9964 35309 10004 35848
rect 10059 35848 10060 35888
rect 10100 35848 10101 35888
rect 10059 35839 10101 35848
rect 10156 35888 10196 35897
rect 10060 35754 10100 35839
rect 10156 35645 10196 35848
rect 10252 35888 10292 36259
rect 10348 35897 10388 36856
rect 10444 36737 10484 37360
rect 10443 36728 10485 36737
rect 10443 36688 10444 36728
rect 10484 36688 10485 36728
rect 10443 36679 10485 36688
rect 10540 36728 10580 37603
rect 10540 36485 10580 36688
rect 10636 36728 10676 38032
rect 10732 37988 10772 37997
rect 10732 37829 10772 37948
rect 10731 37820 10773 37829
rect 10731 37780 10732 37820
rect 10772 37780 10773 37820
rect 10731 37771 10773 37780
rect 10731 37484 10773 37493
rect 10731 37444 10732 37484
rect 10772 37444 10773 37484
rect 10731 37435 10773 37444
rect 10732 36989 10772 37435
rect 10731 36980 10773 36989
rect 10731 36940 10732 36980
rect 10772 36940 10773 36980
rect 10731 36931 10773 36940
rect 10636 36679 10676 36688
rect 10539 36476 10581 36485
rect 10539 36436 10540 36476
rect 10580 36436 10581 36476
rect 10539 36427 10581 36436
rect 10539 36056 10581 36065
rect 10539 36016 10540 36056
rect 10580 36016 10581 36056
rect 10539 36007 10581 36016
rect 10155 35636 10197 35645
rect 10155 35596 10156 35636
rect 10196 35596 10197 35636
rect 10155 35587 10197 35596
rect 10252 35309 10292 35848
rect 10347 35888 10389 35897
rect 10347 35848 10348 35888
rect 10388 35848 10389 35888
rect 10347 35839 10389 35848
rect 10540 35888 10580 36007
rect 10540 35839 10580 35848
rect 10348 35754 10388 35839
rect 10828 35309 10868 42928
rect 10923 42020 10965 42029
rect 10923 41980 10924 42020
rect 10964 41980 10965 42020
rect 10923 41971 10965 41980
rect 10924 39677 10964 41971
rect 11020 41609 11060 42928
rect 11115 42188 11157 42197
rect 11115 42148 11116 42188
rect 11156 42148 11157 42188
rect 11115 42139 11157 42148
rect 11019 41600 11061 41609
rect 11019 41560 11020 41600
rect 11060 41560 11061 41600
rect 11019 41551 11061 41560
rect 11116 40004 11156 42139
rect 11020 39964 11156 40004
rect 10923 39668 10965 39677
rect 10923 39628 10924 39668
rect 10964 39628 10965 39668
rect 10923 39619 10965 39628
rect 10923 37988 10965 37997
rect 10923 37948 10924 37988
rect 10964 37948 10965 37988
rect 10923 37939 10965 37948
rect 10924 37854 10964 37939
rect 10923 36140 10965 36149
rect 10923 36100 10924 36140
rect 10964 36100 10965 36140
rect 10923 36091 10965 36100
rect 9963 35300 10005 35309
rect 9963 35260 9964 35300
rect 10004 35260 10005 35300
rect 9963 35251 10005 35260
rect 10251 35300 10293 35309
rect 10251 35260 10252 35300
rect 10292 35260 10293 35300
rect 10251 35251 10293 35260
rect 10827 35300 10869 35309
rect 10827 35260 10828 35300
rect 10868 35260 10869 35300
rect 10827 35251 10869 35260
rect 9484 35216 9524 35225
rect 9524 35176 9812 35216
rect 9484 35167 9524 35176
rect 9676 34964 9716 34973
rect 9580 34924 9676 34964
rect 9580 34460 9620 34924
rect 9676 34915 9716 34924
rect 9772 34964 9812 35176
rect 10060 35195 10100 35204
rect 10060 35048 10100 35155
rect 9964 35008 10100 35048
rect 9964 34964 10004 35008
rect 9772 34924 10004 34964
rect 9532 34420 9620 34460
rect 9532 34418 9572 34420
rect 9532 34369 9572 34378
rect 9676 34208 9716 34217
rect 9579 33872 9621 33881
rect 9579 33832 9580 33872
rect 9620 33832 9621 33872
rect 9579 33823 9621 33832
rect 9387 31184 9429 31193
rect 9387 31144 9388 31184
rect 9428 31144 9429 31184
rect 9387 31135 9429 31144
rect 9580 30848 9620 33823
rect 9676 31529 9716 34168
rect 9772 33629 9812 34924
rect 10924 34805 10964 36091
rect 10923 34796 10965 34805
rect 10923 34756 10924 34796
rect 10964 34756 10965 34796
rect 10923 34747 10965 34756
rect 10059 34628 10101 34637
rect 10059 34588 10060 34628
rect 10100 34588 10101 34628
rect 10059 34579 10101 34588
rect 10060 34469 10100 34579
rect 11020 34544 11060 39964
rect 11116 38240 11156 38249
rect 11116 37325 11156 38200
rect 11115 37316 11157 37325
rect 11115 37276 11116 37316
rect 11156 37276 11157 37316
rect 11115 37267 11157 37276
rect 11116 36728 11156 36737
rect 11116 36233 11156 36688
rect 11115 36224 11157 36233
rect 11115 36184 11116 36224
rect 11156 36184 11157 36224
rect 11115 36175 11157 36184
rect 11212 36149 11252 42928
rect 11404 41693 11444 42928
rect 11403 41684 11445 41693
rect 11403 41644 11404 41684
rect 11444 41644 11445 41684
rect 11403 41635 11445 41644
rect 11596 41609 11636 42928
rect 11788 41609 11828 42928
rect 11980 42533 12020 42928
rect 11979 42524 12021 42533
rect 11979 42484 11980 42524
rect 12020 42484 12021 42524
rect 11979 42475 12021 42484
rect 11595 41600 11637 41609
rect 11595 41560 11596 41600
rect 11636 41560 11637 41600
rect 11595 41551 11637 41560
rect 11787 41600 11829 41609
rect 12172 41600 12212 42928
rect 12364 41609 12404 42928
rect 12556 42197 12596 42928
rect 12555 42188 12597 42197
rect 12555 42148 12556 42188
rect 12596 42148 12597 42188
rect 12555 42139 12597 42148
rect 11787 41560 11788 41600
rect 11828 41560 11829 41600
rect 11787 41551 11829 41560
rect 12076 41560 12212 41600
rect 12363 41600 12405 41609
rect 12363 41560 12364 41600
rect 12404 41560 12405 41600
rect 11980 41264 12020 41273
rect 11404 41224 11980 41264
rect 11307 39920 11349 39929
rect 11307 39880 11308 39920
rect 11348 39880 11349 39920
rect 11307 39871 11349 39880
rect 11211 36140 11253 36149
rect 11211 36100 11212 36140
rect 11252 36100 11253 36140
rect 11211 36091 11253 36100
rect 11308 36065 11348 39871
rect 11115 36056 11157 36065
rect 11115 36016 11116 36056
rect 11156 36016 11157 36056
rect 11115 36007 11157 36016
rect 11307 36056 11349 36065
rect 11307 36016 11308 36056
rect 11348 36016 11349 36056
rect 11307 36007 11349 36016
rect 11116 34805 11156 36007
rect 11211 35384 11253 35393
rect 11211 35344 11212 35384
rect 11252 35344 11253 35384
rect 11211 35335 11253 35344
rect 11115 34796 11157 34805
rect 11115 34756 11116 34796
rect 11156 34756 11157 34796
rect 11115 34747 11157 34756
rect 11020 34504 11156 34544
rect 10059 34460 10101 34469
rect 10059 34420 10060 34460
rect 10100 34420 10101 34460
rect 10059 34411 10101 34420
rect 9964 34376 10004 34385
rect 9868 34208 9908 34217
rect 9771 33620 9813 33629
rect 9771 33580 9772 33620
rect 9812 33580 9813 33620
rect 9771 33571 9813 33580
rect 9868 32957 9908 34168
rect 9867 32948 9909 32957
rect 9867 32908 9868 32948
rect 9908 32908 9909 32948
rect 9867 32899 9909 32908
rect 9964 32369 10004 34336
rect 10060 34376 10100 34411
rect 10060 34325 10100 34336
rect 10156 34376 10196 34385
rect 10059 34208 10101 34217
rect 10059 34168 10060 34208
rect 10100 34168 10101 34208
rect 10059 34159 10101 34168
rect 10060 32864 10100 34159
rect 10156 33881 10196 34336
rect 10348 34376 10388 34385
rect 10348 34217 10388 34336
rect 10444 34376 10484 34385
rect 10347 34208 10389 34217
rect 10347 34168 10348 34208
rect 10388 34168 10389 34208
rect 10347 34159 10389 34168
rect 10444 33881 10484 34336
rect 10540 34376 10580 34385
rect 10540 34049 10580 34336
rect 10923 34376 10965 34385
rect 10923 34336 10924 34376
rect 10964 34336 10965 34376
rect 10923 34327 10965 34336
rect 11020 34376 11060 34387
rect 10924 34217 10964 34327
rect 11020 34301 11060 34336
rect 11019 34292 11061 34301
rect 11019 34252 11020 34292
rect 11060 34252 11061 34292
rect 11019 34243 11061 34252
rect 10636 34208 10676 34217
rect 10923 34208 10965 34217
rect 10676 34168 10772 34208
rect 10636 34159 10676 34168
rect 10539 34040 10581 34049
rect 10539 34000 10540 34040
rect 10580 34000 10581 34040
rect 10539 33991 10581 34000
rect 10155 33872 10197 33881
rect 10155 33832 10156 33872
rect 10196 33832 10197 33872
rect 10155 33823 10197 33832
rect 10443 33872 10485 33881
rect 10443 33832 10444 33872
rect 10484 33832 10485 33872
rect 10443 33823 10485 33832
rect 10635 33872 10677 33881
rect 10635 33832 10636 33872
rect 10676 33832 10677 33872
rect 10635 33823 10677 33832
rect 10156 33704 10196 33715
rect 10156 33629 10196 33664
rect 10155 33620 10197 33629
rect 10155 33580 10156 33620
rect 10196 33580 10197 33620
rect 10155 33571 10197 33580
rect 10347 33452 10389 33461
rect 10347 33412 10348 33452
rect 10388 33412 10389 33452
rect 10347 33403 10389 33412
rect 10348 33318 10388 33403
rect 10444 33116 10484 33823
rect 10539 33704 10581 33713
rect 10539 33664 10540 33704
rect 10580 33664 10581 33704
rect 10539 33655 10581 33664
rect 10540 33570 10580 33655
rect 10444 33067 10484 33076
rect 10636 33032 10676 33823
rect 10540 32992 10676 33032
rect 10252 32864 10292 32873
rect 10060 32824 10252 32864
rect 9963 32360 10005 32369
rect 9963 32320 9964 32360
rect 10004 32320 10005 32360
rect 9963 32311 10005 32320
rect 10156 32192 10196 32824
rect 10252 32815 10292 32824
rect 10444 32705 10484 32790
rect 10443 32696 10485 32705
rect 10443 32656 10444 32696
rect 10484 32656 10485 32696
rect 10443 32647 10485 32656
rect 10540 32528 10580 32992
rect 10635 32864 10677 32873
rect 10635 32824 10636 32864
rect 10676 32824 10677 32864
rect 10635 32815 10677 32824
rect 10636 32730 10676 32815
rect 10444 32488 10580 32528
rect 10348 32192 10388 32201
rect 10156 32152 10348 32192
rect 10059 32108 10101 32117
rect 10059 32068 10060 32108
rect 10100 32068 10101 32108
rect 10059 32059 10101 32068
rect 9675 31520 9717 31529
rect 9675 31480 9676 31520
rect 9716 31480 9717 31520
rect 9675 31471 9717 31480
rect 9580 30808 9908 30848
rect 9140 30640 9236 30680
rect 9388 30680 9428 30689
rect 9100 30631 9140 30640
rect 9003 30428 9045 30437
rect 9003 30388 9004 30428
rect 9044 30388 9045 30428
rect 9003 30379 9045 30388
rect 9388 30260 9428 30640
rect 9772 30680 9812 30689
rect 9004 30220 9428 30260
rect 9484 30596 9524 30605
rect 8907 29924 8949 29933
rect 8907 29884 8908 29924
rect 8948 29884 8949 29924
rect 8907 29875 8949 29884
rect 8812 29840 8852 29849
rect 8812 29681 8852 29800
rect 8907 29756 8949 29765
rect 8907 29716 8908 29756
rect 8948 29716 8949 29756
rect 8907 29707 8949 29716
rect 8236 29632 8756 29672
rect 8811 29672 8853 29681
rect 8811 29632 8812 29672
rect 8852 29632 8853 29672
rect 8139 29252 8181 29261
rect 8139 29212 8140 29252
rect 8180 29212 8181 29252
rect 8139 29203 8181 29212
rect 8140 29168 8180 29203
rect 8140 29117 8180 29128
rect 8236 29168 8276 29632
rect 8811 29623 8853 29632
rect 8908 29622 8948 29707
rect 8427 29420 8469 29429
rect 8427 29380 8428 29420
rect 8468 29380 8469 29420
rect 8427 29371 8469 29380
rect 8428 29261 8468 29371
rect 8427 29252 8469 29261
rect 8427 29212 8428 29252
rect 8468 29212 8469 29252
rect 8427 29203 8469 29212
rect 8236 29119 8276 29128
rect 8428 29168 8468 29203
rect 8428 29118 8468 29128
rect 8620 29168 8660 29177
rect 8235 28916 8277 28925
rect 8235 28876 8236 28916
rect 8276 28876 8277 28916
rect 8235 28867 8277 28876
rect 8428 28916 8468 28925
rect 8140 27656 8180 27665
rect 8140 26825 8180 27616
rect 8236 26830 8276 28867
rect 8331 27068 8373 27077
rect 8331 27028 8332 27068
rect 8372 27028 8373 27068
rect 8331 27019 8373 27028
rect 8139 26816 8181 26825
rect 8139 26776 8140 26816
rect 8180 26776 8181 26816
rect 8236 26781 8276 26790
rect 8139 26767 8181 26776
rect 8043 26060 8085 26069
rect 8043 26020 8044 26060
rect 8084 26020 8085 26060
rect 8043 26011 8085 26020
rect 8043 25892 8085 25901
rect 8043 25852 8044 25892
rect 8084 25852 8085 25892
rect 8043 25843 8085 25852
rect 7700 25264 7988 25304
rect 8044 25304 8084 25843
rect 7660 24464 7700 25264
rect 8044 25255 8084 25264
rect 7852 25136 7892 25145
rect 7892 25096 7988 25136
rect 7852 25087 7892 25096
rect 7948 24627 7988 25096
rect 7948 24578 7988 24587
rect 8140 24716 8180 24725
rect 8140 24473 8180 24676
rect 8139 24464 8181 24473
rect 7660 24424 8084 24464
rect 7659 23960 7701 23969
rect 7659 23920 7660 23960
rect 7700 23920 7701 23960
rect 7659 23911 7701 23920
rect 7947 23960 7989 23969
rect 7947 23920 7948 23960
rect 7988 23920 7989 23960
rect 7947 23911 7989 23920
rect 7660 23806 7700 23911
rect 7660 23757 7700 23766
rect 7563 23624 7605 23633
rect 7563 23584 7564 23624
rect 7604 23584 7605 23624
rect 7563 23575 7605 23584
rect 7852 23624 7892 23633
rect 7467 23120 7509 23129
rect 7467 23080 7468 23120
rect 7508 23080 7509 23120
rect 7467 23071 7509 23080
rect 7852 22793 7892 23584
rect 7948 23036 7988 23911
rect 8044 23120 8084 24424
rect 8139 24424 8140 24464
rect 8180 24424 8181 24464
rect 8139 24415 8181 24424
rect 8332 23381 8372 27019
rect 8428 26816 8468 28876
rect 8620 28757 8660 29128
rect 9004 29000 9044 30220
rect 9484 30176 9524 30556
rect 9676 30596 9716 30605
rect 9580 30512 9620 30521
rect 9580 30353 9620 30472
rect 9579 30344 9621 30353
rect 9579 30304 9580 30344
rect 9620 30304 9621 30344
rect 9579 30295 9621 30304
rect 8812 28960 9044 29000
rect 9100 30136 9524 30176
rect 8619 28748 8661 28757
rect 8619 28708 8620 28748
rect 8660 28708 8661 28748
rect 8619 28699 8661 28708
rect 8523 28328 8565 28337
rect 8523 28288 8524 28328
rect 8564 28288 8565 28328
rect 8523 28279 8565 28288
rect 8524 28194 8564 28279
rect 8716 28160 8756 28169
rect 8716 27656 8756 28120
rect 8812 27908 8852 28960
rect 9004 28337 9044 28422
rect 9003 28328 9045 28337
rect 9003 28288 9004 28328
rect 9044 28288 9045 28328
rect 9003 28279 9045 28288
rect 8908 28160 8948 28169
rect 8948 28120 9044 28160
rect 8908 28111 8948 28120
rect 8812 27868 8948 27908
rect 8668 27646 8756 27656
rect 8708 27616 8756 27646
rect 8812 27740 8852 27749
rect 8668 27597 8708 27606
rect 8812 27329 8852 27700
rect 8811 27320 8853 27329
rect 8811 27280 8812 27320
rect 8852 27280 8853 27320
rect 8811 27271 8853 27280
rect 8716 27068 8756 27077
rect 8908 27068 8948 27868
rect 9004 27833 9044 28120
rect 9003 27824 9045 27833
rect 9003 27784 9004 27824
rect 9044 27784 9045 27824
rect 9003 27775 9045 27784
rect 9100 27740 9140 30136
rect 9579 30092 9621 30101
rect 9484 30052 9580 30092
rect 9620 30052 9621 30092
rect 9196 30008 9236 30017
rect 9387 30008 9429 30017
rect 9236 29968 9332 30008
rect 9196 29959 9236 29968
rect 9195 29420 9237 29429
rect 9195 29380 9196 29420
rect 9236 29380 9237 29420
rect 9195 29371 9237 29380
rect 9196 28589 9236 29371
rect 9195 28580 9237 28589
rect 9195 28540 9196 28580
rect 9236 28540 9237 28580
rect 9195 28531 9237 28540
rect 9195 28412 9237 28421
rect 9195 28372 9196 28412
rect 9236 28372 9237 28412
rect 9195 28363 9237 28372
rect 9196 28328 9236 28363
rect 9196 28277 9236 28288
rect 9100 27691 9140 27700
rect 9003 27656 9045 27665
rect 9003 27616 9004 27656
rect 9044 27616 9045 27656
rect 9003 27607 9045 27616
rect 9196 27656 9236 27665
rect 8756 27028 8948 27068
rect 8716 27019 8756 27028
rect 8716 26816 8756 26825
rect 8428 26776 8716 26816
rect 8716 26767 8756 26776
rect 9004 26816 9044 27607
rect 9099 27572 9141 27581
rect 9099 27532 9100 27572
rect 9140 27532 9141 27572
rect 9099 27523 9141 27532
rect 9100 26909 9140 27523
rect 9196 27488 9236 27616
rect 9292 27656 9332 29968
rect 9387 29968 9388 30008
rect 9428 29968 9429 30008
rect 9387 29959 9429 29968
rect 9388 29668 9428 29959
rect 9388 29619 9428 29628
rect 9484 29840 9524 30052
rect 9579 30043 9621 30052
rect 9579 29924 9621 29933
rect 9579 29884 9580 29924
rect 9620 29884 9621 29924
rect 9579 29875 9621 29884
rect 9387 29252 9429 29261
rect 9387 29212 9388 29252
rect 9428 29212 9429 29252
rect 9387 29203 9429 29212
rect 9292 27607 9332 27616
rect 9388 27488 9428 29203
rect 9484 29000 9524 29800
rect 9580 29840 9620 29875
rect 9580 29789 9620 29800
rect 9676 29000 9716 30556
rect 9772 30092 9812 30640
rect 9868 30260 9908 30808
rect 9964 30680 10004 30689
rect 9964 30521 10004 30640
rect 9963 30512 10005 30521
rect 9963 30472 9964 30512
rect 10004 30472 10005 30512
rect 9963 30463 10005 30472
rect 9868 30220 10004 30260
rect 9868 30092 9908 30101
rect 9772 30052 9868 30092
rect 9868 30043 9908 30052
rect 9964 29840 10004 30220
rect 10060 30017 10100 32059
rect 10156 31277 10196 32152
rect 10348 32143 10388 32152
rect 10251 31436 10293 31445
rect 10251 31396 10252 31436
rect 10292 31396 10293 31436
rect 10251 31387 10293 31396
rect 10155 31268 10197 31277
rect 10155 31228 10156 31268
rect 10196 31228 10197 31268
rect 10155 31219 10197 31228
rect 10059 30008 10101 30017
rect 10059 29968 10060 30008
rect 10100 29968 10101 30008
rect 10059 29959 10101 29968
rect 10156 29840 10196 29849
rect 9964 29800 10156 29840
rect 9867 29756 9909 29765
rect 9867 29716 9868 29756
rect 9908 29716 9909 29756
rect 9867 29707 9909 29716
rect 9868 29429 9908 29707
rect 9867 29420 9909 29429
rect 9867 29380 9868 29420
rect 9908 29380 9909 29420
rect 9867 29371 9909 29380
rect 9868 29168 9908 29177
rect 9484 28960 9620 29000
rect 9676 28960 9812 29000
rect 9483 27656 9525 27665
rect 9483 27616 9484 27656
rect 9524 27616 9525 27656
rect 9483 27607 9525 27616
rect 9580 27656 9620 28960
rect 9772 27740 9812 28960
rect 9772 27691 9812 27700
rect 9484 27522 9524 27607
rect 9196 27448 9428 27488
rect 9196 27077 9236 27162
rect 9195 27068 9237 27077
rect 9195 27028 9196 27068
rect 9236 27028 9237 27068
rect 9195 27019 9237 27028
rect 9099 26900 9141 26909
rect 9099 26860 9100 26900
rect 9140 26860 9141 26900
rect 9099 26851 9141 26860
rect 9004 26767 9044 26776
rect 9196 26816 9236 26825
rect 9292 26816 9332 27448
rect 9387 26900 9429 26909
rect 9387 26860 9388 26900
rect 9428 26860 9429 26900
rect 9387 26851 9429 26860
rect 9236 26776 9332 26816
rect 9388 26816 9428 26851
rect 9196 26767 9236 26776
rect 9388 26765 9428 26776
rect 9484 26816 9524 26825
rect 9580 26816 9620 27616
rect 9676 27656 9716 27665
rect 9676 27077 9716 27616
rect 9675 27068 9717 27077
rect 9675 27028 9676 27068
rect 9716 27028 9717 27068
rect 9675 27019 9717 27028
rect 9772 26993 9812 27078
rect 9771 26984 9813 26993
rect 9771 26944 9772 26984
rect 9812 26944 9813 26984
rect 9676 26909 9716 26940
rect 9771 26935 9813 26944
rect 9675 26900 9717 26909
rect 9675 26860 9676 26900
rect 9716 26860 9717 26900
rect 9675 26851 9717 26860
rect 9524 26776 9620 26816
rect 9676 26816 9716 26851
rect 9484 26767 9524 26776
rect 8427 26648 8469 26657
rect 9676 26648 9716 26776
rect 9771 26816 9813 26825
rect 9771 26776 9772 26816
rect 9812 26776 9813 26816
rect 9771 26767 9813 26776
rect 8427 26608 8428 26648
rect 8468 26608 8469 26648
rect 8427 26599 8469 26608
rect 9484 26608 9716 26648
rect 8428 26514 8468 26599
rect 9291 26564 9333 26573
rect 9291 26524 9292 26564
rect 9332 26524 9333 26564
rect 9291 26515 9333 26524
rect 8619 26480 8661 26489
rect 8619 26440 8620 26480
rect 8660 26440 8661 26480
rect 8619 26431 8661 26440
rect 8811 26480 8853 26489
rect 8811 26440 8812 26480
rect 8852 26440 8853 26480
rect 8811 26431 8853 26440
rect 9099 26480 9141 26489
rect 9099 26440 9100 26480
rect 9140 26440 9141 26480
rect 9099 26431 9141 26440
rect 8620 23801 8660 26431
rect 8715 26144 8757 26153
rect 8715 26104 8716 26144
rect 8756 26104 8757 26144
rect 8715 26095 8757 26104
rect 8716 26010 8756 26095
rect 8715 25808 8757 25817
rect 8715 25768 8716 25808
rect 8756 25768 8757 25808
rect 8715 25759 8757 25768
rect 8716 25481 8756 25759
rect 8715 25472 8757 25481
rect 8715 25432 8716 25472
rect 8756 25432 8757 25472
rect 8715 25423 8757 25432
rect 8716 24632 8756 25423
rect 8619 23792 8661 23801
rect 8619 23752 8620 23792
rect 8660 23752 8661 23792
rect 8619 23743 8661 23752
rect 8331 23372 8373 23381
rect 8331 23332 8332 23372
rect 8372 23332 8373 23372
rect 8331 23323 8373 23332
rect 8332 23120 8372 23129
rect 8044 23080 8332 23120
rect 7948 22996 8084 23036
rect 7851 22784 7893 22793
rect 7851 22744 7852 22784
rect 7892 22744 7988 22784
rect 7851 22735 7893 22744
rect 7275 22700 7317 22709
rect 7275 22660 7276 22700
rect 7316 22660 7317 22700
rect 7275 22651 7317 22660
rect 7755 22700 7797 22709
rect 7755 22660 7756 22700
rect 7796 22660 7797 22700
rect 7755 22651 7797 22660
rect 7371 22532 7413 22541
rect 7371 22492 7372 22532
rect 7412 22492 7413 22532
rect 7371 22483 7413 22492
rect 7275 22448 7317 22457
rect 7275 22408 7276 22448
rect 7316 22408 7317 22448
rect 7275 22399 7317 22408
rect 7276 22364 7316 22399
rect 7276 22313 7316 22324
rect 7180 22196 7220 22240
rect 7180 22156 7316 22196
rect 7179 21608 7221 21617
rect 7179 21568 7180 21608
rect 7220 21568 7221 21608
rect 7179 21559 7221 21568
rect 7180 21474 7220 21559
rect 7276 21533 7316 22156
rect 7275 21524 7317 21533
rect 7275 21484 7276 21524
rect 7316 21484 7317 21524
rect 7275 21475 7317 21484
rect 7083 21356 7125 21365
rect 7083 21316 7084 21356
rect 7124 21316 7125 21356
rect 7083 21307 7125 21316
rect 6891 21188 6933 21197
rect 6891 21148 6892 21188
rect 6932 21148 6933 21188
rect 6891 21139 6933 21148
rect 6796 20971 6836 20980
rect 6892 20180 6932 20220
rect 6700 20140 6836 20180
rect 6700 20082 6740 20091
rect 6700 19937 6740 20042
rect 6699 19928 6741 19937
rect 6699 19888 6700 19928
rect 6740 19888 6741 19928
rect 6699 19879 6741 19888
rect 6796 19760 6836 20140
rect 6892 20105 6932 20140
rect 7084 20180 7124 20189
rect 7372 20180 7412 22483
rect 7756 22280 7796 22651
rect 7659 22112 7701 22121
rect 7659 22072 7660 22112
rect 7700 22072 7701 22112
rect 7659 22063 7701 22072
rect 7660 21603 7700 22063
rect 7756 21617 7796 22240
rect 7852 21692 7892 21701
rect 7660 21554 7700 21563
rect 7755 21608 7797 21617
rect 7755 21568 7756 21608
rect 7796 21568 7797 21608
rect 7755 21559 7797 21568
rect 7467 21524 7509 21533
rect 7467 21484 7468 21524
rect 7508 21484 7509 21524
rect 7467 21475 7509 21484
rect 6891 20096 6933 20105
rect 6891 20056 6892 20096
rect 6932 20056 6933 20096
rect 6891 20047 6933 20056
rect 6892 20045 6932 20047
rect 6891 19928 6933 19937
rect 6891 19888 6892 19928
rect 6932 19888 6933 19928
rect 6891 19879 6933 19888
rect 6700 19720 6836 19760
rect 6700 17828 6740 19720
rect 6796 18584 6836 18593
rect 6796 18425 6836 18544
rect 6795 18416 6837 18425
rect 6795 18376 6796 18416
rect 6836 18376 6837 18416
rect 6795 18367 6837 18376
rect 6795 17996 6837 18005
rect 6795 17956 6796 17996
rect 6836 17956 6837 17996
rect 6795 17947 6837 17956
rect 6700 17165 6740 17788
rect 6796 17828 6836 17947
rect 6796 17779 6836 17788
rect 6892 17333 6932 19879
rect 7084 19601 7124 20140
rect 7180 20140 7412 20180
rect 7083 19592 7125 19601
rect 7083 19552 7084 19592
rect 7124 19552 7125 19592
rect 7083 19543 7125 19552
rect 6988 19256 7028 19267
rect 7180 19256 7220 20140
rect 7276 20082 7316 20091
rect 7276 19508 7316 20042
rect 7372 19508 7412 19517
rect 7276 19468 7372 19508
rect 7372 19459 7412 19468
rect 6988 19181 7028 19216
rect 7084 19216 7220 19256
rect 7371 19256 7413 19265
rect 7371 19216 7372 19256
rect 7412 19216 7413 19256
rect 6987 19172 7029 19181
rect 6987 19132 6988 19172
rect 7028 19132 7029 19172
rect 6987 19123 7029 19132
rect 6987 18752 7029 18761
rect 6987 18712 6988 18752
rect 7028 18712 7029 18752
rect 6987 18703 7029 18712
rect 6988 18618 7028 18703
rect 7084 18593 7124 19216
rect 7371 19207 7413 19216
rect 7180 19088 7220 19097
rect 7083 18584 7125 18593
rect 7083 18544 7084 18584
rect 7124 18544 7125 18584
rect 7083 18535 7125 18544
rect 6891 17324 6933 17333
rect 6891 17284 6892 17324
rect 6932 17284 6933 17324
rect 6891 17275 6933 17284
rect 6699 17156 6741 17165
rect 6699 17116 6700 17156
rect 6740 17116 6741 17156
rect 6699 17107 6741 17116
rect 6699 16988 6741 16997
rect 6699 16948 6700 16988
rect 6740 16948 6741 16988
rect 6699 16939 6741 16948
rect 6796 16988 6836 16997
rect 6700 16854 6740 16939
rect 6796 16829 6836 16948
rect 6795 16820 6837 16829
rect 6795 16780 6796 16820
rect 6836 16780 6837 16820
rect 6795 16771 6837 16780
rect 6603 16568 6645 16577
rect 6603 16528 6604 16568
rect 6644 16528 6645 16568
rect 6603 16519 6645 16528
rect 6411 16400 6453 16409
rect 6411 16360 6412 16400
rect 6452 16360 6453 16400
rect 6411 16351 6453 16360
rect 6311 16241 6351 16326
rect 6310 16232 6352 16241
rect 6310 16192 6311 16232
rect 6351 16192 6352 16232
rect 6310 16183 6352 16192
rect 6411 16232 6453 16241
rect 6411 16192 6412 16232
rect 6452 16192 6453 16232
rect 6411 16183 6453 16192
rect 6508 16232 6548 16241
rect 6700 16232 6740 16241
rect 6412 16098 6452 16183
rect 6316 16064 6356 16073
rect 6124 15772 6260 15812
rect 6220 14804 6260 15772
rect 6316 15056 6356 16024
rect 6508 15149 6548 16192
rect 6604 16192 6700 16232
rect 6604 15485 6644 16192
rect 6700 16183 6740 16192
rect 6796 16232 6836 16241
rect 6699 15560 6741 15569
rect 6699 15520 6700 15560
rect 6740 15520 6741 15560
rect 6699 15511 6741 15520
rect 6603 15476 6645 15485
rect 6603 15436 6604 15476
rect 6644 15436 6645 15476
rect 6603 15427 6645 15436
rect 6700 15426 6740 15511
rect 6699 15308 6741 15317
rect 6699 15268 6700 15308
rect 6740 15268 6741 15308
rect 6699 15259 6741 15268
rect 6507 15140 6549 15149
rect 6507 15100 6508 15140
rect 6548 15100 6549 15140
rect 6507 15091 6549 15100
rect 6316 15016 6452 15056
rect 6412 14972 6452 15016
rect 6412 14932 6644 14972
rect 6220 14755 6260 14764
rect 6316 14888 6356 14897
rect 6027 14720 6069 14729
rect 6027 14680 6028 14720
rect 6068 14680 6069 14720
rect 6027 14671 6069 14680
rect 6124 14720 6164 14729
rect 5972 14008 6068 14048
rect 5548 13999 5588 14008
rect 5932 13999 5972 14008
rect 5260 13924 5396 13964
rect 5260 13217 5300 13924
rect 5452 13796 5492 13805
rect 5356 13756 5452 13796
rect 5259 13208 5301 13217
rect 5259 13168 5260 13208
rect 5300 13168 5301 13208
rect 5259 13159 5301 13168
rect 5163 13040 5205 13049
rect 5163 13000 5164 13040
rect 5204 13000 5205 13040
rect 5163 12991 5205 13000
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4779 11780 4821 11789
rect 4779 11740 4780 11780
rect 4820 11740 4821 11780
rect 4779 11731 4821 11740
rect 5259 11780 5301 11789
rect 5259 11740 5260 11780
rect 5300 11740 5301 11780
rect 5259 11731 5301 11740
rect 4395 11696 4437 11705
rect 4395 11656 4396 11696
rect 4436 11656 4437 11696
rect 4395 11647 4437 11656
rect 4587 11696 4629 11705
rect 4587 11656 4588 11696
rect 4628 11656 4629 11696
rect 4587 11647 4629 11656
rect 4875 11696 4917 11705
rect 4875 11656 4876 11696
rect 4916 11656 4917 11696
rect 4875 11647 4917 11656
rect 5260 11696 5300 11731
rect 4396 11562 4436 11647
rect 4779 11612 4821 11621
rect 4779 11572 4780 11612
rect 4820 11572 4821 11612
rect 4779 11563 4821 11572
rect 4587 11528 4629 11537
rect 4587 11488 4588 11528
rect 4628 11488 4629 11528
rect 4587 11479 4629 11488
rect 4491 11444 4533 11453
rect 4491 11404 4492 11444
rect 4532 11404 4533 11444
rect 4491 11395 4533 11404
rect 3723 11276 3765 11285
rect 3723 11236 3724 11276
rect 3764 11236 3765 11276
rect 3723 11227 3765 11236
rect 3249 11068 3380 11108
rect 3531 11108 3573 11117
rect 3531 11068 3532 11108
rect 3572 11068 3573 11108
rect 3147 11024 3189 11033
rect 3147 10984 3148 11024
rect 3188 10984 3189 11024
rect 3147 10975 3189 10984
rect 3249 11014 3289 11068
rect 3531 11059 3573 11068
rect 3148 10890 3188 10975
rect 3249 10949 3289 10974
rect 3243 10940 3289 10949
rect 3243 10900 3244 10940
rect 3284 10900 3289 10940
rect 3724 11024 3764 11227
rect 3243 10891 3285 10900
rect 3724 10865 3764 10984
rect 4395 10940 4437 10949
rect 4395 10900 4396 10940
rect 4436 10900 4437 10940
rect 4395 10891 4437 10900
rect 3435 10856 3477 10865
rect 3435 10816 3436 10856
rect 3476 10816 3477 10856
rect 3435 10807 3477 10816
rect 3723 10856 3765 10865
rect 3723 10816 3724 10856
rect 3764 10816 3765 10856
rect 3723 10807 3765 10816
rect 4107 10856 4149 10865
rect 4107 10816 4108 10856
rect 4148 10816 4149 10856
rect 4107 10807 4149 10816
rect 3339 10520 3381 10529
rect 3339 10480 3340 10520
rect 3380 10480 3381 10520
rect 3339 10471 3381 10480
rect 3243 10184 3285 10193
rect 3340 10184 3380 10471
rect 3243 10144 3244 10184
rect 3284 10144 3380 10184
rect 3243 10135 3285 10144
rect 3148 10100 3188 10109
rect 3051 10016 3093 10025
rect 3051 9976 3052 10016
rect 3092 9976 3093 10016
rect 3051 9967 3093 9976
rect 2955 9764 2997 9773
rect 2955 9724 2956 9764
rect 2996 9724 2997 9764
rect 2955 9715 2997 9724
rect 3148 9689 3188 10060
rect 3244 10050 3284 10135
rect 3243 9848 3285 9857
rect 3243 9808 3244 9848
rect 3284 9808 3285 9848
rect 3243 9799 3285 9808
rect 3147 9680 3189 9689
rect 3147 9640 3148 9680
rect 3188 9640 3189 9680
rect 3147 9631 3189 9640
rect 3244 9680 3284 9799
rect 3244 9631 3284 9640
rect 3436 9521 3476 10807
rect 3532 10772 3572 10781
rect 3532 10361 3572 10732
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 3531 10352 3573 10361
rect 3531 10312 3532 10352
rect 3572 10312 3573 10352
rect 3531 10303 3573 10312
rect 4011 10352 4053 10361
rect 4011 10312 4012 10352
rect 4052 10312 4053 10352
rect 4011 10303 4053 10312
rect 4012 10198 4052 10303
rect 3532 10184 3572 10195
rect 4012 10149 4052 10158
rect 3532 10109 3572 10144
rect 3531 10100 3573 10109
rect 3531 10060 3532 10100
rect 3572 10060 3573 10100
rect 3531 10051 3573 10060
rect 3820 10100 3860 10109
rect 4108 10100 4148 10807
rect 4203 10688 4245 10697
rect 4203 10648 4204 10688
rect 4244 10648 4245 10688
rect 4203 10639 4245 10648
rect 4204 10361 4244 10639
rect 4203 10352 4245 10361
rect 4203 10312 4204 10352
rect 4244 10312 4245 10352
rect 4203 10303 4245 10312
rect 3860 10060 4148 10100
rect 3820 10051 3860 10060
rect 3531 9596 3573 9605
rect 3531 9556 3532 9596
rect 3572 9556 3573 9596
rect 3531 9547 3573 9556
rect 3723 9596 3765 9605
rect 3723 9556 3724 9596
rect 3764 9556 3765 9596
rect 3723 9547 3765 9556
rect 3051 9512 3093 9521
rect 3051 9472 3052 9512
rect 3092 9472 3093 9512
rect 3051 9463 3093 9472
rect 3435 9512 3477 9521
rect 3435 9472 3436 9512
rect 3476 9472 3477 9512
rect 3435 9463 3477 9472
rect 3052 9378 3092 9463
rect 3339 9260 3381 9269
rect 3339 9220 3340 9260
rect 3380 9220 3381 9260
rect 3339 9211 3381 9220
rect 3436 9260 3476 9269
rect 3243 8924 3285 8933
rect 3243 8884 3244 8924
rect 3284 8884 3285 8924
rect 3243 8875 3285 8884
rect 3244 8790 3284 8875
rect 2860 8707 2900 8716
rect 2955 8588 2997 8597
rect 2955 8548 2956 8588
rect 2996 8548 2997 8588
rect 2955 8539 2997 8548
rect 2956 8168 2996 8539
rect 3052 8504 3092 8513
rect 3092 8464 3284 8504
rect 3052 8455 3092 8464
rect 2956 8119 2996 8128
rect 2188 6439 2228 6448
rect 2764 6434 2804 6443
rect 2860 7990 3140 8000
rect 2860 7960 3100 7990
rect 2187 6236 2229 6245
rect 2187 6196 2188 6236
rect 2228 6196 2229 6236
rect 2187 6187 2229 6196
rect 2667 6236 2709 6245
rect 2667 6196 2668 6236
rect 2708 6196 2709 6236
rect 2667 6187 2709 6196
rect 2091 6068 2133 6077
rect 2091 6028 2092 6068
rect 2132 6028 2133 6068
rect 2091 6019 2133 6028
rect 1996 5599 2036 5608
rect 1899 5480 1941 5489
rect 1899 5440 1900 5480
rect 1940 5440 1941 5480
rect 1899 5431 1941 5440
rect 1612 5104 1748 5144
rect 1612 4976 1652 4985
rect 1612 4649 1652 4936
rect 1611 4640 1653 4649
rect 1611 4600 1612 4640
rect 1652 4600 1653 4640
rect 1611 4591 1653 4600
rect 1708 4397 1748 5104
rect 1803 4472 1845 4481
rect 1803 4432 1804 4472
rect 1844 4432 1845 4472
rect 1803 4423 1845 4432
rect 1707 4388 1749 4397
rect 1707 4348 1708 4388
rect 1748 4348 1749 4388
rect 1707 4339 1749 4348
rect 1516 4087 1556 4096
rect 1612 4136 1652 4145
rect 1612 3968 1652 4096
rect 1324 3928 1652 3968
rect 1708 4136 1748 4145
rect 1227 3919 1269 3928
rect 844 2500 1076 2540
rect 844 953 884 2500
rect 1228 1868 1268 3919
rect 1708 3809 1748 4096
rect 1804 4136 1844 4423
rect 1804 4087 1844 4096
rect 1515 3800 1557 3809
rect 1515 3760 1516 3800
rect 1556 3760 1557 3800
rect 1515 3751 1557 3760
rect 1707 3800 1749 3809
rect 1900 3800 1940 5431
rect 2092 5396 2132 6019
rect 2188 5648 2228 6187
rect 2283 5816 2325 5825
rect 2283 5776 2284 5816
rect 2324 5776 2325 5816
rect 2283 5767 2325 5776
rect 2380 5816 2420 5825
rect 2284 5732 2324 5767
rect 2284 5681 2324 5692
rect 2380 5657 2420 5776
rect 2476 5732 2516 5741
rect 2188 5573 2228 5608
rect 2379 5648 2421 5657
rect 2379 5608 2380 5648
rect 2420 5608 2421 5648
rect 2379 5599 2421 5608
rect 2187 5564 2229 5573
rect 2187 5524 2188 5564
rect 2228 5524 2229 5564
rect 2187 5515 2229 5524
rect 2188 5484 2228 5515
rect 2092 5356 2420 5396
rect 2091 5228 2133 5237
rect 2091 5188 2092 5228
rect 2132 5188 2133 5228
rect 2091 5179 2133 5188
rect 1995 5060 2037 5069
rect 1995 5020 1996 5060
rect 2036 5020 2037 5060
rect 1995 5011 2037 5020
rect 1996 4136 2036 5011
rect 1996 4087 2036 4096
rect 1995 3968 2037 3977
rect 1995 3928 1996 3968
rect 2036 3928 2037 3968
rect 1995 3919 2037 3928
rect 1707 3760 1708 3800
rect 1748 3760 1749 3800
rect 1707 3751 1749 3760
rect 1804 3760 1940 3800
rect 1419 3632 1461 3641
rect 1419 3592 1420 3632
rect 1460 3592 1461 3632
rect 1419 3583 1461 3592
rect 1323 2792 1365 2801
rect 1323 2752 1324 2792
rect 1364 2752 1365 2792
rect 1323 2743 1365 2752
rect 1228 1819 1268 1828
rect 1324 1280 1364 2743
rect 1420 2624 1460 3583
rect 1516 2885 1556 3751
rect 1611 3716 1653 3725
rect 1611 3676 1612 3716
rect 1652 3676 1653 3716
rect 1611 3667 1653 3676
rect 1515 2876 1557 2885
rect 1515 2836 1516 2876
rect 1556 2836 1557 2876
rect 1515 2827 1557 2836
rect 1612 2801 1652 3667
rect 1708 3296 1748 3305
rect 1611 2792 1653 2801
rect 1611 2752 1612 2792
rect 1652 2752 1653 2792
rect 1611 2743 1653 2752
rect 1612 2658 1652 2743
rect 1420 2120 1460 2584
rect 1708 2297 1748 3256
rect 1707 2288 1749 2297
rect 1707 2248 1708 2288
rect 1748 2248 1749 2288
rect 1707 2239 1749 2248
rect 1612 2120 1652 2129
rect 1420 2080 1612 2120
rect 1612 2071 1652 2080
rect 1708 1784 1748 1793
rect 1420 1700 1460 1709
rect 1420 1457 1460 1660
rect 1419 1448 1461 1457
rect 1419 1408 1420 1448
rect 1460 1408 1461 1448
rect 1419 1399 1461 1408
rect 1708 1373 1748 1744
rect 1707 1364 1749 1373
rect 1707 1324 1708 1364
rect 1748 1324 1749 1364
rect 1707 1315 1749 1324
rect 1324 1231 1364 1240
rect 1515 1196 1557 1205
rect 1515 1156 1516 1196
rect 1556 1156 1557 1196
rect 1515 1147 1557 1156
rect 1516 1062 1556 1147
rect 843 944 885 953
rect 843 904 844 944
rect 884 904 885 944
rect 843 895 885 904
rect 1708 944 1748 953
rect 1708 533 1748 904
rect 1707 524 1749 533
rect 1707 484 1708 524
rect 1748 484 1749 524
rect 1707 475 1749 484
rect 1804 80 1844 3760
rect 1899 3632 1941 3641
rect 1899 3592 1900 3632
rect 1940 3592 1941 3632
rect 1899 3583 1941 3592
rect 1900 2792 1940 3583
rect 1996 3464 2036 3919
rect 1996 3415 2036 3424
rect 2092 3221 2132 5179
rect 2283 4220 2325 4229
rect 2283 4180 2284 4220
rect 2324 4180 2325 4220
rect 2283 4171 2325 4180
rect 2187 4136 2229 4145
rect 2187 4096 2188 4136
rect 2228 4096 2229 4136
rect 2187 4087 2229 4096
rect 2188 3893 2228 4087
rect 2187 3884 2229 3893
rect 2187 3844 2188 3884
rect 2228 3844 2229 3884
rect 2187 3835 2229 3844
rect 2091 3212 2133 3221
rect 2091 3172 2092 3212
rect 2132 3172 2133 3212
rect 2091 3163 2133 3172
rect 1900 2204 1940 2752
rect 2092 2372 2132 3163
rect 2188 2633 2228 2718
rect 2187 2624 2229 2633
rect 2187 2584 2188 2624
rect 2228 2584 2229 2624
rect 2187 2575 2229 2584
rect 2092 2332 2228 2372
rect 1900 2164 2132 2204
rect 1900 2120 1940 2164
rect 1900 2071 1940 2080
rect 1995 2036 2037 2045
rect 1995 1996 1996 2036
rect 2036 1996 2037 2036
rect 1995 1987 2037 1996
rect 1996 1112 2036 1987
rect 2092 1121 2132 2164
rect 2188 1952 2228 2332
rect 2188 1903 2228 1912
rect 2187 1616 2229 1625
rect 2187 1576 2188 1616
rect 2228 1576 2229 1616
rect 2187 1567 2229 1576
rect 1996 1063 2036 1072
rect 2091 1112 2133 1121
rect 2091 1072 2092 1112
rect 2132 1072 2133 1112
rect 2091 1063 2133 1072
rect 2092 978 2132 1063
rect 1995 944 2037 953
rect 1995 904 1996 944
rect 2036 904 2037 944
rect 1995 895 2037 904
rect 1996 80 2036 895
rect 2188 80 2228 1567
rect 2284 1289 2324 4171
rect 2283 1280 2325 1289
rect 2283 1240 2284 1280
rect 2324 1240 2325 1280
rect 2283 1231 2325 1240
rect 2380 80 2420 5356
rect 2476 3137 2516 5692
rect 2571 5648 2613 5657
rect 2571 5608 2572 5648
rect 2612 5608 2613 5648
rect 2571 5599 2613 5608
rect 2572 5514 2612 5599
rect 2475 3128 2517 3137
rect 2475 3088 2476 3128
rect 2516 3088 2517 3128
rect 2475 3079 2517 3088
rect 2475 1280 2517 1289
rect 2475 1240 2476 1280
rect 2516 1240 2517 1280
rect 2475 1231 2517 1240
rect 2476 1196 2516 1231
rect 2476 1145 2516 1156
rect 2571 1196 2613 1205
rect 2571 1156 2572 1196
rect 2612 1156 2613 1196
rect 2571 1147 2613 1156
rect 2572 1062 2612 1147
rect 2668 944 2708 6187
rect 2764 5900 2804 5909
rect 2860 5900 2900 7960
rect 3100 7941 3140 7950
rect 2955 7832 2997 7841
rect 2955 7792 2956 7832
rect 2996 7792 2997 7832
rect 2955 7783 2997 7792
rect 2956 6161 2996 7783
rect 3244 6917 3284 8464
rect 3243 6908 3285 6917
rect 3243 6868 3244 6908
rect 3284 6868 3285 6908
rect 3243 6859 3285 6868
rect 3244 6488 3284 6497
rect 3051 6236 3093 6245
rect 3051 6196 3052 6236
rect 3092 6196 3093 6236
rect 3051 6187 3093 6196
rect 2955 6152 2997 6161
rect 2955 6112 2956 6152
rect 2996 6112 2997 6152
rect 2955 6103 2997 6112
rect 2804 5860 2900 5900
rect 2764 5851 2804 5860
rect 2956 5648 2996 5657
rect 3052 5648 3092 6187
rect 3244 6161 3284 6448
rect 3243 6152 3285 6161
rect 3243 6112 3244 6152
rect 3284 6112 3285 6152
rect 3243 6103 3285 6112
rect 2996 5608 3092 5648
rect 2956 5599 2996 5608
rect 2860 4976 2900 4985
rect 3147 4976 3189 4985
rect 2900 4936 3148 4976
rect 3188 4936 3189 4976
rect 2860 4927 2900 4936
rect 3147 4927 3189 4936
rect 3244 4976 3284 4985
rect 2859 4724 2901 4733
rect 2859 4684 2860 4724
rect 2900 4684 2901 4724
rect 2859 4675 2901 4684
rect 3052 4724 3092 4733
rect 2860 1709 2900 4675
rect 3052 3305 3092 4684
rect 3148 4136 3188 4927
rect 3244 4733 3284 4936
rect 3243 4724 3285 4733
rect 3243 4684 3244 4724
rect 3284 4684 3285 4724
rect 3243 4675 3285 4684
rect 3244 4136 3284 4145
rect 3148 4096 3244 4136
rect 3051 3296 3093 3305
rect 3051 3256 3052 3296
rect 3092 3256 3093 3296
rect 3051 3247 3093 3256
rect 3148 2465 3188 4096
rect 3244 4087 3284 4096
rect 3340 4052 3380 9211
rect 3436 7337 3476 9220
rect 3532 8840 3572 9547
rect 3724 9462 3764 9547
rect 3819 9512 3861 9521
rect 3819 9472 3820 9512
rect 3860 9472 3861 9512
rect 3819 9463 3861 9472
rect 4108 9512 4148 9521
rect 4204 9512 4244 10303
rect 4148 9472 4244 9512
rect 4299 9512 4341 9521
rect 4299 9472 4300 9512
rect 4340 9472 4341 9512
rect 3820 9378 3860 9463
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3532 8800 3764 8840
rect 3724 8756 3764 8800
rect 3724 8716 3860 8756
rect 3531 8672 3573 8681
rect 3531 8632 3532 8672
rect 3572 8632 3573 8672
rect 3531 8623 3573 8632
rect 3628 8672 3668 8681
rect 3668 8632 3764 8672
rect 3628 8623 3668 8632
rect 3532 8538 3572 8623
rect 3724 8345 3764 8632
rect 3723 8336 3765 8345
rect 3723 8296 3724 8336
rect 3764 8296 3765 8336
rect 3723 8287 3765 8296
rect 3724 8093 3764 8287
rect 3723 8084 3765 8093
rect 3723 8044 3724 8084
rect 3764 8044 3765 8084
rect 3723 8035 3765 8044
rect 3628 8000 3668 8009
rect 3628 7757 3668 7960
rect 3820 7757 3860 8716
rect 3916 8672 3956 8681
rect 4108 8672 4148 9472
rect 4299 9463 4341 9472
rect 4396 9512 4436 10891
rect 4492 10184 4532 11395
rect 4588 11394 4628 11479
rect 4780 11478 4820 11563
rect 4876 11562 4916 11647
rect 5260 11645 5300 11656
rect 5068 11537 5108 11622
rect 5067 11528 5109 11537
rect 5067 11488 5068 11528
rect 5108 11488 5109 11528
rect 5067 11479 5109 11488
rect 4779 11360 4821 11369
rect 4779 11320 4780 11360
rect 4820 11320 4821 11360
rect 4779 11311 4821 11320
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4780 10277 4820 11311
rect 5067 11192 5109 11201
rect 5067 11152 5068 11192
rect 5108 11152 5109 11192
rect 5067 11143 5109 11152
rect 4971 11108 5013 11117
rect 4971 11068 4972 11108
rect 5012 11068 5013 11108
rect 4971 11059 5013 11068
rect 4972 11024 5012 11059
rect 4972 10973 5012 10984
rect 4779 10268 4821 10277
rect 4779 10228 4780 10268
rect 4820 10228 4821 10268
rect 4779 10219 4821 10228
rect 5068 10268 5108 11143
rect 5164 11024 5204 11035
rect 5164 10949 5204 10984
rect 5163 10940 5205 10949
rect 5163 10900 5164 10940
rect 5204 10900 5205 10940
rect 5163 10891 5205 10900
rect 5068 10219 5108 10228
rect 4492 9857 4532 10144
rect 4683 10100 4725 10109
rect 4683 10060 4684 10100
rect 4724 10060 4725 10100
rect 4683 10051 4725 10060
rect 4587 10016 4629 10025
rect 4587 9976 4588 10016
rect 4628 9976 4629 10016
rect 4587 9967 4629 9976
rect 4491 9848 4533 9857
rect 4491 9808 4492 9848
rect 4532 9808 4533 9848
rect 4491 9799 4533 9808
rect 4491 9680 4533 9689
rect 4491 9640 4492 9680
rect 4532 9640 4533 9680
rect 4491 9631 4533 9640
rect 4492 9546 4532 9631
rect 4396 9463 4436 9472
rect 4588 9512 4628 9967
rect 4588 9463 4628 9472
rect 4684 9512 4724 10051
rect 4684 9463 4724 9472
rect 4300 8933 4340 9463
rect 4780 9344 4820 10219
rect 4972 10184 5012 10193
rect 4972 10100 5012 10144
rect 5067 10100 5109 10109
rect 4972 10060 5068 10100
rect 5108 10060 5109 10100
rect 5067 10051 5109 10060
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4875 9680 4917 9689
rect 5356 9680 5396 13756
rect 5452 13747 5492 13756
rect 5740 13796 5780 13805
rect 5780 13756 5972 13796
rect 5740 13747 5780 13756
rect 5547 13208 5589 13217
rect 5547 13168 5548 13208
rect 5588 13168 5589 13208
rect 5547 13159 5589 13168
rect 5451 12788 5493 12797
rect 5451 12748 5452 12788
rect 5492 12748 5493 12788
rect 5451 12739 5493 12748
rect 5452 12536 5492 12739
rect 5452 10352 5492 12496
rect 5548 11033 5588 13159
rect 5739 13040 5781 13049
rect 5739 13000 5740 13040
rect 5780 13000 5781 13040
rect 5739 12991 5781 13000
rect 5643 12620 5685 12629
rect 5643 12580 5644 12620
rect 5684 12580 5685 12620
rect 5643 12571 5685 12580
rect 5644 12486 5684 12571
rect 5547 11024 5589 11033
rect 5547 10984 5548 11024
rect 5588 10984 5589 11024
rect 5547 10975 5589 10984
rect 5740 10361 5780 12991
rect 5835 12704 5877 12713
rect 5835 12664 5836 12704
rect 5876 12664 5877 12704
rect 5835 12655 5877 12664
rect 5836 12570 5876 12655
rect 5932 12536 5972 13756
rect 6028 12797 6068 14008
rect 6124 13469 6164 14680
rect 6219 14552 6261 14561
rect 6219 14512 6220 14552
rect 6260 14512 6261 14552
rect 6219 14503 6261 14512
rect 6123 13460 6165 13469
rect 6123 13420 6124 13460
rect 6164 13420 6165 13460
rect 6123 13411 6165 13420
rect 6123 13208 6165 13217
rect 6123 13168 6124 13208
rect 6164 13168 6165 13208
rect 6123 13159 6165 13168
rect 6124 13074 6164 13159
rect 6027 12788 6069 12797
rect 6027 12748 6028 12788
rect 6068 12748 6069 12788
rect 6027 12739 6069 12748
rect 5932 12526 6020 12536
rect 5932 12496 5980 12526
rect 5980 12477 6020 12486
rect 5835 12452 5877 12461
rect 5835 12412 5836 12452
rect 5876 12412 5877 12452
rect 5835 12403 5877 12412
rect 5739 10352 5781 10361
rect 5452 10312 5684 10352
rect 4875 9640 4876 9680
rect 4916 9640 4917 9680
rect 4875 9631 4917 9640
rect 5260 9640 5396 9680
rect 5452 10184 5492 10193
rect 4876 9512 4916 9631
rect 4876 9463 4916 9472
rect 4588 9304 4820 9344
rect 4299 8924 4341 8933
rect 4299 8884 4300 8924
rect 4340 8884 4341 8924
rect 4299 8875 4341 8884
rect 4588 8840 4628 9304
rect 4971 9092 5013 9101
rect 4971 9052 4972 9092
rect 5012 9052 5013 9092
rect 4971 9043 5013 9052
rect 4683 8924 4725 8933
rect 4683 8884 4684 8924
rect 4724 8884 4725 8924
rect 4683 8875 4725 8884
rect 4492 8800 4628 8840
rect 3956 8632 4148 8672
rect 4203 8672 4245 8681
rect 4203 8632 4204 8672
rect 4244 8632 4245 8672
rect 3916 8623 3956 8632
rect 4203 8623 4245 8632
rect 4300 8672 4340 8681
rect 4107 7916 4149 7925
rect 4107 7876 4108 7916
rect 4148 7876 4149 7916
rect 4107 7867 4149 7876
rect 4204 7916 4244 8623
rect 4108 7782 4148 7867
rect 4204 7841 4244 7876
rect 4203 7832 4245 7841
rect 4203 7792 4204 7832
rect 4244 7792 4245 7832
rect 4203 7783 4245 7792
rect 3627 7748 3669 7757
rect 3627 7708 3628 7748
rect 3668 7708 3669 7748
rect 3627 7699 3669 7708
rect 3819 7748 3861 7757
rect 3819 7708 3820 7748
rect 3860 7708 3861 7748
rect 3819 7699 3861 7708
rect 4300 7673 4340 8632
rect 4396 8672 4436 8681
rect 4396 8429 4436 8632
rect 4395 8420 4437 8429
rect 4395 8380 4396 8420
rect 4436 8380 4437 8420
rect 4395 8371 4437 8380
rect 4395 7916 4437 7925
rect 4395 7876 4396 7916
rect 4436 7876 4437 7916
rect 4395 7867 4437 7876
rect 3531 7664 3573 7673
rect 3531 7624 3532 7664
rect 3572 7624 3573 7664
rect 3531 7615 3573 7624
rect 4299 7664 4341 7673
rect 4299 7624 4300 7664
rect 4340 7624 4341 7664
rect 4299 7615 4341 7624
rect 3532 7412 3572 7615
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3628 7412 3668 7421
rect 3532 7372 3628 7412
rect 3628 7363 3668 7372
rect 3819 7412 3861 7421
rect 3819 7372 3820 7412
rect 3860 7372 3861 7412
rect 3819 7363 3861 7372
rect 3435 7328 3477 7337
rect 3435 7288 3436 7328
rect 3476 7288 3477 7328
rect 3435 7279 3477 7288
rect 3436 7160 3476 7169
rect 3436 6245 3476 7120
rect 3820 7160 3860 7363
rect 4107 7328 4149 7337
rect 4107 7288 4108 7328
rect 4148 7288 4149 7328
rect 4107 7279 4149 7288
rect 4011 7244 4053 7253
rect 4011 7204 4012 7244
rect 4052 7204 4053 7244
rect 4011 7195 4053 7204
rect 3820 7111 3860 7120
rect 4012 7160 4052 7195
rect 4012 7109 4052 7120
rect 3915 6992 3957 7001
rect 3915 6952 3916 6992
rect 3956 6952 3957 6992
rect 3915 6943 3957 6952
rect 3916 6858 3956 6943
rect 3723 6488 3765 6497
rect 3723 6448 3724 6488
rect 3764 6448 3765 6488
rect 3723 6439 3765 6448
rect 3820 6488 3860 6497
rect 4108 6488 4148 7279
rect 4396 7244 4436 7867
rect 4492 7421 4532 8800
rect 4684 8420 4724 8875
rect 4972 8765 5012 9043
rect 4971 8756 5013 8765
rect 4971 8716 4972 8756
rect 5012 8716 5013 8756
rect 4971 8707 5013 8716
rect 4780 8672 4820 8683
rect 4780 8597 4820 8632
rect 4875 8672 4917 8681
rect 4875 8632 4876 8672
rect 4916 8632 4917 8672
rect 4875 8623 4917 8632
rect 4779 8588 4821 8597
rect 4779 8548 4780 8588
rect 4820 8548 4821 8588
rect 4779 8539 4821 8548
rect 4876 8538 4916 8623
rect 5260 8504 5300 9640
rect 5356 8681 5396 8766
rect 5355 8672 5397 8681
rect 5355 8632 5356 8672
rect 5396 8632 5397 8672
rect 5355 8623 5397 8632
rect 5452 8513 5492 10144
rect 5547 10184 5589 10193
rect 5547 10144 5548 10184
rect 5588 10144 5589 10184
rect 5547 10135 5589 10144
rect 5548 10050 5588 10135
rect 5644 9932 5684 10312
rect 5739 10312 5740 10352
rect 5780 10312 5781 10352
rect 5739 10303 5781 10312
rect 5739 10100 5781 10109
rect 5739 10060 5740 10100
rect 5780 10060 5781 10100
rect 5739 10051 5781 10060
rect 5548 9892 5684 9932
rect 5451 8504 5493 8513
rect 5260 8464 5396 8504
rect 4684 8380 4820 8420
rect 4588 8000 4628 8009
rect 4588 7589 4628 7960
rect 4684 8000 4724 8009
rect 4587 7580 4629 7589
rect 4587 7540 4588 7580
rect 4628 7540 4629 7580
rect 4587 7531 4629 7540
rect 4491 7412 4533 7421
rect 4491 7372 4492 7412
rect 4532 7372 4533 7412
rect 4491 7363 4533 7372
rect 4396 7204 4532 7244
rect 4203 7160 4245 7169
rect 4203 7120 4204 7160
rect 4244 7120 4245 7160
rect 4203 7111 4245 7120
rect 4204 7026 4244 7111
rect 3860 6448 4148 6488
rect 4204 6488 4244 6497
rect 3820 6439 3860 6448
rect 3724 6354 3764 6439
rect 3435 6236 3477 6245
rect 3435 6196 3436 6236
rect 3476 6196 3477 6236
rect 3435 6187 3477 6196
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 4204 5993 4244 6448
rect 4300 6488 4340 6497
rect 4340 6448 4436 6488
rect 4300 6439 4340 6448
rect 4203 5984 4245 5993
rect 4203 5944 4204 5984
rect 4244 5944 4245 5984
rect 4203 5935 4245 5944
rect 3531 5816 3573 5825
rect 3531 5776 3532 5816
rect 3572 5776 3573 5816
rect 3531 5767 3573 5776
rect 3435 4472 3477 4481
rect 3435 4432 3436 4472
rect 3476 4432 3477 4472
rect 3435 4423 3477 4432
rect 3436 4388 3476 4423
rect 3436 4337 3476 4348
rect 3532 4220 3572 5767
rect 4204 5648 4244 5657
rect 4204 5489 4244 5608
rect 4203 5480 4245 5489
rect 4203 5440 4204 5480
rect 4244 5440 4245 5480
rect 4203 5431 4245 5440
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 3532 4180 3764 4220
rect 3628 4052 3668 4061
rect 3340 4012 3628 4052
rect 3628 4003 3668 4012
rect 3627 3800 3669 3809
rect 3627 3760 3628 3800
rect 3668 3760 3669 3800
rect 3627 3751 3669 3760
rect 3339 3632 3381 3641
rect 3339 3592 3340 3632
rect 3380 3592 3381 3632
rect 3339 3583 3381 3592
rect 3531 3632 3573 3641
rect 3531 3592 3532 3632
rect 3572 3592 3573 3632
rect 3531 3583 3573 3592
rect 3628 3632 3668 3751
rect 3724 3641 3764 4180
rect 3820 4141 3860 4150
rect 3820 4061 3860 4101
rect 4299 4136 4341 4145
rect 4299 4096 4300 4136
rect 4340 4096 4341 4136
rect 4299 4087 4341 4096
rect 3819 4052 3861 4061
rect 3819 4012 3820 4052
rect 3860 4012 3861 4052
rect 3819 4003 3861 4012
rect 3820 3716 3860 4003
rect 4300 4002 4340 4087
rect 4396 3893 4436 6448
rect 4492 6320 4532 7204
rect 4587 6740 4629 6749
rect 4587 6700 4588 6740
rect 4628 6700 4629 6740
rect 4587 6691 4629 6700
rect 4588 6488 4628 6691
rect 4684 6581 4724 7960
rect 4683 6572 4725 6581
rect 4683 6532 4684 6572
rect 4724 6532 4725 6572
rect 4683 6523 4725 6532
rect 4588 6439 4628 6448
rect 4492 6280 4628 6320
rect 4491 6152 4533 6161
rect 4491 6112 4492 6152
rect 4532 6112 4533 6152
rect 4491 6103 4533 6112
rect 4492 5648 4532 6103
rect 4492 5599 4532 5608
rect 4491 4976 4533 4985
rect 4491 4936 4492 4976
rect 4532 4936 4533 4976
rect 4491 4927 4533 4936
rect 4492 4842 4532 4927
rect 4588 4724 4628 6280
rect 4780 6077 4820 8380
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4971 8168 5013 8177
rect 4971 8128 4972 8168
rect 5012 8128 5013 8168
rect 4971 8119 5013 8128
rect 5164 8168 5204 8177
rect 4972 8000 5012 8119
rect 4972 7951 5012 7960
rect 5067 8000 5109 8009
rect 5067 7960 5068 8000
rect 5108 7960 5109 8000
rect 5067 7951 5109 7960
rect 5068 7866 5108 7951
rect 5164 7841 5204 8128
rect 5260 8000 5300 8009
rect 5163 7832 5205 7841
rect 5163 7792 5164 7832
rect 5204 7792 5205 7832
rect 5163 7783 5205 7792
rect 5260 7505 5300 7960
rect 5356 8000 5396 8464
rect 5451 8464 5452 8504
rect 5492 8464 5493 8504
rect 5451 8455 5493 8464
rect 5456 8252 5498 8261
rect 5456 8212 5457 8252
rect 5497 8212 5498 8252
rect 5456 8203 5498 8212
rect 5356 7951 5396 7960
rect 5457 8000 5497 8203
rect 5457 7951 5497 7960
rect 5259 7496 5301 7505
rect 5259 7456 5260 7496
rect 5300 7456 5301 7496
rect 5259 7447 5301 7456
rect 5452 7160 5492 7169
rect 5548 7160 5588 9892
rect 5643 9512 5685 9521
rect 5643 9472 5644 9512
rect 5684 9472 5685 9512
rect 5643 9463 5685 9472
rect 5644 8336 5684 9463
rect 5740 8933 5780 10051
rect 5836 9008 5876 12403
rect 6220 12293 6260 14503
rect 6316 13385 6356 14848
rect 6412 14804 6452 14813
rect 6315 13376 6357 13385
rect 6315 13336 6316 13376
rect 6356 13336 6357 13376
rect 6315 13327 6357 13336
rect 6315 13040 6357 13049
rect 6315 13000 6316 13040
rect 6356 13000 6357 13040
rect 6315 12991 6357 13000
rect 6316 12906 6356 12991
rect 6412 12545 6452 14764
rect 6508 14720 6548 14729
rect 6508 13721 6548 14680
rect 6507 13712 6549 13721
rect 6507 13672 6508 13712
rect 6548 13672 6549 13712
rect 6507 13663 6549 13672
rect 6604 13553 6644 14932
rect 6700 14552 6740 15259
rect 6796 14888 6836 16192
rect 6892 16157 6932 17275
rect 7084 16997 7124 18535
rect 7180 17753 7220 19048
rect 7372 18425 7412 19207
rect 7371 18416 7413 18425
rect 7371 18376 7372 18416
rect 7412 18376 7413 18416
rect 7371 18367 7413 18376
rect 7179 17744 7221 17753
rect 7179 17704 7180 17744
rect 7220 17704 7221 17744
rect 7179 17695 7221 17704
rect 7276 17744 7316 17753
rect 7276 17240 7316 17704
rect 7180 17200 7316 17240
rect 7083 16988 7125 16997
rect 7083 16948 7084 16988
rect 7124 16948 7125 16988
rect 7083 16939 7125 16948
rect 7180 16325 7220 17200
rect 7276 17072 7316 17081
rect 7179 16316 7221 16325
rect 7179 16276 7180 16316
rect 7220 16276 7221 16316
rect 7179 16267 7221 16276
rect 7084 16232 7124 16241
rect 6891 16148 6933 16157
rect 6891 16108 6892 16148
rect 6932 16108 6933 16148
rect 6891 16099 6933 16108
rect 7084 16073 7124 16192
rect 7083 16064 7125 16073
rect 7083 16024 7084 16064
rect 7124 16024 7125 16064
rect 7083 16015 7125 16024
rect 7180 15896 7220 16267
rect 7276 15989 7316 17032
rect 7371 16652 7413 16661
rect 7371 16612 7372 16652
rect 7412 16612 7413 16652
rect 7371 16603 7413 16612
rect 7275 15980 7317 15989
rect 7275 15940 7276 15980
rect 7316 15940 7317 15980
rect 7275 15931 7317 15940
rect 7084 15856 7220 15896
rect 6891 15644 6933 15653
rect 6891 15604 6892 15644
rect 6932 15604 6933 15644
rect 6891 15595 6933 15604
rect 6892 15510 6932 15595
rect 6987 15476 7029 15485
rect 6987 15436 6988 15476
rect 7028 15436 7029 15476
rect 6987 15427 7029 15436
rect 6892 14888 6932 14897
rect 6796 14848 6892 14888
rect 6892 14839 6932 14848
rect 6796 14720 6836 14729
rect 6988 14720 7028 15427
rect 7084 15392 7124 15856
rect 7179 15644 7221 15653
rect 7179 15604 7180 15644
rect 7220 15604 7221 15644
rect 7179 15595 7221 15604
rect 7180 15560 7220 15595
rect 7180 15509 7220 15520
rect 7275 15560 7317 15569
rect 7275 15520 7276 15560
rect 7316 15520 7317 15560
rect 7275 15511 7317 15520
rect 7276 15426 7316 15511
rect 7084 15352 7220 15392
rect 6836 14680 6932 14720
rect 6796 14671 6836 14680
rect 6892 14561 6932 14680
rect 6988 14671 7028 14680
rect 7083 14720 7125 14729
rect 7083 14680 7084 14720
rect 7124 14680 7125 14720
rect 7083 14671 7125 14680
rect 7084 14586 7124 14671
rect 6891 14552 6933 14561
rect 6700 14512 6836 14552
rect 6603 13544 6645 13553
rect 6508 13504 6604 13544
rect 6644 13504 6645 13544
rect 6411 12536 6453 12545
rect 6411 12496 6412 12536
rect 6452 12496 6453 12536
rect 6411 12487 6453 12496
rect 6508 12536 6548 13504
rect 6603 13495 6645 13504
rect 6604 13410 6644 13495
rect 6604 13208 6644 13217
rect 6604 13049 6644 13168
rect 6699 13208 6741 13217
rect 6699 13168 6700 13208
rect 6740 13168 6741 13208
rect 6699 13159 6741 13168
rect 6700 13074 6740 13159
rect 6603 13040 6645 13049
rect 6603 13000 6604 13040
rect 6644 13000 6645 13040
rect 6603 12991 6645 13000
rect 6508 12487 6548 12496
rect 6027 12284 6069 12293
rect 6027 12244 6028 12284
rect 6068 12244 6069 12284
rect 6027 12235 6069 12244
rect 6219 12284 6261 12293
rect 6219 12244 6220 12284
rect 6260 12244 6261 12284
rect 6219 12235 6261 12244
rect 5931 11360 5973 11369
rect 5931 11320 5932 11360
rect 5972 11320 5973 11360
rect 5931 11311 5973 11320
rect 5932 10268 5972 11311
rect 6028 11033 6068 12235
rect 6220 11360 6260 12235
rect 6603 11780 6645 11789
rect 6508 11740 6604 11780
rect 6644 11740 6645 11780
rect 6508 11696 6548 11740
rect 6603 11731 6645 11740
rect 6508 11647 6548 11656
rect 6700 11696 6740 11705
rect 6796 11696 6836 14512
rect 6891 14512 6892 14552
rect 6932 14512 6933 14552
rect 6891 14503 6933 14512
rect 6892 13637 6932 14503
rect 7180 14468 7220 15352
rect 7084 14428 7220 14468
rect 6891 13628 6933 13637
rect 6891 13588 6892 13628
rect 6932 13588 6933 13628
rect 6891 13579 6933 13588
rect 7084 13460 7124 14428
rect 7179 14300 7221 14309
rect 7179 14260 7180 14300
rect 7220 14260 7221 14300
rect 7179 14251 7221 14260
rect 7180 14048 7220 14251
rect 7180 13999 7220 14008
rect 6892 13420 7124 13460
rect 6892 12377 6932 13420
rect 6987 13292 7029 13301
rect 6987 13252 6988 13292
rect 7028 13252 7029 13292
rect 6987 13243 7029 13252
rect 7179 13292 7221 13301
rect 7179 13252 7180 13292
rect 7220 13252 7221 13292
rect 7179 13243 7221 13252
rect 6988 12536 7028 13243
rect 7084 13208 7124 13217
rect 7084 12620 7124 13168
rect 7180 13158 7220 13243
rect 7084 12580 7316 12620
rect 6891 12368 6933 12377
rect 6891 12328 6892 12368
rect 6932 12328 6933 12368
rect 6891 12319 6933 12328
rect 6988 11873 7028 12496
rect 7084 12452 7124 12461
rect 7124 12412 7220 12452
rect 7084 12403 7124 12412
rect 7083 12284 7125 12293
rect 7083 12244 7084 12284
rect 7124 12244 7125 12284
rect 7083 12235 7125 12244
rect 6987 11864 7029 11873
rect 6987 11824 6988 11864
rect 7028 11824 7029 11864
rect 6987 11815 7029 11824
rect 6740 11656 6836 11696
rect 6987 11696 7029 11705
rect 6987 11656 6988 11696
rect 7028 11656 7029 11696
rect 6700 11647 6740 11656
rect 6987 11647 7029 11656
rect 6891 11360 6933 11369
rect 6220 11320 6548 11360
rect 6219 11108 6261 11117
rect 6219 11068 6220 11108
rect 6260 11068 6261 11108
rect 6219 11059 6261 11068
rect 6411 11108 6453 11117
rect 6411 11068 6412 11108
rect 6452 11068 6453 11108
rect 6411 11059 6453 11068
rect 6027 11024 6069 11033
rect 6027 10984 6028 11024
rect 6068 10984 6069 11024
rect 6027 10975 6069 10984
rect 6027 10268 6069 10277
rect 5932 10228 6028 10268
rect 6068 10228 6069 10268
rect 5932 10184 5972 10228
rect 6027 10219 6069 10228
rect 5932 10135 5972 10144
rect 6220 10109 6260 11059
rect 6412 11024 6452 11059
rect 6412 10973 6452 10984
rect 6219 10100 6261 10109
rect 6219 10060 6220 10100
rect 6260 10060 6261 10100
rect 6219 10051 6261 10060
rect 6124 9521 6164 9606
rect 6123 9512 6165 9521
rect 6123 9472 6124 9512
rect 6164 9472 6165 9512
rect 6123 9463 6165 9472
rect 6220 9344 6260 10051
rect 6508 9512 6548 11320
rect 6891 11320 6892 11360
rect 6932 11320 6933 11360
rect 6891 11311 6933 11320
rect 6603 11276 6645 11285
rect 6603 11236 6604 11276
rect 6644 11236 6740 11276
rect 6603 11227 6645 11236
rect 6603 11108 6645 11117
rect 6603 11068 6604 11108
rect 6644 11068 6645 11108
rect 6603 11059 6645 11068
rect 6604 10974 6644 11059
rect 6508 9463 6548 9472
rect 6124 9304 6260 9344
rect 5836 8968 5972 9008
rect 5739 8924 5781 8933
rect 5739 8884 5740 8924
rect 5780 8884 5781 8924
rect 5739 8875 5781 8884
rect 5836 8677 5876 8686
rect 5639 8296 5684 8336
rect 5740 8637 5836 8677
rect 5639 8084 5679 8296
rect 5740 8261 5780 8637
rect 5836 8628 5876 8637
rect 5932 8420 5972 8968
rect 6027 8840 6069 8849
rect 6027 8800 6028 8840
rect 6068 8800 6069 8840
rect 6027 8791 6069 8800
rect 6028 8588 6068 8791
rect 6028 8539 6068 8548
rect 5932 8380 6068 8420
rect 5739 8252 5781 8261
rect 5739 8212 5740 8252
rect 5780 8212 5781 8252
rect 5739 8203 5781 8212
rect 6028 8168 6068 8380
rect 5836 8128 6068 8168
rect 5836 8126 5876 8128
rect 5639 8044 5780 8084
rect 5836 8077 5876 8086
rect 5643 7412 5685 7421
rect 5643 7372 5644 7412
rect 5684 7372 5685 7412
rect 5643 7363 5685 7372
rect 5644 7278 5684 7363
rect 5492 7120 5588 7160
rect 5452 7111 5492 7120
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5548 6245 5588 7120
rect 5643 7076 5685 7085
rect 5643 7036 5644 7076
rect 5684 7036 5685 7076
rect 5643 7027 5685 7036
rect 5547 6236 5589 6245
rect 5547 6196 5548 6236
rect 5588 6196 5589 6236
rect 5547 6187 5589 6196
rect 4779 6068 4821 6077
rect 4779 6028 4780 6068
rect 4820 6028 4821 6068
rect 4779 6019 4821 6028
rect 5355 5984 5397 5993
rect 5355 5944 5356 5984
rect 5396 5944 5397 5984
rect 5355 5935 5397 5944
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 5356 5144 5396 5935
rect 5260 5104 5396 5144
rect 4876 4976 4916 4985
rect 4780 4936 4876 4976
rect 4492 4684 4628 4724
rect 4684 4724 4724 4733
rect 4395 3884 4437 3893
rect 4395 3844 4396 3884
rect 4436 3844 4437 3884
rect 4395 3835 4437 3844
rect 3820 3676 4052 3716
rect 3628 3583 3668 3592
rect 3723 3632 3765 3641
rect 3723 3592 3724 3632
rect 3764 3592 3956 3632
rect 3723 3583 3765 3592
rect 3244 3464 3284 3473
rect 3244 2969 3284 3424
rect 3340 3221 3380 3583
rect 3436 3548 3476 3557
rect 3436 3389 3476 3508
rect 3435 3380 3477 3389
rect 3435 3340 3436 3380
rect 3476 3340 3477 3380
rect 3435 3331 3477 3340
rect 3339 3212 3381 3221
rect 3339 3172 3340 3212
rect 3380 3172 3381 3212
rect 3339 3163 3381 3172
rect 3243 2960 3285 2969
rect 3243 2920 3244 2960
rect 3284 2920 3285 2960
rect 3243 2911 3285 2920
rect 3147 2456 3189 2465
rect 3147 2416 3148 2456
rect 3188 2416 3189 2456
rect 3147 2407 3189 2416
rect 2955 2288 2997 2297
rect 2955 2248 2956 2288
rect 2996 2248 2997 2288
rect 2955 2239 2997 2248
rect 2859 1700 2901 1709
rect 2859 1660 2860 1700
rect 2900 1660 2901 1700
rect 2859 1651 2901 1660
rect 2763 1280 2805 1289
rect 2763 1240 2764 1280
rect 2804 1240 2805 1280
rect 2763 1231 2805 1240
rect 2572 904 2708 944
rect 2572 80 2612 904
rect 2764 80 2804 1231
rect 2956 80 2996 2239
rect 3340 1448 3380 3163
rect 3435 2960 3477 2969
rect 3435 2920 3436 2960
rect 3476 2920 3477 2960
rect 3435 2911 3477 2920
rect 3436 2624 3476 2911
rect 3532 2876 3572 3583
rect 3723 3464 3765 3473
rect 3723 3424 3724 3464
rect 3764 3424 3765 3464
rect 3723 3415 3765 3424
rect 3820 3464 3860 3473
rect 3724 3330 3764 3415
rect 3820 3212 3860 3424
rect 3916 3464 3956 3592
rect 3916 3415 3956 3424
rect 4012 3389 4052 3676
rect 4492 3641 4532 4684
rect 4587 4388 4629 4397
rect 4587 4348 4588 4388
rect 4628 4348 4629 4388
rect 4587 4339 4629 4348
rect 4588 4145 4628 4339
rect 4587 4136 4629 4145
rect 4587 4096 4588 4136
rect 4628 4096 4629 4136
rect 4587 4087 4629 4096
rect 4491 3632 4533 3641
rect 4491 3592 4492 3632
rect 4532 3592 4533 3632
rect 4491 3583 4533 3592
rect 4107 3548 4149 3557
rect 4107 3508 4108 3548
rect 4148 3508 4149 3548
rect 4107 3499 4149 3508
rect 4011 3380 4053 3389
rect 4011 3340 4012 3380
rect 4052 3340 4053 3380
rect 4011 3331 4053 3340
rect 4108 3212 4148 3499
rect 4588 3464 4628 4087
rect 4684 3548 4724 4684
rect 4780 4397 4820 4936
rect 4876 4927 4916 4936
rect 4971 4892 5013 4901
rect 4971 4852 4972 4892
rect 5012 4852 5013 4892
rect 4971 4843 5013 4852
rect 4875 4724 4917 4733
rect 4875 4684 4876 4724
rect 4916 4684 4917 4724
rect 4875 4675 4917 4684
rect 4779 4388 4821 4397
rect 4779 4348 4780 4388
rect 4820 4348 4821 4388
rect 4779 4339 4821 4348
rect 4779 4220 4821 4229
rect 4779 4180 4780 4220
rect 4820 4180 4821 4220
rect 4779 4171 4821 4180
rect 4876 4220 4916 4675
rect 4876 4171 4916 4180
rect 4780 4086 4820 4171
rect 4972 3968 5012 4843
rect 5260 4136 5300 5104
rect 5355 4556 5397 4565
rect 5355 4516 5356 4556
rect 5396 4516 5397 4556
rect 5355 4507 5397 4516
rect 5356 4145 5396 4507
rect 5260 4087 5300 4096
rect 5355 4136 5397 4145
rect 5355 4096 5356 4136
rect 5396 4096 5397 4136
rect 5355 4087 5397 4096
rect 5356 4002 5396 4087
rect 4780 3928 5012 3968
rect 4780 3632 4820 3928
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 5451 3716 5493 3725
rect 5451 3676 5452 3716
rect 5492 3676 5493 3716
rect 5451 3667 5493 3676
rect 4971 3632 5013 3641
rect 4780 3592 4916 3632
rect 4684 3508 4820 3548
rect 4588 3415 4628 3424
rect 4684 3445 4724 3454
rect 4491 3380 4533 3389
rect 4491 3340 4492 3380
rect 4532 3340 4533 3380
rect 4491 3331 4533 3340
rect 4300 3296 4340 3305
rect 4340 3256 4436 3296
rect 4300 3247 4340 3256
rect 3820 3172 4148 3212
rect 4203 3128 4245 3137
rect 4203 3088 4204 3128
rect 4244 3088 4245 3128
rect 4203 3079 4245 3088
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 3628 2876 3668 2885
rect 3532 2836 3628 2876
rect 3531 2708 3573 2717
rect 3531 2668 3532 2708
rect 3572 2668 3573 2708
rect 3531 2659 3573 2668
rect 3436 2575 3476 2584
rect 3435 2456 3477 2465
rect 3435 2416 3436 2456
rect 3476 2416 3477 2456
rect 3435 2407 3477 2416
rect 3436 1952 3476 2407
rect 3436 1903 3476 1912
rect 3340 1408 3476 1448
rect 3051 1364 3093 1373
rect 3051 1324 3052 1364
rect 3092 1324 3093 1364
rect 3051 1315 3093 1324
rect 3052 1112 3092 1315
rect 3339 1280 3381 1289
rect 3339 1240 3340 1280
rect 3380 1240 3381 1280
rect 3436 1280 3476 1408
rect 3532 1364 3572 2659
rect 3628 2633 3668 2836
rect 3627 2624 3669 2633
rect 3627 2584 3628 2624
rect 3668 2584 3669 2624
rect 3627 2575 3669 2584
rect 4012 2540 4052 2549
rect 4012 2213 4052 2500
rect 4204 2456 4244 3079
rect 4204 2407 4244 2416
rect 4396 2624 4436 3256
rect 4107 2288 4149 2297
rect 4107 2248 4108 2288
rect 4148 2248 4149 2288
rect 4107 2239 4149 2248
rect 4011 2204 4053 2213
rect 4011 2164 4012 2204
rect 4052 2164 4053 2204
rect 4011 2155 4053 2164
rect 4011 1952 4053 1961
rect 4011 1912 4012 1952
rect 4052 1912 4053 1952
rect 4011 1903 4053 1912
rect 4108 1952 4148 2239
rect 4396 2213 4436 2584
rect 4492 2624 4532 3331
rect 4684 3221 4724 3405
rect 4683 3212 4725 3221
rect 4683 3172 4684 3212
rect 4724 3172 4725 3212
rect 4683 3163 4725 3172
rect 4780 2717 4820 3508
rect 4876 2792 4916 3592
rect 4971 3592 4972 3632
rect 5012 3592 5013 3632
rect 4971 3583 5013 3592
rect 4972 3221 5012 3583
rect 5068 3380 5108 3389
rect 4971 3212 5013 3221
rect 4971 3172 4972 3212
rect 5012 3172 5013 3212
rect 4971 3163 5013 3172
rect 4972 2885 5012 3163
rect 5068 2960 5108 3340
rect 5164 3380 5204 3389
rect 5204 3340 5396 3380
rect 5164 3331 5204 3340
rect 5068 2920 5204 2960
rect 4971 2876 5013 2885
rect 4971 2836 4972 2876
rect 5012 2836 5013 2876
rect 4971 2827 5013 2836
rect 4876 2743 4916 2752
rect 5067 2792 5109 2801
rect 5067 2752 5068 2792
rect 5108 2752 5109 2792
rect 5067 2743 5109 2752
rect 4779 2708 4821 2717
rect 4779 2668 4780 2708
rect 4820 2668 4821 2708
rect 4779 2659 4821 2668
rect 5068 2708 5108 2743
rect 5068 2657 5108 2668
rect 4492 2575 4532 2584
rect 4780 2540 4820 2549
rect 4587 2456 4629 2465
rect 4587 2416 4588 2456
rect 4628 2416 4629 2456
rect 4587 2407 4629 2416
rect 4491 2372 4533 2381
rect 4491 2332 4492 2372
rect 4532 2332 4533 2372
rect 4491 2323 4533 2332
rect 4203 2204 4245 2213
rect 4203 2164 4204 2204
rect 4244 2164 4245 2204
rect 4203 2155 4245 2164
rect 4395 2204 4437 2213
rect 4395 2164 4396 2204
rect 4436 2164 4437 2204
rect 4395 2155 4437 2164
rect 4108 1903 4148 1912
rect 3628 1793 3668 1878
rect 4012 1818 4052 1903
rect 3627 1784 3669 1793
rect 3627 1744 3628 1784
rect 3668 1744 3669 1784
rect 3627 1735 3669 1744
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 4011 1364 4053 1373
rect 3532 1324 3764 1364
rect 3436 1240 3668 1280
rect 3339 1231 3381 1240
rect 3052 1063 3092 1072
rect 3147 1112 3189 1121
rect 3147 1072 3148 1112
rect 3188 1072 3189 1112
rect 3147 1063 3189 1072
rect 3148 80 3188 1063
rect 3340 80 3380 1231
rect 3532 1117 3572 1126
rect 3436 1077 3532 1112
rect 3436 1072 3572 1077
rect 3436 869 3476 1072
rect 3532 1068 3572 1072
rect 3531 944 3573 953
rect 3531 904 3532 944
rect 3572 904 3573 944
rect 3531 895 3573 904
rect 3435 860 3477 869
rect 3435 820 3436 860
rect 3476 820 3477 860
rect 3435 811 3477 820
rect 3532 80 3572 895
rect 3628 860 3668 1240
rect 3724 1028 3764 1324
rect 4011 1324 4012 1364
rect 4052 1324 4053 1364
rect 4011 1315 4053 1324
rect 3915 1280 3957 1289
rect 3915 1240 3916 1280
rect 3956 1240 3957 1280
rect 3915 1231 3957 1240
rect 3916 1146 3956 1231
rect 3724 979 3764 988
rect 3628 820 3764 860
rect 3724 80 3764 820
rect 4012 776 4052 1315
rect 4204 1289 4244 2155
rect 4492 1952 4532 2323
rect 4492 1903 4532 1912
rect 4588 1868 4628 2407
rect 4299 1532 4341 1541
rect 4299 1492 4300 1532
rect 4340 1492 4341 1532
rect 4299 1483 4341 1492
rect 4203 1280 4245 1289
rect 4203 1240 4204 1280
rect 4244 1240 4245 1280
rect 4203 1231 4245 1240
rect 4204 1146 4244 1231
rect 4107 1112 4149 1121
rect 4107 1072 4108 1112
rect 4148 1072 4149 1112
rect 4107 1063 4149 1072
rect 3916 736 4052 776
rect 3916 80 3956 736
rect 4108 80 4148 1063
rect 4300 80 4340 1483
rect 4588 1448 4628 1828
rect 4492 1408 4628 1448
rect 4492 80 4532 1408
rect 4780 1289 4820 2500
rect 5164 2465 5204 2920
rect 5260 2549 5300 2580
rect 5259 2540 5301 2549
rect 5259 2500 5260 2540
rect 5300 2500 5301 2540
rect 5259 2491 5301 2500
rect 5163 2456 5205 2465
rect 5163 2416 5164 2456
rect 5204 2416 5205 2456
rect 5163 2407 5205 2416
rect 5260 2456 5300 2491
rect 5260 2405 5300 2416
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5067 2120 5109 2129
rect 5067 2080 5068 2120
rect 5108 2080 5109 2120
rect 5067 2071 5109 2080
rect 5068 1952 5108 2071
rect 5068 1903 5108 1912
rect 4684 1280 4724 1289
rect 4779 1280 4821 1289
rect 4724 1240 4780 1280
rect 4820 1240 4821 1280
rect 4684 1231 4724 1240
rect 4779 1231 4821 1240
rect 4780 1146 4820 1231
rect 4876 1196 4916 1205
rect 4683 1112 4725 1121
rect 4683 1072 4684 1112
rect 4724 1072 4725 1112
rect 4683 1063 4725 1072
rect 4684 80 4724 1063
rect 4876 1037 4916 1156
rect 5259 1196 5301 1205
rect 5259 1156 5260 1196
rect 5300 1156 5301 1196
rect 5259 1147 5301 1156
rect 5260 1062 5300 1147
rect 5356 1121 5396 3340
rect 5452 2624 5492 3667
rect 5548 3296 5588 6187
rect 5644 5480 5684 7027
rect 5740 5741 5780 8044
rect 5836 7990 6020 8000
rect 5836 7960 5980 7990
rect 5836 7412 5876 7960
rect 5980 7941 6020 7950
rect 5836 7363 5876 7372
rect 6028 7160 6068 7169
rect 6124 7160 6164 9304
rect 6316 9260 6356 9269
rect 6356 9220 6644 9260
rect 6316 9211 6356 9220
rect 6315 9092 6357 9101
rect 6315 9052 6316 9092
rect 6356 9052 6357 9092
rect 6315 9043 6357 9052
rect 6219 8840 6261 8849
rect 6219 8800 6220 8840
rect 6260 8800 6261 8840
rect 6219 8791 6261 8800
rect 6220 8706 6260 8791
rect 6219 8336 6261 8345
rect 6219 8296 6220 8336
rect 6260 8296 6261 8336
rect 6219 8287 6261 8296
rect 5932 7120 6028 7160
rect 6068 7120 6164 7160
rect 5836 6488 5876 6497
rect 5932 6488 5972 7120
rect 6028 7111 6068 7120
rect 6027 6656 6069 6665
rect 6027 6616 6028 6656
rect 6068 6616 6069 6656
rect 6027 6607 6069 6616
rect 6028 6522 6068 6607
rect 5876 6448 5972 6488
rect 5836 6439 5876 6448
rect 5931 5900 5973 5909
rect 5931 5860 5932 5900
rect 5972 5860 5973 5900
rect 5931 5851 5973 5860
rect 5932 5766 5972 5851
rect 6123 5816 6165 5825
rect 6123 5776 6124 5816
rect 6164 5776 6165 5816
rect 6123 5767 6165 5776
rect 5739 5732 5781 5741
rect 5739 5692 5740 5732
rect 5780 5692 5781 5732
rect 5739 5683 5781 5692
rect 5740 5648 5780 5683
rect 5740 5564 5780 5608
rect 6124 5648 6164 5767
rect 6124 5599 6164 5608
rect 6027 5564 6069 5573
rect 5740 5524 5972 5564
rect 5644 5440 5780 5480
rect 5643 4892 5685 4901
rect 5643 4852 5644 4892
rect 5684 4852 5685 4892
rect 5643 4843 5685 4852
rect 5644 4304 5684 4843
rect 5644 4255 5684 4264
rect 5740 4136 5780 5440
rect 5835 5144 5877 5153
rect 5835 5104 5836 5144
rect 5876 5104 5877 5144
rect 5835 5095 5877 5104
rect 5644 4096 5780 4136
rect 5644 3464 5684 4096
rect 5644 3415 5684 3424
rect 5739 3464 5781 3473
rect 5739 3424 5740 3464
rect 5780 3424 5781 3464
rect 5739 3415 5781 3424
rect 5548 3256 5684 3296
rect 5644 2801 5684 3256
rect 5740 2876 5780 3415
rect 5740 2827 5780 2836
rect 5643 2792 5685 2801
rect 5643 2752 5644 2792
rect 5684 2752 5685 2792
rect 5643 2743 5685 2752
rect 5548 2633 5588 2718
rect 5836 2708 5876 5095
rect 5932 4985 5972 5524
rect 6027 5524 6028 5564
rect 6068 5524 6069 5564
rect 6027 5515 6069 5524
rect 5931 4976 5973 4985
rect 5931 4936 5932 4976
rect 5972 4936 5973 4976
rect 5931 4927 5973 4936
rect 5931 4304 5973 4313
rect 5931 4264 5932 4304
rect 5972 4264 5973 4304
rect 5931 4255 5973 4264
rect 5932 4170 5972 4255
rect 5931 3800 5973 3809
rect 5931 3760 5932 3800
rect 5972 3760 5973 3800
rect 5931 3751 5973 3760
rect 5740 2668 5876 2708
rect 5452 2575 5492 2584
rect 5547 2624 5589 2633
rect 5547 2584 5548 2624
rect 5588 2584 5589 2624
rect 5547 2575 5589 2584
rect 5740 2624 5780 2668
rect 5932 2633 5972 3751
rect 6028 2708 6068 5515
rect 6123 4976 6165 4985
rect 6123 4936 6124 4976
rect 6164 4936 6165 4976
rect 6123 4927 6165 4936
rect 6124 4842 6164 4927
rect 6220 4472 6260 8287
rect 6316 6152 6356 9043
rect 6604 8672 6644 9220
rect 6700 9101 6740 11236
rect 6796 11108 6836 11117
rect 6699 9092 6741 9101
rect 6699 9052 6700 9092
rect 6740 9052 6741 9092
rect 6699 9043 6741 9052
rect 6604 8623 6644 8632
rect 6700 8672 6740 8681
rect 6700 8429 6740 8632
rect 6699 8420 6741 8429
rect 6699 8380 6700 8420
rect 6740 8380 6741 8420
rect 6699 8371 6741 8380
rect 6699 8252 6741 8261
rect 6699 8212 6700 8252
rect 6740 8212 6741 8252
rect 6699 8203 6741 8212
rect 6508 8000 6548 8009
rect 6508 7673 6548 7960
rect 6507 7664 6549 7673
rect 6507 7624 6508 7664
rect 6548 7624 6549 7664
rect 6507 7615 6549 7624
rect 6507 7412 6549 7421
rect 6507 7372 6508 7412
rect 6548 7372 6549 7412
rect 6507 7363 6549 7372
rect 6508 6665 6548 7363
rect 6700 7085 6740 8203
rect 6796 7253 6836 11068
rect 6795 7244 6837 7253
rect 6795 7204 6796 7244
rect 6836 7204 6837 7244
rect 6795 7195 6837 7204
rect 6699 7076 6741 7085
rect 6699 7036 6700 7076
rect 6740 7036 6741 7076
rect 6699 7027 6741 7036
rect 6507 6656 6549 6665
rect 6507 6616 6508 6656
rect 6548 6616 6549 6656
rect 6507 6607 6549 6616
rect 6412 6572 6452 6581
rect 6412 6329 6452 6532
rect 6604 6474 6644 6483
rect 6604 6329 6644 6434
rect 6411 6320 6453 6329
rect 6411 6280 6412 6320
rect 6452 6280 6453 6320
rect 6411 6271 6453 6280
rect 6603 6320 6645 6329
rect 6603 6280 6604 6320
rect 6644 6280 6645 6320
rect 6603 6271 6645 6280
rect 6316 6112 6452 6152
rect 6315 5312 6357 5321
rect 6315 5272 6316 5312
rect 6356 5272 6357 5312
rect 6315 5263 6357 5272
rect 6316 5060 6356 5263
rect 6316 5011 6356 5020
rect 6412 4808 6452 6112
rect 6892 5069 6932 11311
rect 6988 11019 7028 11647
rect 6988 10970 7028 10979
rect 6987 9596 7029 9605
rect 6987 9556 6988 9596
rect 7028 9556 7029 9596
rect 6987 9547 7029 9556
rect 6988 8000 7028 9547
rect 7084 8849 7124 12235
rect 7180 11201 7220 12412
rect 7276 11537 7316 12580
rect 7372 12293 7412 16603
rect 7468 14216 7508 21475
rect 7755 21188 7797 21197
rect 7755 21148 7756 21188
rect 7796 21148 7797 21188
rect 7755 21139 7797 21148
rect 7756 20180 7796 21139
rect 7660 20140 7796 20180
rect 7563 19256 7605 19265
rect 7563 19216 7564 19256
rect 7604 19216 7605 19256
rect 7563 19207 7605 19216
rect 7564 19122 7604 19207
rect 7563 18584 7605 18593
rect 7563 18544 7564 18584
rect 7604 18544 7605 18584
rect 7563 18535 7605 18544
rect 7564 15065 7604 18535
rect 7660 16409 7700 20140
rect 7756 20096 7796 20140
rect 7756 20047 7796 20056
rect 7852 19853 7892 21652
rect 7851 19844 7893 19853
rect 7851 19804 7852 19844
rect 7892 19804 7893 19844
rect 7851 19795 7893 19804
rect 7755 18164 7797 18173
rect 7755 18124 7756 18164
rect 7796 18124 7797 18164
rect 7755 18115 7797 18124
rect 7756 17912 7796 18115
rect 7852 17996 7892 19795
rect 7948 18173 7988 22744
rect 8044 21608 8084 22996
rect 8140 22205 8180 23080
rect 8332 23071 8372 23080
rect 8524 22868 8564 22877
rect 8332 22828 8524 22868
rect 8332 22364 8372 22828
rect 8524 22819 8564 22828
rect 8620 22700 8660 23743
rect 8284 22324 8372 22364
rect 8524 22660 8660 22700
rect 8284 22322 8324 22324
rect 8284 22273 8324 22282
rect 8139 22196 8181 22205
rect 8139 22156 8140 22196
rect 8180 22156 8181 22196
rect 8139 22147 8181 22156
rect 8427 22112 8469 22121
rect 8427 22072 8428 22112
rect 8468 22072 8469 22112
rect 8427 22063 8469 22072
rect 8084 21568 8180 21608
rect 8044 21559 8084 21568
rect 8044 20768 8084 20777
rect 8044 19349 8084 20728
rect 8043 19340 8085 19349
rect 8043 19300 8044 19340
rect 8084 19300 8085 19340
rect 8043 19291 8085 19300
rect 8043 18584 8085 18593
rect 8043 18544 8044 18584
rect 8084 18544 8085 18584
rect 8043 18535 8085 18544
rect 8044 18450 8084 18535
rect 7947 18164 7989 18173
rect 7947 18124 7948 18164
rect 7988 18124 7989 18164
rect 7947 18115 7989 18124
rect 7852 17956 7988 17996
rect 7948 17912 7988 17956
rect 7756 17872 7892 17912
rect 7948 17872 8084 17912
rect 7756 17749 7796 17758
rect 7756 17669 7796 17709
rect 7755 17660 7797 17669
rect 7755 17620 7756 17660
rect 7796 17620 7797 17660
rect 7755 17611 7797 17620
rect 7756 17067 7796 17611
rect 7756 17018 7796 17027
rect 7659 16400 7701 16409
rect 7659 16360 7660 16400
rect 7700 16360 7701 16400
rect 7659 16351 7701 16360
rect 7660 15476 7700 15485
rect 7660 15233 7700 15436
rect 7755 15476 7797 15485
rect 7755 15436 7756 15476
rect 7796 15436 7797 15476
rect 7755 15427 7797 15436
rect 7756 15342 7796 15427
rect 7659 15224 7701 15233
rect 7659 15184 7660 15224
rect 7700 15184 7701 15224
rect 7659 15175 7701 15184
rect 7563 15056 7605 15065
rect 7563 15016 7564 15056
rect 7604 15016 7605 15056
rect 7563 15007 7605 15016
rect 7564 14720 7604 14731
rect 7564 14645 7604 14680
rect 7563 14636 7605 14645
rect 7563 14596 7564 14636
rect 7604 14596 7605 14636
rect 7563 14587 7605 14596
rect 7468 14176 7604 14216
rect 7467 14048 7509 14057
rect 7467 14008 7468 14048
rect 7508 14008 7509 14048
rect 7467 13999 7509 14008
rect 7468 13914 7508 13999
rect 7467 13796 7509 13805
rect 7564 13796 7604 14176
rect 7467 13756 7468 13796
rect 7508 13756 7604 13796
rect 7467 13747 7509 13756
rect 7659 13544 7701 13553
rect 7659 13504 7660 13544
rect 7700 13504 7701 13544
rect 7659 13495 7701 13504
rect 7467 13208 7509 13217
rect 7467 13168 7468 13208
rect 7508 13168 7509 13208
rect 7467 13159 7509 13168
rect 7660 13208 7700 13495
rect 7852 13301 7892 17872
rect 7948 17669 7988 17754
rect 7947 17660 7989 17669
rect 7947 17620 7948 17660
rect 7988 17620 7989 17660
rect 7947 17611 7989 17620
rect 7947 17492 7989 17501
rect 7947 17452 7948 17492
rect 7988 17452 7989 17492
rect 7947 17443 7989 17452
rect 7948 17240 7988 17443
rect 7948 17191 7988 17200
rect 7947 14384 7989 14393
rect 8044 14384 8084 17872
rect 8140 17837 8180 21568
rect 8236 20012 8276 20021
rect 8236 19769 8276 19972
rect 8331 20012 8373 20021
rect 8331 19972 8332 20012
rect 8372 19972 8373 20012
rect 8331 19963 8373 19972
rect 8332 19878 8372 19963
rect 8235 19760 8277 19769
rect 8235 19720 8236 19760
rect 8276 19720 8277 19760
rect 8235 19711 8277 19720
rect 8139 17828 8181 17837
rect 8139 17788 8140 17828
rect 8180 17788 8181 17828
rect 8139 17779 8181 17788
rect 8236 17744 8276 17753
rect 8236 17240 8276 17704
rect 8428 17324 8468 22063
rect 8524 21533 8564 22660
rect 8716 22616 8756 24592
rect 8620 22576 8756 22616
rect 8523 21524 8565 21533
rect 8523 21484 8524 21524
rect 8564 21484 8565 21524
rect 8523 21475 8565 21484
rect 8524 18593 8564 21475
rect 8620 19265 8660 22576
rect 8812 20945 8852 26431
rect 8907 25892 8949 25901
rect 8907 25852 8908 25892
rect 8948 25852 8949 25892
rect 8907 25843 8949 25852
rect 8908 25758 8948 25843
rect 9003 23792 9045 23801
rect 9003 23752 9004 23792
rect 9044 23752 9045 23792
rect 9003 23743 9045 23752
rect 8907 23204 8949 23213
rect 8907 23164 8908 23204
rect 8948 23164 8949 23204
rect 8907 23155 8949 23164
rect 8811 20936 8853 20945
rect 8811 20896 8812 20936
rect 8852 20896 8853 20936
rect 8811 20887 8853 20896
rect 8908 20180 8948 23155
rect 9004 21440 9044 23743
rect 9100 21617 9140 26431
rect 9195 26228 9237 26237
rect 9195 26188 9196 26228
rect 9236 26188 9237 26228
rect 9195 26179 9237 26188
rect 9196 26144 9236 26179
rect 9196 26093 9236 26104
rect 9292 26144 9332 26515
rect 9292 26095 9332 26104
rect 9387 26144 9429 26153
rect 9387 26104 9388 26144
rect 9428 26104 9429 26144
rect 9387 26095 9429 26104
rect 9195 25388 9237 25397
rect 9195 25348 9196 25388
rect 9236 25348 9237 25388
rect 9195 25339 9237 25348
rect 9196 22625 9236 25339
rect 9388 25313 9428 26095
rect 9484 25397 9524 26608
rect 9579 26480 9621 26489
rect 9772 26480 9812 26767
rect 9579 26440 9580 26480
rect 9620 26440 9621 26480
rect 9579 26431 9621 26440
rect 9676 26440 9812 26480
rect 9483 25388 9525 25397
rect 9483 25348 9484 25388
rect 9524 25348 9525 25388
rect 9483 25339 9525 25348
rect 9292 25304 9332 25313
rect 9387 25304 9429 25313
rect 9332 25264 9388 25304
rect 9428 25264 9429 25304
rect 9292 25255 9332 25264
rect 9387 25255 9429 25264
rect 9484 25136 9524 25145
rect 9292 25096 9484 25136
rect 9292 23792 9332 25096
rect 9484 25087 9524 25096
rect 9292 23743 9332 23752
rect 9387 23792 9429 23801
rect 9387 23752 9388 23792
rect 9428 23752 9429 23792
rect 9387 23743 9429 23752
rect 9388 23658 9428 23743
rect 9483 23708 9525 23717
rect 9483 23668 9484 23708
rect 9524 23668 9525 23708
rect 9483 23659 9525 23668
rect 9484 23120 9524 23659
rect 9484 23071 9524 23080
rect 9195 22616 9237 22625
rect 9195 22576 9196 22616
rect 9236 22576 9237 22616
rect 9195 22567 9237 22576
rect 9196 22280 9236 22289
rect 9196 21776 9236 22240
rect 9292 22280 9332 22289
rect 9292 22037 9332 22240
rect 9291 22028 9333 22037
rect 9291 21988 9292 22028
rect 9332 21988 9333 22028
rect 9291 21979 9333 21988
rect 9484 21776 9524 21785
rect 9196 21736 9484 21776
rect 9484 21727 9524 21736
rect 9099 21608 9141 21617
rect 9099 21568 9100 21608
rect 9140 21568 9141 21608
rect 9099 21559 9141 21568
rect 9292 21608 9332 21617
rect 9004 21400 9140 21440
rect 9003 21272 9045 21281
rect 9003 21232 9004 21272
rect 9044 21232 9045 21272
rect 9003 21223 9045 21232
rect 9004 20945 9044 21223
rect 9003 20936 9045 20945
rect 9003 20896 9004 20936
rect 9044 20896 9045 20936
rect 9003 20887 9045 20896
rect 8908 20140 9044 20180
rect 8716 20096 8756 20105
rect 8619 19256 8661 19265
rect 8619 19216 8620 19256
rect 8660 19216 8661 19256
rect 8619 19207 8661 19216
rect 8523 18584 8565 18593
rect 8523 18544 8524 18584
rect 8564 18544 8565 18584
rect 8523 18535 8565 18544
rect 8524 17744 8564 17753
rect 8524 17585 8564 17704
rect 8716 17669 8756 20056
rect 8812 20096 8852 20105
rect 8852 20056 8948 20096
rect 8812 20047 8852 20056
rect 8811 19256 8853 19265
rect 8811 19216 8812 19256
rect 8852 19216 8853 19256
rect 8811 19207 8853 19216
rect 8812 19122 8852 19207
rect 8908 18761 8948 20056
rect 8907 18752 8949 18761
rect 8907 18712 8908 18752
rect 8948 18712 8949 18752
rect 8907 18703 8949 18712
rect 8908 17912 8948 17921
rect 8620 17660 8660 17669
rect 8523 17576 8565 17585
rect 8523 17536 8524 17576
rect 8564 17536 8565 17576
rect 8523 17527 8565 17536
rect 8620 17501 8660 17620
rect 8715 17660 8757 17669
rect 8715 17620 8716 17660
rect 8756 17620 8757 17660
rect 8715 17611 8757 17620
rect 8619 17492 8661 17501
rect 8619 17452 8620 17492
rect 8660 17452 8661 17492
rect 8619 17443 8661 17452
rect 8428 17284 8660 17324
rect 8236 17200 8564 17240
rect 8235 17072 8277 17081
rect 8235 17032 8236 17072
rect 8276 17032 8277 17072
rect 8235 17023 8277 17032
rect 8236 16938 8276 17023
rect 8140 16820 8180 16829
rect 8140 16241 8180 16780
rect 8235 16820 8277 16829
rect 8235 16780 8236 16820
rect 8276 16780 8277 16820
rect 8235 16771 8277 16780
rect 8139 16232 8181 16241
rect 8139 16192 8140 16232
rect 8180 16192 8181 16232
rect 8139 16183 8181 16192
rect 8236 15560 8276 16771
rect 8427 16568 8469 16577
rect 8427 16528 8428 16568
rect 8468 16528 8469 16568
rect 8427 16519 8469 16528
rect 8236 15511 8276 15520
rect 8332 16232 8372 16241
rect 8332 14897 8372 16192
rect 8331 14888 8373 14897
rect 8331 14848 8332 14888
rect 8372 14848 8373 14888
rect 8331 14839 8373 14848
rect 8332 14561 8372 14839
rect 8331 14552 8373 14561
rect 8331 14512 8332 14552
rect 8372 14512 8373 14552
rect 8331 14503 8373 14512
rect 7947 14344 7948 14384
rect 7988 14344 8084 14384
rect 7947 14335 7989 14344
rect 7851 13292 7893 13301
rect 7851 13252 7852 13292
rect 7892 13252 7893 13292
rect 7851 13243 7893 13252
rect 7660 13159 7700 13168
rect 7468 12536 7508 13159
rect 7563 12620 7605 12629
rect 7563 12580 7564 12620
rect 7604 12580 7605 12620
rect 7563 12571 7605 12580
rect 7371 12284 7413 12293
rect 7371 12244 7372 12284
rect 7412 12244 7413 12284
rect 7371 12235 7413 12244
rect 7371 11696 7413 11705
rect 7371 11656 7372 11696
rect 7412 11656 7413 11696
rect 7371 11647 7413 11656
rect 7275 11528 7317 11537
rect 7275 11488 7276 11528
rect 7316 11488 7317 11528
rect 7275 11479 7317 11488
rect 7275 11276 7317 11285
rect 7275 11236 7276 11276
rect 7316 11236 7317 11276
rect 7275 11227 7317 11236
rect 7179 11192 7221 11201
rect 7179 11152 7180 11192
rect 7220 11152 7221 11192
rect 7179 11143 7221 11152
rect 7180 10184 7220 10195
rect 7180 10109 7220 10144
rect 7179 10100 7221 10109
rect 7179 10060 7180 10100
rect 7220 10060 7221 10100
rect 7179 10051 7221 10060
rect 7276 9773 7316 11227
rect 7372 10100 7412 11647
rect 7468 11369 7508 12496
rect 7564 12536 7604 12571
rect 7852 12536 7892 12545
rect 7564 12485 7604 12496
rect 7756 12496 7852 12536
rect 7563 11612 7605 11621
rect 7563 11572 7564 11612
rect 7604 11572 7605 11612
rect 7563 11563 7605 11572
rect 7467 11360 7509 11369
rect 7467 11320 7468 11360
rect 7508 11320 7509 11360
rect 7467 11311 7509 11320
rect 7468 11024 7508 11033
rect 7468 10613 7508 10984
rect 7467 10604 7509 10613
rect 7467 10564 7468 10604
rect 7508 10564 7509 10604
rect 7467 10555 7509 10564
rect 7275 9764 7317 9773
rect 7275 9724 7276 9764
rect 7316 9724 7317 9764
rect 7275 9715 7317 9724
rect 7083 8840 7125 8849
rect 7083 8800 7084 8840
rect 7124 8800 7125 8840
rect 7083 8791 7125 8800
rect 7084 8672 7124 8681
rect 7084 8597 7124 8632
rect 7180 8672 7220 8681
rect 7276 8672 7316 9715
rect 7220 8632 7316 8672
rect 7180 8623 7220 8632
rect 7083 8588 7125 8597
rect 7083 8548 7084 8588
rect 7124 8548 7125 8588
rect 7083 8539 7125 8548
rect 7084 8345 7124 8539
rect 7179 8504 7221 8513
rect 7179 8464 7180 8504
rect 7220 8464 7221 8504
rect 7179 8455 7221 8464
rect 7083 8336 7125 8345
rect 7083 8296 7084 8336
rect 7124 8296 7125 8336
rect 7083 8287 7125 8296
rect 7083 8168 7125 8177
rect 7083 8128 7084 8168
rect 7124 8128 7125 8168
rect 7083 8119 7125 8128
rect 6988 7951 7028 7960
rect 7084 8000 7124 8119
rect 7084 7951 7124 7960
rect 7083 7832 7125 7841
rect 7083 7792 7084 7832
rect 7124 7792 7125 7832
rect 7083 7783 7125 7792
rect 7084 6488 7124 7783
rect 7084 6439 7124 6448
rect 7180 5153 7220 8455
rect 7276 7580 7316 8632
rect 7372 7757 7412 10060
rect 7564 8504 7604 11563
rect 7659 11276 7701 11285
rect 7659 11236 7660 11276
rect 7700 11236 7701 11276
rect 7659 11227 7701 11236
rect 7660 10697 7700 11227
rect 7659 10688 7701 10697
rect 7659 10648 7660 10688
rect 7700 10648 7701 10688
rect 7659 10639 7701 10648
rect 7660 9344 7700 10639
rect 7756 10184 7796 12496
rect 7852 12487 7892 12496
rect 7852 12284 7892 12293
rect 7852 10352 7892 12244
rect 7948 11873 7988 14335
rect 8188 13217 8228 13226
rect 8228 13177 8276 13208
rect 8188 13168 8276 13177
rect 8044 12536 8084 12545
rect 7947 11864 7989 11873
rect 7947 11824 7948 11864
rect 7988 11824 7989 11864
rect 7947 11815 7989 11824
rect 7947 11696 7989 11705
rect 7947 11656 7948 11696
rect 7988 11656 7989 11696
rect 7947 11647 7989 11656
rect 7948 11562 7988 11647
rect 7947 11276 7989 11285
rect 7947 11236 7948 11276
rect 7988 11236 7989 11276
rect 7947 11227 7989 11236
rect 7948 11024 7988 11227
rect 8044 11117 8084 12496
rect 8140 12536 8180 12545
rect 8140 12377 8180 12496
rect 8139 12368 8181 12377
rect 8139 12328 8140 12368
rect 8180 12328 8181 12368
rect 8139 12319 8181 12328
rect 8140 11864 8180 11873
rect 8236 11864 8276 13168
rect 8331 13124 8373 13133
rect 8331 13084 8332 13124
rect 8372 13084 8373 13124
rect 8331 13075 8373 13084
rect 8332 12990 8372 13075
rect 8428 12956 8468 16519
rect 8524 16400 8564 17200
rect 8524 16351 8564 16360
rect 8620 16232 8660 17284
rect 8715 17156 8757 17165
rect 8715 17116 8716 17156
rect 8756 17116 8757 17156
rect 8715 17107 8757 17116
rect 8716 17072 8756 17107
rect 8716 17021 8756 17032
rect 8908 16745 8948 17872
rect 9004 17417 9044 20140
rect 9100 17912 9140 21400
rect 9292 20768 9332 21568
rect 9387 21608 9429 21617
rect 9387 21568 9388 21608
rect 9428 21568 9429 21608
rect 9387 21559 9429 21568
rect 9195 20516 9237 20525
rect 9195 20476 9196 20516
rect 9236 20476 9237 20516
rect 9195 20467 9237 20476
rect 9196 20105 9236 20467
rect 9195 20096 9237 20105
rect 9195 20056 9196 20096
rect 9236 20056 9237 20096
rect 9195 20047 9237 20056
rect 9196 18929 9236 20047
rect 9195 18920 9237 18929
rect 9195 18880 9196 18920
rect 9236 18880 9237 18920
rect 9195 18871 9237 18880
rect 9292 18593 9332 20728
rect 9388 19601 9428 21559
rect 9580 21365 9620 26431
rect 9676 26144 9716 26440
rect 9868 26153 9908 29128
rect 9964 28757 10004 29800
rect 10156 29791 10196 29800
rect 10252 29252 10292 31387
rect 10348 31352 10388 31363
rect 10444 31352 10484 32488
rect 10539 32360 10581 32369
rect 10539 32320 10540 32360
rect 10580 32320 10581 32360
rect 10539 32311 10581 32320
rect 10540 32117 10580 32311
rect 10539 32108 10581 32117
rect 10539 32068 10540 32108
rect 10580 32068 10581 32108
rect 10539 32059 10581 32068
rect 10635 32024 10677 32033
rect 10635 31984 10636 32024
rect 10676 31984 10677 32024
rect 10635 31975 10677 31984
rect 10540 31520 10580 31529
rect 10636 31520 10676 31975
rect 10732 31529 10772 34168
rect 10923 34168 10924 34208
rect 10964 34168 10965 34208
rect 10923 34159 10965 34168
rect 10924 33461 10964 34159
rect 10923 33452 10965 33461
rect 10923 33412 10924 33452
rect 10964 33412 10965 33452
rect 10923 33403 10965 33412
rect 10827 32696 10869 32705
rect 10827 32656 10828 32696
rect 10868 32656 10869 32696
rect 10827 32647 10869 32656
rect 10828 32285 10868 32647
rect 11116 32528 11156 34504
rect 11212 32537 11252 35335
rect 11308 35216 11348 35225
rect 11308 34973 11348 35176
rect 11307 34964 11349 34973
rect 11307 34924 11308 34964
rect 11348 34924 11349 34964
rect 11307 34915 11349 34924
rect 11308 33881 11348 34915
rect 11404 34805 11444 41224
rect 11980 41215 12020 41224
rect 11979 41096 12021 41105
rect 11979 41056 11980 41096
rect 12020 41056 12021 41096
rect 11979 41047 12021 41056
rect 11499 40844 11541 40853
rect 11499 40804 11500 40844
rect 11540 40804 11541 40844
rect 11499 40795 11541 40804
rect 11500 37661 11540 40795
rect 11980 40424 12020 41047
rect 11884 39752 11924 39761
rect 11980 39752 12020 40384
rect 12076 40181 12116 41560
rect 12363 41551 12405 41560
rect 12364 41264 12404 41273
rect 12172 41012 12212 41021
rect 12212 40972 12308 41012
rect 12172 40963 12212 40972
rect 12171 40676 12213 40685
rect 12171 40636 12172 40676
rect 12212 40636 12213 40676
rect 12171 40627 12213 40636
rect 12172 40542 12212 40627
rect 12075 40172 12117 40181
rect 12075 40132 12076 40172
rect 12116 40132 12117 40172
rect 12075 40123 12117 40132
rect 12171 40004 12213 40013
rect 12171 39964 12172 40004
rect 12212 39964 12213 40004
rect 12171 39955 12213 39964
rect 12075 39836 12117 39845
rect 12075 39796 12076 39836
rect 12116 39796 12117 39836
rect 12075 39787 12117 39796
rect 11924 39712 12020 39752
rect 11595 39164 11637 39173
rect 11595 39124 11596 39164
rect 11636 39124 11637 39164
rect 11595 39115 11637 39124
rect 11499 37652 11541 37661
rect 11499 37612 11500 37652
rect 11540 37612 11541 37652
rect 11499 37603 11541 37612
rect 11499 37400 11541 37409
rect 11499 37360 11500 37400
rect 11540 37360 11541 37400
rect 11499 37351 11541 37360
rect 11500 36569 11540 37351
rect 11596 36989 11636 39115
rect 11788 38912 11828 38921
rect 11884 38912 11924 39712
rect 12076 39702 12116 39787
rect 11979 39500 12021 39509
rect 11979 39460 11980 39500
rect 12020 39460 12021 39500
rect 11979 39451 12021 39460
rect 11828 38872 11924 38912
rect 11691 38240 11733 38249
rect 11691 38200 11692 38240
rect 11732 38200 11733 38240
rect 11691 38191 11733 38200
rect 11692 37400 11732 38191
rect 11595 36980 11637 36989
rect 11595 36940 11596 36980
rect 11636 36940 11637 36980
rect 11595 36931 11637 36940
rect 11596 36714 11636 36723
rect 11499 36560 11541 36569
rect 11499 36520 11500 36560
rect 11540 36520 11541 36560
rect 11499 36511 11541 36520
rect 11596 36149 11636 36674
rect 11595 36140 11637 36149
rect 11595 36100 11596 36140
rect 11636 36100 11637 36140
rect 11595 36091 11637 36100
rect 11692 36056 11732 37360
rect 11788 37064 11828 38872
rect 11980 38828 12020 39451
rect 12172 39341 12212 39955
rect 12171 39332 12213 39341
rect 12171 39292 12172 39332
rect 12212 39292 12213 39332
rect 12171 39283 12213 39292
rect 11980 38501 12020 38788
rect 12172 38744 12212 38753
rect 11979 38492 12021 38501
rect 11979 38452 11980 38492
rect 12020 38452 12021 38492
rect 11979 38443 12021 38452
rect 11884 37232 11924 37241
rect 12076 37232 12116 37241
rect 11924 37192 12020 37232
rect 11884 37183 11924 37192
rect 11788 37024 11924 37064
rect 11788 36821 11828 36906
rect 11787 36812 11829 36821
rect 11787 36772 11788 36812
rect 11828 36772 11829 36812
rect 11787 36763 11829 36772
rect 11787 36056 11829 36065
rect 11692 36016 11788 36056
rect 11828 36016 11829 36056
rect 11787 36007 11829 36016
rect 11788 35888 11828 36007
rect 11788 35839 11828 35848
rect 11596 35216 11636 35225
rect 11403 34796 11445 34805
rect 11403 34756 11404 34796
rect 11444 34756 11445 34796
rect 11403 34747 11445 34756
rect 11499 34712 11541 34721
rect 11499 34672 11500 34712
rect 11540 34672 11541 34712
rect 11499 34663 11541 34672
rect 11500 34469 11540 34663
rect 11499 34460 11541 34469
rect 11499 34420 11500 34460
rect 11540 34420 11541 34460
rect 11499 34411 11541 34420
rect 11403 34376 11445 34385
rect 11403 34336 11404 34376
rect 11444 34336 11445 34376
rect 11403 34327 11445 34336
rect 11404 34242 11444 34327
rect 11500 34326 11540 34411
rect 11307 33872 11349 33881
rect 11307 33832 11308 33872
rect 11348 33832 11349 33872
rect 11307 33823 11349 33832
rect 11596 33704 11636 35176
rect 11691 34040 11733 34049
rect 11691 34000 11692 34040
rect 11732 34000 11733 34040
rect 11691 33991 11733 34000
rect 11404 33664 11636 33704
rect 11404 33620 11444 33664
rect 11308 33580 11444 33620
rect 11308 33116 11348 33580
rect 11308 33067 11348 33076
rect 11595 32864 11637 32873
rect 11595 32824 11596 32864
rect 11636 32824 11637 32864
rect 11595 32815 11637 32824
rect 11596 32730 11636 32815
rect 11020 32488 11156 32528
rect 11211 32528 11253 32537
rect 11211 32488 11212 32528
rect 11252 32488 11253 32528
rect 10827 32276 10869 32285
rect 10827 32236 10828 32276
rect 10868 32236 10869 32276
rect 10827 32227 10869 32236
rect 10828 32192 10868 32227
rect 10828 32141 10868 32152
rect 10580 31480 10676 31520
rect 10731 31520 10773 31529
rect 10731 31480 10732 31520
rect 10772 31480 10773 31520
rect 10540 31471 10580 31480
rect 10731 31471 10773 31480
rect 10924 31352 10964 31363
rect 10444 31312 10676 31352
rect 10348 31277 10388 31312
rect 10347 31268 10389 31277
rect 10347 31228 10348 31268
rect 10388 31228 10389 31268
rect 10347 31219 10389 31228
rect 10348 30605 10388 31219
rect 10443 31184 10485 31193
rect 10443 31144 10444 31184
rect 10484 31144 10485 31184
rect 10443 31135 10485 31144
rect 10347 30596 10389 30605
rect 10347 30556 10348 30596
rect 10388 30556 10389 30596
rect 10347 30547 10389 30556
rect 10156 29212 10292 29252
rect 10060 28916 10100 28925
rect 9963 28748 10005 28757
rect 9963 28708 9964 28748
rect 10004 28708 10005 28748
rect 9963 28699 10005 28708
rect 9963 27320 10005 27329
rect 9963 27280 9964 27320
rect 10004 27280 10005 27320
rect 9963 27271 10005 27280
rect 9676 26095 9716 26104
rect 9867 26144 9909 26153
rect 9867 26104 9868 26144
rect 9908 26104 9909 26144
rect 9867 26095 9909 26104
rect 9772 26060 9812 26069
rect 9772 25892 9812 26020
rect 9676 25852 9812 25892
rect 9676 24473 9716 25852
rect 9964 25808 10004 27271
rect 10060 26816 10100 28876
rect 10156 27656 10196 29212
rect 10252 29168 10292 29212
rect 10348 29168 10388 29177
rect 10252 29128 10348 29168
rect 10348 29119 10388 29128
rect 10444 29000 10484 31135
rect 10539 30428 10581 30437
rect 10539 30388 10540 30428
rect 10580 30388 10581 30428
rect 10539 30379 10581 30388
rect 10348 28960 10484 29000
rect 10348 28001 10388 28960
rect 10444 28328 10484 28337
rect 10347 27992 10389 28001
rect 10347 27952 10348 27992
rect 10388 27952 10389 27992
rect 10347 27943 10389 27952
rect 10444 27824 10484 28288
rect 10156 26993 10196 27616
rect 10252 27784 10484 27824
rect 10155 26984 10197 26993
rect 10155 26944 10156 26984
rect 10196 26944 10197 26984
rect 10155 26935 10197 26944
rect 10060 26767 10100 26776
rect 10156 26816 10196 26825
rect 9772 25768 10004 25808
rect 9675 24464 9717 24473
rect 9675 24424 9676 24464
rect 9716 24424 9717 24464
rect 9675 24415 9717 24424
rect 9772 23885 9812 25768
rect 10059 25724 10101 25733
rect 10059 25684 10060 25724
rect 10100 25684 10101 25724
rect 10059 25675 10101 25684
rect 9963 25304 10005 25313
rect 9963 25264 9964 25304
rect 10004 25264 10005 25304
rect 9963 25255 10005 25264
rect 9964 24632 10004 25255
rect 10060 24641 10100 25675
rect 10156 24725 10196 26776
rect 10252 26573 10292 27784
rect 10540 27572 10580 30379
rect 10636 29000 10676 31312
rect 10924 31277 10964 31312
rect 10923 31268 10965 31277
rect 10923 31228 10924 31268
rect 10964 31228 10965 31268
rect 10923 31219 10965 31228
rect 10924 31109 10964 31219
rect 11020 31193 11060 32488
rect 11211 32479 11253 32488
rect 11403 32444 11445 32453
rect 11692 32444 11732 33991
rect 11788 33713 11828 33778
rect 11884 33713 11924 37024
rect 11980 36728 12020 37192
rect 12076 36905 12116 37192
rect 12075 36896 12117 36905
rect 12075 36856 12076 36896
rect 12116 36856 12117 36896
rect 12172 36896 12212 38704
rect 12268 38333 12308 40972
rect 12364 40181 12404 41224
rect 12748 40853 12788 42928
rect 12747 40844 12789 40853
rect 12747 40804 12748 40844
rect 12788 40804 12789 40844
rect 12747 40795 12789 40804
rect 12460 40424 12500 40433
rect 12363 40172 12405 40181
rect 12363 40132 12364 40172
rect 12404 40132 12405 40172
rect 12363 40123 12405 40132
rect 12364 40013 12404 40123
rect 12363 40004 12405 40013
rect 12363 39964 12364 40004
rect 12404 39964 12405 40004
rect 12363 39955 12405 39964
rect 12364 39752 12404 39761
rect 12364 39173 12404 39712
rect 12460 39509 12500 40384
rect 12748 40424 12788 40433
rect 12555 40004 12597 40013
rect 12555 39964 12556 40004
rect 12596 39964 12597 40004
rect 12555 39955 12597 39964
rect 12556 39761 12596 39955
rect 12748 39920 12788 40384
rect 12844 40340 12884 40349
rect 12844 40181 12884 40300
rect 12843 40172 12885 40181
rect 12843 40132 12844 40172
rect 12884 40132 12885 40172
rect 12843 40123 12885 40132
rect 12940 40004 12980 42928
rect 13132 40760 13172 42928
rect 13324 42197 13364 42928
rect 13323 42188 13365 42197
rect 13323 42148 13324 42188
rect 13364 42148 13365 42188
rect 13323 42139 13365 42148
rect 13516 42113 13556 42928
rect 13515 42104 13557 42113
rect 13515 42064 13516 42104
rect 13556 42064 13557 42104
rect 13515 42055 13557 42064
rect 13708 42029 13748 42928
rect 13900 42281 13940 42928
rect 13899 42272 13941 42281
rect 13899 42232 13900 42272
rect 13940 42232 13941 42272
rect 13899 42223 13941 42232
rect 13707 42020 13749 42029
rect 13707 41980 13708 42020
rect 13748 41980 13749 42020
rect 13707 41971 13749 41980
rect 13612 41264 13652 41273
rect 13996 41264 14036 41273
rect 13132 40720 13268 40760
rect 13131 40592 13173 40601
rect 13131 40552 13132 40592
rect 13172 40552 13173 40592
rect 13131 40543 13173 40552
rect 13132 40458 13172 40543
rect 12940 39964 13172 40004
rect 12748 39880 12980 39920
rect 12555 39752 12597 39761
rect 12555 39712 12556 39752
rect 12596 39712 12597 39752
rect 12555 39703 12597 39712
rect 12652 39752 12692 39761
rect 12459 39500 12501 39509
rect 12459 39460 12460 39500
rect 12500 39460 12501 39500
rect 12459 39451 12501 39460
rect 12555 39332 12597 39341
rect 12555 39292 12556 39332
rect 12596 39292 12597 39332
rect 12555 39283 12597 39292
rect 12363 39164 12405 39173
rect 12363 39124 12364 39164
rect 12404 39124 12405 39164
rect 12363 39115 12405 39124
rect 12364 38912 12404 38921
rect 12364 38828 12404 38872
rect 12556 38828 12596 39283
rect 12364 38788 12596 38828
rect 12267 38324 12309 38333
rect 12267 38284 12268 38324
rect 12308 38284 12309 38324
rect 12267 38275 12309 38284
rect 12363 38240 12405 38249
rect 12363 38200 12364 38240
rect 12404 38200 12405 38240
rect 12363 38191 12405 38200
rect 12555 38240 12597 38249
rect 12555 38200 12556 38240
rect 12596 38200 12597 38240
rect 12555 38191 12597 38200
rect 12364 38106 12404 38191
rect 12556 38106 12596 38191
rect 12363 37988 12405 37997
rect 12363 37948 12364 37988
rect 12404 37948 12405 37988
rect 12363 37939 12405 37948
rect 12267 37400 12309 37409
rect 12267 37360 12268 37400
rect 12308 37360 12309 37400
rect 12267 37351 12309 37360
rect 12268 37266 12308 37351
rect 12172 36856 12308 36896
rect 12075 36847 12117 36856
rect 12076 36728 12116 36737
rect 11980 36688 12076 36728
rect 12076 36679 12116 36688
rect 12171 36728 12213 36737
rect 12171 36688 12172 36728
rect 12212 36688 12213 36728
rect 12171 36679 12213 36688
rect 12172 36594 12212 36679
rect 12075 36560 12117 36569
rect 12075 36520 12076 36560
rect 12116 36520 12117 36560
rect 12075 36511 12117 36520
rect 11979 36140 12021 36149
rect 11979 36100 11980 36140
rect 12020 36100 12021 36140
rect 11979 36091 12021 36100
rect 11980 36006 12020 36091
rect 11979 34628 12021 34637
rect 11979 34588 11980 34628
rect 12020 34588 12021 34628
rect 11979 34579 12021 34588
rect 11980 34385 12020 34579
rect 11979 34376 12021 34385
rect 11979 34336 11980 34376
rect 12020 34336 12021 34376
rect 11979 34327 12021 34336
rect 12076 34376 12116 36511
rect 12171 36392 12213 36401
rect 12171 36352 12172 36392
rect 12212 36352 12213 36392
rect 12171 36343 12213 36352
rect 12172 34637 12212 36343
rect 12171 34628 12213 34637
rect 12171 34588 12172 34628
rect 12212 34588 12213 34628
rect 12171 34579 12213 34588
rect 12268 34553 12308 36856
rect 12364 36737 12404 37939
rect 12459 37736 12501 37745
rect 12459 37696 12460 37736
rect 12500 37696 12501 37736
rect 12459 37687 12501 37696
rect 12363 36728 12405 36737
rect 12363 36688 12364 36728
rect 12404 36688 12405 36728
rect 12363 36679 12405 36688
rect 12363 36224 12405 36233
rect 12363 36184 12364 36224
rect 12404 36184 12405 36224
rect 12363 36175 12405 36184
rect 12364 35888 12404 36175
rect 12364 35839 12404 35848
rect 12460 35300 12500 37687
rect 12652 37325 12692 39712
rect 12748 39752 12788 39761
rect 12748 38417 12788 39712
rect 12940 39080 12980 39880
rect 13035 39752 13077 39761
rect 13035 39712 13036 39752
rect 13076 39712 13077 39752
rect 13035 39703 13077 39712
rect 13036 39584 13076 39703
rect 13036 39535 13076 39544
rect 12940 39040 13076 39080
rect 12747 38408 12789 38417
rect 12747 38368 12748 38408
rect 12788 38368 12789 38408
rect 12747 38359 12789 38368
rect 12748 38240 12788 38249
rect 12940 38240 12980 38249
rect 12788 38200 12884 38240
rect 12748 38191 12788 38200
rect 12747 38072 12789 38081
rect 12747 38032 12748 38072
rect 12788 38032 12789 38072
rect 12747 38023 12789 38032
rect 12748 37938 12788 38023
rect 12844 37661 12884 38200
rect 12843 37652 12885 37661
rect 12843 37612 12844 37652
rect 12884 37612 12885 37652
rect 12843 37603 12885 37612
rect 12940 37493 12980 38200
rect 12939 37484 12981 37493
rect 12939 37444 12940 37484
rect 12980 37444 12981 37484
rect 12939 37435 12981 37444
rect 12651 37316 12693 37325
rect 12651 37276 12652 37316
rect 12692 37276 12693 37316
rect 12651 37267 12693 37276
rect 12651 37148 12693 37157
rect 12651 37108 12652 37148
rect 12692 37108 12693 37148
rect 12651 37099 12693 37108
rect 12555 36728 12597 36737
rect 12555 36688 12556 36728
rect 12596 36688 12597 36728
rect 12555 36679 12597 36688
rect 12556 36594 12596 36679
rect 12652 36644 12692 37099
rect 13036 36980 13076 39040
rect 13132 38921 13172 39964
rect 13131 38912 13173 38921
rect 13131 38872 13132 38912
rect 13172 38872 13173 38912
rect 13131 38863 13173 38872
rect 13132 37997 13172 38863
rect 13131 37988 13173 37997
rect 13131 37948 13132 37988
rect 13172 37948 13173 37988
rect 13131 37939 13173 37948
rect 13131 37400 13173 37409
rect 13131 37360 13132 37400
rect 13172 37360 13173 37400
rect 13131 37351 13173 37360
rect 12555 36392 12597 36401
rect 12652 36392 12692 36604
rect 12555 36352 12556 36392
rect 12596 36352 12692 36392
rect 12844 36940 13076 36980
rect 12555 36343 12597 36352
rect 12844 36149 12884 36940
rect 13132 36896 13172 37351
rect 12940 36856 13172 36896
rect 12843 36140 12885 36149
rect 12843 36100 12844 36140
rect 12884 36100 12885 36140
rect 12843 36091 12885 36100
rect 12555 36056 12597 36065
rect 12555 36016 12556 36056
rect 12596 36016 12597 36056
rect 12555 36007 12597 36016
rect 12460 35251 12500 35260
rect 12267 34544 12309 34553
rect 12267 34504 12268 34544
rect 12308 34504 12309 34544
rect 12267 34495 12309 34504
rect 12460 34381 12500 34390
rect 12076 34341 12460 34376
rect 12076 34336 12500 34341
rect 11980 34242 12020 34327
rect 12076 33881 12116 34336
rect 12460 34332 12500 34336
rect 12363 34040 12405 34049
rect 12363 34000 12364 34040
rect 12404 34000 12405 34040
rect 12363 33991 12405 34000
rect 11980 33872 12020 33881
rect 12075 33872 12117 33881
rect 12020 33832 12076 33872
rect 12116 33832 12117 33872
rect 11980 33823 12020 33832
rect 12075 33823 12117 33832
rect 12076 33738 12116 33823
rect 11787 33704 11829 33713
rect 11787 33655 11788 33704
rect 11828 33655 11829 33704
rect 11883 33704 11925 33713
rect 11883 33664 11884 33704
rect 11924 33664 11925 33704
rect 11883 33655 11925 33664
rect 12364 33704 12404 33991
rect 11788 33634 11828 33643
rect 12364 33209 12404 33664
rect 12363 33200 12405 33209
rect 12363 33160 12364 33200
rect 12404 33160 12405 33200
rect 12363 33151 12405 33160
rect 12364 33032 12404 33041
rect 11403 32404 11404 32444
rect 11444 32404 11445 32444
rect 11403 32395 11445 32404
rect 11596 32404 11732 32444
rect 11788 32992 12364 33032
rect 11115 32360 11157 32369
rect 11115 32320 11116 32360
rect 11156 32320 11157 32360
rect 11115 32311 11157 32320
rect 11116 32192 11156 32311
rect 11116 32143 11156 32152
rect 11212 32192 11252 32201
rect 11212 31613 11252 32152
rect 11211 31604 11253 31613
rect 11211 31564 11212 31604
rect 11252 31564 11253 31604
rect 11211 31555 11253 31564
rect 11307 31352 11349 31361
rect 11307 31312 11308 31352
rect 11348 31312 11349 31352
rect 11307 31303 11349 31312
rect 11019 31184 11061 31193
rect 11019 31144 11020 31184
rect 11060 31144 11061 31184
rect 11019 31135 11061 31144
rect 10923 31100 10965 31109
rect 10923 31060 10924 31100
rect 10964 31060 10965 31100
rect 10923 31051 10965 31060
rect 11115 30764 11157 30773
rect 11115 30724 11116 30764
rect 11156 30724 11157 30764
rect 11115 30715 11157 30724
rect 11116 29681 11156 30715
rect 11212 30680 11252 30691
rect 11212 30605 11252 30640
rect 11211 30596 11253 30605
rect 11211 30556 11212 30596
rect 11252 30556 11253 30596
rect 11211 30547 11253 30556
rect 11212 30269 11252 30547
rect 11211 30260 11253 30269
rect 11211 30220 11212 30260
rect 11252 30220 11253 30260
rect 11211 30211 11253 30220
rect 11115 29672 11157 29681
rect 11115 29632 11116 29672
rect 11156 29632 11157 29672
rect 11115 29623 11157 29632
rect 11308 29000 11348 31303
rect 11404 30689 11444 32395
rect 11499 32192 11541 32201
rect 11499 32152 11500 32192
rect 11540 32152 11541 32192
rect 11499 32143 11541 32152
rect 11500 32024 11540 32143
rect 11500 31975 11540 31984
rect 11596 31940 11636 32404
rect 11692 32192 11732 32203
rect 11692 32117 11732 32152
rect 11691 32108 11733 32117
rect 11691 32068 11692 32108
rect 11732 32068 11733 32108
rect 11691 32059 11733 32068
rect 11692 31940 11732 31949
rect 11596 31900 11692 31940
rect 11692 31891 11732 31900
rect 11788 31772 11828 32992
rect 12364 32983 12404 32992
rect 12556 32875 12596 36007
rect 12843 35888 12885 35897
rect 12843 35848 12844 35888
rect 12884 35848 12885 35888
rect 12843 35839 12885 35848
rect 12844 35216 12884 35839
rect 12844 35167 12884 35176
rect 12652 34292 12692 34301
rect 12940 34292 12980 36856
rect 13132 36728 13172 36737
rect 13132 36401 13172 36688
rect 13131 36392 13173 36401
rect 13131 36352 13132 36392
rect 13172 36352 13173 36392
rect 13131 36343 13173 36352
rect 13035 35636 13077 35645
rect 13035 35596 13036 35636
rect 13076 35596 13077 35636
rect 13035 35587 13077 35596
rect 13036 34544 13076 35587
rect 13228 35384 13268 40720
rect 13324 40508 13364 40517
rect 13364 40468 13460 40508
rect 13324 40459 13364 40468
rect 13324 39752 13364 39761
rect 13324 37241 13364 39712
rect 13323 37232 13365 37241
rect 13323 37192 13324 37232
rect 13364 37192 13365 37232
rect 13323 37183 13365 37192
rect 13420 35645 13460 40468
rect 13612 40349 13652 41224
rect 13900 41224 13996 41264
rect 13803 41012 13845 41021
rect 13803 40972 13804 41012
rect 13844 40972 13845 41012
rect 13803 40963 13845 40972
rect 13804 40878 13844 40963
rect 13708 40424 13748 40433
rect 13611 40340 13653 40349
rect 13611 40300 13612 40340
rect 13652 40300 13653 40340
rect 13611 40291 13653 40300
rect 13516 40256 13556 40265
rect 13516 39593 13556 40216
rect 13515 39584 13557 39593
rect 13515 39544 13516 39584
rect 13556 39544 13557 39584
rect 13515 39535 13557 39544
rect 13708 39089 13748 40384
rect 13900 40097 13940 41224
rect 13996 41215 14036 41224
rect 14092 40517 14132 42928
rect 14091 40508 14133 40517
rect 14091 40468 14092 40508
rect 14132 40468 14133 40508
rect 14091 40459 14133 40468
rect 14284 40433 14324 42928
rect 14476 41693 14516 42928
rect 14667 42904 14668 42928
rect 14708 42928 14728 42944
rect 14840 42928 14920 43008
rect 15032 42928 15112 43008
rect 15224 42928 15304 43008
rect 15416 42928 15496 43008
rect 15608 42928 15688 43008
rect 15800 42928 15880 43008
rect 15992 42928 16072 43008
rect 16184 42928 16264 43008
rect 16376 42928 16456 43008
rect 16568 42928 16648 43008
rect 16760 42928 16840 43008
rect 16952 42928 17032 43008
rect 17144 42928 17224 43008
rect 17336 42928 17416 43008
rect 17528 42928 17608 43008
rect 17720 42928 17800 43008
rect 17912 42928 17992 43008
rect 18104 42928 18184 43008
rect 18296 42928 18376 43008
rect 18488 42928 18568 43008
rect 18680 42928 18760 43008
rect 18872 42928 18952 43008
rect 19064 42928 19144 43008
rect 19256 42944 19336 43008
rect 19256 42928 19276 42944
rect 14708 42904 14709 42928
rect 14667 42895 14709 42904
rect 14475 41684 14517 41693
rect 14475 41644 14476 41684
rect 14516 41644 14517 41684
rect 14475 41635 14517 41644
rect 14475 41180 14517 41189
rect 14475 41140 14476 41180
rect 14516 41140 14517 41180
rect 14475 41131 14517 41140
rect 14283 40424 14325 40433
rect 14283 40384 14284 40424
rect 14324 40384 14325 40424
rect 14283 40375 14325 40384
rect 13995 40340 14037 40349
rect 13995 40300 13996 40340
rect 14036 40300 14037 40340
rect 13995 40291 14037 40300
rect 13899 40088 13941 40097
rect 13899 40048 13900 40088
rect 13940 40048 13941 40088
rect 13899 40039 13941 40048
rect 13897 39089 13937 39146
rect 13707 39080 13749 39089
rect 13707 39040 13708 39080
rect 13748 39040 13749 39080
rect 13707 39031 13749 39040
rect 13896 39080 13938 39089
rect 13896 39040 13897 39080
rect 13937 39054 13940 39080
rect 13896 39031 13900 39040
rect 13900 39005 13940 39014
rect 13515 38996 13557 39005
rect 13515 38956 13516 38996
rect 13556 38956 13557 38996
rect 13515 38947 13557 38956
rect 13516 38501 13556 38947
rect 13612 38912 13652 38921
rect 13900 38904 13940 38913
rect 13612 38669 13652 38872
rect 13804 38864 13900 38904
rect 13611 38660 13653 38669
rect 13611 38620 13612 38660
rect 13652 38620 13653 38660
rect 13611 38611 13653 38620
rect 13515 38492 13557 38501
rect 13515 38452 13516 38492
rect 13556 38452 13557 38492
rect 13515 38443 13557 38452
rect 13516 37997 13556 38443
rect 13515 37988 13557 37997
rect 13515 37948 13516 37988
rect 13556 37948 13557 37988
rect 13515 37939 13557 37948
rect 13707 37652 13749 37661
rect 13707 37612 13708 37652
rect 13748 37612 13749 37652
rect 13707 37603 13749 37612
rect 13708 37518 13748 37603
rect 13515 37484 13557 37493
rect 13515 37444 13516 37484
rect 13556 37444 13557 37484
rect 13515 37435 13557 37444
rect 13516 37400 13556 37435
rect 13516 37349 13556 37360
rect 13707 37400 13749 37409
rect 13707 37360 13708 37400
rect 13748 37360 13749 37400
rect 13707 37351 13749 37360
rect 13708 37266 13748 37351
rect 13804 37157 13844 38864
rect 13900 38855 13940 38864
rect 13996 38744 14036 40291
rect 14187 40004 14229 40013
rect 14187 39964 14188 40004
rect 14228 39964 14229 40004
rect 14187 39955 14229 39964
rect 13900 38704 14036 38744
rect 14092 38744 14132 38753
rect 13900 37661 13940 38704
rect 14092 38501 14132 38704
rect 14091 38492 14133 38501
rect 14091 38452 14092 38492
rect 14132 38452 14133 38492
rect 14091 38443 14133 38452
rect 14188 38240 14228 39955
rect 14476 39509 14516 41131
rect 14860 40853 14900 42928
rect 15052 41945 15092 42928
rect 15051 41936 15093 41945
rect 15051 41896 15052 41936
rect 15092 41896 15093 41936
rect 15051 41887 15093 41896
rect 15244 41525 15284 42928
rect 15243 41516 15285 41525
rect 15243 41476 15244 41516
rect 15284 41476 15285 41516
rect 15243 41467 15285 41476
rect 15244 41264 15284 41273
rect 14859 40844 14901 40853
rect 14859 40804 14860 40844
rect 14900 40804 14901 40844
rect 14859 40795 14901 40804
rect 14859 40424 14901 40433
rect 14859 40384 14860 40424
rect 14900 40384 14901 40424
rect 14859 40375 14901 40384
rect 14956 40424 14996 40433
rect 14667 40340 14709 40349
rect 14667 40300 14668 40340
rect 14708 40300 14709 40340
rect 14667 40291 14709 40300
rect 14571 40004 14613 40013
rect 14571 39964 14572 40004
rect 14612 39964 14613 40004
rect 14571 39955 14613 39964
rect 14572 39752 14612 39955
rect 14572 39703 14612 39712
rect 14475 39500 14517 39509
rect 14475 39460 14476 39500
rect 14516 39460 14517 39500
rect 14475 39451 14517 39460
rect 14571 39416 14613 39425
rect 14571 39376 14572 39416
rect 14612 39376 14613 39416
rect 14571 39367 14613 39376
rect 14283 39332 14325 39341
rect 14283 39292 14284 39332
rect 14324 39292 14325 39332
rect 14283 39283 14325 39292
rect 14284 39173 14324 39283
rect 14283 39164 14325 39173
rect 14283 39124 14284 39164
rect 14324 39124 14325 39164
rect 14283 39115 14325 39124
rect 14284 38912 14324 39115
rect 14284 38863 14324 38872
rect 14380 38912 14420 38923
rect 14380 38837 14420 38872
rect 14476 38912 14516 38921
rect 14379 38828 14421 38837
rect 14379 38788 14380 38828
rect 14420 38788 14421 38828
rect 14379 38779 14421 38788
rect 14476 38501 14516 38872
rect 14572 38912 14612 39367
rect 14668 38921 14708 40291
rect 14764 39500 14804 39509
rect 14764 39425 14804 39460
rect 14764 39416 14806 39425
rect 14764 39376 14765 39416
rect 14805 39376 14806 39416
rect 14764 39367 14806 39376
rect 14763 39164 14805 39173
rect 14763 39124 14764 39164
rect 14804 39124 14805 39164
rect 14763 39115 14805 39124
rect 14572 38863 14612 38872
rect 14667 38912 14709 38921
rect 14667 38872 14668 38912
rect 14708 38872 14709 38912
rect 14667 38863 14709 38872
rect 14764 38912 14804 39115
rect 14860 39080 14900 40375
rect 14956 40013 14996 40384
rect 15147 40256 15189 40265
rect 15147 40216 15148 40256
rect 15188 40216 15189 40256
rect 15147 40207 15189 40216
rect 15148 40122 15188 40207
rect 14955 40004 14997 40013
rect 14955 39964 14956 40004
rect 14996 39964 14997 40004
rect 14955 39955 14997 39964
rect 15244 39920 15284 41224
rect 15436 41189 15476 42928
rect 15628 41609 15668 42928
rect 15627 41600 15669 41609
rect 15627 41560 15628 41600
rect 15668 41560 15669 41600
rect 15627 41551 15669 41560
rect 15531 41432 15573 41441
rect 15531 41392 15532 41432
rect 15572 41392 15573 41432
rect 15531 41383 15573 41392
rect 15435 41180 15477 41189
rect 15435 41140 15436 41180
rect 15476 41140 15477 41180
rect 15435 41131 15477 41140
rect 15435 41012 15477 41021
rect 15435 40972 15436 41012
rect 15476 40972 15477 41012
rect 15435 40963 15477 40972
rect 15436 40878 15476 40963
rect 15532 40844 15572 41383
rect 15628 41264 15668 41273
rect 15628 41105 15668 41224
rect 15627 41096 15669 41105
rect 15627 41056 15628 41096
rect 15668 41056 15669 41096
rect 15627 41047 15669 41056
rect 15532 40804 15668 40844
rect 15148 39880 15284 39920
rect 15340 40424 15380 40433
rect 15051 39836 15093 39845
rect 15051 39796 15052 39836
rect 15092 39796 15093 39836
rect 15051 39787 15093 39796
rect 14955 39752 14997 39761
rect 14955 39712 14956 39752
rect 14996 39712 14997 39752
rect 14955 39703 14997 39712
rect 15052 39752 15092 39787
rect 14956 39618 14996 39703
rect 14860 39040 14996 39080
rect 14764 38660 14804 38872
rect 14859 38912 14901 38921
rect 14859 38872 14860 38912
rect 14900 38872 14901 38912
rect 14859 38863 14901 38872
rect 14860 38778 14900 38863
rect 14956 38828 14996 39040
rect 15052 38912 15092 39712
rect 15052 38863 15092 38872
rect 14956 38779 14996 38788
rect 15051 38744 15093 38753
rect 15051 38704 15052 38744
rect 15092 38704 15093 38744
rect 15051 38695 15093 38704
rect 14764 38620 14996 38660
rect 14475 38492 14517 38501
rect 14475 38452 14476 38492
rect 14516 38452 14517 38492
rect 14475 38443 14517 38452
rect 14859 38492 14901 38501
rect 14859 38452 14860 38492
rect 14900 38452 14901 38492
rect 14859 38443 14901 38452
rect 14667 38408 14709 38417
rect 14667 38368 14668 38408
rect 14708 38368 14709 38408
rect 14667 38359 14709 38368
rect 14860 38408 14900 38443
rect 14380 38324 14420 38333
rect 14092 38200 14188 38240
rect 13899 37652 13941 37661
rect 13899 37612 13900 37652
rect 13940 37612 13941 37652
rect 13899 37603 13941 37612
rect 14092 37568 14132 38200
rect 14188 38191 14228 38200
rect 14283 38240 14325 38249
rect 14283 38200 14284 38240
rect 14324 38200 14325 38240
rect 14380 38240 14420 38284
rect 14571 38240 14613 38249
rect 14380 38200 14572 38240
rect 14612 38200 14613 38240
rect 14283 38191 14325 38200
rect 14571 38191 14613 38200
rect 14668 38240 14708 38359
rect 14860 38357 14900 38368
rect 14668 38191 14708 38200
rect 14764 38240 14804 38249
rect 14187 38072 14229 38081
rect 14187 38032 14188 38072
rect 14228 38032 14229 38072
rect 14187 38023 14229 38032
rect 13996 37528 14132 37568
rect 13900 37400 13940 37409
rect 13803 37148 13845 37157
rect 13803 37108 13804 37148
rect 13844 37108 13845 37148
rect 13803 37099 13845 37108
rect 13804 36812 13844 36821
rect 13516 36772 13804 36812
rect 13419 35636 13461 35645
rect 13419 35596 13420 35636
rect 13460 35596 13461 35636
rect 13419 35587 13461 35596
rect 13516 35393 13556 36772
rect 13804 36763 13844 36772
rect 13660 36686 13700 36695
rect 13660 36644 13700 36646
rect 13660 36604 13844 36644
rect 13707 36140 13749 36149
rect 13707 36100 13708 36140
rect 13748 36100 13749 36140
rect 13707 36091 13749 36100
rect 13804 36140 13844 36604
rect 13900 36233 13940 37360
rect 13899 36224 13941 36233
rect 13899 36184 13900 36224
rect 13940 36184 13941 36224
rect 13899 36175 13941 36184
rect 13804 36091 13844 36100
rect 13611 36056 13653 36065
rect 13611 36016 13612 36056
rect 13652 36016 13653 36056
rect 13611 36007 13653 36016
rect 13612 35888 13652 36007
rect 13612 35839 13652 35848
rect 13611 35636 13653 35645
rect 13611 35596 13612 35636
rect 13652 35596 13653 35636
rect 13611 35587 13653 35596
rect 13515 35384 13557 35393
rect 13228 35344 13460 35384
rect 13132 35216 13172 35227
rect 13132 35141 13172 35176
rect 13227 35216 13269 35225
rect 13227 35176 13228 35216
rect 13268 35176 13269 35216
rect 13227 35167 13269 35176
rect 13131 35132 13173 35141
rect 13131 35092 13132 35132
rect 13172 35092 13173 35132
rect 13131 35083 13173 35092
rect 13036 34504 13172 34544
rect 13036 34376 13076 34387
rect 13036 34301 13076 34336
rect 12692 34252 12980 34292
rect 13035 34292 13077 34301
rect 13035 34252 13036 34292
rect 13076 34252 13077 34292
rect 12652 34243 12692 34252
rect 13035 34243 13077 34252
rect 12651 33284 12693 33293
rect 12651 33244 12652 33284
rect 12692 33244 12693 33284
rect 12651 33235 12693 33244
rect 11980 32864 12020 32873
rect 11884 32638 11924 32647
rect 11884 32453 11924 32598
rect 11883 32444 11925 32453
rect 11883 32404 11884 32444
rect 11924 32404 11925 32444
rect 11883 32395 11925 32404
rect 11980 32285 12020 32824
rect 12075 32864 12117 32873
rect 12075 32824 12076 32864
rect 12116 32824 12117 32864
rect 12075 32815 12117 32824
rect 12267 32864 12309 32873
rect 12267 32824 12268 32864
rect 12308 32824 12309 32864
rect 12267 32815 12309 32824
rect 12460 32835 12596 32875
rect 12076 32730 12116 32815
rect 12171 32780 12213 32789
rect 12171 32740 12172 32780
rect 12212 32740 12213 32780
rect 12171 32731 12213 32740
rect 12172 32360 12212 32731
rect 12076 32320 12212 32360
rect 12268 32360 12308 32815
rect 12363 32696 12405 32705
rect 12363 32656 12364 32696
rect 12404 32656 12405 32696
rect 12363 32647 12405 32656
rect 11979 32276 12021 32285
rect 11979 32236 11980 32276
rect 12020 32236 12021 32276
rect 11979 32227 12021 32236
rect 11596 31732 11828 31772
rect 11884 32192 11924 32201
rect 11499 31268 11541 31277
rect 11499 31228 11500 31268
rect 11540 31228 11541 31268
rect 11499 31219 11541 31228
rect 11500 30773 11540 31219
rect 11499 30764 11541 30773
rect 11499 30724 11500 30764
rect 11540 30724 11541 30764
rect 11499 30715 11541 30724
rect 11403 30680 11445 30689
rect 11403 30640 11404 30680
rect 11444 30640 11445 30680
rect 11403 30631 11445 30640
rect 11596 30680 11636 31732
rect 11691 31520 11733 31529
rect 11691 31480 11692 31520
rect 11732 31480 11733 31520
rect 11691 31471 11733 31480
rect 11596 30631 11636 30640
rect 11692 30596 11732 31471
rect 11884 31109 11924 32152
rect 11980 32192 12020 32227
rect 11980 32141 12020 32152
rect 11883 31100 11925 31109
rect 11883 31060 11884 31100
rect 11924 31060 11925 31100
rect 11883 31051 11925 31060
rect 12076 30932 12116 32320
rect 12268 32311 12308 32320
rect 12172 32192 12212 32203
rect 12172 32117 12212 32152
rect 12364 32192 12404 32647
rect 12460 32360 12500 32835
rect 12556 32705 12596 32790
rect 12555 32696 12597 32705
rect 12555 32656 12556 32696
rect 12596 32656 12597 32696
rect 12555 32647 12597 32656
rect 12652 32360 12692 33235
rect 12843 33032 12885 33041
rect 13132 33032 13172 34504
rect 13228 34133 13268 35167
rect 13323 35132 13365 35141
rect 13323 35092 13324 35132
rect 13364 35092 13365 35132
rect 13323 35083 13365 35092
rect 13227 34124 13269 34133
rect 13227 34084 13228 34124
rect 13268 34084 13269 34124
rect 13227 34075 13269 34084
rect 13324 33293 13364 35083
rect 13420 34040 13460 35344
rect 13515 35344 13516 35384
rect 13556 35344 13557 35384
rect 13515 35335 13557 35344
rect 13515 34964 13557 34973
rect 13515 34924 13516 34964
rect 13556 34924 13557 34964
rect 13515 34915 13557 34924
rect 13516 34830 13556 34915
rect 13612 34637 13652 35587
rect 13708 35393 13748 36091
rect 13996 36056 14036 37528
rect 14091 37400 14133 37409
rect 14091 37360 14092 37400
rect 14132 37360 14133 37400
rect 14091 37351 14133 37360
rect 14188 37400 14228 38023
rect 14284 37409 14324 38191
rect 14572 38106 14612 38191
rect 14667 38072 14709 38081
rect 14667 38032 14668 38072
rect 14708 38032 14709 38072
rect 14667 38023 14709 38032
rect 14571 37988 14613 37997
rect 14571 37948 14572 37988
rect 14612 37948 14613 37988
rect 14571 37939 14613 37948
rect 14379 37652 14421 37661
rect 14379 37612 14380 37652
rect 14420 37612 14421 37652
rect 14379 37603 14421 37612
rect 14380 37518 14420 37603
rect 14188 37351 14228 37360
rect 14283 37400 14325 37409
rect 14283 37360 14284 37400
rect 14324 37360 14325 37400
rect 14283 37351 14325 37360
rect 14380 37400 14420 37409
rect 14092 37266 14132 37351
rect 14380 37241 14420 37360
rect 14572 37400 14612 37939
rect 14668 37652 14708 38023
rect 14668 37603 14708 37612
rect 14764 37493 14804 38200
rect 14956 38081 14996 38620
rect 15052 38249 15092 38695
rect 15148 38417 15188 39880
rect 15243 39752 15285 39761
rect 15243 39712 15244 39752
rect 15284 39712 15285 39752
rect 15243 39703 15285 39712
rect 15244 39618 15284 39703
rect 15243 39500 15285 39509
rect 15243 39460 15244 39500
rect 15284 39460 15285 39500
rect 15243 39451 15285 39460
rect 15244 39366 15284 39451
rect 15340 39341 15380 40384
rect 15436 40424 15476 40435
rect 15532 40433 15572 40518
rect 15436 40349 15476 40384
rect 15531 40424 15573 40433
rect 15531 40384 15532 40424
rect 15572 40384 15573 40424
rect 15531 40375 15573 40384
rect 15628 40424 15668 40804
rect 15820 40433 15860 42928
rect 16012 41105 16052 42928
rect 16204 42533 16244 42928
rect 16203 42524 16245 42533
rect 16203 42484 16204 42524
rect 16244 42484 16245 42524
rect 16203 42475 16245 42484
rect 16396 42365 16436 42928
rect 16395 42356 16437 42365
rect 16395 42316 16396 42356
rect 16436 42316 16437 42356
rect 16395 42307 16437 42316
rect 16491 41348 16533 41357
rect 16491 41308 16492 41348
rect 16532 41308 16533 41348
rect 16491 41299 16533 41308
rect 16299 41264 16341 41273
rect 16299 41224 16300 41264
rect 16340 41224 16341 41264
rect 16299 41215 16341 41224
rect 16011 41096 16053 41105
rect 16011 41056 16012 41096
rect 16052 41056 16053 41096
rect 16011 41047 16053 41056
rect 16107 41012 16149 41021
rect 16107 40972 16108 41012
rect 16148 40972 16149 41012
rect 16107 40963 16149 40972
rect 15628 40375 15668 40384
rect 15819 40424 15861 40433
rect 15819 40384 15820 40424
rect 15860 40384 15861 40424
rect 15819 40375 15861 40384
rect 15916 40424 15956 40433
rect 15435 40340 15477 40349
rect 15435 40300 15436 40340
rect 15476 40300 15477 40340
rect 15435 40291 15477 40300
rect 15531 40256 15573 40265
rect 15820 40256 15860 40265
rect 15531 40216 15532 40256
rect 15572 40216 15573 40256
rect 15531 40207 15573 40216
rect 15724 40216 15820 40256
rect 15435 40004 15477 40013
rect 15435 39964 15436 40004
rect 15476 39964 15477 40004
rect 15435 39955 15477 39964
rect 15339 39332 15381 39341
rect 15339 39292 15340 39332
rect 15380 39292 15381 39332
rect 15339 39283 15381 39292
rect 15340 39089 15380 39174
rect 15339 39080 15381 39089
rect 15339 39040 15340 39080
rect 15380 39040 15381 39080
rect 15339 39031 15381 39040
rect 15340 38912 15380 38921
rect 15244 38872 15340 38912
rect 15147 38408 15189 38417
rect 15147 38368 15148 38408
rect 15188 38368 15189 38408
rect 15147 38359 15189 38368
rect 15051 38240 15093 38249
rect 15148 38240 15188 38249
rect 15051 38200 15052 38240
rect 15092 38200 15148 38240
rect 15051 38191 15093 38200
rect 15148 38191 15188 38200
rect 15052 38106 15092 38191
rect 14955 38072 14997 38081
rect 14955 38032 14956 38072
rect 14996 38032 14997 38072
rect 14955 38023 14997 38032
rect 15244 37745 15284 38872
rect 15340 38863 15380 38872
rect 15436 38744 15476 39955
rect 15532 39752 15572 40207
rect 15532 39703 15572 39712
rect 15628 39752 15668 39761
rect 15724 39752 15764 40216
rect 15820 40207 15860 40216
rect 15916 40013 15956 40384
rect 16012 40424 16052 40435
rect 16012 40349 16052 40384
rect 16108 40403 16148 40963
rect 16300 40685 16340 41215
rect 16299 40676 16341 40685
rect 16299 40636 16300 40676
rect 16340 40636 16341 40676
rect 16299 40627 16341 40636
rect 16300 40508 16340 40627
rect 16492 40592 16532 41299
rect 16588 41021 16628 42928
rect 16587 41012 16629 41021
rect 16587 40972 16588 41012
rect 16628 40972 16629 41012
rect 16587 40963 16629 40972
rect 16780 40592 16820 42928
rect 16875 41432 16917 41441
rect 16875 41392 16876 41432
rect 16916 41392 16917 41432
rect 16875 41383 16917 41392
rect 16876 41264 16916 41383
rect 16876 41215 16916 41224
rect 16972 40769 17012 42928
rect 17164 41525 17204 42928
rect 17356 42701 17396 42928
rect 17548 42869 17588 42928
rect 17547 42860 17589 42869
rect 17547 42820 17548 42860
rect 17588 42820 17589 42860
rect 17547 42811 17589 42820
rect 17355 42692 17397 42701
rect 17355 42652 17356 42692
rect 17396 42652 17397 42692
rect 17355 42643 17397 42652
rect 17643 42188 17685 42197
rect 17643 42148 17644 42188
rect 17684 42148 17685 42188
rect 17643 42139 17685 42148
rect 17163 41516 17205 41525
rect 17163 41476 17164 41516
rect 17204 41476 17205 41516
rect 17163 41467 17205 41476
rect 17068 41273 17108 41358
rect 17259 41348 17301 41357
rect 17259 41308 17260 41348
rect 17300 41308 17301 41348
rect 17259 41299 17301 41308
rect 17067 41264 17109 41273
rect 17067 41224 17068 41264
rect 17108 41224 17109 41264
rect 17067 41215 17109 41224
rect 17260 41264 17300 41299
rect 17260 41213 17300 41224
rect 17356 41264 17396 41273
rect 17067 41012 17109 41021
rect 17067 40972 17068 41012
rect 17108 40972 17109 41012
rect 17067 40963 17109 40972
rect 17068 40878 17108 40963
rect 16971 40760 17013 40769
rect 16971 40720 16972 40760
rect 17012 40720 17013 40760
rect 16971 40711 17013 40720
rect 17356 40601 17396 41224
rect 17644 41180 17684 42139
rect 17740 41441 17780 42928
rect 17835 42776 17877 42785
rect 17835 42736 17836 42776
rect 17876 42736 17877 42776
rect 17835 42727 17877 42736
rect 17739 41432 17781 41441
rect 17739 41392 17740 41432
rect 17780 41392 17781 41432
rect 17739 41383 17781 41392
rect 17740 41180 17780 41189
rect 17644 41140 17740 41180
rect 17740 41131 17780 41140
rect 17836 41096 17876 42727
rect 17932 41525 17972 42928
rect 18124 42617 18164 42928
rect 18123 42608 18165 42617
rect 18123 42568 18124 42608
rect 18164 42568 18165 42608
rect 18123 42559 18165 42568
rect 18027 41684 18069 41693
rect 18027 41644 18028 41684
rect 18068 41644 18069 41684
rect 18027 41635 18069 41644
rect 17931 41516 17973 41525
rect 17931 41476 17932 41516
rect 17972 41476 17973 41516
rect 17931 41467 17973 41476
rect 17932 41096 17972 41105
rect 17836 41056 17932 41096
rect 17932 41047 17972 41056
rect 17547 41012 17589 41021
rect 17547 40972 17548 41012
rect 17588 40972 17589 41012
rect 17547 40963 17589 40972
rect 17548 40878 17588 40963
rect 17355 40592 17397 40601
rect 16492 40552 16628 40592
rect 16780 40552 17204 40592
rect 16300 40468 16435 40508
rect 16395 40464 16435 40468
rect 16395 40424 16436 40464
rect 16396 40375 16436 40384
rect 16492 40424 16532 40433
rect 16108 40354 16148 40363
rect 16011 40340 16053 40349
rect 16011 40300 16012 40340
rect 16052 40300 16053 40340
rect 16011 40291 16053 40300
rect 16300 40256 16340 40265
rect 16300 40088 16340 40216
rect 16204 40048 16340 40088
rect 15915 40004 15957 40013
rect 15915 39964 15916 40004
rect 15956 39964 15957 40004
rect 15915 39955 15957 39964
rect 16204 39761 16244 40048
rect 16299 39920 16341 39929
rect 16299 39880 16300 39920
rect 16340 39880 16341 39920
rect 16299 39871 16341 39880
rect 15668 39712 15764 39752
rect 15820 39752 15860 39761
rect 16203 39752 16245 39761
rect 15860 39712 15956 39752
rect 15628 39703 15668 39712
rect 15820 39703 15860 39712
rect 15819 39500 15861 39509
rect 15819 39460 15820 39500
rect 15860 39460 15861 39500
rect 15819 39451 15861 39460
rect 15627 39416 15669 39425
rect 15627 39376 15628 39416
rect 15668 39376 15669 39416
rect 15627 39367 15669 39376
rect 15531 39080 15573 39089
rect 15531 39040 15532 39080
rect 15572 39040 15573 39080
rect 15531 39031 15573 39040
rect 15532 38946 15572 39031
rect 15340 38704 15476 38744
rect 15243 37736 15285 37745
rect 15243 37696 15244 37736
rect 15284 37696 15285 37736
rect 15243 37687 15285 37696
rect 15340 37661 15380 38704
rect 15435 38240 15477 38249
rect 15435 38200 15436 38240
rect 15476 38200 15477 38240
rect 15435 38191 15477 38200
rect 15532 38240 15572 38249
rect 15436 38106 15476 38191
rect 15532 37997 15572 38200
rect 15628 38165 15668 39367
rect 15820 39366 15860 39451
rect 15916 39248 15956 39712
rect 16203 39712 16204 39752
rect 16244 39712 16245 39752
rect 16203 39703 16245 39712
rect 16300 39752 16340 39871
rect 16300 39703 16340 39712
rect 16011 39668 16053 39677
rect 16011 39628 16012 39668
rect 16052 39628 16053 39668
rect 16011 39619 16053 39628
rect 16012 39534 16052 39619
rect 16492 39509 16532 40384
rect 16588 40424 16628 40552
rect 16588 39845 16628 40384
rect 16683 40424 16725 40433
rect 16683 40384 16684 40424
rect 16724 40384 16725 40424
rect 16683 40375 16725 40384
rect 16876 40424 16916 40433
rect 16587 39836 16629 39845
rect 16587 39796 16588 39836
rect 16628 39796 16629 39836
rect 16587 39787 16629 39796
rect 16491 39500 16533 39509
rect 16491 39460 16492 39500
rect 16532 39460 16533 39500
rect 16491 39451 16533 39460
rect 15916 39208 16340 39248
rect 15724 39124 16052 39164
rect 15724 39080 15764 39124
rect 16012 39080 16052 39124
rect 16012 39040 16244 39080
rect 15724 39031 15764 39040
rect 15724 38912 15764 38921
rect 15724 38501 15764 38872
rect 15915 38912 15957 38921
rect 15915 38872 15916 38912
rect 15956 38872 15957 38912
rect 15915 38863 15957 38872
rect 16012 38912 16052 38921
rect 16204 38912 16244 39040
rect 16300 38996 16340 39208
rect 16300 38947 16340 38956
rect 16052 38872 16148 38912
rect 16012 38863 16052 38872
rect 15916 38778 15956 38863
rect 15723 38492 15765 38501
rect 15723 38452 15724 38492
rect 15764 38452 15765 38492
rect 15723 38443 15765 38452
rect 16108 38324 16148 38872
rect 16204 38863 16244 38872
rect 16396 38912 16436 38921
rect 16588 38912 16628 38921
rect 16436 38872 16532 38912
rect 16396 38863 16436 38872
rect 16395 38660 16437 38669
rect 16395 38620 16396 38660
rect 16436 38620 16437 38660
rect 16395 38611 16437 38620
rect 16108 38284 16340 38324
rect 15627 38156 15669 38165
rect 15627 38116 15628 38156
rect 15668 38116 15669 38156
rect 15627 38107 15669 38116
rect 16012 38156 16052 38165
rect 16203 38156 16245 38165
rect 16052 38116 16148 38156
rect 16012 38107 16052 38116
rect 15819 38072 15861 38081
rect 15819 38032 15820 38072
rect 15860 38032 15861 38072
rect 15819 38023 15861 38032
rect 15531 37988 15573 37997
rect 15531 37948 15532 37988
rect 15572 37948 15573 37988
rect 15531 37939 15573 37948
rect 15820 37938 15860 38023
rect 16011 37988 16053 37997
rect 16011 37948 16012 37988
rect 16052 37948 16053 37988
rect 16011 37939 16053 37948
rect 15339 37652 15381 37661
rect 15339 37612 15340 37652
rect 15380 37612 15381 37652
rect 15339 37603 15381 37612
rect 15531 37652 15573 37661
rect 15531 37612 15532 37652
rect 15572 37612 15573 37652
rect 15531 37603 15573 37612
rect 14763 37484 14805 37493
rect 14763 37444 14764 37484
rect 14804 37444 14805 37484
rect 14763 37435 14805 37444
rect 14572 37351 14612 37360
rect 14667 37400 14709 37409
rect 14667 37360 14668 37400
rect 14708 37360 14709 37400
rect 14667 37351 14709 37360
rect 14187 37232 14229 37241
rect 14187 37192 14188 37232
rect 14228 37192 14229 37232
rect 14187 37183 14229 37192
rect 14379 37232 14421 37241
rect 14379 37192 14380 37232
rect 14420 37192 14421 37232
rect 14379 37183 14421 37192
rect 14091 37064 14133 37073
rect 14091 37024 14092 37064
rect 14132 37024 14133 37064
rect 14091 37015 14133 37024
rect 14092 36728 14132 37015
rect 14092 36679 14132 36688
rect 13900 36016 14036 36056
rect 13707 35384 13749 35393
rect 13707 35344 13708 35384
rect 13748 35344 13749 35384
rect 13707 35335 13749 35344
rect 13708 35216 13748 35225
rect 13611 34628 13653 34637
rect 13611 34588 13612 34628
rect 13652 34588 13653 34628
rect 13611 34579 13653 34588
rect 13708 34553 13748 35176
rect 13707 34544 13749 34553
rect 13707 34504 13708 34544
rect 13748 34504 13749 34544
rect 13707 34495 13749 34504
rect 13708 34301 13748 34495
rect 13707 34292 13749 34301
rect 13707 34252 13708 34292
rect 13748 34252 13749 34292
rect 13707 34243 13749 34252
rect 13420 34000 13556 34040
rect 13419 33872 13461 33881
rect 13419 33832 13420 33872
rect 13460 33832 13461 33872
rect 13419 33823 13461 33832
rect 13323 33284 13365 33293
rect 13323 33244 13324 33284
rect 13364 33244 13365 33284
rect 13323 33235 13365 33244
rect 12843 32992 12844 33032
rect 12884 32992 12885 33032
rect 12843 32983 12885 32992
rect 12940 32992 13172 33032
rect 12748 32864 12788 32873
rect 12748 32537 12788 32824
rect 12844 32864 12884 32983
rect 12844 32815 12884 32824
rect 12747 32528 12789 32537
rect 12747 32488 12748 32528
rect 12788 32488 12789 32528
rect 12747 32479 12789 32488
rect 12940 32453 12980 32992
rect 13035 32864 13077 32873
rect 13324 32864 13364 32873
rect 13035 32824 13036 32864
rect 13076 32824 13077 32864
rect 13035 32815 13077 32824
rect 13228 32824 13324 32864
rect 13036 32730 13076 32815
rect 13131 32780 13173 32789
rect 13131 32740 13132 32780
rect 13172 32740 13173 32780
rect 13131 32731 13173 32740
rect 13132 32646 13172 32731
rect 13035 32528 13077 32537
rect 13035 32488 13036 32528
rect 13076 32488 13077 32528
rect 13035 32479 13077 32488
rect 12939 32444 12981 32453
rect 12939 32404 12940 32444
rect 12980 32404 12981 32444
rect 12939 32395 12981 32404
rect 12460 32320 12596 32360
rect 12652 32320 12884 32360
rect 12364 32143 12404 32152
rect 12460 32192 12500 32201
rect 12171 32108 12213 32117
rect 12171 32068 12172 32108
rect 12212 32068 12213 32108
rect 12171 32059 12213 32068
rect 12460 31781 12500 32152
rect 12459 31772 12501 31781
rect 12459 31732 12460 31772
rect 12500 31732 12501 31772
rect 12459 31723 12501 31732
rect 12556 31445 12596 32320
rect 12651 32192 12693 32201
rect 12651 32152 12652 32192
rect 12692 32152 12693 32192
rect 12651 32143 12693 32152
rect 12748 32192 12788 32203
rect 12652 32058 12692 32143
rect 12748 32117 12788 32152
rect 12747 32108 12789 32117
rect 12747 32068 12748 32108
rect 12788 32068 12789 32108
rect 12747 32059 12789 32068
rect 12171 31436 12213 31445
rect 12171 31396 12172 31436
rect 12212 31396 12213 31436
rect 12171 31387 12213 31396
rect 12555 31436 12597 31445
rect 12555 31396 12556 31436
rect 12596 31396 12597 31436
rect 12555 31387 12597 31396
rect 12172 31352 12212 31387
rect 12172 31301 12212 31312
rect 12652 31352 12692 31361
rect 12364 31268 12404 31277
rect 12652 31268 12692 31312
rect 12747 31352 12789 31361
rect 12747 31312 12748 31352
rect 12788 31312 12789 31352
rect 12747 31303 12789 31312
rect 12404 31228 12692 31268
rect 12364 31219 12404 31228
rect 12748 31218 12788 31303
rect 12267 31100 12309 31109
rect 12267 31060 12268 31100
rect 12308 31060 12309 31100
rect 12267 31051 12309 31060
rect 11980 30892 12116 30932
rect 12171 30932 12213 30941
rect 12171 30892 12172 30932
rect 12212 30892 12213 30932
rect 11884 30605 11924 30690
rect 11980 30680 12020 30892
rect 12171 30883 12213 30892
rect 11980 30631 12020 30640
rect 11692 30547 11732 30556
rect 11883 30596 11925 30605
rect 11883 30556 11884 30596
rect 11924 30556 11925 30596
rect 11883 30547 11925 30556
rect 12172 30596 12212 30883
rect 12172 30547 12212 30556
rect 11404 30437 11444 30522
rect 11788 30512 11828 30521
rect 11403 30428 11445 30437
rect 11403 30388 11404 30428
rect 11444 30388 11445 30428
rect 11403 30379 11445 30388
rect 11788 30269 11828 30472
rect 11979 30428 12021 30437
rect 11979 30388 11980 30428
rect 12020 30388 12021 30428
rect 12268 30428 12308 31051
rect 12363 30848 12405 30857
rect 12363 30808 12364 30848
rect 12404 30808 12405 30848
rect 12363 30799 12405 30808
rect 12364 30714 12404 30799
rect 12555 30764 12597 30773
rect 12555 30724 12556 30764
rect 12596 30724 12597 30764
rect 12555 30715 12597 30724
rect 12556 30680 12596 30715
rect 12556 30629 12596 30640
rect 12459 30428 12501 30437
rect 12268 30388 12404 30428
rect 11979 30379 12021 30388
rect 11403 30260 11445 30269
rect 11403 30220 11404 30260
rect 11444 30220 11445 30260
rect 11403 30211 11445 30220
rect 11787 30260 11829 30269
rect 11787 30220 11788 30260
rect 11828 30220 11829 30260
rect 11787 30211 11829 30220
rect 11404 29840 11444 30211
rect 11788 30008 11828 30017
rect 11404 29177 11444 29800
rect 11692 29968 11788 30008
rect 11595 29672 11637 29681
rect 11595 29632 11596 29672
rect 11636 29632 11637 29672
rect 11595 29623 11637 29632
rect 11596 29538 11636 29623
rect 11403 29168 11445 29177
rect 11403 29128 11404 29168
rect 11444 29128 11445 29168
rect 11403 29119 11445 29128
rect 11595 29168 11637 29177
rect 11595 29128 11596 29168
rect 11636 29128 11637 29168
rect 11595 29119 11637 29128
rect 11596 29034 11636 29119
rect 10636 28960 10868 29000
rect 11308 28960 11540 29000
rect 10636 28160 10676 28169
rect 10676 28120 10772 28160
rect 10636 28111 10676 28120
rect 10635 27992 10677 28001
rect 10635 27952 10636 27992
rect 10676 27952 10677 27992
rect 10635 27943 10677 27952
rect 10444 27532 10580 27572
rect 10347 27152 10389 27161
rect 10347 27112 10348 27152
rect 10388 27112 10389 27152
rect 10347 27103 10389 27112
rect 10251 26564 10293 26573
rect 10251 26524 10252 26564
rect 10292 26524 10293 26564
rect 10251 26515 10293 26524
rect 10252 26321 10292 26515
rect 10251 26312 10293 26321
rect 10251 26272 10252 26312
rect 10292 26272 10293 26312
rect 10251 26263 10293 26272
rect 10252 26144 10292 26153
rect 10155 24716 10197 24725
rect 10155 24676 10156 24716
rect 10196 24676 10197 24716
rect 10155 24667 10197 24676
rect 9868 24592 9964 24632
rect 9868 23969 9908 24592
rect 9964 24583 10004 24592
rect 10059 24632 10101 24641
rect 10059 24592 10060 24632
rect 10100 24592 10101 24632
rect 10059 24583 10101 24592
rect 9963 24464 10005 24473
rect 9963 24424 9964 24464
rect 10004 24424 10005 24464
rect 9963 24415 10005 24424
rect 9867 23960 9909 23969
rect 9867 23920 9868 23960
rect 9908 23920 9909 23960
rect 9867 23911 9909 23920
rect 9771 23876 9813 23885
rect 9771 23836 9772 23876
rect 9812 23836 9813 23876
rect 9771 23827 9813 23836
rect 9772 23742 9812 23827
rect 9868 23792 9908 23801
rect 9675 22784 9717 22793
rect 9675 22744 9676 22784
rect 9716 22744 9717 22784
rect 9675 22735 9717 22744
rect 9676 22364 9716 22735
rect 9676 22315 9716 22324
rect 9772 22280 9812 22289
rect 9675 21608 9717 21617
rect 9675 21568 9676 21608
rect 9716 21568 9717 21608
rect 9675 21559 9717 21568
rect 9676 21474 9716 21559
rect 9579 21356 9621 21365
rect 9579 21316 9580 21356
rect 9620 21316 9621 21356
rect 9579 21307 9621 21316
rect 9675 21272 9717 21281
rect 9675 21232 9676 21272
rect 9716 21232 9717 21272
rect 9675 21223 9717 21232
rect 9676 20777 9716 21223
rect 9675 20768 9717 20777
rect 9675 20728 9676 20768
rect 9716 20728 9717 20768
rect 9675 20719 9717 20728
rect 9676 20634 9716 20719
rect 9484 20600 9524 20609
rect 9524 20560 9620 20600
rect 9484 20551 9524 20560
rect 9483 20432 9525 20441
rect 9483 20392 9484 20432
rect 9524 20392 9525 20432
rect 9483 20383 9525 20392
rect 9387 19592 9429 19601
rect 9387 19552 9388 19592
rect 9428 19552 9429 19592
rect 9387 19543 9429 19552
rect 9484 19424 9524 20383
rect 9580 20105 9620 20560
rect 9579 20096 9621 20105
rect 9579 20056 9580 20096
rect 9620 20056 9621 20096
rect 9579 20047 9621 20056
rect 9772 19685 9812 22240
rect 9771 19676 9813 19685
rect 9771 19636 9772 19676
rect 9812 19636 9813 19676
rect 9771 19627 9813 19636
rect 9771 19508 9813 19517
rect 9771 19468 9772 19508
rect 9812 19468 9813 19508
rect 9771 19459 9813 19468
rect 9388 19384 9524 19424
rect 9291 18584 9333 18593
rect 9291 18544 9292 18584
rect 9332 18544 9333 18584
rect 9388 18584 9428 19384
rect 9676 19256 9716 19265
rect 9484 19216 9676 19256
rect 9484 18752 9524 19216
rect 9676 19207 9716 19216
rect 9772 19256 9812 19459
rect 9484 18703 9524 18712
rect 9676 18584 9716 18593
rect 9388 18544 9676 18584
rect 9291 18535 9333 18544
rect 9676 18535 9716 18544
rect 9292 18450 9332 18535
rect 9100 17872 9332 17912
rect 9195 17744 9237 17753
rect 9195 17704 9196 17744
rect 9236 17704 9237 17744
rect 9195 17695 9237 17704
rect 9196 17610 9236 17695
rect 9099 17576 9141 17585
rect 9099 17536 9100 17576
rect 9140 17536 9141 17576
rect 9099 17527 9141 17536
rect 9100 17442 9140 17527
rect 9003 17408 9045 17417
rect 9003 17368 9004 17408
rect 9044 17368 9045 17408
rect 9003 17359 9045 17368
rect 9003 17072 9045 17081
rect 9003 17032 9004 17072
rect 9044 17032 9045 17072
rect 9003 17023 9045 17032
rect 9100 17072 9140 17081
rect 9004 16938 9044 17023
rect 8907 16736 8949 16745
rect 8907 16696 8908 16736
rect 8948 16696 8949 16736
rect 8907 16687 8949 16696
rect 9100 16409 9140 17032
rect 9292 16913 9332 17872
rect 9579 17744 9621 17753
rect 9579 17704 9580 17744
rect 9620 17704 9621 17744
rect 9579 17695 9621 17704
rect 9580 17610 9620 17695
rect 9483 17576 9525 17585
rect 9483 17536 9484 17576
rect 9524 17536 9525 17576
rect 9483 17527 9525 17536
rect 9291 16904 9333 16913
rect 9291 16864 9292 16904
rect 9332 16864 9333 16904
rect 9291 16855 9333 16864
rect 9292 16484 9332 16855
rect 9388 16820 9428 16829
rect 9388 16661 9428 16780
rect 9387 16652 9429 16661
rect 9387 16612 9388 16652
rect 9428 16612 9429 16652
rect 9387 16603 9429 16612
rect 9292 16444 9428 16484
rect 9099 16400 9141 16409
rect 9099 16360 9100 16400
rect 9140 16360 9141 16400
rect 9099 16351 9141 16360
rect 8716 16232 8756 16241
rect 8620 16192 8716 16232
rect 8523 13208 8565 13217
rect 8523 13168 8524 13208
rect 8564 13168 8565 13208
rect 8523 13159 8565 13168
rect 8524 13074 8564 13159
rect 8428 12916 8564 12956
rect 8332 12536 8372 12545
rect 8372 12496 8468 12536
rect 8332 12487 8372 12496
rect 8331 12368 8373 12377
rect 8331 12328 8332 12368
rect 8372 12328 8373 12368
rect 8331 12319 8373 12328
rect 8332 11948 8372 12319
rect 8332 11899 8372 11908
rect 8180 11824 8276 11864
rect 8140 11815 8180 11824
rect 8331 11528 8373 11537
rect 8428 11528 8468 12496
rect 8331 11488 8332 11528
rect 8372 11488 8468 11528
rect 8331 11479 8373 11488
rect 8524 11444 8564 12916
rect 8620 11705 8660 16192
rect 8716 16183 8756 16192
rect 8908 16232 8948 16241
rect 9099 16232 9141 16241
rect 8948 16192 9044 16232
rect 8908 16183 8948 16192
rect 8812 16064 8852 16073
rect 8716 15546 8756 15555
rect 8716 14645 8756 15506
rect 8812 14897 8852 16024
rect 8907 15644 8949 15653
rect 8907 15604 8908 15644
rect 8948 15604 8949 15644
rect 8907 15595 8949 15604
rect 8908 15510 8948 15595
rect 8907 15392 8949 15401
rect 8907 15352 8908 15392
rect 8948 15352 8949 15392
rect 8907 15343 8949 15352
rect 8811 14888 8853 14897
rect 8811 14848 8812 14888
rect 8852 14848 8853 14888
rect 8811 14839 8853 14848
rect 8812 14720 8852 14729
rect 8715 14636 8757 14645
rect 8715 14596 8716 14636
rect 8756 14596 8757 14636
rect 8715 14587 8757 14596
rect 8812 14561 8852 14680
rect 8811 14552 8853 14561
rect 8811 14512 8812 14552
rect 8852 14512 8853 14552
rect 8811 14503 8853 14512
rect 8908 14384 8948 15343
rect 9004 15233 9044 16192
rect 9099 16192 9100 16232
rect 9140 16192 9141 16232
rect 9099 16183 9141 16192
rect 9196 16232 9236 16241
rect 9100 15401 9140 16183
rect 9196 15560 9236 16192
rect 9292 16232 9332 16241
rect 9388 16232 9428 16444
rect 9332 16192 9428 16232
rect 9292 16183 9332 16192
rect 9291 15644 9333 15653
rect 9291 15604 9292 15644
rect 9332 15604 9333 15644
rect 9291 15595 9333 15604
rect 9099 15392 9141 15401
rect 9099 15352 9100 15392
rect 9140 15352 9141 15392
rect 9099 15343 9141 15352
rect 9003 15224 9045 15233
rect 9003 15184 9004 15224
rect 9044 15184 9045 15224
rect 9003 15175 9045 15184
rect 9004 14972 9044 14981
rect 9196 14972 9236 15520
rect 9292 15560 9332 15595
rect 9292 15509 9332 15520
rect 9387 15560 9429 15569
rect 9387 15520 9388 15560
rect 9428 15520 9429 15560
rect 9387 15511 9429 15520
rect 9044 14932 9236 14972
rect 9004 14923 9044 14932
rect 9195 14720 9237 14729
rect 9195 14680 9196 14720
rect 9236 14680 9237 14720
rect 9195 14671 9237 14680
rect 9292 14720 9332 14729
rect 9196 14586 9236 14671
rect 8812 14344 8948 14384
rect 9195 14384 9237 14393
rect 9195 14344 9196 14384
rect 9236 14344 9237 14384
rect 8715 14216 8757 14225
rect 8715 14176 8716 14216
rect 8756 14176 8757 14216
rect 8715 14167 8757 14176
rect 8716 14048 8756 14167
rect 8716 12125 8756 14008
rect 8715 12116 8757 12125
rect 8715 12076 8716 12116
rect 8756 12076 8757 12116
rect 8715 12067 8757 12076
rect 8715 11948 8757 11957
rect 8715 11908 8716 11948
rect 8756 11908 8757 11948
rect 8715 11899 8757 11908
rect 8619 11696 8661 11705
rect 8619 11656 8620 11696
rect 8660 11656 8661 11696
rect 8619 11647 8661 11656
rect 8716 11696 8756 11899
rect 8620 11562 8660 11647
rect 8428 11404 8564 11444
rect 8428 11360 8468 11404
rect 8332 11320 8468 11360
rect 8619 11360 8661 11369
rect 8619 11320 8620 11360
rect 8660 11320 8661 11360
rect 8043 11108 8085 11117
rect 8043 11068 8044 11108
rect 8084 11068 8085 11108
rect 8043 11059 8085 11068
rect 7948 10975 7988 10984
rect 8235 11024 8277 11033
rect 8235 10984 8236 11024
rect 8276 10984 8277 11024
rect 8235 10975 8277 10984
rect 8043 10940 8085 10949
rect 8043 10900 8044 10940
rect 8084 10900 8085 10940
rect 8043 10891 8085 10900
rect 8044 10806 8084 10891
rect 7852 10312 8180 10352
rect 7756 10135 7796 10144
rect 7851 10184 7893 10193
rect 7851 10144 7852 10184
rect 7892 10144 7893 10184
rect 7851 10135 7893 10144
rect 7948 10184 7988 10193
rect 7852 10050 7892 10135
rect 7755 10016 7797 10025
rect 7755 9976 7756 10016
rect 7796 9976 7797 10016
rect 7755 9967 7797 9976
rect 7756 9521 7796 9967
rect 7755 9512 7797 9521
rect 7755 9472 7756 9512
rect 7796 9472 7797 9512
rect 7755 9463 7797 9472
rect 7948 9428 7988 10144
rect 8043 10184 8085 10193
rect 8043 10144 8044 10184
rect 8084 10144 8085 10184
rect 8043 10135 8085 10144
rect 8044 10050 8084 10135
rect 8140 10016 8180 10312
rect 8236 10184 8276 10975
rect 8236 10135 8276 10144
rect 8140 9976 8276 10016
rect 7852 9388 7988 9428
rect 7660 9304 7796 9344
rect 7660 8681 7700 8766
rect 7659 8672 7701 8681
rect 7659 8632 7660 8672
rect 7700 8632 7701 8672
rect 7659 8623 7701 8632
rect 7564 8464 7700 8504
rect 7467 8252 7509 8261
rect 7467 8212 7468 8252
rect 7508 8212 7509 8252
rect 7467 8203 7509 8212
rect 7468 8000 7508 8203
rect 7468 7951 7508 7960
rect 7564 8000 7604 8009
rect 7371 7748 7413 7757
rect 7371 7708 7372 7748
rect 7412 7708 7413 7748
rect 7371 7699 7413 7708
rect 7276 7540 7412 7580
rect 7276 7169 7316 7254
rect 7372 7244 7412 7540
rect 7564 7421 7604 7960
rect 7563 7412 7605 7421
rect 7563 7372 7564 7412
rect 7604 7372 7605 7412
rect 7563 7363 7605 7372
rect 7372 7204 7604 7244
rect 7275 7160 7317 7169
rect 7275 7120 7276 7160
rect 7316 7120 7317 7160
rect 7275 7111 7317 7120
rect 7275 6992 7317 7001
rect 7275 6952 7276 6992
rect 7316 6952 7317 6992
rect 7275 6943 7317 6952
rect 7467 6992 7509 7001
rect 7467 6952 7468 6992
rect 7508 6952 7509 6992
rect 7467 6943 7509 6952
rect 7179 5144 7221 5153
rect 7179 5104 7180 5144
rect 7220 5104 7221 5144
rect 7179 5095 7221 5104
rect 6891 5060 6933 5069
rect 6891 5020 6892 5060
rect 6932 5020 6933 5060
rect 6891 5011 6933 5020
rect 6795 4976 6837 4985
rect 6795 4936 6796 4976
rect 6836 4936 6837 4976
rect 6795 4927 6837 4936
rect 6507 4892 6549 4901
rect 6507 4852 6508 4892
rect 6548 4852 6644 4892
rect 6507 4843 6549 4852
rect 6124 4432 6260 4472
rect 6316 4768 6452 4808
rect 6124 4052 6164 4432
rect 6219 4304 6261 4313
rect 6219 4264 6220 4304
rect 6260 4264 6261 4304
rect 6219 4255 6261 4264
rect 6220 4170 6260 4255
rect 6124 4012 6260 4052
rect 6124 3450 6164 3475
rect 6124 3389 6164 3410
rect 6123 3380 6165 3389
rect 6123 3340 6124 3380
rect 6164 3340 6165 3380
rect 6123 3331 6165 3340
rect 6220 3053 6260 4012
rect 6316 3725 6356 4768
rect 6508 4758 6548 4843
rect 6508 4136 6548 4145
rect 6412 4096 6508 4136
rect 6412 3809 6452 4096
rect 6508 4087 6548 4096
rect 6604 4136 6644 4852
rect 6796 4304 6836 4927
rect 6987 4892 7029 4901
rect 6987 4852 6988 4892
rect 7028 4852 7029 4892
rect 6987 4843 7029 4852
rect 6988 4758 7028 4843
rect 7180 4724 7220 4733
rect 6988 4397 7028 4482
rect 6987 4388 7029 4397
rect 6987 4348 6988 4388
rect 7028 4348 7029 4388
rect 6987 4339 7029 4348
rect 6796 4264 6932 4304
rect 6796 4136 6836 4145
rect 6892 4136 6932 4264
rect 6604 3884 6644 4096
rect 6700 4115 6740 4124
rect 6836 4096 6932 4136
rect 7083 4136 7125 4145
rect 7083 4096 7084 4136
rect 7124 4096 7125 4136
rect 6796 4087 6836 4096
rect 7083 4087 7125 4096
rect 6700 3977 6740 4075
rect 7084 4002 7124 4087
rect 6699 3968 6741 3977
rect 6699 3928 6700 3968
rect 6740 3928 6741 3968
rect 6699 3919 6741 3928
rect 6508 3844 6644 3884
rect 6411 3800 6453 3809
rect 6411 3760 6412 3800
rect 6452 3760 6453 3800
rect 6411 3751 6453 3760
rect 6315 3716 6357 3725
rect 6315 3676 6316 3716
rect 6356 3676 6357 3716
rect 6315 3667 6357 3676
rect 6508 3632 6548 3844
rect 6315 3548 6357 3557
rect 6315 3508 6316 3548
rect 6356 3508 6357 3548
rect 6315 3499 6357 3508
rect 6316 3414 6356 3499
rect 6411 3296 6453 3305
rect 6411 3256 6412 3296
rect 6452 3256 6453 3296
rect 6411 3247 6453 3256
rect 6219 3044 6261 3053
rect 6219 3004 6220 3044
rect 6260 3004 6261 3044
rect 6219 2995 6261 3004
rect 6123 2792 6165 2801
rect 6123 2752 6124 2792
rect 6164 2752 6165 2792
rect 6123 2743 6165 2752
rect 6028 2659 6068 2668
rect 6124 2658 6164 2743
rect 6220 2708 6260 2995
rect 6220 2659 6260 2668
rect 6316 2633 6356 2718
rect 5740 2575 5780 2584
rect 5931 2624 5973 2633
rect 5931 2584 5932 2624
rect 5972 2584 5973 2624
rect 5931 2575 5973 2584
rect 6315 2624 6357 2633
rect 6315 2584 6316 2624
rect 6356 2584 6357 2624
rect 6315 2575 6357 2584
rect 5835 2540 5877 2549
rect 5835 2500 5836 2540
rect 5876 2500 5877 2540
rect 5835 2491 5877 2500
rect 6027 2540 6069 2549
rect 6027 2500 6028 2540
rect 6068 2500 6069 2540
rect 6027 2491 6069 2500
rect 5451 2456 5493 2465
rect 5451 2416 5452 2456
rect 5492 2416 5493 2456
rect 5451 2407 5493 2416
rect 5452 1205 5492 2407
rect 5739 2288 5781 2297
rect 5739 2248 5740 2288
rect 5780 2248 5781 2288
rect 5739 2239 5781 2248
rect 5547 2120 5589 2129
rect 5547 2080 5548 2120
rect 5588 2080 5589 2120
rect 5547 2071 5589 2080
rect 5740 2120 5780 2239
rect 5740 2071 5780 2080
rect 5548 1947 5588 2071
rect 5548 1898 5588 1907
rect 5643 1280 5685 1289
rect 5643 1240 5644 1280
rect 5684 1240 5685 1280
rect 5643 1231 5685 1240
rect 5451 1196 5493 1205
rect 5451 1156 5452 1196
rect 5492 1156 5493 1196
rect 5451 1147 5493 1156
rect 5644 1196 5684 1231
rect 5644 1145 5684 1156
rect 5355 1112 5397 1121
rect 5836 1112 5876 2491
rect 5931 2204 5973 2213
rect 5931 2164 5932 2204
rect 5972 2164 5973 2204
rect 5931 2155 5973 2164
rect 5932 1868 5972 2155
rect 5932 1819 5972 1828
rect 5355 1072 5356 1112
rect 5396 1072 5397 1112
rect 5355 1063 5397 1072
rect 5740 1072 5876 1112
rect 6028 1112 6068 2491
rect 6412 1952 6452 3247
rect 6508 2792 6548 3592
rect 6795 3632 6837 3641
rect 7180 3632 7220 4684
rect 7276 4136 7316 6943
rect 7371 6236 7413 6245
rect 7371 6196 7372 6236
rect 7412 6196 7413 6236
rect 7371 6187 7413 6196
rect 7372 5741 7412 6187
rect 7371 5732 7413 5741
rect 7371 5692 7372 5732
rect 7412 5692 7413 5732
rect 7371 5683 7413 5692
rect 7372 5648 7412 5683
rect 7372 5597 7412 5608
rect 7371 5228 7413 5237
rect 7371 5188 7372 5228
rect 7412 5188 7413 5228
rect 7371 5179 7413 5188
rect 7372 5060 7412 5179
rect 7372 5011 7412 5020
rect 7276 4087 7316 4096
rect 7468 4136 7508 6943
rect 7564 6908 7604 7204
rect 7660 7160 7700 8464
rect 7660 7111 7700 7120
rect 7756 7160 7796 9304
rect 7852 8588 7892 9388
rect 8140 9344 8180 9353
rect 7948 9260 7988 9269
rect 7948 8849 7988 9220
rect 8140 9092 8180 9304
rect 8044 9052 8180 9092
rect 7947 8840 7989 8849
rect 7947 8800 7948 8840
rect 7988 8800 7989 8840
rect 7947 8791 7989 8800
rect 7852 8548 7988 8588
rect 7756 7111 7796 7120
rect 7851 7160 7893 7169
rect 7851 7120 7852 7160
rect 7892 7120 7893 7160
rect 7851 7111 7893 7120
rect 7948 7160 7988 8548
rect 8044 8513 8084 9052
rect 8139 8840 8181 8849
rect 8139 8800 8140 8840
rect 8180 8800 8181 8840
rect 8139 8791 8181 8800
rect 8140 8686 8180 8791
rect 8140 8637 8180 8646
rect 8043 8504 8085 8513
rect 8043 8464 8044 8504
rect 8084 8464 8085 8504
rect 8043 8455 8085 8464
rect 8043 8000 8085 8009
rect 8043 7960 8044 8000
rect 8084 7960 8085 8000
rect 8043 7951 8085 7960
rect 8044 7866 8084 7951
rect 8236 7421 8276 9976
rect 8332 9512 8372 11320
rect 8619 11311 8661 11320
rect 8523 11108 8565 11117
rect 8523 11068 8524 11108
rect 8564 11068 8565 11108
rect 8523 11059 8565 11068
rect 8428 11024 8468 11033
rect 8428 10445 8468 10984
rect 8524 11024 8564 11059
rect 8427 10436 8469 10445
rect 8427 10396 8428 10436
rect 8468 10396 8469 10436
rect 8427 10387 8469 10396
rect 8524 10193 8564 10984
rect 8523 10184 8565 10193
rect 8523 10144 8524 10184
rect 8564 10144 8565 10184
rect 8523 10135 8565 10144
rect 8372 9472 8468 9512
rect 8332 9463 8372 9472
rect 8331 8504 8373 8513
rect 8331 8464 8332 8504
rect 8372 8464 8373 8504
rect 8428 8504 8468 9472
rect 8523 9428 8565 9437
rect 8523 9388 8524 9428
rect 8564 9388 8565 9428
rect 8523 9379 8565 9388
rect 8524 9017 8564 9379
rect 8620 9185 8660 11311
rect 8619 9176 8661 9185
rect 8619 9136 8620 9176
rect 8660 9136 8661 9176
rect 8619 9127 8661 9136
rect 8523 9008 8565 9017
rect 8523 8968 8524 9008
rect 8564 8968 8565 9008
rect 8523 8959 8565 8968
rect 8524 8672 8564 8959
rect 8619 8756 8661 8765
rect 8619 8716 8620 8756
rect 8660 8716 8661 8756
rect 8619 8707 8661 8716
rect 8524 8623 8564 8632
rect 8428 8464 8564 8504
rect 8331 8455 8373 8464
rect 8332 8370 8372 8455
rect 8331 7748 8373 7757
rect 8331 7708 8332 7748
rect 8372 7708 8373 7748
rect 8331 7699 8373 7708
rect 8235 7412 8277 7421
rect 8235 7372 8236 7412
rect 8276 7372 8277 7412
rect 8235 7363 8277 7372
rect 8140 7328 8180 7337
rect 8044 7288 8140 7328
rect 8044 7169 8084 7288
rect 8140 7279 8180 7288
rect 8332 7302 8372 7699
rect 8427 7496 8469 7505
rect 8427 7456 8428 7496
rect 8468 7456 8469 7496
rect 8427 7447 8469 7456
rect 8332 7253 8372 7262
rect 7948 7111 7988 7120
rect 8043 7160 8085 7169
rect 8043 7120 8044 7160
rect 8084 7120 8085 7160
rect 8043 7111 8085 7120
rect 8332 7152 8372 7161
rect 7852 7026 7892 7111
rect 8332 7076 8372 7112
rect 8236 7036 8372 7076
rect 8236 6908 8276 7036
rect 7564 6868 8276 6908
rect 8331 6908 8373 6917
rect 8331 6868 8332 6908
rect 8372 6868 8373 6908
rect 8331 6859 8373 6868
rect 8332 6740 8372 6859
rect 8236 6700 8372 6740
rect 8043 6656 8085 6665
rect 8043 6616 8044 6656
rect 8084 6616 8085 6656
rect 8043 6607 8085 6616
rect 7564 6497 7604 6582
rect 7563 6488 7605 6497
rect 7563 6448 7564 6488
rect 7604 6448 7605 6488
rect 7563 6439 7605 6448
rect 8044 6488 8084 6607
rect 8044 6439 8084 6448
rect 8140 6488 8180 6497
rect 7659 6404 7701 6413
rect 7659 6364 7660 6404
rect 7700 6364 7701 6404
rect 7659 6355 7701 6364
rect 7563 6320 7605 6329
rect 7563 6280 7564 6320
rect 7604 6280 7605 6320
rect 7563 6271 7605 6280
rect 7564 5900 7604 6271
rect 7660 6270 7700 6355
rect 8043 6320 8085 6329
rect 8043 6280 8044 6320
rect 8084 6280 8085 6320
rect 8043 6271 8085 6280
rect 7564 5851 7604 5860
rect 7948 5653 7988 5662
rect 7756 5480 7796 5489
rect 7468 4087 7508 4096
rect 7564 5440 7756 5480
rect 7372 3968 7412 3979
rect 7564 3968 7604 5440
rect 7756 5431 7796 5440
rect 7948 5153 7988 5613
rect 7947 5144 7989 5153
rect 7947 5104 7948 5144
rect 7988 5104 7989 5144
rect 7947 5095 7989 5104
rect 7756 4985 7796 5070
rect 7660 4976 7700 4985
rect 7660 4472 7700 4936
rect 7755 4976 7797 4985
rect 7755 4936 7756 4976
rect 7796 4936 7797 4976
rect 7755 4927 7797 4936
rect 7948 4976 7988 4985
rect 7755 4808 7797 4817
rect 7755 4768 7756 4808
rect 7796 4768 7797 4808
rect 7755 4759 7797 4768
rect 7756 4674 7796 4759
rect 7948 4565 7988 4936
rect 7947 4556 7989 4565
rect 7947 4516 7948 4556
rect 7988 4516 7989 4556
rect 7947 4507 7989 4516
rect 7660 4432 7796 4472
rect 7659 4304 7701 4313
rect 7659 4264 7660 4304
rect 7700 4264 7701 4304
rect 7659 4255 7701 4264
rect 7660 4136 7700 4255
rect 7660 4087 7700 4096
rect 7564 3928 7700 3968
rect 7372 3893 7412 3928
rect 7371 3884 7413 3893
rect 7371 3844 7372 3884
rect 7412 3844 7413 3884
rect 7371 3835 7413 3844
rect 6795 3592 6796 3632
rect 6836 3592 6837 3632
rect 6795 3583 6837 3592
rect 7084 3592 7220 3632
rect 6796 3464 6836 3583
rect 6796 3415 6836 3424
rect 6508 2743 6548 2752
rect 6988 2633 7028 2718
rect 6892 2624 6932 2633
rect 6892 2036 6932 2584
rect 6987 2624 7029 2633
rect 6987 2584 6988 2624
rect 7028 2584 7029 2624
rect 6987 2575 7029 2584
rect 6796 1996 6932 2036
rect 6412 1903 6452 1912
rect 6507 1952 6549 1961
rect 6507 1912 6508 1952
rect 6548 1912 6549 1952
rect 6507 1903 6549 1912
rect 6508 1818 6548 1903
rect 6796 1793 6836 1996
rect 6987 1952 7029 1961
rect 6987 1912 6988 1952
rect 7028 1912 7029 1952
rect 6987 1903 7029 1912
rect 6891 1868 6933 1877
rect 6891 1828 6892 1868
rect 6932 1828 6933 1868
rect 6891 1819 6933 1828
rect 6795 1784 6837 1793
rect 6795 1744 6796 1784
rect 6836 1744 6837 1784
rect 6795 1735 6837 1744
rect 6892 1734 6932 1819
rect 6988 1818 7028 1903
rect 6123 1700 6165 1709
rect 6123 1660 6124 1700
rect 6164 1660 6165 1700
rect 6123 1651 6165 1660
rect 6124 1566 6164 1651
rect 6219 1280 6261 1289
rect 6219 1240 6220 1280
rect 6260 1240 6261 1280
rect 6219 1231 6261 1240
rect 6603 1280 6645 1289
rect 6603 1240 6604 1280
rect 6644 1240 6645 1280
rect 6603 1231 6645 1240
rect 6795 1280 6837 1289
rect 6795 1240 6796 1280
rect 6836 1240 6837 1280
rect 6795 1231 6837 1240
rect 6987 1280 7029 1289
rect 6987 1240 6988 1280
rect 7028 1240 7029 1280
rect 6987 1231 7029 1240
rect 6123 1196 6165 1205
rect 6123 1156 6124 1196
rect 6164 1156 6165 1196
rect 6123 1147 6165 1156
rect 4875 1028 4917 1037
rect 5740 1028 5780 1072
rect 6028 1063 6068 1072
rect 4875 988 4876 1028
rect 4916 988 4917 1028
rect 4875 979 4917 988
rect 5644 988 5780 1028
rect 5068 944 5108 953
rect 5452 944 5492 953
rect 5108 904 5396 944
rect 5068 895 5108 904
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 4875 608 4917 617
rect 4875 568 4876 608
rect 4916 568 4917 608
rect 4875 559 4917 568
rect 5259 608 5301 617
rect 5259 568 5260 608
rect 5300 568 5301 608
rect 5259 559 5301 568
rect 4876 80 4916 559
rect 5067 104 5109 113
rect 5067 80 5068 104
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 64 5068 80
rect 5108 80 5109 104
rect 5260 80 5300 559
rect 5356 281 5396 904
rect 5492 904 5588 944
rect 5452 895 5492 904
rect 5451 692 5493 701
rect 5451 652 5452 692
rect 5492 652 5493 692
rect 5451 643 5493 652
rect 5355 272 5397 281
rect 5355 232 5356 272
rect 5396 232 5397 272
rect 5355 223 5397 232
rect 5452 80 5492 643
rect 5548 449 5588 904
rect 5547 440 5589 449
rect 5547 400 5548 440
rect 5588 400 5589 440
rect 5547 391 5589 400
rect 5644 80 5684 988
rect 5836 944 5876 953
rect 6027 944 6069 953
rect 5876 904 5972 944
rect 5836 895 5876 904
rect 5835 692 5877 701
rect 5835 652 5836 692
rect 5876 652 5877 692
rect 5835 643 5877 652
rect 5836 80 5876 643
rect 5932 533 5972 904
rect 6027 904 6028 944
rect 6068 904 6069 944
rect 6027 895 6069 904
rect 5931 524 5973 533
rect 5931 484 5932 524
rect 5972 484 5973 524
rect 5931 475 5973 484
rect 6028 80 6068 895
rect 6124 197 6164 1147
rect 6123 188 6165 197
rect 6123 148 6124 188
rect 6164 148 6165 188
rect 6123 139 6165 148
rect 6220 80 6260 1231
rect 6411 608 6453 617
rect 6411 568 6412 608
rect 6452 568 6453 608
rect 6411 559 6453 568
rect 6412 80 6452 559
rect 6604 80 6644 1231
rect 6796 80 6836 1231
rect 6988 80 7028 1231
rect 7084 1121 7124 3592
rect 7467 3044 7509 3053
rect 7467 3004 7468 3044
rect 7508 3004 7509 3044
rect 7467 2995 7509 3004
rect 7371 2960 7413 2969
rect 7371 2920 7372 2960
rect 7412 2920 7413 2960
rect 7371 2911 7413 2920
rect 7372 2708 7412 2911
rect 7372 2659 7412 2668
rect 7468 2708 7508 2995
rect 7468 2659 7508 2668
rect 7563 2540 7605 2549
rect 7563 2500 7564 2540
rect 7604 2500 7605 2540
rect 7563 2491 7605 2500
rect 7467 2372 7509 2381
rect 7467 2332 7468 2372
rect 7508 2332 7509 2372
rect 7467 2323 7509 2332
rect 7468 1952 7508 2323
rect 7468 1903 7508 1912
rect 7275 1364 7317 1373
rect 7275 1324 7276 1364
rect 7316 1324 7317 1364
rect 7275 1315 7317 1324
rect 7179 1280 7221 1289
rect 7179 1240 7180 1280
rect 7220 1240 7221 1280
rect 7179 1231 7221 1240
rect 7083 1112 7125 1121
rect 7083 1072 7084 1112
rect 7124 1072 7125 1112
rect 7083 1063 7125 1072
rect 7180 80 7220 1231
rect 7276 1112 7316 1315
rect 7468 1280 7508 1291
rect 7468 1205 7508 1240
rect 7467 1196 7509 1205
rect 7467 1156 7468 1196
rect 7508 1156 7509 1196
rect 7467 1147 7509 1156
rect 7564 1112 7604 2491
rect 7660 2213 7700 3928
rect 7756 2801 7796 4432
rect 8044 3968 8084 6271
rect 8140 5909 8180 6448
rect 8139 5900 8181 5909
rect 8139 5860 8140 5900
rect 8180 5860 8181 5900
rect 8139 5851 8181 5860
rect 8236 5312 8276 6700
rect 8428 6665 8468 7447
rect 8524 7253 8564 8464
rect 8620 8093 8660 8707
rect 8716 8681 8756 11656
rect 8812 11024 8852 14344
rect 9195 14335 9237 14344
rect 8907 14132 8949 14141
rect 8907 14092 8908 14132
rect 8948 14092 8949 14132
rect 8907 14083 8949 14092
rect 8908 13998 8948 14083
rect 9100 14006 9140 14015
rect 9196 14006 9236 14335
rect 9140 13966 9236 14006
rect 9100 13957 9140 13966
rect 9004 11696 9044 11707
rect 9004 11621 9044 11656
rect 9196 11621 9236 13966
rect 9292 12209 9332 14680
rect 9388 13889 9428 15511
rect 9484 15308 9524 17527
rect 9772 17324 9812 19216
rect 9868 19088 9908 23752
rect 9964 22280 10004 24415
rect 10156 24389 10196 24474
rect 10155 24380 10197 24389
rect 10155 24340 10156 24380
rect 10196 24340 10197 24380
rect 10155 24331 10197 24340
rect 10059 22952 10101 22961
rect 10059 22912 10060 22952
rect 10100 22912 10101 22952
rect 10059 22903 10101 22912
rect 10060 22709 10100 22903
rect 10252 22793 10292 26104
rect 10348 25388 10388 27103
rect 10444 26825 10484 27532
rect 10636 27488 10676 27943
rect 10540 27448 10676 27488
rect 10540 26900 10580 27448
rect 10635 27320 10677 27329
rect 10635 27280 10636 27320
rect 10676 27280 10677 27320
rect 10635 27271 10677 27280
rect 10636 26909 10676 27271
rect 10443 26816 10485 26825
rect 10443 26776 10444 26816
rect 10484 26776 10485 26816
rect 10443 26767 10485 26776
rect 10443 25892 10485 25901
rect 10443 25852 10444 25892
rect 10484 25852 10485 25892
rect 10443 25843 10485 25852
rect 10348 25339 10388 25348
rect 10444 24632 10484 25843
rect 10540 25733 10580 26860
rect 10635 26900 10677 26909
rect 10635 26860 10636 26900
rect 10676 26860 10677 26900
rect 10635 26851 10677 26860
rect 10636 26766 10676 26851
rect 10732 26139 10772 28120
rect 10732 26090 10772 26099
rect 10635 25976 10677 25985
rect 10635 25936 10636 25976
rect 10676 25936 10677 25976
rect 10635 25927 10677 25936
rect 10539 25724 10581 25733
rect 10539 25684 10540 25724
rect 10580 25684 10581 25724
rect 10539 25675 10581 25684
rect 10539 25556 10581 25565
rect 10539 25516 10540 25556
rect 10580 25516 10581 25556
rect 10539 25507 10581 25516
rect 10540 25422 10580 25507
rect 10444 24583 10484 24592
rect 10540 24632 10580 24641
rect 10348 23792 10388 23801
rect 10348 23633 10388 23752
rect 10540 23717 10580 24592
rect 10539 23708 10581 23717
rect 10539 23668 10540 23708
rect 10580 23668 10581 23708
rect 10539 23659 10581 23668
rect 10347 23624 10389 23633
rect 10347 23584 10348 23624
rect 10388 23584 10389 23624
rect 10347 23575 10389 23584
rect 10347 23456 10389 23465
rect 10347 23416 10348 23456
rect 10388 23416 10389 23456
rect 10347 23407 10389 23416
rect 10251 22784 10293 22793
rect 10251 22744 10252 22784
rect 10292 22744 10293 22784
rect 10251 22735 10293 22744
rect 10059 22700 10101 22709
rect 10059 22660 10060 22700
rect 10100 22660 10101 22700
rect 10059 22651 10101 22660
rect 10251 22616 10293 22625
rect 10251 22576 10252 22616
rect 10292 22576 10293 22616
rect 10251 22567 10293 22576
rect 10059 22280 10101 22289
rect 9964 22240 10060 22280
rect 10100 22240 10101 22280
rect 10059 22231 10101 22240
rect 10252 22280 10292 22567
rect 10252 22231 10292 22240
rect 10060 22028 10100 22231
rect 10060 21988 10196 22028
rect 9963 20096 10005 20105
rect 9963 20056 9964 20096
rect 10004 20056 10005 20096
rect 9963 20047 10005 20056
rect 10060 20096 10100 20105
rect 9964 19962 10004 20047
rect 10060 19844 10100 20056
rect 9964 19804 10100 19844
rect 9964 19517 10004 19804
rect 10059 19676 10101 19685
rect 10059 19636 10060 19676
rect 10100 19636 10101 19676
rect 10059 19627 10101 19636
rect 9963 19508 10005 19517
rect 9963 19468 9964 19508
rect 10004 19468 10005 19508
rect 9963 19459 10005 19468
rect 9868 19048 10004 19088
rect 9867 18920 9909 18929
rect 9867 18880 9868 18920
rect 9908 18880 9909 18920
rect 9867 18871 9909 18880
rect 9676 17284 9812 17324
rect 9579 17156 9621 17165
rect 9579 17116 9580 17156
rect 9620 17116 9621 17156
rect 9579 17107 9621 17116
rect 9580 17022 9620 17107
rect 9676 16325 9716 17284
rect 9771 17156 9813 17165
rect 9771 17116 9772 17156
rect 9812 17116 9813 17156
rect 9771 17107 9813 17116
rect 9772 17072 9812 17107
rect 9772 17021 9812 17032
rect 9675 16316 9717 16325
rect 9675 16276 9676 16316
rect 9716 16276 9717 16316
rect 9675 16267 9717 16276
rect 9676 16182 9716 16267
rect 9772 16232 9812 16241
rect 9772 16073 9812 16192
rect 9771 16064 9813 16073
rect 9771 16024 9772 16064
rect 9812 16024 9813 16064
rect 9771 16015 9813 16024
rect 9675 15896 9717 15905
rect 9675 15856 9676 15896
rect 9716 15856 9717 15896
rect 9675 15847 9717 15856
rect 9676 15560 9716 15847
rect 9772 15560 9812 15569
rect 9868 15560 9908 18871
rect 9964 17249 10004 19048
rect 9963 17240 10005 17249
rect 9963 17200 9964 17240
rect 10004 17200 10005 17240
rect 9963 17191 10005 17200
rect 9964 16241 10004 17191
rect 9963 16232 10005 16241
rect 9963 16192 9964 16232
rect 10004 16192 10005 16232
rect 9963 16183 10005 16192
rect 9963 15980 10005 15989
rect 10060 15980 10100 19627
rect 9963 15940 9964 15980
rect 10004 15940 10100 15980
rect 10156 19256 10196 21988
rect 9963 15931 10005 15940
rect 9676 15511 9716 15520
rect 9769 15520 9772 15545
rect 9812 15520 9908 15560
rect 9769 15505 9812 15520
rect 9769 15401 9809 15505
rect 9769 15392 9813 15401
rect 9769 15352 9772 15392
rect 9812 15352 9813 15392
rect 9771 15343 9813 15352
rect 9484 15268 9620 15308
rect 9483 15140 9525 15149
rect 9483 15100 9484 15140
rect 9524 15100 9525 15140
rect 9483 15091 9525 15100
rect 9484 14552 9524 15091
rect 9484 14503 9524 14512
rect 9387 13880 9429 13889
rect 9387 13840 9388 13880
rect 9428 13840 9429 13880
rect 9387 13831 9429 13840
rect 9580 12704 9620 15268
rect 9771 15224 9813 15233
rect 9771 15184 9772 15224
rect 9812 15184 9813 15224
rect 9771 15175 9813 15184
rect 9675 14720 9717 14729
rect 9675 14680 9676 14720
rect 9716 14680 9717 14720
rect 9675 14671 9717 14680
rect 9772 14720 9812 15175
rect 9964 14981 10004 15931
rect 10156 15905 10196 19216
rect 10252 19256 10292 19265
rect 10252 19181 10292 19216
rect 10250 19172 10292 19181
rect 10250 19132 10251 19172
rect 10291 19132 10292 19172
rect 10250 19123 10292 19132
rect 10251 16232 10293 16241
rect 10251 16192 10252 16232
rect 10292 16192 10293 16232
rect 10251 16183 10293 16192
rect 10252 16098 10292 16183
rect 10155 15896 10197 15905
rect 10155 15856 10156 15896
rect 10196 15856 10197 15896
rect 10155 15847 10197 15856
rect 10252 15560 10292 15569
rect 10060 15520 10252 15560
rect 9963 14972 10005 14981
rect 9963 14932 9964 14972
rect 10004 14932 10005 14972
rect 9963 14923 10005 14932
rect 9963 14804 10005 14813
rect 9963 14764 9964 14804
rect 10004 14764 10005 14804
rect 9963 14755 10005 14764
rect 9676 14477 9716 14671
rect 9675 14468 9717 14477
rect 9675 14428 9676 14468
rect 9716 14428 9717 14468
rect 9675 14419 9717 14428
rect 9675 13628 9717 13637
rect 9675 13588 9676 13628
rect 9716 13588 9717 13628
rect 9675 13579 9717 13588
rect 9676 13292 9716 13579
rect 9772 13469 9812 14680
rect 9868 14720 9908 14729
rect 9771 13460 9813 13469
rect 9771 13420 9772 13460
rect 9812 13420 9813 13460
rect 9771 13411 9813 13420
rect 9676 13252 9812 13292
rect 9772 13250 9812 13252
rect 9772 13201 9812 13210
rect 9771 12704 9813 12713
rect 9580 12664 9716 12704
rect 9580 12536 9620 12545
rect 9291 12200 9333 12209
rect 9291 12160 9292 12200
rect 9332 12160 9333 12200
rect 9291 12151 9333 12160
rect 9580 12125 9620 12496
rect 9676 12461 9716 12664
rect 9771 12664 9772 12704
rect 9812 12664 9813 12704
rect 9771 12655 9813 12664
rect 9772 12570 9812 12655
rect 9675 12452 9717 12461
rect 9675 12412 9676 12452
rect 9716 12412 9717 12452
rect 9675 12403 9717 12412
rect 9868 12368 9908 14680
rect 9964 14720 10004 14755
rect 9964 14669 10004 14680
rect 9963 14552 10005 14561
rect 9963 14512 9964 14552
rect 10004 14512 10005 14552
rect 9963 14503 10005 14512
rect 9964 14393 10004 14503
rect 9963 14384 10005 14393
rect 9963 14344 9964 14384
rect 10004 14344 10005 14384
rect 9963 14335 10005 14344
rect 9963 14216 10005 14225
rect 9963 14176 9964 14216
rect 10004 14176 10005 14216
rect 9963 14167 10005 14176
rect 9964 13460 10004 14167
rect 10060 14048 10100 15520
rect 10252 15511 10292 15520
rect 10348 15149 10388 23407
rect 10443 23120 10485 23129
rect 10443 23080 10444 23120
rect 10484 23080 10485 23120
rect 10443 23071 10485 23080
rect 10444 21617 10484 23071
rect 10539 22700 10581 22709
rect 10539 22660 10540 22700
rect 10580 22660 10581 22700
rect 10539 22651 10581 22660
rect 10540 21944 10580 22651
rect 10636 22112 10676 25927
rect 10731 25388 10773 25397
rect 10731 25348 10732 25388
rect 10772 25348 10773 25388
rect 10731 25339 10773 25348
rect 10732 25304 10772 25339
rect 10828 25313 10868 28960
rect 11307 28748 11349 28757
rect 11307 28708 11308 28748
rect 11348 28708 11349 28748
rect 11307 28699 11349 28708
rect 11211 28664 11253 28673
rect 11211 28624 11212 28664
rect 11252 28624 11253 28664
rect 11211 28615 11253 28624
rect 11019 28496 11061 28505
rect 11019 28456 11020 28496
rect 11060 28456 11061 28496
rect 11019 28447 11061 28456
rect 10923 28328 10965 28337
rect 10923 28288 10924 28328
rect 10964 28288 10965 28328
rect 10923 28279 10965 28288
rect 11020 28328 11060 28447
rect 11020 28279 11060 28288
rect 11116 28328 11156 28337
rect 11212 28328 11252 28615
rect 11308 28580 11348 28699
rect 11308 28531 11348 28540
rect 11308 28337 11348 28422
rect 11156 28288 11252 28328
rect 11307 28328 11349 28337
rect 11307 28288 11308 28328
rect 11348 28288 11349 28328
rect 11116 28279 11156 28288
rect 11307 28279 11349 28288
rect 11500 28328 11540 28960
rect 11692 28505 11732 29968
rect 11788 29959 11828 29968
rect 11980 29168 12020 30379
rect 12364 29933 12404 30388
rect 12459 30388 12460 30428
rect 12500 30388 12501 30428
rect 12459 30379 12501 30388
rect 12363 29924 12405 29933
rect 12363 29884 12364 29924
rect 12404 29884 12405 29924
rect 12363 29875 12405 29884
rect 12172 29840 12212 29849
rect 12075 29756 12117 29765
rect 12075 29716 12076 29756
rect 12116 29716 12117 29756
rect 12075 29707 12117 29716
rect 12076 29622 12116 29707
rect 12076 29168 12116 29177
rect 11980 29128 12076 29168
rect 11787 29000 11829 29009
rect 11787 28960 11788 29000
rect 11828 28960 11829 29000
rect 11787 28951 11829 28960
rect 11788 28866 11828 28951
rect 11691 28496 11733 28505
rect 11691 28456 11692 28496
rect 11732 28456 11733 28496
rect 11691 28447 11733 28456
rect 11979 28496 12021 28505
rect 11979 28456 11980 28496
rect 12020 28456 12021 28496
rect 11979 28447 12021 28456
rect 10924 26480 10964 28279
rect 11403 27656 11445 27665
rect 11403 27616 11404 27656
rect 11444 27616 11445 27656
rect 11403 27607 11445 27616
rect 11116 26816 11156 26827
rect 11116 26741 11156 26776
rect 11115 26732 11157 26741
rect 11115 26692 11116 26732
rect 11156 26692 11348 26732
rect 11115 26683 11157 26692
rect 10924 26440 11060 26480
rect 10923 26312 10965 26321
rect 10923 26272 10924 26312
rect 10964 26272 10965 26312
rect 10923 26263 10965 26272
rect 10924 26178 10964 26263
rect 10732 25253 10772 25264
rect 10827 25304 10869 25313
rect 10827 25264 10828 25304
rect 10868 25264 10869 25304
rect 10827 25255 10869 25264
rect 11020 24716 11060 26440
rect 11116 26144 11156 26155
rect 11116 26069 11156 26104
rect 11211 26144 11253 26153
rect 11211 26104 11212 26144
rect 11252 26104 11253 26144
rect 11211 26095 11253 26104
rect 11115 26060 11157 26069
rect 11115 26020 11116 26060
rect 11156 26020 11157 26060
rect 11115 26011 11157 26020
rect 11020 24676 11156 24716
rect 11116 24557 11156 24676
rect 10923 24548 10965 24557
rect 10923 24508 10924 24548
rect 10964 24508 10965 24548
rect 10923 24499 10965 24508
rect 11020 24548 11060 24557
rect 10924 24414 10964 24499
rect 10827 24380 10869 24389
rect 10827 24340 10828 24380
rect 10868 24340 10869 24380
rect 10827 24331 10869 24340
rect 10731 23960 10773 23969
rect 10731 23920 10732 23960
rect 10772 23920 10773 23960
rect 10731 23911 10773 23920
rect 10732 23129 10772 23911
rect 10828 23806 10868 24331
rect 11020 23876 11060 24508
rect 11115 24548 11157 24557
rect 11115 24508 11116 24548
rect 11156 24508 11157 24548
rect 11115 24499 11157 24508
rect 11212 24044 11252 26095
rect 10828 23757 10868 23766
rect 10924 23836 11060 23876
rect 11115 24004 11252 24044
rect 10924 23549 10964 23836
rect 11020 23708 11060 23717
rect 11115 23708 11155 24004
rect 11308 23960 11348 26692
rect 11404 25901 11444 27607
rect 11500 27161 11540 28288
rect 11595 28328 11637 28337
rect 11595 28288 11596 28328
rect 11636 28288 11637 28328
rect 11595 28279 11637 28288
rect 11692 28328 11732 28337
rect 11732 28288 11924 28328
rect 11692 28279 11732 28288
rect 11596 28194 11636 28279
rect 11787 28160 11829 28169
rect 11787 28120 11788 28160
rect 11828 28120 11829 28160
rect 11787 28111 11829 28120
rect 11788 28026 11828 28111
rect 11691 27908 11733 27917
rect 11691 27868 11692 27908
rect 11732 27868 11733 27908
rect 11691 27859 11733 27868
rect 11596 27404 11636 27413
rect 11499 27152 11541 27161
rect 11499 27112 11500 27152
rect 11540 27112 11541 27152
rect 11499 27103 11541 27112
rect 11499 26984 11541 26993
rect 11499 26944 11500 26984
rect 11540 26944 11541 26984
rect 11499 26935 11541 26944
rect 11500 26573 11540 26935
rect 11596 26830 11636 27364
rect 11596 26781 11636 26790
rect 11499 26564 11541 26573
rect 11499 26524 11500 26564
rect 11540 26524 11541 26564
rect 11499 26515 11541 26524
rect 11403 25892 11445 25901
rect 11403 25852 11404 25892
rect 11444 25852 11445 25892
rect 11403 25843 11445 25852
rect 11595 25388 11637 25397
rect 11595 25348 11596 25388
rect 11636 25348 11637 25388
rect 11595 25339 11637 25348
rect 11060 23668 11155 23708
rect 11212 23920 11348 23960
rect 11500 24632 11540 24641
rect 11020 23659 11060 23668
rect 10923 23540 10965 23549
rect 10923 23500 10924 23540
rect 10964 23500 10965 23540
rect 10923 23491 10965 23500
rect 10731 23120 10773 23129
rect 10731 23080 10732 23120
rect 10772 23080 10773 23120
rect 10731 23071 10773 23080
rect 10732 22986 10772 23071
rect 11212 22952 11252 23920
rect 11308 23792 11348 23801
rect 11348 23752 11360 23792
rect 11308 23743 11360 23752
rect 11320 23708 11360 23743
rect 11403 23708 11445 23717
rect 11320 23668 11404 23708
rect 11444 23668 11445 23708
rect 11403 23659 11445 23668
rect 11404 23120 11444 23129
rect 11212 22912 11348 22952
rect 10924 22868 10964 22877
rect 10964 22828 11252 22868
rect 10924 22819 10964 22828
rect 10780 22289 10820 22298
rect 11212 22280 11252 22828
rect 11308 22457 11348 22912
rect 11404 22877 11444 23080
rect 11403 22868 11445 22877
rect 11403 22828 11404 22868
rect 11444 22828 11445 22868
rect 11403 22819 11445 22828
rect 11403 22616 11445 22625
rect 11403 22576 11404 22616
rect 11444 22576 11445 22616
rect 11403 22567 11445 22576
rect 11307 22448 11349 22457
rect 11307 22408 11308 22448
rect 11348 22408 11349 22448
rect 11307 22399 11349 22408
rect 10820 22249 11156 22280
rect 10780 22240 11156 22249
rect 10924 22112 10964 22121
rect 10636 22072 10924 22112
rect 10924 22063 10964 22072
rect 10540 21904 11060 21944
rect 10731 21776 10773 21785
rect 10731 21736 10732 21776
rect 10772 21736 10773 21776
rect 10731 21727 10773 21736
rect 10443 21608 10485 21617
rect 10443 21568 10444 21608
rect 10484 21568 10485 21608
rect 10443 21559 10485 21568
rect 10444 20012 10484 20021
rect 10444 19853 10484 19972
rect 10540 20012 10580 20021
rect 10443 19844 10485 19853
rect 10443 19804 10444 19844
rect 10484 19804 10485 19844
rect 10443 19795 10485 19804
rect 10540 19685 10580 19972
rect 10539 19676 10581 19685
rect 10539 19636 10540 19676
rect 10580 19636 10581 19676
rect 10539 19627 10581 19636
rect 10732 19256 10772 21727
rect 10923 21608 10965 21617
rect 10923 21568 10924 21608
rect 10964 21568 10965 21608
rect 10923 21559 10965 21568
rect 10636 19216 10732 19256
rect 10443 19172 10485 19181
rect 10443 19132 10444 19172
rect 10484 19132 10485 19172
rect 10443 19123 10485 19132
rect 10444 18845 10484 19123
rect 10443 18836 10485 18845
rect 10443 18796 10444 18836
rect 10484 18796 10485 18836
rect 10443 18787 10485 18796
rect 10444 15569 10484 18787
rect 10636 15989 10676 19216
rect 10732 19207 10772 19216
rect 10924 20768 10964 21559
rect 10924 18593 10964 20728
rect 11020 20096 11060 21904
rect 11116 21776 11156 22240
rect 11212 22231 11252 22240
rect 11308 22280 11348 22289
rect 11308 22037 11348 22240
rect 11307 22028 11349 22037
rect 11307 21988 11308 22028
rect 11348 21988 11349 22028
rect 11307 21979 11349 21988
rect 11116 21727 11156 21736
rect 11404 20777 11444 22567
rect 11308 20768 11348 20777
rect 11403 20768 11445 20777
rect 11348 20728 11404 20768
rect 11444 20728 11445 20768
rect 11308 20719 11348 20728
rect 11403 20719 11445 20728
rect 11404 20634 11444 20719
rect 11116 20600 11156 20609
rect 11116 20105 11156 20560
rect 11500 20525 11540 24592
rect 11596 23717 11636 25339
rect 11595 23708 11637 23717
rect 11595 23668 11596 23708
rect 11636 23668 11637 23708
rect 11595 23659 11637 23668
rect 11596 22037 11636 23659
rect 11692 22541 11732 27859
rect 11884 27824 11924 28288
rect 11980 28169 12020 28447
rect 12076 28337 12116 29128
rect 12172 28841 12212 29800
rect 12460 29840 12500 30379
rect 12555 30260 12597 30269
rect 12555 30220 12556 30260
rect 12596 30220 12597 30260
rect 12555 30211 12597 30220
rect 12460 29791 12500 29800
rect 12363 29504 12405 29513
rect 12363 29464 12364 29504
rect 12404 29464 12405 29504
rect 12363 29455 12405 29464
rect 12364 29168 12404 29455
rect 12459 29252 12501 29261
rect 12459 29212 12460 29252
rect 12500 29212 12501 29252
rect 12459 29203 12501 29212
rect 12364 29119 12404 29128
rect 12460 29118 12500 29203
rect 12267 29084 12309 29093
rect 12267 29044 12268 29084
rect 12308 29044 12309 29084
rect 12267 29035 12309 29044
rect 12171 28832 12213 28841
rect 12171 28792 12172 28832
rect 12212 28792 12213 28832
rect 12171 28783 12213 28792
rect 12268 28337 12308 29035
rect 12556 29000 12596 30211
rect 12747 29924 12789 29933
rect 12747 29884 12748 29924
rect 12788 29884 12789 29924
rect 12747 29875 12789 29884
rect 12748 29790 12788 29875
rect 12844 29840 12884 32320
rect 12940 32192 12980 32203
rect 13036 32192 13076 32479
rect 13131 32444 13173 32453
rect 13131 32404 13132 32444
rect 13172 32404 13173 32444
rect 13131 32395 13173 32404
rect 13132 32360 13172 32395
rect 13132 32309 13172 32320
rect 13036 32152 13172 32192
rect 12940 32117 12980 32152
rect 12939 32108 12981 32117
rect 12939 32068 12940 32108
rect 12980 32068 12981 32108
rect 12939 32059 12981 32068
rect 12940 31940 12980 31949
rect 12940 30605 12980 31900
rect 13035 31520 13077 31529
rect 13035 31480 13036 31520
rect 13076 31480 13077 31520
rect 13035 31471 13077 31480
rect 12939 30596 12981 30605
rect 12939 30556 12940 30596
rect 12980 30556 12981 30596
rect 12939 30547 12981 30556
rect 12940 30092 12980 30101
rect 13036 30092 13076 31471
rect 13132 31436 13172 32152
rect 13228 32117 13268 32824
rect 13324 32815 13364 32824
rect 13324 32201 13364 32286
rect 13323 32192 13365 32201
rect 13323 32152 13324 32192
rect 13364 32152 13365 32192
rect 13323 32143 13365 32152
rect 13227 32108 13269 32117
rect 13227 32068 13228 32108
rect 13268 32068 13269 32108
rect 13227 32059 13269 32068
rect 13324 32024 13364 32033
rect 13420 32024 13460 33823
rect 13364 31984 13460 32024
rect 13324 31975 13364 31984
rect 13516 31520 13556 34000
rect 13611 33704 13653 33713
rect 13611 33664 13612 33704
rect 13652 33664 13653 33704
rect 13611 33655 13653 33664
rect 13612 33570 13652 33655
rect 13804 33452 13844 33461
rect 13708 33412 13804 33452
rect 13708 32873 13748 33412
rect 13804 33403 13844 33412
rect 13803 33116 13845 33125
rect 13803 33076 13804 33116
rect 13844 33076 13845 33116
rect 13803 33067 13845 33076
rect 13707 32864 13749 32873
rect 13707 32824 13708 32864
rect 13748 32824 13749 32864
rect 13707 32815 13749 32824
rect 13804 32864 13844 33067
rect 13804 32815 13844 32824
rect 13708 32730 13748 32815
rect 13708 32192 13748 32201
rect 13612 32152 13708 32192
rect 13612 31613 13652 32152
rect 13708 32143 13748 32152
rect 13707 32024 13749 32033
rect 13707 31984 13708 32024
rect 13748 31984 13749 32024
rect 13707 31975 13749 31984
rect 13611 31604 13653 31613
rect 13611 31564 13612 31604
rect 13652 31564 13653 31604
rect 13611 31555 13653 31564
rect 13132 31387 13172 31396
rect 13420 31480 13556 31520
rect 13228 31352 13268 31363
rect 13228 31277 13268 31312
rect 13227 31268 13269 31277
rect 13227 31228 13228 31268
rect 13268 31228 13269 31268
rect 13227 31219 13269 31228
rect 13228 30941 13268 31219
rect 13227 30932 13269 30941
rect 13227 30892 13228 30932
rect 13268 30892 13269 30932
rect 13227 30883 13269 30892
rect 13420 30521 13460 31480
rect 13515 31352 13557 31361
rect 13515 31312 13516 31352
rect 13556 31312 13557 31352
rect 13515 31303 13557 31312
rect 13419 30512 13461 30521
rect 13419 30472 13420 30512
rect 13460 30472 13461 30512
rect 13419 30463 13461 30472
rect 12980 30052 13076 30092
rect 12940 30043 12980 30052
rect 13132 29840 13172 29849
rect 12844 29800 13132 29840
rect 13172 29800 13460 29840
rect 13132 29791 13172 29800
rect 13131 29672 13173 29681
rect 13131 29632 13132 29672
rect 13172 29632 13173 29672
rect 13131 29623 13173 29632
rect 12364 28960 12596 29000
rect 12940 29168 12980 29177
rect 12075 28328 12117 28337
rect 12075 28288 12076 28328
rect 12116 28288 12117 28328
rect 12075 28279 12117 28288
rect 12267 28328 12309 28337
rect 12267 28288 12268 28328
rect 12308 28288 12309 28328
rect 12267 28279 12309 28288
rect 12364 28328 12404 28960
rect 12748 28916 12788 28925
rect 12652 28876 12748 28916
rect 12364 28279 12404 28288
rect 12555 28328 12597 28337
rect 12555 28288 12556 28328
rect 12596 28288 12597 28328
rect 12555 28279 12597 28288
rect 11979 28160 12021 28169
rect 11979 28120 11980 28160
rect 12020 28120 12021 28160
rect 11979 28111 12021 28120
rect 11884 27775 11924 27784
rect 11979 27824 12021 27833
rect 11979 27784 11980 27824
rect 12020 27784 12021 27824
rect 11979 27775 12021 27784
rect 11787 27740 11829 27749
rect 11787 27700 11788 27740
rect 11828 27700 11829 27740
rect 11787 27691 11829 27700
rect 11788 27656 11828 27691
rect 11788 27605 11828 27616
rect 11980 27656 12020 27775
rect 11787 27404 11829 27413
rect 11787 27364 11788 27404
rect 11828 27364 11829 27404
rect 11787 27355 11829 27364
rect 11788 26732 11828 27355
rect 11883 27236 11925 27245
rect 11883 27196 11884 27236
rect 11924 27196 11925 27236
rect 11883 27187 11925 27196
rect 11788 26683 11828 26692
rect 11787 26564 11829 26573
rect 11787 26524 11788 26564
rect 11828 26524 11829 26564
rect 11787 26515 11829 26524
rect 11788 24725 11828 26515
rect 11787 24716 11829 24725
rect 11787 24676 11788 24716
rect 11828 24676 11829 24716
rect 11787 24667 11829 24676
rect 11788 22709 11828 24667
rect 11787 22700 11829 22709
rect 11787 22660 11788 22700
rect 11828 22660 11829 22700
rect 11787 22651 11829 22660
rect 11691 22532 11733 22541
rect 11691 22492 11692 22532
rect 11732 22492 11733 22532
rect 11691 22483 11733 22492
rect 11884 22373 11924 27187
rect 11980 27077 12020 27616
rect 12076 27656 12116 28279
rect 12460 28244 12500 28253
rect 12363 28160 12405 28169
rect 12363 28120 12364 28160
rect 12404 28120 12405 28160
rect 12363 28111 12405 28120
rect 12267 28076 12309 28085
rect 12267 28036 12268 28076
rect 12308 28036 12309 28076
rect 12267 28027 12309 28036
rect 12076 27607 12116 27616
rect 12075 27320 12117 27329
rect 12075 27280 12076 27320
rect 12116 27280 12117 27320
rect 12075 27271 12117 27280
rect 11979 27068 12021 27077
rect 11979 27028 11980 27068
rect 12020 27028 12021 27068
rect 11979 27019 12021 27028
rect 11979 26816 12021 26825
rect 11979 26776 11980 26816
rect 12020 26776 12021 26816
rect 11979 26767 12021 26776
rect 11980 26682 12020 26767
rect 11979 25892 12021 25901
rect 11979 25852 11980 25892
rect 12020 25852 12021 25892
rect 11979 25843 12021 25852
rect 11980 25304 12020 25843
rect 12076 25649 12116 27271
rect 12075 25640 12117 25649
rect 12075 25600 12076 25640
rect 12116 25600 12117 25640
rect 12075 25591 12117 25600
rect 12268 25481 12308 28027
rect 12364 27488 12404 28111
rect 12460 27917 12500 28204
rect 12556 28169 12596 28279
rect 12555 28160 12597 28169
rect 12555 28120 12556 28160
rect 12596 28120 12597 28160
rect 12555 28111 12597 28120
rect 12459 27908 12501 27917
rect 12459 27868 12460 27908
rect 12500 27868 12501 27908
rect 12459 27859 12501 27868
rect 12459 27740 12501 27749
rect 12459 27700 12460 27740
rect 12500 27700 12501 27740
rect 12459 27691 12501 27700
rect 12460 27656 12500 27691
rect 12460 27605 12500 27616
rect 12556 27656 12596 27665
rect 12652 27656 12692 28876
rect 12748 28867 12788 28876
rect 12940 28757 12980 29128
rect 13036 29084 13076 29093
rect 12939 28748 12981 28757
rect 12939 28708 12940 28748
rect 12980 28708 12981 28748
rect 12939 28699 12981 28708
rect 12940 28580 12980 28589
rect 13036 28580 13076 29044
rect 13132 29000 13172 29623
rect 13324 29168 13364 29177
rect 13132 28951 13172 28960
rect 13228 29084 13268 29093
rect 13131 28664 13173 28673
rect 13131 28624 13132 28664
rect 13172 28624 13173 28664
rect 13131 28615 13173 28624
rect 12980 28540 13076 28580
rect 12940 28531 12980 28540
rect 12748 28496 12788 28505
rect 12788 28456 12884 28496
rect 12748 28447 12788 28456
rect 12844 28160 12884 28456
rect 12940 28337 12980 28422
rect 12939 28328 12981 28337
rect 12939 28288 12940 28328
rect 12980 28288 12981 28328
rect 12939 28279 12981 28288
rect 13132 28328 13172 28615
rect 13228 28505 13268 29044
rect 13227 28496 13269 28505
rect 13227 28456 13228 28496
rect 13268 28456 13269 28496
rect 13227 28447 13269 28456
rect 13132 28279 13172 28288
rect 13228 28328 13268 28337
rect 13228 28160 13268 28288
rect 12844 28120 13268 28160
rect 13324 28076 13364 29128
rect 13420 28841 13460 29800
rect 13419 28832 13461 28841
rect 13419 28792 13420 28832
rect 13460 28792 13461 28832
rect 13419 28783 13461 28792
rect 13419 28664 13461 28673
rect 13419 28624 13420 28664
rect 13460 28624 13461 28664
rect 13419 28615 13461 28624
rect 12748 28036 13364 28076
rect 13420 28328 13460 28615
rect 13516 28496 13556 31303
rect 13612 29000 13652 31555
rect 13708 31529 13748 31975
rect 13707 31520 13749 31529
rect 13707 31480 13708 31520
rect 13748 31480 13749 31520
rect 13707 31471 13749 31480
rect 13708 31352 13748 31363
rect 13708 31277 13748 31312
rect 13707 31268 13749 31277
rect 13707 31228 13708 31268
rect 13748 31228 13749 31268
rect 13707 31219 13749 31228
rect 13803 30764 13845 30773
rect 13803 30724 13804 30764
rect 13844 30724 13845 30764
rect 13803 30715 13845 30724
rect 13804 30680 13844 30715
rect 13900 30680 13940 36016
rect 13996 35888 14036 35897
rect 14188 35888 14228 37183
rect 14379 36896 14421 36905
rect 14379 36856 14380 36896
rect 14420 36856 14421 36896
rect 14379 36847 14421 36856
rect 14283 35972 14325 35981
rect 14283 35932 14284 35972
rect 14324 35932 14325 35972
rect 14283 35923 14325 35932
rect 14036 35848 14228 35888
rect 13996 34049 14036 35848
rect 14284 35729 14324 35923
rect 14283 35720 14325 35729
rect 14283 35680 14284 35720
rect 14324 35680 14325 35720
rect 14283 35671 14325 35680
rect 14187 34376 14229 34385
rect 14187 34336 14188 34376
rect 14228 34336 14229 34376
rect 14187 34327 14229 34336
rect 14284 34376 14324 34385
rect 14091 34292 14133 34301
rect 14091 34252 14092 34292
rect 14132 34252 14133 34292
rect 14091 34243 14133 34252
rect 13995 34040 14037 34049
rect 13995 34000 13996 34040
rect 14036 34000 14037 34040
rect 13995 33991 14037 34000
rect 13996 33704 14036 33713
rect 14092 33704 14132 34243
rect 14036 33664 14132 33704
rect 13996 33655 14036 33664
rect 14188 33545 14228 34327
rect 14284 33965 14324 34336
rect 14283 33956 14325 33965
rect 14283 33916 14284 33956
rect 14324 33916 14325 33956
rect 14283 33907 14325 33916
rect 14284 33713 14324 33907
rect 14283 33704 14325 33713
rect 14283 33664 14284 33704
rect 14324 33664 14325 33704
rect 14283 33655 14325 33664
rect 14187 33536 14229 33545
rect 14187 33496 14188 33536
rect 14228 33496 14229 33536
rect 14187 33487 14229 33496
rect 14187 33116 14229 33125
rect 14187 33076 14188 33116
rect 14228 33076 14229 33116
rect 14187 33067 14229 33076
rect 13995 32864 14037 32873
rect 13995 32824 13996 32864
rect 14036 32824 14037 32864
rect 13995 32815 14037 32824
rect 14188 32864 14228 33067
rect 14283 32948 14325 32957
rect 14283 32908 14284 32948
rect 14324 32908 14325 32948
rect 14283 32899 14325 32908
rect 13996 32201 14036 32815
rect 14188 32789 14228 32824
rect 14284 32814 14324 32899
rect 14187 32780 14229 32789
rect 14187 32740 14188 32780
rect 14228 32740 14229 32780
rect 14187 32731 14229 32740
rect 14380 32453 14420 36847
rect 14475 35636 14517 35645
rect 14475 35596 14476 35636
rect 14516 35596 14517 35636
rect 14475 35587 14517 35596
rect 14476 34637 14516 35587
rect 14571 35300 14613 35309
rect 14571 35260 14572 35300
rect 14612 35260 14613 35300
rect 14571 35251 14613 35260
rect 14475 34628 14517 34637
rect 14475 34588 14476 34628
rect 14516 34588 14517 34628
rect 14475 34579 14517 34588
rect 14572 34376 14612 35251
rect 14668 34628 14708 37351
rect 14764 37241 14804 37435
rect 14860 37400 14900 37409
rect 14763 37232 14805 37241
rect 14763 37192 14764 37232
rect 14804 37192 14805 37232
rect 14763 37183 14805 37192
rect 14860 35645 14900 37360
rect 14956 37400 14996 37409
rect 14859 35636 14901 35645
rect 14859 35596 14860 35636
rect 14900 35596 14901 35636
rect 14859 35587 14901 35596
rect 14956 35384 14996 37360
rect 15052 37400 15092 37409
rect 15052 37157 15092 37360
rect 15435 37400 15477 37409
rect 15435 37360 15436 37400
rect 15476 37360 15477 37400
rect 15435 37351 15477 37360
rect 15532 37400 15572 37603
rect 15723 37568 15765 37577
rect 15723 37528 15724 37568
rect 15764 37528 15765 37568
rect 15723 37519 15765 37528
rect 15532 37351 15572 37360
rect 15628 37484 15668 37493
rect 15148 37232 15188 37241
rect 15051 37148 15093 37157
rect 15051 37108 15052 37148
rect 15092 37108 15093 37148
rect 15051 37099 15093 37108
rect 15052 36569 15092 37099
rect 15051 36560 15093 36569
rect 15051 36520 15052 36560
rect 15092 36520 15093 36560
rect 15051 36511 15093 36520
rect 15148 35645 15188 37192
rect 15340 36728 15380 36737
rect 15244 36688 15340 36728
rect 15436 36728 15476 37351
rect 15628 37241 15668 37444
rect 15724 37434 15764 37519
rect 15820 37484 15860 37493
rect 15627 37232 15669 37241
rect 15627 37192 15628 37232
rect 15668 37192 15669 37232
rect 15627 37183 15669 37192
rect 15532 36896 15572 36905
rect 15820 36896 15860 37444
rect 15572 36856 15860 36896
rect 15532 36847 15572 36856
rect 15436 36688 15668 36728
rect 15244 36233 15284 36688
rect 15340 36679 15380 36688
rect 15435 36560 15477 36569
rect 15340 36520 15436 36560
rect 15476 36520 15477 36560
rect 15243 36224 15285 36233
rect 15243 36184 15244 36224
rect 15284 36184 15285 36224
rect 15243 36175 15285 36184
rect 15244 35888 15284 36175
rect 15340 35972 15380 36520
rect 15435 36511 15477 36520
rect 15436 36149 15476 36234
rect 15435 36140 15477 36149
rect 15435 36100 15436 36140
rect 15476 36100 15477 36140
rect 15435 36091 15477 36100
rect 15340 35932 15476 35972
rect 15147 35636 15189 35645
rect 15147 35596 15148 35636
rect 15188 35596 15189 35636
rect 15147 35587 15189 35596
rect 14668 34579 14708 34588
rect 14764 35344 14996 35384
rect 14668 34376 14708 34385
rect 14572 34336 14668 34376
rect 14668 34327 14708 34336
rect 14764 34208 14804 35344
rect 14956 35216 14996 35227
rect 14956 35141 14996 35176
rect 15244 35141 15284 35848
rect 15339 35636 15381 35645
rect 15339 35596 15340 35636
rect 15380 35596 15381 35636
rect 15339 35587 15381 35596
rect 15340 35216 15380 35587
rect 15340 35167 15380 35176
rect 14955 35132 14997 35141
rect 14955 35092 14956 35132
rect 14996 35092 14997 35132
rect 14955 35083 14997 35092
rect 15243 35132 15285 35141
rect 15243 35092 15244 35132
rect 15284 35092 15285 35132
rect 15243 35083 15285 35092
rect 14955 34964 14997 34973
rect 14955 34924 14956 34964
rect 14996 34924 14997 34964
rect 14955 34915 14997 34924
rect 15147 34964 15189 34973
rect 15147 34924 15148 34964
rect 15188 34924 15189 34964
rect 15147 34915 15189 34924
rect 15340 34964 15380 34973
rect 14956 34544 14996 34915
rect 15148 34830 15188 34915
rect 15051 34628 15093 34637
rect 15051 34588 15052 34628
rect 15092 34588 15093 34628
rect 15051 34579 15093 34588
rect 14955 34504 14996 34544
rect 14955 34460 14995 34504
rect 14955 34420 14996 34460
rect 14860 34376 14900 34385
rect 14860 34217 14900 34336
rect 14956 34376 14996 34420
rect 14956 34327 14996 34336
rect 14476 34168 14804 34208
rect 14859 34208 14901 34217
rect 14859 34168 14860 34208
rect 14900 34168 14901 34208
rect 14379 32444 14421 32453
rect 14379 32404 14380 32444
rect 14420 32404 14421 32444
rect 14379 32395 14421 32404
rect 14476 32360 14516 34168
rect 14859 34159 14901 34168
rect 15052 34040 15092 34579
rect 15148 34217 15188 34302
rect 15147 34208 15189 34217
rect 15147 34168 15148 34208
rect 15188 34168 15189 34208
rect 15147 34159 15189 34168
rect 15052 34000 15188 34040
rect 14763 33704 14805 33713
rect 14763 33664 14764 33704
rect 14804 33664 14805 33704
rect 14763 33655 14805 33664
rect 14667 33536 14709 33545
rect 14667 33496 14668 33536
rect 14708 33496 14709 33536
rect 14667 33487 14709 33496
rect 14668 32537 14708 33487
rect 14764 32864 14804 33655
rect 15148 33536 15188 34000
rect 15243 33956 15285 33965
rect 15243 33916 15244 33956
rect 15284 33916 15285 33956
rect 15243 33907 15285 33916
rect 15244 33704 15284 33907
rect 15244 33655 15284 33664
rect 15148 33496 15284 33536
rect 15147 33284 15189 33293
rect 15147 33244 15148 33284
rect 15188 33244 15189 33284
rect 15147 33235 15189 33244
rect 14667 32528 14709 32537
rect 14667 32488 14668 32528
rect 14708 32488 14709 32528
rect 14667 32479 14709 32488
rect 14476 32311 14516 32320
rect 14284 32236 14420 32276
rect 13995 32192 14037 32201
rect 13995 32152 13996 32192
rect 14036 32152 14037 32192
rect 13995 32143 14037 32152
rect 14284 32117 14324 32236
rect 14380 32192 14420 32236
rect 14380 32143 14420 32152
rect 14571 32192 14613 32201
rect 14571 32152 14572 32192
rect 14612 32152 14613 32192
rect 14571 32143 14613 32152
rect 14668 32192 14708 32479
rect 14764 32369 14804 32824
rect 14955 32696 14997 32705
rect 14955 32656 14956 32696
rect 14996 32656 14997 32696
rect 14955 32647 14997 32656
rect 14763 32360 14805 32369
rect 14763 32320 14764 32360
rect 14804 32320 14805 32360
rect 14763 32311 14805 32320
rect 14764 32201 14804 32311
rect 14668 32143 14708 32152
rect 14763 32192 14805 32201
rect 14763 32152 14764 32192
rect 14804 32152 14805 32192
rect 14763 32143 14805 32152
rect 14283 32108 14325 32117
rect 14283 32068 14284 32108
rect 14324 32068 14325 32108
rect 14283 32059 14325 32068
rect 14572 32058 14612 32143
rect 14956 32033 14996 32647
rect 15051 32192 15093 32201
rect 15051 32152 15052 32192
rect 15092 32152 15093 32192
rect 15051 32143 15093 32152
rect 15148 32192 15188 33235
rect 15244 32878 15284 33496
rect 15340 32957 15380 34924
rect 15436 34460 15476 35932
rect 15532 35216 15572 35225
rect 15532 34637 15572 35176
rect 15628 34973 15668 36688
rect 15820 36644 15860 36856
rect 15916 37400 15956 37409
rect 15916 36812 15956 37360
rect 16012 37232 16052 37939
rect 16108 37829 16148 38116
rect 16203 38116 16204 38156
rect 16244 38116 16245 38156
rect 16203 38107 16245 38116
rect 16204 38072 16244 38107
rect 16204 38021 16244 38032
rect 16107 37820 16149 37829
rect 16107 37780 16108 37820
rect 16148 37780 16149 37820
rect 16107 37771 16149 37780
rect 16107 37652 16149 37661
rect 16107 37612 16108 37652
rect 16148 37612 16149 37652
rect 16107 37603 16149 37612
rect 16108 37518 16148 37603
rect 16300 37577 16340 38284
rect 16396 38240 16436 38611
rect 16396 37997 16436 38200
rect 16395 37988 16437 37997
rect 16395 37948 16396 37988
rect 16436 37948 16437 37988
rect 16395 37939 16437 37948
rect 16299 37568 16341 37577
rect 16299 37528 16300 37568
rect 16340 37528 16341 37568
rect 16299 37519 16341 37528
rect 16108 37400 16148 37409
rect 16299 37400 16341 37409
rect 16148 37360 16244 37400
rect 16108 37351 16148 37360
rect 16012 37192 16148 37232
rect 15916 36763 15956 36772
rect 16011 36728 16053 36737
rect 15916 36705 15956 36714
rect 16011 36688 16012 36728
rect 16052 36688 16053 36728
rect 16011 36679 16053 36688
rect 15916 36644 15956 36665
rect 15820 36604 15956 36644
rect 16012 36594 16052 36679
rect 15723 36560 15765 36569
rect 15723 36520 15724 36560
rect 15764 36520 15765 36560
rect 15723 36511 15765 36520
rect 15724 36149 15764 36511
rect 16108 36476 16148 37192
rect 16204 36896 16244 37360
rect 16299 37360 16300 37400
rect 16340 37360 16341 37400
rect 16299 37351 16341 37360
rect 16396 37400 16436 37409
rect 16300 37266 16340 37351
rect 16396 36980 16436 37360
rect 16492 37232 16532 38872
rect 16588 38585 16628 38872
rect 16587 38576 16629 38585
rect 16587 38536 16588 38576
rect 16628 38536 16629 38576
rect 16587 38527 16629 38536
rect 16684 37442 16724 40375
rect 16684 37393 16724 37402
rect 16780 40256 16820 40265
rect 16780 37400 16820 40216
rect 16876 39089 16916 40384
rect 16972 40424 17012 40433
rect 16972 39929 17012 40384
rect 17068 40424 17108 40435
rect 17068 40349 17108 40384
rect 17067 40340 17109 40349
rect 17067 40300 17068 40340
rect 17108 40300 17109 40340
rect 17067 40291 17109 40300
rect 16971 39920 17013 39929
rect 16971 39880 16972 39920
rect 17012 39880 17013 39920
rect 16971 39871 17013 39880
rect 17068 39089 17108 40291
rect 16875 39080 16917 39089
rect 16875 39040 16876 39080
rect 16916 39040 16917 39080
rect 16875 39031 16917 39040
rect 17067 39080 17109 39089
rect 17067 39040 17068 39080
rect 17108 39040 17109 39080
rect 17067 39031 17109 39040
rect 16875 37484 16917 37493
rect 16875 37444 16876 37484
rect 16916 37444 16917 37484
rect 16875 37435 16917 37444
rect 16780 37351 16820 37360
rect 16876 37400 16916 37435
rect 16876 37349 16916 37360
rect 17068 37325 17108 39031
rect 17164 37652 17204 40552
rect 17355 40552 17356 40592
rect 17396 40552 17397 40592
rect 17355 40543 17397 40552
rect 17932 40508 17972 40517
rect 18028 40508 18068 41635
rect 18316 41357 18356 42928
rect 18508 42272 18548 42928
rect 18412 42232 18548 42272
rect 18315 41348 18357 41357
rect 18315 41308 18316 41348
rect 18356 41308 18357 41348
rect 18315 41299 18357 41308
rect 18124 41180 18164 41189
rect 18164 41140 18260 41180
rect 18124 41131 18164 41140
rect 18123 40592 18165 40601
rect 18123 40552 18124 40592
rect 18164 40552 18165 40592
rect 18123 40543 18165 40552
rect 17972 40468 18068 40508
rect 17932 40459 17972 40468
rect 18124 40458 18164 40543
rect 17259 40424 17301 40433
rect 17259 40384 17260 40424
rect 17300 40384 17301 40424
rect 17259 40375 17301 40384
rect 17452 40424 17492 40433
rect 17260 40290 17300 40375
rect 17355 40256 17397 40265
rect 17355 40216 17356 40256
rect 17396 40216 17397 40256
rect 17355 40207 17397 40216
rect 17356 40122 17396 40207
rect 17452 40004 17492 40384
rect 17356 39964 17492 40004
rect 17548 40424 17588 40433
rect 17356 39341 17396 39964
rect 17548 39920 17588 40384
rect 17740 40256 17780 40265
rect 17780 40216 17876 40256
rect 17740 40207 17780 40216
rect 17452 39880 17588 39920
rect 17355 39332 17397 39341
rect 17355 39292 17356 39332
rect 17396 39292 17397 39332
rect 17355 39283 17397 39292
rect 17356 37820 17396 39283
rect 17452 38081 17492 39880
rect 17739 39836 17781 39845
rect 17739 39796 17740 39836
rect 17780 39796 17781 39836
rect 17739 39787 17781 39796
rect 17548 39752 17588 39761
rect 17548 38828 17588 39712
rect 17740 39702 17780 39787
rect 17836 39080 17876 40216
rect 18123 39752 18165 39761
rect 18123 39712 18124 39752
rect 18164 39712 18165 39752
rect 18123 39703 18165 39712
rect 17931 39668 17973 39677
rect 17931 39628 17932 39668
rect 17972 39628 17973 39668
rect 17931 39619 17973 39628
rect 17932 39534 17972 39619
rect 18124 39584 18164 39703
rect 18124 39535 18164 39544
rect 18220 39080 18260 41140
rect 18315 41012 18357 41021
rect 18315 40972 18316 41012
rect 18356 40972 18357 41012
rect 18315 40963 18357 40972
rect 18316 40878 18356 40963
rect 18315 40508 18357 40517
rect 18315 40468 18316 40508
rect 18356 40468 18357 40508
rect 18315 40459 18357 40468
rect 18316 40374 18356 40459
rect 18412 40349 18452 42232
rect 18507 42104 18549 42113
rect 18507 42064 18508 42104
rect 18548 42064 18549 42104
rect 18507 42055 18549 42064
rect 18508 41180 18548 42055
rect 18700 41945 18740 42928
rect 18892 42701 18932 42928
rect 18891 42692 18933 42701
rect 18891 42652 18892 42692
rect 18932 42652 18933 42692
rect 18891 42643 18933 42652
rect 18699 41936 18741 41945
rect 18699 41896 18700 41936
rect 18740 41896 18741 41936
rect 18699 41887 18741 41896
rect 19084 41861 19124 42928
rect 19275 42904 19276 42928
rect 19316 42928 19336 42944
rect 19448 42928 19528 43008
rect 19316 42904 19317 42928
rect 19275 42895 19317 42904
rect 19275 42272 19317 42281
rect 19275 42232 19276 42272
rect 19316 42232 19317 42272
rect 19275 42223 19317 42232
rect 19083 41852 19125 41861
rect 19083 41812 19084 41852
rect 19124 41812 19125 41852
rect 19083 41803 19125 41812
rect 18508 41131 18548 41140
rect 18891 41180 18933 41189
rect 18891 41140 18892 41180
rect 18932 41140 18933 41180
rect 18891 41131 18933 41140
rect 19276 41180 19316 42223
rect 19468 41693 19508 42928
rect 19563 42524 19605 42533
rect 19563 42484 19564 42524
rect 19604 42484 19605 42524
rect 19563 42475 19605 42484
rect 19467 41684 19509 41693
rect 19467 41644 19468 41684
rect 19508 41644 19509 41684
rect 19467 41635 19509 41644
rect 19371 41600 19413 41609
rect 19371 41560 19372 41600
rect 19412 41560 19413 41600
rect 19371 41551 19413 41560
rect 19276 41131 19316 41140
rect 18892 41046 18932 41131
rect 19084 41021 19124 41106
rect 18700 41012 18740 41021
rect 18604 40972 18700 41012
rect 18507 40676 18549 40685
rect 18507 40636 18508 40676
rect 18548 40636 18549 40676
rect 18507 40627 18549 40636
rect 18508 40542 18548 40627
rect 18411 40340 18453 40349
rect 18411 40300 18412 40340
rect 18452 40300 18453 40340
rect 18411 40291 18453 40300
rect 18507 40088 18549 40097
rect 18507 40048 18508 40088
rect 18548 40048 18549 40088
rect 18507 40039 18549 40048
rect 18508 39668 18548 40039
rect 18508 39619 18548 39628
rect 18316 39500 18356 39509
rect 18316 39341 18356 39460
rect 18315 39332 18357 39341
rect 18315 39292 18316 39332
rect 18356 39292 18357 39332
rect 18315 39283 18357 39292
rect 17836 39040 17972 39080
rect 17836 38912 17876 38923
rect 17836 38837 17876 38872
rect 17643 38828 17685 38837
rect 17548 38788 17644 38828
rect 17684 38788 17685 38828
rect 17643 38779 17685 38788
rect 17835 38828 17877 38837
rect 17835 38788 17836 38828
rect 17876 38788 17877 38828
rect 17835 38779 17877 38788
rect 17644 38240 17684 38779
rect 17835 38660 17877 38669
rect 17835 38620 17836 38660
rect 17876 38620 17877 38660
rect 17835 38611 17877 38620
rect 17739 38576 17781 38585
rect 17739 38536 17740 38576
rect 17780 38536 17781 38576
rect 17739 38527 17781 38536
rect 17740 38249 17780 38527
rect 17836 38408 17876 38611
rect 17836 38359 17876 38368
rect 17548 38200 17644 38240
rect 17451 38072 17493 38081
rect 17451 38032 17452 38072
rect 17492 38032 17493 38072
rect 17451 38023 17493 38032
rect 17548 37820 17588 38200
rect 17644 38191 17684 38200
rect 17739 38240 17781 38249
rect 17739 38200 17740 38240
rect 17780 38200 17781 38240
rect 17739 38191 17781 38200
rect 17164 37603 17204 37612
rect 17260 37780 17396 37820
rect 17452 37780 17588 37820
rect 17260 37493 17300 37780
rect 17259 37484 17301 37493
rect 17259 37444 17260 37484
rect 17300 37444 17301 37484
rect 17259 37435 17301 37444
rect 17356 37484 17396 37493
rect 17067 37316 17109 37325
rect 17067 37276 17068 37316
rect 17108 37276 17109 37316
rect 17067 37267 17109 37276
rect 16588 37232 16628 37241
rect 16492 37192 16588 37232
rect 16588 37183 16628 37192
rect 16875 37232 16917 37241
rect 16875 37192 16876 37232
rect 16916 37192 16917 37232
rect 16875 37183 16917 37192
rect 17163 37232 17205 37241
rect 17163 37192 17164 37232
rect 17204 37192 17205 37232
rect 17163 37183 17205 37192
rect 16491 36980 16533 36989
rect 16396 36940 16492 36980
rect 16532 36940 16533 36980
rect 16491 36931 16533 36940
rect 16204 36856 16435 36896
rect 16395 36821 16435 36856
rect 16395 36812 16437 36821
rect 16395 36772 16396 36812
rect 16436 36772 16437 36812
rect 16395 36763 16437 36772
rect 16299 36728 16341 36737
rect 16204 36713 16244 36722
rect 16299 36688 16300 36728
rect 16340 36688 16341 36728
rect 16684 36728 16724 36737
rect 16299 36679 16341 36688
rect 16457 36713 16497 36722
rect 16204 36653 16244 36673
rect 16203 36644 16245 36653
rect 16203 36604 16204 36644
rect 16244 36604 16245 36644
rect 16203 36595 16245 36604
rect 16204 36578 16244 36595
rect 16300 36594 16340 36679
rect 16108 36436 16244 36476
rect 15915 36392 15957 36401
rect 15915 36352 15916 36392
rect 15956 36352 15957 36392
rect 15915 36343 15957 36352
rect 15723 36140 15765 36149
rect 15723 36100 15724 36140
rect 15764 36100 15765 36140
rect 15723 36091 15765 36100
rect 15724 35888 15764 36091
rect 15724 35839 15764 35848
rect 15724 35216 15764 35225
rect 15627 34964 15669 34973
rect 15627 34924 15628 34964
rect 15668 34924 15669 34964
rect 15627 34915 15669 34924
rect 15531 34628 15573 34637
rect 15531 34588 15532 34628
rect 15572 34588 15573 34628
rect 15531 34579 15573 34588
rect 15436 34420 15572 34460
rect 15436 34334 15476 34343
rect 15435 34294 15436 34301
rect 15476 34294 15477 34301
rect 15435 34292 15477 34294
rect 15435 34252 15436 34292
rect 15476 34252 15477 34292
rect 15435 34243 15477 34252
rect 15436 34199 15476 34243
rect 15436 33872 15476 33881
rect 15532 33872 15572 34420
rect 15476 33832 15572 33872
rect 15436 33823 15476 33832
rect 15627 33788 15669 33797
rect 15627 33748 15628 33788
rect 15668 33748 15669 33788
rect 15627 33739 15669 33748
rect 15628 33704 15668 33739
rect 15435 33536 15477 33545
rect 15435 33496 15436 33536
rect 15476 33496 15477 33536
rect 15435 33487 15477 33496
rect 15339 32948 15381 32957
rect 15339 32908 15340 32948
rect 15380 32908 15381 32948
rect 15339 32899 15381 32908
rect 15244 32789 15284 32838
rect 15243 32780 15285 32789
rect 15243 32740 15244 32780
rect 15284 32740 15285 32780
rect 15243 32731 15285 32740
rect 15436 32780 15476 33487
rect 15628 33377 15668 33664
rect 15627 33368 15669 33377
rect 15627 33328 15628 33368
rect 15668 33328 15669 33368
rect 15627 33319 15669 33328
rect 15724 33032 15764 35176
rect 15916 33461 15956 36343
rect 16011 36308 16053 36317
rect 16011 36268 16012 36308
rect 16052 36268 16053 36308
rect 16011 36259 16053 36268
rect 16012 35888 16052 36259
rect 16012 35309 16052 35848
rect 16107 35804 16149 35813
rect 16107 35764 16108 35804
rect 16148 35764 16149 35804
rect 16107 35755 16149 35764
rect 16108 35670 16148 35755
rect 16011 35300 16053 35309
rect 16011 35260 16012 35300
rect 16052 35260 16053 35300
rect 16011 35251 16053 35260
rect 16107 34628 16149 34637
rect 16107 34588 16108 34628
rect 16148 34588 16149 34628
rect 16107 34579 16149 34588
rect 15915 33452 15957 33461
rect 15915 33412 15916 33452
rect 15956 33412 15957 33452
rect 15915 33403 15957 33412
rect 15819 33284 15861 33293
rect 15819 33244 15820 33284
rect 15860 33244 15861 33284
rect 15819 33235 15861 33244
rect 15436 32731 15476 32740
rect 15532 32992 15764 33032
rect 15244 32714 15284 32731
rect 15532 32360 15572 32992
rect 15820 32948 15860 33235
rect 16108 33116 16148 34579
rect 16108 33067 16148 33076
rect 15724 32908 15860 32948
rect 15627 32864 15669 32873
rect 15627 32824 15628 32864
rect 15668 32824 15669 32864
rect 15627 32815 15669 32824
rect 15724 32864 15764 32908
rect 15916 32864 15956 32873
rect 16108 32864 16148 32873
rect 15724 32815 15764 32824
rect 15820 32843 15860 32852
rect 15628 32730 15668 32815
rect 15956 32824 16108 32864
rect 15916 32815 15956 32824
rect 16108 32815 16148 32824
rect 15820 32789 15860 32803
rect 15819 32780 15861 32789
rect 15819 32740 15820 32780
rect 15860 32740 15861 32780
rect 15819 32731 15861 32740
rect 15820 32708 15860 32731
rect 15819 32528 15861 32537
rect 15819 32488 15820 32528
rect 15860 32488 15861 32528
rect 15819 32479 15861 32488
rect 15532 32320 15668 32360
rect 13995 32024 14037 32033
rect 13995 31984 13996 32024
rect 14036 31984 14037 32024
rect 13995 31975 14037 31984
rect 14379 32024 14421 32033
rect 14379 31984 14380 32024
rect 14420 31984 14421 32024
rect 14379 31975 14421 31984
rect 14955 32024 14997 32033
rect 14955 31984 14956 32024
rect 14996 31984 14997 32024
rect 14955 31975 14997 31984
rect 13996 31890 14036 31975
rect 14188 31357 14228 31366
rect 13996 30848 14036 30857
rect 14188 30848 14228 31317
rect 14380 31268 14420 31975
rect 14667 31940 14709 31949
rect 14667 31900 14668 31940
rect 14708 31900 14709 31940
rect 14667 31891 14709 31900
rect 14475 31856 14517 31865
rect 14475 31816 14476 31856
rect 14516 31816 14517 31856
rect 14475 31807 14517 31816
rect 14380 31219 14420 31228
rect 14036 30808 14228 30848
rect 13996 30799 14036 30808
rect 14476 30689 14516 31807
rect 14187 30680 14229 30689
rect 13900 30640 14132 30680
rect 13804 29933 13844 30640
rect 13803 29924 13845 29933
rect 13803 29884 13804 29924
rect 13844 29884 13845 29924
rect 13803 29875 13845 29884
rect 13708 29177 13748 29262
rect 13707 29168 13749 29177
rect 13707 29128 13708 29168
rect 13748 29128 13749 29168
rect 13707 29119 13749 29128
rect 13612 28960 13844 29000
rect 13516 28456 13748 28496
rect 13516 28328 13556 28337
rect 13420 28288 13516 28328
rect 12748 27824 12788 28036
rect 12748 27775 12788 27784
rect 13035 27824 13077 27833
rect 13035 27784 13036 27824
rect 13076 27784 13077 27824
rect 13035 27775 13077 27784
rect 12596 27616 12692 27656
rect 12556 27607 12596 27616
rect 12940 27572 12980 27583
rect 12940 27497 12980 27532
rect 12939 27488 12981 27497
rect 12364 27448 12500 27488
rect 12364 26144 12404 26153
rect 12364 25901 12404 26104
rect 12363 25892 12405 25901
rect 12363 25852 12364 25892
rect 12404 25852 12405 25892
rect 12363 25843 12405 25852
rect 12267 25472 12309 25481
rect 12267 25432 12268 25472
rect 12308 25432 12309 25472
rect 12267 25423 12309 25432
rect 12363 25388 12405 25397
rect 12363 25348 12364 25388
rect 12404 25348 12405 25388
rect 12363 25339 12405 25348
rect 11980 25229 12020 25264
rect 12364 25254 12404 25339
rect 11979 25220 12021 25229
rect 11979 25180 11980 25220
rect 12020 25180 12021 25220
rect 11979 25171 12021 25180
rect 12172 25136 12212 25145
rect 12076 25096 12172 25136
rect 12076 24622 12116 25096
rect 12172 25087 12212 25096
rect 12363 25136 12405 25145
rect 12363 25096 12364 25136
rect 12404 25096 12405 25136
rect 12363 25087 12405 25096
rect 12364 24968 12404 25087
rect 12172 24928 12404 24968
rect 12172 24800 12212 24928
rect 12172 24751 12212 24760
rect 12028 24590 12116 24622
rect 12068 24582 12116 24590
rect 12460 24632 12500 27448
rect 12939 27448 12940 27488
rect 12980 27448 12981 27488
rect 12939 27439 12981 27448
rect 12651 27152 12693 27161
rect 12651 27112 12652 27152
rect 12692 27112 12693 27152
rect 12651 27103 12693 27112
rect 12555 26228 12597 26237
rect 12555 26188 12556 26228
rect 12596 26188 12597 26228
rect 12555 26179 12597 26188
rect 12556 26094 12596 26179
rect 12555 25556 12597 25565
rect 12555 25516 12556 25556
rect 12596 25516 12597 25556
rect 12555 25507 12597 25516
rect 12556 25422 12596 25507
rect 12555 25220 12597 25229
rect 12555 25180 12556 25220
rect 12596 25180 12597 25220
rect 12555 25171 12597 25180
rect 12460 24583 12500 24592
rect 12028 24541 12068 24550
rect 12363 24548 12405 24557
rect 12363 24508 12364 24548
rect 12404 24508 12405 24548
rect 12363 24499 12405 24508
rect 12364 24414 12404 24499
rect 12556 23885 12596 25171
rect 12555 23876 12597 23885
rect 12555 23836 12556 23876
rect 12596 23836 12597 23876
rect 12555 23827 12597 23836
rect 12556 23792 12596 23827
rect 12652 23801 12692 27103
rect 12939 27068 12981 27077
rect 12939 27028 12940 27068
rect 12980 27028 12981 27068
rect 12939 27019 12981 27028
rect 12747 26816 12789 26825
rect 12747 26776 12748 26816
rect 12788 26776 12789 26816
rect 12747 26767 12789 26776
rect 12748 25817 12788 26767
rect 12843 26228 12885 26237
rect 12843 26188 12844 26228
rect 12884 26188 12885 26228
rect 12843 26179 12885 26188
rect 12844 26144 12884 26179
rect 12844 26093 12884 26104
rect 12940 26144 12980 27019
rect 13036 26480 13076 27775
rect 13420 27740 13460 28288
rect 13516 28279 13556 28288
rect 13324 27700 13460 27740
rect 13131 27656 13173 27665
rect 13131 27616 13132 27656
rect 13172 27616 13173 27656
rect 13131 27607 13173 27616
rect 13132 27488 13172 27607
rect 13132 27439 13172 27448
rect 13324 26825 13364 27700
rect 13516 27656 13556 27665
rect 13420 27637 13460 27646
rect 13420 27068 13460 27597
rect 13420 27019 13460 27028
rect 13228 26816 13268 26825
rect 13228 26573 13268 26776
rect 13323 26816 13365 26825
rect 13323 26776 13324 26816
rect 13364 26776 13365 26816
rect 13323 26767 13365 26776
rect 13227 26564 13269 26573
rect 13227 26524 13228 26564
rect 13268 26524 13269 26564
rect 13227 26515 13269 26524
rect 13036 26440 13172 26480
rect 13132 26144 13172 26440
rect 13324 26144 13364 26153
rect 13132 26104 13324 26144
rect 12747 25808 12789 25817
rect 12747 25768 12748 25808
rect 12788 25768 12789 25808
rect 12747 25759 12789 25768
rect 12940 25397 12980 26104
rect 13324 26095 13364 26104
rect 13420 26144 13460 26153
rect 12939 25388 12981 25397
rect 12939 25348 12940 25388
rect 12980 25348 12981 25388
rect 12939 25339 12981 25348
rect 12747 25304 12789 25313
rect 12747 25264 12748 25304
rect 12788 25264 12789 25304
rect 12747 25255 12789 25264
rect 12748 24800 12788 25255
rect 13420 25061 13460 26104
rect 13419 25052 13461 25061
rect 13419 25012 13420 25052
rect 13460 25012 13461 25052
rect 13419 25003 13461 25012
rect 12748 24760 13076 24800
rect 12748 24632 12788 24641
rect 12748 24044 12788 24592
rect 12844 24632 12884 24641
rect 12884 24592 12980 24632
rect 12844 24583 12884 24592
rect 12748 23995 12788 24004
rect 12075 23204 12117 23213
rect 12075 23164 12076 23204
rect 12116 23164 12117 23204
rect 12075 23155 12117 23164
rect 11883 22364 11925 22373
rect 11883 22324 11884 22364
rect 11924 22324 11925 22364
rect 11883 22315 11925 22324
rect 11692 22280 11732 22289
rect 11692 22121 11732 22240
rect 11788 22280 11828 22291
rect 11788 22205 11828 22240
rect 11787 22196 11829 22205
rect 11787 22156 11788 22196
rect 11828 22156 11829 22196
rect 11787 22147 11829 22156
rect 11691 22112 11733 22121
rect 11691 22072 11692 22112
rect 11732 22072 11733 22112
rect 11691 22063 11733 22072
rect 11595 22028 11637 22037
rect 11595 21988 11596 22028
rect 11636 21988 11637 22028
rect 11595 21979 11637 21988
rect 11692 21449 11732 22063
rect 11884 21785 11924 22315
rect 11883 21776 11925 21785
rect 11883 21736 11884 21776
rect 11924 21736 11925 21776
rect 11883 21727 11925 21736
rect 11691 21440 11733 21449
rect 11691 21400 11692 21440
rect 11732 21400 11733 21440
rect 11691 21391 11733 21400
rect 12076 20609 12116 23155
rect 12556 23120 12596 23752
rect 12651 23792 12693 23801
rect 12651 23752 12652 23792
rect 12692 23752 12693 23792
rect 12651 23743 12693 23752
rect 12652 23120 12692 23129
rect 12556 23080 12652 23120
rect 12652 23071 12692 23080
rect 12844 22868 12884 22877
rect 12651 22784 12693 22793
rect 12651 22744 12652 22784
rect 12692 22744 12693 22784
rect 12651 22735 12693 22744
rect 12267 22364 12309 22373
rect 12267 22324 12268 22364
rect 12308 22324 12309 22364
rect 12267 22315 12309 22324
rect 12268 22280 12308 22315
rect 12268 22229 12308 22240
rect 12267 21608 12309 21617
rect 12267 21568 12268 21608
rect 12308 21568 12309 21608
rect 12267 21559 12309 21568
rect 12268 21474 12308 21559
rect 12652 21365 12692 22735
rect 12844 22448 12884 22828
rect 12748 22408 12884 22448
rect 12748 22294 12788 22408
rect 12940 22373 12980 24592
rect 13036 23969 13076 24760
rect 13227 24548 13269 24557
rect 13227 24508 13228 24548
rect 13268 24508 13269 24548
rect 13227 24499 13269 24508
rect 13324 24548 13364 24557
rect 13516 24548 13556 27616
rect 13611 27488 13653 27497
rect 13611 27448 13612 27488
rect 13652 27448 13653 27488
rect 13611 27439 13653 27448
rect 13612 26816 13652 27439
rect 13612 26767 13652 26776
rect 13611 26564 13653 26573
rect 13611 26524 13612 26564
rect 13652 26524 13653 26564
rect 13611 26515 13653 26524
rect 13364 24508 13556 24548
rect 13228 24305 13268 24499
rect 13227 24296 13269 24305
rect 13227 24256 13228 24296
rect 13268 24256 13269 24296
rect 13227 24247 13269 24256
rect 13227 24044 13269 24053
rect 13227 24004 13228 24044
rect 13268 24004 13269 24044
rect 13227 23995 13269 24004
rect 13035 23960 13077 23969
rect 13035 23920 13036 23960
rect 13076 23920 13077 23960
rect 13035 23911 13077 23920
rect 13036 23876 13076 23911
rect 13228 23910 13268 23995
rect 13036 23825 13076 23836
rect 13324 23708 13364 24508
rect 13612 24305 13652 26515
rect 13611 24296 13653 24305
rect 13611 24256 13612 24296
rect 13652 24256 13653 24296
rect 13611 24247 13653 24256
rect 13612 24044 13652 24053
rect 13708 24044 13748 28456
rect 13804 25061 13844 28960
rect 13900 27572 13940 27581
rect 13900 26909 13940 27532
rect 13996 27572 14036 27581
rect 13899 26900 13941 26909
rect 13899 26860 13900 26900
rect 13940 26860 13941 26900
rect 13899 26851 13941 26860
rect 13996 26657 14036 27532
rect 13995 26648 14037 26657
rect 13995 26608 13996 26648
rect 14036 26608 14037 26648
rect 13995 26599 14037 26608
rect 13899 26480 13941 26489
rect 13899 26440 13900 26480
rect 13940 26440 13941 26480
rect 13899 26431 13941 26440
rect 13900 26144 13940 26431
rect 13995 26228 14037 26237
rect 13995 26188 13996 26228
rect 14036 26188 14037 26228
rect 13995 26179 14037 26188
rect 13900 25733 13940 26104
rect 13899 25724 13941 25733
rect 13899 25684 13900 25724
rect 13940 25684 13941 25724
rect 13899 25675 13941 25684
rect 13899 25472 13941 25481
rect 13899 25432 13900 25472
rect 13940 25432 13941 25472
rect 13899 25423 13941 25432
rect 13803 25052 13845 25061
rect 13803 25012 13804 25052
rect 13844 25012 13845 25052
rect 13803 25003 13845 25012
rect 13652 24004 13748 24044
rect 13804 24632 13844 24641
rect 13804 24044 13844 24592
rect 13900 24473 13940 25423
rect 13996 25304 14036 26179
rect 13996 25229 14036 25264
rect 13995 25220 14037 25229
rect 13995 25180 13996 25220
rect 14036 25180 14037 25220
rect 13995 25171 14037 25180
rect 13899 24464 13941 24473
rect 13899 24424 13900 24464
rect 13940 24424 13941 24464
rect 13899 24415 13941 24424
rect 13995 24044 14037 24053
rect 13804 24004 13940 24044
rect 13612 23995 13652 24004
rect 13420 23876 13460 23885
rect 13420 23792 13460 23836
rect 13803 23876 13845 23885
rect 13803 23836 13804 23876
rect 13844 23836 13845 23876
rect 13803 23827 13845 23836
rect 13420 23752 13652 23792
rect 13324 23668 13460 23708
rect 13323 23288 13365 23297
rect 13323 23248 13324 23288
rect 13364 23248 13365 23288
rect 13323 23239 13365 23248
rect 13324 23154 13364 23239
rect 13131 23036 13173 23045
rect 13131 22996 13132 23036
rect 13172 22996 13173 23036
rect 13131 22987 13173 22996
rect 13132 22902 13172 22987
rect 13227 22700 13269 22709
rect 13227 22660 13228 22700
rect 13268 22660 13269 22700
rect 13227 22651 13269 22660
rect 12939 22364 12981 22373
rect 12939 22324 12940 22364
rect 12980 22324 12981 22364
rect 12939 22315 12981 22324
rect 13131 22364 13173 22373
rect 13131 22324 13132 22364
rect 13172 22324 13173 22364
rect 13131 22315 13173 22324
rect 12748 22245 12788 22254
rect 12939 22112 12981 22121
rect 12939 22072 12940 22112
rect 12980 22072 12981 22112
rect 12939 22063 12981 22072
rect 12940 21978 12980 22063
rect 12843 21860 12885 21869
rect 12843 21820 12844 21860
rect 12884 21820 12885 21860
rect 12843 21811 12885 21820
rect 12651 21356 12693 21365
rect 12651 21316 12652 21356
rect 12692 21316 12693 21356
rect 12651 21307 12693 21316
rect 12652 20861 12692 21307
rect 12651 20852 12693 20861
rect 12651 20812 12652 20852
rect 12692 20812 12693 20852
rect 12651 20803 12693 20812
rect 12556 20768 12596 20777
rect 12556 20609 12596 20728
rect 12747 20684 12789 20693
rect 12747 20644 12748 20684
rect 12788 20644 12789 20684
rect 12747 20635 12789 20644
rect 11691 20600 11733 20609
rect 11691 20560 11692 20600
rect 11732 20560 11733 20600
rect 11691 20551 11733 20560
rect 12075 20600 12117 20609
rect 12075 20560 12076 20600
rect 12116 20560 12117 20600
rect 12075 20551 12117 20560
rect 12555 20600 12597 20609
rect 12555 20560 12556 20600
rect 12596 20560 12597 20600
rect 12555 20551 12597 20560
rect 11499 20516 11541 20525
rect 11499 20476 11500 20516
rect 11540 20476 11541 20516
rect 11499 20467 11541 20476
rect 11692 20180 11732 20551
rect 12748 20550 12788 20635
rect 12652 20273 12692 20358
rect 12651 20264 12693 20273
rect 12651 20224 12652 20264
rect 12692 20224 12693 20264
rect 12651 20215 12693 20224
rect 11692 20131 11732 20140
rect 11020 20047 11060 20056
rect 11115 20096 11157 20105
rect 11115 20056 11116 20096
rect 11156 20056 11157 20096
rect 11115 20047 11157 20056
rect 11499 20096 11541 20105
rect 11499 20051 11500 20096
rect 11540 20051 11541 20096
rect 11499 20047 11541 20051
rect 11979 20096 12021 20105
rect 11979 20056 11980 20096
rect 12020 20056 12021 20096
rect 11979 20047 12021 20056
rect 12172 20096 12212 20105
rect 11500 19961 11540 20047
rect 11211 19844 11253 19853
rect 11211 19804 11212 19844
rect 11252 19804 11253 19844
rect 11211 19795 11253 19804
rect 11691 19844 11733 19853
rect 11691 19804 11692 19844
rect 11732 19804 11733 19844
rect 11691 19795 11733 19804
rect 11212 19517 11252 19795
rect 11499 19760 11541 19769
rect 11499 19720 11500 19760
rect 11540 19720 11541 19760
rect 11499 19711 11541 19720
rect 11211 19508 11253 19517
rect 11211 19468 11212 19508
rect 11252 19468 11253 19508
rect 11211 19459 11253 19468
rect 11212 19261 11252 19270
rect 11116 18752 11156 18761
rect 11212 18752 11252 19221
rect 11404 19172 11444 19181
rect 11500 19172 11540 19711
rect 11692 19601 11732 19795
rect 11691 19592 11733 19601
rect 11691 19552 11692 19592
rect 11732 19552 11733 19592
rect 11691 19543 11733 19552
rect 11595 19340 11637 19349
rect 11595 19300 11596 19340
rect 11636 19300 11637 19340
rect 11595 19291 11637 19300
rect 11596 19256 11636 19291
rect 11596 19205 11636 19216
rect 11444 19132 11540 19172
rect 11404 19123 11444 19132
rect 11156 18712 11252 18752
rect 11116 18703 11156 18712
rect 10923 18584 10965 18593
rect 11308 18584 11348 18593
rect 10923 18544 10924 18584
rect 10964 18544 11156 18584
rect 10923 18535 10965 18544
rect 10924 18450 10964 18535
rect 10828 17753 10868 17838
rect 10923 17828 10965 17837
rect 10923 17788 10924 17828
rect 10964 17788 10965 17828
rect 10923 17779 10965 17788
rect 10827 17744 10869 17753
rect 10732 17704 10828 17744
rect 10868 17704 10869 17744
rect 10732 17165 10772 17704
rect 10827 17695 10869 17704
rect 10827 17576 10869 17585
rect 10827 17536 10828 17576
rect 10868 17536 10869 17576
rect 10827 17527 10869 17536
rect 10731 17156 10773 17165
rect 10731 17116 10732 17156
rect 10772 17116 10773 17156
rect 10731 17107 10773 17116
rect 10828 16484 10868 17527
rect 10924 17240 10964 17779
rect 11019 17576 11061 17585
rect 11019 17536 11020 17576
rect 11060 17536 11061 17576
rect 11019 17527 11061 17536
rect 11020 17442 11060 17527
rect 10924 17200 11060 17240
rect 10923 17072 10965 17081
rect 10923 17032 10924 17072
rect 10964 17032 10965 17072
rect 10923 17023 10965 17032
rect 11020 17072 11060 17200
rect 10732 16444 10868 16484
rect 10732 16246 10772 16444
rect 10635 15980 10677 15989
rect 10635 15940 10636 15980
rect 10676 15940 10677 15980
rect 10635 15931 10677 15940
rect 10443 15560 10485 15569
rect 10443 15520 10444 15560
rect 10484 15520 10485 15560
rect 10443 15511 10485 15520
rect 10347 15140 10389 15149
rect 10347 15100 10348 15140
rect 10388 15100 10389 15140
rect 10347 15091 10389 15100
rect 10539 15140 10581 15149
rect 10539 15100 10540 15140
rect 10580 15100 10581 15140
rect 10539 15091 10581 15100
rect 10347 14888 10389 14897
rect 10347 14848 10348 14888
rect 10388 14848 10389 14888
rect 10347 14839 10389 14848
rect 10156 14720 10196 14729
rect 10156 14225 10196 14680
rect 10348 14720 10388 14839
rect 10348 14671 10388 14680
rect 10444 14720 10484 14731
rect 10444 14645 10484 14680
rect 10443 14636 10485 14645
rect 10443 14596 10444 14636
rect 10484 14596 10485 14636
rect 10443 14587 10485 14596
rect 10252 14552 10292 14561
rect 10155 14216 10197 14225
rect 10155 14176 10156 14216
rect 10196 14176 10197 14216
rect 10155 14167 10197 14176
rect 10060 14008 10196 14048
rect 10059 13880 10101 13889
rect 10059 13840 10060 13880
rect 10100 13840 10101 13880
rect 10059 13831 10101 13840
rect 9964 13411 10004 13420
rect 9964 13040 10004 13049
rect 9964 12545 10004 13000
rect 9963 12536 10005 12545
rect 9963 12496 9964 12536
rect 10004 12496 10005 12536
rect 9963 12487 10005 12496
rect 9964 12368 10004 12377
rect 9868 12328 9964 12368
rect 9964 12319 10004 12328
rect 9675 12284 9717 12293
rect 9675 12244 9676 12284
rect 9716 12244 9717 12284
rect 9675 12235 9717 12244
rect 9579 12116 9621 12125
rect 9579 12076 9580 12116
rect 9620 12076 9621 12116
rect 9579 12067 9621 12076
rect 9676 12041 9716 12235
rect 9675 12032 9717 12041
rect 9675 11992 9676 12032
rect 9716 11992 9717 12032
rect 9675 11983 9717 11992
rect 9580 11864 9620 11873
rect 9292 11824 9524 11864
rect 9003 11612 9045 11621
rect 9003 11572 9004 11612
rect 9044 11572 9045 11612
rect 9003 11563 9045 11572
rect 9195 11612 9237 11621
rect 9195 11572 9196 11612
rect 9236 11572 9237 11612
rect 9195 11563 9237 11572
rect 9292 11276 9332 11824
rect 9484 11780 9524 11824
rect 9484 11731 9524 11740
rect 9196 11236 9332 11276
rect 9388 11696 9428 11705
rect 9099 11108 9141 11117
rect 9099 11068 9100 11108
rect 9140 11068 9141 11108
rect 9099 11059 9141 11068
rect 8812 10781 8852 10984
rect 9100 11024 9140 11059
rect 9100 10973 9140 10984
rect 8811 10772 8853 10781
rect 8811 10732 8812 10772
rect 8852 10732 8853 10772
rect 8811 10723 8853 10732
rect 9099 10772 9141 10781
rect 9099 10732 9100 10772
rect 9140 10732 9141 10772
rect 9099 10723 9141 10732
rect 9100 10638 9140 10723
rect 9003 10436 9045 10445
rect 9003 10396 9004 10436
rect 9044 10396 9045 10436
rect 9003 10387 9045 10396
rect 9004 10193 9044 10387
rect 9196 10352 9236 11236
rect 9291 11108 9333 11117
rect 9291 11068 9292 11108
rect 9332 11068 9333 11108
rect 9291 11059 9333 11068
rect 9292 10974 9332 11059
rect 9100 10312 9236 10352
rect 9003 10184 9045 10193
rect 9003 10144 9004 10184
rect 9044 10144 9045 10184
rect 9003 10135 9045 10144
rect 8811 9428 8853 9437
rect 8811 9388 8812 9428
rect 8852 9388 8853 9428
rect 8811 9379 8853 9388
rect 8715 8672 8757 8681
rect 8715 8632 8716 8672
rect 8756 8632 8757 8672
rect 8715 8623 8757 8632
rect 8715 8252 8757 8261
rect 8715 8212 8716 8252
rect 8756 8212 8757 8252
rect 8715 8203 8757 8212
rect 8619 8084 8661 8093
rect 8619 8044 8620 8084
rect 8660 8044 8661 8084
rect 8619 8035 8661 8044
rect 8716 7757 8756 8203
rect 8715 7748 8757 7757
rect 8715 7708 8716 7748
rect 8756 7708 8757 7748
rect 8715 7699 8757 7708
rect 8715 7328 8757 7337
rect 8715 7288 8716 7328
rect 8756 7288 8757 7328
rect 8715 7279 8757 7288
rect 8523 7244 8565 7253
rect 8523 7204 8524 7244
rect 8564 7204 8565 7244
rect 8523 7195 8565 7204
rect 8716 7160 8756 7279
rect 8716 7111 8756 7120
rect 8620 7076 8660 7085
rect 8524 7036 8620 7076
rect 8427 6656 8469 6665
rect 8427 6616 8428 6656
rect 8468 6616 8469 6656
rect 8427 6607 8469 6616
rect 8331 6572 8373 6581
rect 8331 6532 8332 6572
rect 8372 6532 8373 6572
rect 8331 6523 8373 6532
rect 7852 3928 8084 3968
rect 8140 5272 8276 5312
rect 7852 3137 7892 3928
rect 7947 3800 7989 3809
rect 7947 3760 7948 3800
rect 7988 3760 7989 3800
rect 7947 3751 7989 3760
rect 7948 3221 7988 3751
rect 8043 3464 8085 3473
rect 8043 3424 8044 3464
rect 8084 3424 8085 3464
rect 8043 3415 8085 3424
rect 8044 3330 8084 3415
rect 7947 3212 7989 3221
rect 7947 3172 7948 3212
rect 7988 3172 7989 3212
rect 7947 3163 7989 3172
rect 7851 3128 7893 3137
rect 7851 3088 7852 3128
rect 7892 3088 7893 3128
rect 7851 3079 7893 3088
rect 7755 2792 7797 2801
rect 7755 2752 7756 2792
rect 7796 2752 7797 2792
rect 7755 2743 7797 2752
rect 7948 2624 7988 3163
rect 8140 2633 8180 5272
rect 8332 5228 8372 6523
rect 8427 6488 8469 6497
rect 8427 6448 8428 6488
rect 8468 6448 8469 6488
rect 8427 6439 8469 6448
rect 8428 6354 8468 6439
rect 8427 6068 8469 6077
rect 8427 6028 8428 6068
rect 8468 6028 8469 6068
rect 8427 6019 8469 6028
rect 8428 5741 8468 6019
rect 8427 5732 8469 5741
rect 8427 5692 8428 5732
rect 8468 5692 8469 5732
rect 8427 5683 8469 5692
rect 8428 5648 8468 5683
rect 8524 5657 8564 7036
rect 8620 7027 8660 7036
rect 8812 6992 8852 9379
rect 9004 8849 9044 10135
rect 9100 9941 9140 10312
rect 9388 10268 9428 11656
rect 9483 11612 9525 11621
rect 9483 11572 9484 11612
rect 9524 11572 9525 11612
rect 9483 11563 9525 11572
rect 9484 11024 9524 11563
rect 9484 10975 9524 10984
rect 9196 10228 9428 10268
rect 9099 9932 9141 9941
rect 9099 9892 9100 9932
rect 9140 9892 9141 9932
rect 9099 9883 9141 9892
rect 9196 9437 9236 10228
rect 9484 10184 9524 10193
rect 9292 10144 9484 10184
rect 9195 9428 9237 9437
rect 9195 9388 9196 9428
rect 9236 9388 9237 9428
rect 9195 9379 9237 9388
rect 9003 8840 9045 8849
rect 9003 8800 9004 8840
rect 9044 8800 9045 8840
rect 9003 8791 9045 8800
rect 9195 8756 9237 8765
rect 9195 8716 9196 8756
rect 9236 8716 9237 8756
rect 9195 8707 9237 8716
rect 9099 8672 9141 8681
rect 9099 8632 9100 8672
rect 9140 8632 9141 8672
rect 9099 8623 9141 8632
rect 9003 8168 9045 8177
rect 9003 8128 9004 8168
rect 9044 8128 9045 8168
rect 9003 8119 9045 8128
rect 8907 8084 8949 8093
rect 8907 8044 8908 8084
rect 8948 8044 8949 8084
rect 8907 8035 8949 8044
rect 8908 7925 8948 8035
rect 8907 7916 8949 7925
rect 8907 7876 8908 7916
rect 8948 7876 8949 7916
rect 8907 7867 8949 7876
rect 9004 7421 9044 8119
rect 9100 7748 9140 8623
rect 9196 7832 9236 8707
rect 9292 8597 9332 10144
rect 9484 10135 9524 10144
rect 9580 9680 9620 11824
rect 9676 11780 9716 11789
rect 9676 10436 9716 11740
rect 9771 11696 9813 11705
rect 9771 11656 9772 11696
rect 9812 11656 9813 11696
rect 9771 11647 9813 11656
rect 9964 11696 10004 11705
rect 9772 11453 9812 11647
rect 9964 11537 10004 11656
rect 9963 11528 10005 11537
rect 9963 11488 9964 11528
rect 10004 11488 10005 11528
rect 9963 11479 10005 11488
rect 9771 11444 9813 11453
rect 9771 11404 9772 11444
rect 9812 11404 9813 11444
rect 9771 11395 9813 11404
rect 9963 11276 10005 11285
rect 9963 11236 9964 11276
rect 10004 11236 10005 11276
rect 9963 11227 10005 11236
rect 9868 10436 9908 10445
rect 9676 10396 9868 10436
rect 9868 10387 9908 10396
rect 9964 10268 10004 11227
rect 9868 10228 10004 10268
rect 9484 9640 9620 9680
rect 9676 10016 9716 10025
rect 9291 8588 9333 8597
rect 9291 8548 9292 8588
rect 9332 8548 9333 8588
rect 9291 8539 9333 8548
rect 9292 8000 9332 8539
rect 9484 8261 9524 9640
rect 9579 9512 9621 9521
rect 9579 9472 9580 9512
rect 9620 9472 9621 9512
rect 9579 9463 9621 9472
rect 9676 9512 9716 9976
rect 9868 9605 9908 10228
rect 10060 10025 10100 13831
rect 10156 13553 10196 14008
rect 10155 13544 10197 13553
rect 10155 13504 10156 13544
rect 10196 13504 10197 13544
rect 10155 13495 10197 13504
rect 10156 12713 10196 13495
rect 10252 13208 10292 14512
rect 10347 14384 10389 14393
rect 10347 14344 10348 14384
rect 10388 14344 10389 14384
rect 10347 14335 10389 14344
rect 10348 14048 10388 14335
rect 10540 14057 10580 15091
rect 10636 14981 10676 15931
rect 10732 15555 10772 16206
rect 10924 16148 10964 17023
rect 11020 16568 11060 17032
rect 11116 16652 11156 18544
rect 11308 16829 11348 18544
rect 11404 18584 11444 18593
rect 11596 18584 11636 18593
rect 11787 18584 11829 18593
rect 11444 18544 11540 18584
rect 11404 18535 11444 18544
rect 11403 18416 11445 18425
rect 11403 18376 11404 18416
rect 11444 18376 11445 18416
rect 11403 18367 11445 18376
rect 11404 17744 11444 18367
rect 11404 17240 11444 17704
rect 11500 17669 11540 18544
rect 11636 18544 11732 18584
rect 11596 18535 11636 18544
rect 11596 18332 11636 18341
rect 11596 17837 11636 18292
rect 11692 18005 11732 18544
rect 11787 18544 11788 18584
rect 11828 18544 11829 18584
rect 11787 18535 11829 18544
rect 11788 18450 11828 18535
rect 11787 18164 11829 18173
rect 11787 18124 11788 18164
rect 11828 18124 11829 18164
rect 11787 18115 11829 18124
rect 11691 17996 11733 18005
rect 11691 17956 11692 17996
rect 11732 17956 11733 17996
rect 11691 17947 11733 17956
rect 11595 17828 11637 17837
rect 11595 17788 11596 17828
rect 11636 17788 11637 17828
rect 11595 17779 11637 17788
rect 11499 17660 11541 17669
rect 11499 17620 11500 17660
rect 11540 17620 11541 17660
rect 11499 17611 11541 17620
rect 11404 17200 11540 17240
rect 11404 17072 11444 17081
rect 11404 16913 11444 17032
rect 11403 16904 11445 16913
rect 11403 16864 11404 16904
rect 11444 16864 11445 16904
rect 11403 16855 11445 16864
rect 11307 16820 11349 16829
rect 11307 16780 11308 16820
rect 11348 16780 11349 16820
rect 11307 16771 11349 16780
rect 11116 16612 11348 16652
rect 11020 16528 11156 16568
rect 11019 16400 11061 16409
rect 11019 16360 11020 16400
rect 11060 16360 11061 16400
rect 11019 16351 11061 16360
rect 10924 16099 10964 16108
rect 10924 15728 10964 15737
rect 11020 15728 11060 16351
rect 10964 15688 11060 15728
rect 10924 15679 10964 15688
rect 11116 15644 11156 16528
rect 10732 15506 10772 15515
rect 11020 15604 11156 15644
rect 10635 14972 10677 14981
rect 10635 14932 10636 14972
rect 10676 14932 10677 14972
rect 10635 14923 10677 14932
rect 11020 14897 11060 15604
rect 11116 15547 11156 15556
rect 11116 15233 11156 15507
rect 11212 15308 11252 15317
rect 11115 15224 11157 15233
rect 11115 15184 11116 15224
rect 11156 15184 11157 15224
rect 11115 15175 11157 15184
rect 10828 14888 10868 14897
rect 10732 14804 10772 14813
rect 10636 14720 10676 14729
rect 10348 13637 10388 14008
rect 10539 14048 10581 14057
rect 10539 14008 10540 14048
rect 10580 14008 10581 14048
rect 10539 13999 10581 14008
rect 10539 13880 10581 13889
rect 10539 13840 10540 13880
rect 10580 13840 10581 13880
rect 10539 13831 10581 13840
rect 10540 13746 10580 13831
rect 10347 13628 10389 13637
rect 10347 13588 10348 13628
rect 10388 13588 10389 13628
rect 10347 13579 10389 13588
rect 10636 13376 10676 14680
rect 10732 14141 10772 14764
rect 10828 14393 10868 14848
rect 11019 14888 11061 14897
rect 11019 14848 11020 14888
rect 11060 14848 11061 14888
rect 11019 14839 11061 14848
rect 10923 14804 10965 14813
rect 10923 14764 10924 14804
rect 10964 14764 10965 14804
rect 10923 14755 10965 14764
rect 10924 14670 10964 14755
rect 11020 14720 11060 14729
rect 10827 14384 10869 14393
rect 10827 14344 10828 14384
rect 10868 14344 10869 14384
rect 10827 14335 10869 14344
rect 10923 14300 10965 14309
rect 11020 14300 11060 14680
rect 11116 14309 11156 15175
rect 11212 14720 11252 15268
rect 11308 14813 11348 16612
rect 11500 16409 11540 17200
rect 11499 16400 11541 16409
rect 11499 16360 11500 16400
rect 11540 16360 11541 16400
rect 11499 16351 11541 16360
rect 11403 16316 11445 16325
rect 11403 16276 11404 16316
rect 11444 16276 11445 16316
rect 11403 16267 11445 16276
rect 11404 15560 11444 16267
rect 11596 16232 11636 16241
rect 11499 15896 11541 15905
rect 11499 15856 11500 15896
rect 11540 15856 11541 15896
rect 11499 15847 11541 15856
rect 11500 15737 11540 15847
rect 11499 15728 11541 15737
rect 11499 15688 11500 15728
rect 11540 15688 11541 15728
rect 11499 15679 11541 15688
rect 11596 15569 11636 16192
rect 11788 15905 11828 18115
rect 11980 17660 12020 20047
rect 12172 18761 12212 20056
rect 12267 20096 12309 20105
rect 12267 20056 12268 20096
rect 12308 20056 12309 20096
rect 12267 20047 12309 20056
rect 12460 20096 12500 20105
rect 12268 19962 12308 20047
rect 12460 19853 12500 20056
rect 12556 20096 12596 20105
rect 12459 19844 12501 19853
rect 12459 19804 12460 19844
rect 12500 19804 12501 19844
rect 12459 19795 12501 19804
rect 12363 19676 12405 19685
rect 12363 19636 12364 19676
rect 12404 19636 12405 19676
rect 12363 19627 12405 19636
rect 12267 18920 12309 18929
rect 12267 18880 12268 18920
rect 12308 18880 12309 18920
rect 12267 18871 12309 18880
rect 12171 18752 12213 18761
rect 12171 18712 12172 18752
rect 12212 18712 12213 18752
rect 12171 18703 12213 18712
rect 11884 17620 12020 17660
rect 11787 15896 11829 15905
rect 11787 15856 11788 15896
rect 11828 15856 11829 15896
rect 11787 15847 11829 15856
rect 11691 15728 11733 15737
rect 11691 15688 11692 15728
rect 11732 15688 11733 15728
rect 11691 15679 11733 15688
rect 11404 15511 11444 15520
rect 11595 15560 11637 15569
rect 11595 15520 11596 15560
rect 11636 15520 11637 15560
rect 11595 15511 11637 15520
rect 11500 15476 11540 15487
rect 11500 15401 11540 15436
rect 11692 15476 11732 15679
rect 11692 15427 11732 15436
rect 11788 15560 11828 15569
rect 11499 15392 11541 15401
rect 11499 15352 11500 15392
rect 11540 15352 11541 15392
rect 11499 15343 11541 15352
rect 11596 15392 11636 15401
rect 11403 14972 11445 14981
rect 11403 14932 11404 14972
rect 11444 14932 11445 14972
rect 11403 14923 11445 14932
rect 11307 14804 11349 14813
rect 11307 14764 11308 14804
rect 11348 14764 11349 14804
rect 11307 14755 11349 14764
rect 10923 14260 10924 14300
rect 10964 14260 10965 14300
rect 10923 14251 10965 14260
rect 11014 14260 11060 14300
rect 11115 14300 11157 14309
rect 11115 14260 11116 14300
rect 11156 14260 11157 14300
rect 10731 14132 10773 14141
rect 10731 14092 10732 14132
rect 10772 14092 10773 14132
rect 10731 14083 10773 14092
rect 10828 14048 10868 14057
rect 10924 14048 10964 14251
rect 11014 14132 11054 14260
rect 11115 14251 11157 14260
rect 11212 14216 11252 14680
rect 11404 14720 11444 14923
rect 11596 14897 11636 15352
rect 11788 15317 11828 15520
rect 11884 15485 11924 17620
rect 12268 16157 12308 18871
rect 12364 17240 12404 19627
rect 12459 18248 12501 18257
rect 12459 18208 12460 18248
rect 12500 18208 12501 18248
rect 12459 18199 12501 18208
rect 12460 17417 12500 18199
rect 12556 18173 12596 20056
rect 12713 20081 12753 20090
rect 12713 19760 12753 20041
rect 12713 19720 12788 19760
rect 12748 18845 12788 19720
rect 12844 19265 12884 21811
rect 13036 20777 13076 20862
rect 13035 20768 13077 20777
rect 13035 20728 13036 20768
rect 13076 20728 13077 20768
rect 13035 20719 13077 20728
rect 13132 20768 13172 22315
rect 13228 21701 13268 22651
rect 13323 22364 13365 22373
rect 13323 22324 13324 22364
rect 13364 22324 13365 22364
rect 13323 22315 13365 22324
rect 13324 22230 13364 22315
rect 13227 21692 13269 21701
rect 13227 21652 13228 21692
rect 13268 21652 13269 21692
rect 13227 21643 13269 21652
rect 13132 20600 13172 20728
rect 12940 20560 13172 20600
rect 12843 19256 12885 19265
rect 12843 19216 12844 19256
rect 12884 19216 12885 19256
rect 12843 19207 12885 19216
rect 12844 19122 12884 19207
rect 12747 18836 12789 18845
rect 12747 18796 12748 18836
rect 12788 18796 12789 18836
rect 12747 18787 12789 18796
rect 12651 18248 12693 18257
rect 12651 18208 12652 18248
rect 12692 18208 12693 18248
rect 12651 18199 12693 18208
rect 12555 18164 12597 18173
rect 12555 18124 12556 18164
rect 12596 18124 12597 18164
rect 12555 18115 12597 18124
rect 12652 17744 12692 18199
rect 12459 17408 12501 17417
rect 12459 17368 12460 17408
rect 12500 17368 12501 17408
rect 12459 17359 12501 17368
rect 12652 17249 12692 17704
rect 12843 17660 12885 17669
rect 12843 17620 12844 17660
rect 12884 17620 12885 17660
rect 12843 17611 12885 17620
rect 12844 17526 12884 17611
rect 12940 17408 12980 20560
rect 13228 20357 13268 21643
rect 13323 21440 13365 21449
rect 13323 21400 13324 21440
rect 13364 21400 13365 21440
rect 13323 21391 13365 21400
rect 13227 20348 13269 20357
rect 13227 20308 13228 20348
rect 13268 20308 13269 20348
rect 13227 20299 13269 20308
rect 13227 20180 13269 20189
rect 13227 20140 13228 20180
rect 13268 20140 13269 20180
rect 13227 20131 13269 20140
rect 13036 20096 13076 20105
rect 13036 19508 13076 20056
rect 13132 20096 13172 20105
rect 13132 19685 13172 20056
rect 13131 19676 13173 19685
rect 13131 19636 13132 19676
rect 13172 19636 13173 19676
rect 13131 19627 13173 19636
rect 13036 19459 13076 19468
rect 13228 18920 13268 20131
rect 13324 20021 13364 21391
rect 13323 20012 13365 20021
rect 13323 19972 13324 20012
rect 13364 19972 13365 20012
rect 13323 19963 13365 19972
rect 13420 19760 13460 23668
rect 13515 23120 13557 23129
rect 13515 23080 13516 23120
rect 13556 23080 13557 23120
rect 13515 23071 13557 23080
rect 13516 22986 13556 23071
rect 13612 22709 13652 23752
rect 13804 23742 13844 23827
rect 13900 23801 13940 24004
rect 13995 24004 13996 24044
rect 14036 24004 14037 24044
rect 13995 23995 14037 24004
rect 13996 23960 14036 23995
rect 13996 23909 14036 23920
rect 13899 23792 13941 23801
rect 13899 23752 13900 23792
rect 13940 23752 13941 23792
rect 13899 23743 13941 23752
rect 13995 23708 14037 23717
rect 13995 23668 13996 23708
rect 14036 23668 14037 23708
rect 13995 23659 14037 23668
rect 13611 22700 13653 22709
rect 13611 22660 13612 22700
rect 13652 22660 13653 22700
rect 13611 22651 13653 22660
rect 13515 22532 13557 22541
rect 13515 22492 13516 22532
rect 13556 22492 13557 22532
rect 13515 22483 13557 22492
rect 13516 22398 13556 22483
rect 13611 22448 13653 22457
rect 13611 22408 13612 22448
rect 13652 22408 13653 22448
rect 13611 22399 13653 22408
rect 13515 21860 13557 21869
rect 13515 21820 13516 21860
rect 13556 21820 13557 21860
rect 13515 21811 13557 21820
rect 13516 21608 13556 21811
rect 13516 21559 13556 21568
rect 13612 21104 13652 22399
rect 13804 22280 13844 22289
rect 13708 21776 13748 21785
rect 13804 21776 13844 22240
rect 13900 22280 13940 22291
rect 13900 22205 13940 22240
rect 13899 22196 13941 22205
rect 13899 22156 13900 22196
rect 13940 22156 13941 22196
rect 13899 22147 13941 22156
rect 13996 21785 14036 23659
rect 13748 21736 13844 21776
rect 13995 21776 14037 21785
rect 13995 21736 13996 21776
rect 14036 21736 14037 21776
rect 13708 21727 13748 21736
rect 13995 21727 14037 21736
rect 13899 21692 13941 21701
rect 13899 21652 13900 21692
rect 13940 21652 13941 21692
rect 13899 21643 13941 21652
rect 13900 21608 13940 21643
rect 13900 21557 13940 21568
rect 14092 21440 14132 30640
rect 14187 30640 14188 30680
rect 14228 30640 14229 30680
rect 14187 30631 14229 30640
rect 14380 30680 14420 30689
rect 14188 25304 14228 30631
rect 14380 30512 14420 30640
rect 14475 30680 14517 30689
rect 14475 30640 14476 30680
rect 14516 30640 14517 30680
rect 14475 30631 14517 30640
rect 14380 30472 14516 30512
rect 14380 29840 14420 29849
rect 14476 29840 14516 30472
rect 14571 29840 14613 29849
rect 14476 29800 14572 29840
rect 14612 29800 14613 29840
rect 14380 29177 14420 29800
rect 14571 29791 14613 29800
rect 14572 29756 14612 29791
rect 14572 29705 14612 29716
rect 14379 29168 14421 29177
rect 14379 29128 14380 29168
rect 14420 29128 14421 29168
rect 14379 29119 14421 29128
rect 14283 28748 14325 28757
rect 14283 28708 14284 28748
rect 14324 28708 14325 28748
rect 14283 28699 14325 28708
rect 14284 27497 14324 28699
rect 14379 28328 14421 28337
rect 14379 28288 14380 28328
rect 14420 28288 14421 28328
rect 14379 28279 14421 28288
rect 14283 27488 14325 27497
rect 14283 27448 14284 27488
rect 14324 27448 14325 27488
rect 14283 27439 14325 27448
rect 14284 25481 14324 27439
rect 14380 26573 14420 28279
rect 14476 27656 14516 27665
rect 14476 27245 14516 27616
rect 14571 27572 14613 27581
rect 14571 27532 14572 27572
rect 14612 27532 14613 27572
rect 14571 27523 14613 27532
rect 14475 27236 14517 27245
rect 14475 27196 14476 27236
rect 14516 27196 14517 27236
rect 14475 27187 14517 27196
rect 14379 26564 14421 26573
rect 14379 26524 14380 26564
rect 14420 26524 14421 26564
rect 14379 26515 14421 26524
rect 14572 26312 14612 27523
rect 14572 26263 14612 26272
rect 14380 26130 14420 26139
rect 14380 25901 14420 26090
rect 14379 25892 14421 25901
rect 14379 25852 14380 25892
rect 14420 25852 14421 25892
rect 14379 25843 14421 25852
rect 14668 25724 14708 31891
rect 14763 31856 14805 31865
rect 14763 31816 14764 31856
rect 14804 31816 14805 31856
rect 14763 31807 14805 31816
rect 14764 30101 14804 31807
rect 14860 31352 14900 31363
rect 14860 31277 14900 31312
rect 14859 31268 14901 31277
rect 14859 31228 14860 31268
rect 14900 31228 14901 31268
rect 14859 31219 14901 31228
rect 14859 30932 14901 30941
rect 14859 30892 14860 30932
rect 14900 30892 14901 30932
rect 14859 30883 14901 30892
rect 14860 30680 14900 30883
rect 14860 30631 14900 30640
rect 14956 30596 14996 30605
rect 14956 30269 14996 30556
rect 14955 30260 14997 30269
rect 14955 30220 14956 30260
rect 14996 30220 14997 30260
rect 14955 30211 14997 30220
rect 14763 30092 14805 30101
rect 14763 30052 14764 30092
rect 14804 30052 14805 30092
rect 14763 30043 14805 30052
rect 14955 29924 14997 29933
rect 14955 29884 14956 29924
rect 14996 29884 14997 29924
rect 14955 29875 14997 29884
rect 14764 29840 14804 29849
rect 14764 29261 14804 29800
rect 14763 29252 14805 29261
rect 14763 29212 14764 29252
rect 14804 29212 14805 29252
rect 14763 29203 14805 29212
rect 14859 29168 14901 29177
rect 14859 29128 14860 29168
rect 14900 29128 14901 29168
rect 14859 29119 14901 29128
rect 14956 29168 14996 29875
rect 15052 29849 15092 32143
rect 15148 31529 15188 32152
rect 15244 32192 15284 32201
rect 15147 31520 15189 31529
rect 15147 31480 15148 31520
rect 15188 31480 15189 31520
rect 15147 31471 15189 31480
rect 15244 31361 15284 32152
rect 15340 32192 15380 32201
rect 15532 32192 15572 32201
rect 15380 32152 15532 32192
rect 15340 32143 15380 32152
rect 15532 32143 15572 32152
rect 15435 32024 15477 32033
rect 15435 31984 15436 32024
rect 15476 31984 15477 32024
rect 15435 31975 15477 31984
rect 15243 31352 15285 31361
rect 15243 31312 15244 31352
rect 15284 31312 15285 31352
rect 15243 31303 15285 31312
rect 15339 31268 15381 31277
rect 15339 31228 15340 31268
rect 15380 31228 15381 31268
rect 15339 31219 15381 31228
rect 15147 30596 15189 30605
rect 15147 30556 15148 30596
rect 15188 30556 15189 30596
rect 15147 30547 15189 30556
rect 15051 29840 15093 29849
rect 15051 29800 15052 29840
rect 15092 29800 15093 29840
rect 15051 29791 15093 29800
rect 15148 29672 15188 30547
rect 14956 29119 14996 29128
rect 15052 29632 15188 29672
rect 14763 28328 14805 28337
rect 14763 28288 14764 28328
rect 14804 28288 14805 28328
rect 14763 28279 14805 28288
rect 14764 28194 14804 28279
rect 14763 27992 14805 28001
rect 14763 27952 14764 27992
rect 14804 27952 14805 27992
rect 14763 27943 14805 27952
rect 14764 26144 14804 27943
rect 14860 26816 14900 29119
rect 15052 28337 15092 29632
rect 15340 29504 15380 31219
rect 15436 30689 15476 31975
rect 15531 31940 15573 31949
rect 15531 31900 15532 31940
rect 15572 31900 15573 31940
rect 15531 31891 15573 31900
rect 15532 31806 15572 31891
rect 15531 31520 15573 31529
rect 15531 31480 15532 31520
rect 15572 31480 15573 31520
rect 15531 31471 15573 31480
rect 15532 31025 15572 31471
rect 15531 31016 15573 31025
rect 15531 30976 15532 31016
rect 15572 30976 15573 31016
rect 15531 30967 15573 30976
rect 15435 30680 15477 30689
rect 15435 30640 15436 30680
rect 15476 30640 15477 30680
rect 15435 30631 15477 30640
rect 15436 30546 15476 30631
rect 15628 30101 15668 32320
rect 15723 32192 15765 32201
rect 15723 32152 15724 32192
rect 15764 32152 15765 32192
rect 15723 32143 15765 32152
rect 15820 32192 15860 32479
rect 16204 32369 16244 36436
rect 16299 36392 16341 36401
rect 16299 36352 16300 36392
rect 16340 36352 16341 36392
rect 16299 36343 16341 36352
rect 16300 36056 16340 36343
rect 16457 36182 16497 36673
rect 16588 36182 16628 36191
rect 16457 36142 16588 36182
rect 16684 36182 16724 36688
rect 16780 36644 16820 36653
rect 16780 36401 16820 36604
rect 16876 36560 16916 37183
rect 16971 36728 17013 36737
rect 16971 36688 16972 36728
rect 17012 36688 17013 36728
rect 16971 36679 17013 36688
rect 17068 36728 17108 36739
rect 16972 36644 17012 36679
rect 17068 36653 17108 36688
rect 16972 36593 17012 36604
rect 17067 36644 17109 36653
rect 17067 36604 17068 36644
rect 17108 36604 17109 36644
rect 17067 36595 17109 36604
rect 16876 36511 16916 36520
rect 16779 36392 16821 36401
rect 16779 36352 16780 36392
rect 16820 36352 16821 36392
rect 16779 36343 16821 36352
rect 17164 36233 17204 37183
rect 17259 37148 17301 37157
rect 17259 37108 17260 37148
rect 17300 37108 17301 37148
rect 17259 37099 17301 37108
rect 17260 36728 17300 37099
rect 17356 36821 17396 37444
rect 17452 37241 17492 37780
rect 17835 37652 17877 37661
rect 17835 37612 17836 37652
rect 17876 37612 17877 37652
rect 17835 37603 17877 37612
rect 17836 37442 17876 37603
rect 17932 37577 17972 39040
rect 18124 39040 18260 39080
rect 18412 39080 18452 39089
rect 18604 39080 18644 40972
rect 18700 40963 18740 40972
rect 19083 41012 19125 41021
rect 19083 40972 19084 41012
rect 19124 40972 19125 41012
rect 19083 40963 19125 40972
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 19179 40676 19221 40685
rect 19179 40636 19180 40676
rect 19220 40636 19221 40676
rect 19179 40627 19221 40636
rect 19372 40676 19412 41551
rect 19467 41432 19509 41441
rect 19467 41392 19468 41432
rect 19508 41392 19509 41432
rect 19467 41383 19509 41392
rect 19468 41298 19508 41383
rect 19564 40676 19604 42475
rect 19755 42356 19797 42365
rect 19755 42316 19756 42356
rect 19796 42316 19797 42356
rect 19755 42307 19797 42316
rect 19756 41264 19796 42307
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 19851 41516 19893 41525
rect 19851 41476 19852 41516
rect 19892 41476 19893 41516
rect 19851 41467 19893 41476
rect 19852 41432 19892 41467
rect 19852 41381 19892 41392
rect 21387 41432 21429 41441
rect 21387 41392 21388 41432
rect 21428 41392 21429 41432
rect 21387 41383 21429 41392
rect 19756 41224 19892 41264
rect 19659 41180 19701 41189
rect 19659 41140 19660 41180
rect 19700 41140 19701 41180
rect 19659 41131 19701 41140
rect 19660 41046 19700 41131
rect 19755 41096 19797 41105
rect 19755 41056 19756 41096
rect 19796 41056 19797 41096
rect 19755 41047 19797 41056
rect 19756 40676 19796 41047
rect 19564 40636 19700 40676
rect 19372 40627 19412 40636
rect 18987 40592 19029 40601
rect 18987 40552 18988 40592
rect 19028 40552 19029 40592
rect 18987 40543 19029 40552
rect 18700 40508 18740 40517
rect 18700 40265 18740 40468
rect 18988 40458 19028 40543
rect 19180 40508 19220 40627
rect 19180 40459 19220 40468
rect 19564 40508 19604 40517
rect 18699 40256 18741 40265
rect 18699 40216 18700 40256
rect 18740 40216 18741 40256
rect 18699 40207 18741 40216
rect 18891 40172 18933 40181
rect 18891 40132 18892 40172
rect 18932 40132 18933 40172
rect 18891 40123 18933 40132
rect 18699 39920 18741 39929
rect 18699 39880 18700 39920
rect 18740 39880 18741 39920
rect 18699 39871 18741 39880
rect 18700 39786 18740 39871
rect 18892 39668 18932 40123
rect 19467 40004 19509 40013
rect 19467 39964 19468 40004
rect 19508 39964 19509 40004
rect 19467 39955 19509 39964
rect 19180 39920 19220 39929
rect 19468 39920 19508 39955
rect 19220 39880 19412 39920
rect 19180 39871 19220 39880
rect 19083 39836 19125 39845
rect 19083 39796 19084 39836
rect 19124 39796 19125 39836
rect 19083 39787 19125 39796
rect 19084 39752 19124 39787
rect 19084 39701 19124 39712
rect 19276 39752 19316 39761
rect 18892 39619 18932 39628
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 18891 39080 18933 39089
rect 18604 39040 18740 39080
rect 18124 39005 18164 39040
rect 18122 38996 18164 39005
rect 18122 38956 18123 38996
rect 18163 38956 18164 38996
rect 18122 38947 18164 38956
rect 18316 38996 18356 39005
rect 18220 38912 18260 38921
rect 18028 38744 18068 38753
rect 18028 37820 18068 38704
rect 18220 38492 18260 38872
rect 18316 38669 18356 38956
rect 18412 38753 18452 39040
rect 18507 38996 18549 39005
rect 18507 38956 18508 38996
rect 18548 38956 18549 38996
rect 18507 38947 18549 38956
rect 18508 38862 18548 38947
rect 18604 38912 18644 38921
rect 18411 38744 18453 38753
rect 18411 38704 18412 38744
rect 18452 38704 18453 38744
rect 18411 38695 18453 38704
rect 18604 38669 18644 38872
rect 18315 38660 18357 38669
rect 18315 38620 18316 38660
rect 18356 38620 18357 38660
rect 18315 38611 18357 38620
rect 18603 38660 18645 38669
rect 18603 38620 18604 38660
rect 18644 38620 18645 38660
rect 18603 38611 18645 38620
rect 18316 38492 18356 38611
rect 18700 38585 18740 39040
rect 18891 39040 18892 39080
rect 18932 39040 18933 39080
rect 18891 39031 18933 39040
rect 18892 38946 18932 39031
rect 19084 38996 19124 39005
rect 18795 38912 18837 38921
rect 18795 38872 18796 38912
rect 18836 38872 18837 38912
rect 18795 38863 18837 38872
rect 18796 38778 18836 38863
rect 18411 38576 18453 38585
rect 18411 38536 18412 38576
rect 18452 38536 18453 38576
rect 18411 38527 18453 38536
rect 18699 38576 18741 38585
rect 18699 38536 18700 38576
rect 18740 38536 18741 38576
rect 18699 38527 18741 38536
rect 18124 38452 18260 38492
rect 18305 38452 18356 38492
rect 18124 38324 18164 38452
rect 18305 38408 18345 38452
rect 18225 38368 18345 38408
rect 18225 38324 18265 38368
rect 18412 38324 18452 38527
rect 18603 38408 18645 38417
rect 18603 38368 18604 38408
rect 18644 38368 18645 38408
rect 18603 38359 18645 38368
rect 18123 38284 18164 38324
rect 18220 38284 18265 38324
rect 18364 38284 18452 38324
rect 18123 38236 18163 38284
rect 18220 38240 18260 38284
rect 18123 38196 18164 38236
rect 18124 37988 18164 38196
rect 18220 38191 18260 38200
rect 18364 38230 18404 38284
rect 18507 38240 18549 38249
rect 18507 38200 18508 38240
rect 18548 38200 18549 38240
rect 18507 38191 18549 38200
rect 18604 38240 18644 38359
rect 19084 38333 19124 38956
rect 19179 38996 19221 39005
rect 19179 38956 19180 38996
rect 19220 38956 19221 38996
rect 19179 38947 19221 38956
rect 18890 38324 18932 38333
rect 18890 38284 18891 38324
rect 18931 38284 18932 38324
rect 18890 38275 18932 38284
rect 19083 38324 19125 38333
rect 19083 38284 19084 38324
rect 19124 38284 19125 38324
rect 19083 38275 19125 38284
rect 18604 38191 18644 38200
rect 18705 38240 18745 38249
rect 18892 38240 18932 38275
rect 18988 38240 19028 38249
rect 18892 38200 18988 38240
rect 18364 38181 18404 38190
rect 18508 38106 18548 38191
rect 18220 37988 18260 37997
rect 18124 37948 18220 37988
rect 18220 37939 18260 37948
rect 18411 37904 18453 37913
rect 18705 37904 18745 38200
rect 18988 38191 19028 38200
rect 19084 38156 19124 38165
rect 19084 37997 19124 38116
rect 19180 38072 19220 38947
rect 19276 38921 19316 39712
rect 19275 38912 19317 38921
rect 19275 38872 19276 38912
rect 19316 38872 19317 38912
rect 19275 38863 19317 38872
rect 19275 38744 19317 38753
rect 19275 38704 19276 38744
rect 19316 38704 19317 38744
rect 19275 38695 19317 38704
rect 19276 38610 19316 38695
rect 19275 38408 19317 38417
rect 19275 38368 19276 38408
rect 19316 38368 19317 38408
rect 19275 38359 19317 38368
rect 19180 38023 19220 38032
rect 19276 38156 19316 38359
rect 19372 38249 19412 39880
rect 19468 39869 19508 39880
rect 19564 39257 19604 40468
rect 19660 39836 19700 40636
rect 19756 40627 19796 40636
rect 19852 39920 19892 41224
rect 20043 41180 20085 41189
rect 20043 41140 20044 41180
rect 20084 41140 20085 41180
rect 20043 41131 20085 41140
rect 20044 41046 20084 41131
rect 19947 40928 19989 40937
rect 19947 40888 19948 40928
rect 19988 40888 19989 40928
rect 19947 40879 19989 40888
rect 19948 40508 19988 40879
rect 19948 40459 19988 40468
rect 20140 40349 20180 40434
rect 20236 40424 20276 40433
rect 21195 40424 21237 40433
rect 20276 40384 20756 40424
rect 20236 40375 20276 40384
rect 20139 40340 20181 40349
rect 20139 40300 20140 40340
rect 20180 40300 20181 40340
rect 20139 40291 20181 40300
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 19852 39871 19892 39880
rect 19660 39796 19796 39836
rect 19659 39668 19701 39677
rect 19659 39628 19660 39668
rect 19700 39628 19701 39668
rect 19659 39619 19701 39628
rect 19660 39534 19700 39619
rect 19563 39248 19605 39257
rect 19563 39208 19564 39248
rect 19604 39208 19605 39248
rect 19563 39199 19605 39208
rect 19756 39080 19796 39796
rect 20043 39668 20085 39677
rect 20043 39628 20044 39668
rect 20084 39628 20085 39668
rect 20043 39619 20085 39628
rect 20044 39534 20084 39619
rect 19852 39080 19892 39089
rect 19756 39040 19852 39080
rect 19852 39031 19892 39040
rect 19467 38996 19509 39005
rect 19467 38956 19468 38996
rect 19508 38956 19509 38996
rect 19467 38947 19509 38956
rect 20044 38996 20084 39005
rect 19468 38862 19508 38947
rect 19563 38912 19605 38921
rect 19563 38872 19564 38912
rect 19604 38872 19605 38912
rect 19563 38863 19605 38872
rect 19564 38417 19604 38863
rect 20044 38837 20084 38956
rect 20043 38828 20085 38837
rect 20043 38788 20044 38828
rect 20084 38788 20085 38828
rect 20043 38779 20085 38788
rect 19660 38744 19700 38753
rect 19700 38704 19796 38744
rect 19660 38695 19700 38704
rect 19563 38408 19605 38417
rect 19563 38368 19564 38408
rect 19604 38368 19605 38408
rect 19563 38359 19605 38368
rect 19371 38240 19413 38249
rect 19371 38200 19372 38240
rect 19412 38200 19413 38240
rect 19756 38240 19796 38704
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 19756 38200 19892 38240
rect 19371 38191 19413 38200
rect 19083 37988 19125 37997
rect 19083 37948 19084 37988
rect 19124 37948 19125 37988
rect 19083 37939 19125 37948
rect 18411 37864 18412 37904
rect 18452 37864 18453 37904
rect 18411 37855 18453 37864
rect 18508 37864 18745 37904
rect 18028 37780 18164 37820
rect 17931 37568 17973 37577
rect 17931 37528 17932 37568
rect 17972 37528 17973 37568
rect 17931 37519 17973 37528
rect 17932 37442 17972 37451
rect 17836 37402 17932 37442
rect 17626 37385 17666 37394
rect 17932 37393 17972 37402
rect 17626 37316 17666 37345
rect 18124 37325 18164 37780
rect 18315 37652 18357 37661
rect 18315 37612 18316 37652
rect 18356 37612 18357 37652
rect 18315 37603 18357 37612
rect 18316 37518 18356 37603
rect 18028 37316 18068 37325
rect 17626 37276 17684 37316
rect 17451 37232 17493 37241
rect 17451 37192 17452 37232
rect 17492 37192 17493 37232
rect 17451 37183 17493 37192
rect 17644 36821 17684 37276
rect 17740 37276 18028 37316
rect 17355 36812 17397 36821
rect 17355 36772 17356 36812
rect 17396 36772 17397 36812
rect 17355 36763 17397 36772
rect 17643 36812 17685 36821
rect 17643 36772 17644 36812
rect 17684 36772 17685 36812
rect 17643 36763 17685 36772
rect 17260 36679 17300 36688
rect 17452 36728 17492 36737
rect 17356 36644 17396 36653
rect 17259 36560 17301 36569
rect 17259 36520 17260 36560
rect 17300 36520 17301 36560
rect 17259 36511 17301 36520
rect 17163 36224 17205 36233
rect 17163 36184 17164 36224
rect 17204 36184 17205 36224
rect 16684 36149 16820 36182
rect 17163 36175 17205 36184
rect 16684 36142 16821 36149
rect 16588 36133 16628 36142
rect 16779 36140 16821 36142
rect 16779 36100 16780 36140
rect 16820 36100 16821 36140
rect 16779 36091 16821 36100
rect 16971 36140 17013 36149
rect 16971 36100 16972 36140
rect 17012 36100 17013 36140
rect 16971 36091 17013 36100
rect 16396 36056 16436 36065
rect 16300 36016 16396 36056
rect 16396 36007 16436 36016
rect 16491 36056 16533 36065
rect 16491 36016 16492 36056
rect 16532 36016 16533 36056
rect 16491 36007 16533 36016
rect 16395 35804 16437 35813
rect 16395 35764 16396 35804
rect 16436 35764 16437 35804
rect 16395 35755 16437 35764
rect 16299 34040 16341 34049
rect 16299 34000 16300 34040
rect 16340 34000 16341 34040
rect 16299 33991 16341 34000
rect 16300 33293 16340 33991
rect 16299 33284 16341 33293
rect 16299 33244 16300 33284
rect 16340 33244 16341 33284
rect 16299 33235 16341 33244
rect 16299 32864 16341 32873
rect 16299 32824 16300 32864
rect 16340 32824 16341 32864
rect 16299 32822 16341 32824
rect 16299 32815 16300 32822
rect 16340 32815 16341 32822
rect 16396 32864 16436 35755
rect 16492 33965 16532 36007
rect 16780 35972 16820 36091
rect 16588 35932 16820 35972
rect 16491 33956 16533 33965
rect 16491 33916 16492 33956
rect 16532 33916 16533 33956
rect 16491 33907 16533 33916
rect 16300 32729 16340 32782
rect 16299 32612 16341 32621
rect 16299 32572 16300 32612
rect 16340 32572 16341 32612
rect 16299 32563 16341 32572
rect 16011 32360 16053 32369
rect 16011 32320 16012 32360
rect 16052 32320 16053 32360
rect 16011 32311 16053 32320
rect 16203 32360 16245 32369
rect 16203 32320 16204 32360
rect 16244 32320 16245 32360
rect 16203 32311 16245 32320
rect 15820 32143 15860 32152
rect 15724 32058 15764 32143
rect 15723 31520 15765 31529
rect 15723 31480 15724 31520
rect 15764 31480 15765 31520
rect 15723 31471 15765 31480
rect 15627 30092 15669 30101
rect 15627 30052 15628 30092
rect 15668 30052 15669 30092
rect 15627 30043 15669 30052
rect 15627 29840 15669 29849
rect 15627 29800 15628 29840
rect 15668 29800 15669 29840
rect 15627 29791 15669 29800
rect 15340 29464 15476 29504
rect 15339 29336 15381 29345
rect 15339 29296 15340 29336
rect 15380 29296 15381 29336
rect 15339 29287 15381 29296
rect 15340 29168 15380 29287
rect 15340 29009 15380 29128
rect 15339 29000 15381 29009
rect 15339 28960 15340 29000
rect 15380 28960 15381 29000
rect 15339 28951 15381 28960
rect 15148 28916 15188 28925
rect 15051 28328 15093 28337
rect 15051 28288 15052 28328
rect 15092 28288 15093 28328
rect 15148 28328 15188 28876
rect 15244 28328 15284 28337
rect 15148 28288 15244 28328
rect 15051 28279 15093 28288
rect 15244 28279 15284 28288
rect 15340 28328 15380 28337
rect 14956 28160 14996 28169
rect 14956 27651 14996 28120
rect 15147 28160 15189 28169
rect 15147 28120 15148 28160
rect 15188 28120 15189 28160
rect 15147 28111 15189 28120
rect 15148 27740 15188 28111
rect 15340 28001 15380 28288
rect 15339 27992 15381 28001
rect 15339 27952 15340 27992
rect 15380 27952 15381 27992
rect 15339 27943 15381 27952
rect 15148 27691 15188 27700
rect 14956 27602 14996 27611
rect 15340 27656 15380 27665
rect 15436 27656 15476 29464
rect 15531 29336 15573 29345
rect 15531 29296 15532 29336
rect 15572 29296 15573 29336
rect 15531 29287 15573 29296
rect 15532 29202 15572 29287
rect 15628 29168 15668 29791
rect 15628 29119 15668 29128
rect 15531 29084 15573 29093
rect 15531 29044 15532 29084
rect 15572 29044 15573 29084
rect 15531 29035 15573 29044
rect 15380 27616 15476 27656
rect 15340 27607 15380 27616
rect 15532 27236 15572 29035
rect 15627 28916 15669 28925
rect 15627 28876 15628 28916
rect 15668 28876 15669 28916
rect 15627 28867 15669 28876
rect 15436 27196 15572 27236
rect 15339 26900 15381 26909
rect 15339 26860 15340 26900
rect 15380 26860 15381 26900
rect 15339 26851 15381 26860
rect 14860 26767 14900 26776
rect 15340 26766 15380 26851
rect 15052 26648 15092 26657
rect 14955 26228 14997 26237
rect 14955 26188 14956 26228
rect 14996 26188 14997 26228
rect 14955 26179 14997 26188
rect 14956 26144 14996 26179
rect 14764 26104 14900 26144
rect 14764 25901 14804 25986
rect 14763 25892 14805 25901
rect 14763 25852 14764 25892
rect 14804 25852 14805 25892
rect 14763 25843 14805 25852
rect 14668 25684 14804 25724
rect 14667 25556 14709 25565
rect 14667 25516 14668 25556
rect 14708 25516 14709 25556
rect 14667 25507 14709 25516
rect 14283 25472 14325 25481
rect 14283 25432 14284 25472
rect 14324 25432 14325 25472
rect 14283 25423 14325 25432
rect 14668 25422 14708 25507
rect 14475 25388 14517 25397
rect 14475 25348 14476 25388
rect 14516 25348 14517 25388
rect 14475 25339 14517 25348
rect 14188 25264 14420 25304
rect 14188 25136 14228 25145
rect 14228 25096 14324 25136
rect 14188 25087 14228 25096
rect 14284 24627 14324 25096
rect 14284 24578 14324 24587
rect 14283 24464 14325 24473
rect 14283 24424 14284 24464
rect 14324 24424 14325 24464
rect 14283 24415 14325 24424
rect 14188 23876 14228 23885
rect 14188 23129 14228 23836
rect 14187 23120 14229 23129
rect 14187 23080 14188 23120
rect 14228 23080 14229 23120
rect 14187 23071 14229 23080
rect 14188 22541 14228 23071
rect 14187 22532 14229 22541
rect 14187 22492 14188 22532
rect 14228 22492 14229 22532
rect 14187 22483 14229 22492
rect 14284 22457 14324 24415
rect 14380 24128 14420 25264
rect 14476 25254 14516 25339
rect 14571 25304 14613 25313
rect 14571 25264 14572 25304
rect 14612 25264 14613 25304
rect 14571 25255 14613 25264
rect 14476 24800 14516 24809
rect 14572 24800 14612 25255
rect 14516 24760 14612 24800
rect 14476 24751 14516 24760
rect 14764 24716 14804 25684
rect 14860 25136 14900 26104
rect 14956 26093 14996 26104
rect 15052 25976 15092 26608
rect 15243 26480 15285 26489
rect 15243 26440 15244 26480
rect 15284 26440 15285 26480
rect 15243 26431 15285 26440
rect 14956 25936 15092 25976
rect 14956 25304 14996 25936
rect 15244 25724 15284 26431
rect 15148 25684 15284 25724
rect 14956 25255 14996 25264
rect 15052 25304 15092 25313
rect 15052 25136 15092 25264
rect 15148 25229 15188 25684
rect 15243 25556 15285 25565
rect 15243 25516 15244 25556
rect 15284 25516 15285 25556
rect 15243 25507 15285 25516
rect 15147 25220 15189 25229
rect 15147 25180 15148 25220
rect 15188 25180 15189 25220
rect 15147 25171 15189 25180
rect 14860 25096 15092 25136
rect 14955 24800 14997 24809
rect 14955 24760 14956 24800
rect 14996 24760 14997 24800
rect 14955 24751 14997 24760
rect 14668 24676 14804 24716
rect 14380 24088 14516 24128
rect 14379 23960 14421 23969
rect 14379 23920 14380 23960
rect 14420 23920 14421 23960
rect 14379 23911 14421 23920
rect 14380 23826 14420 23911
rect 14283 22448 14325 22457
rect 14283 22408 14284 22448
rect 14324 22408 14325 22448
rect 14283 22399 14325 22408
rect 14283 22280 14325 22289
rect 14283 22240 14284 22280
rect 14324 22240 14325 22280
rect 14283 22231 14325 22240
rect 14380 22280 14420 22289
rect 14187 22196 14229 22205
rect 14187 22156 14188 22196
rect 14228 22156 14229 22196
rect 14187 22147 14229 22156
rect 13900 21400 14132 21440
rect 13516 21064 13844 21104
rect 13516 20852 13556 21064
rect 13516 20803 13556 20812
rect 13707 20852 13749 20861
rect 13707 20812 13708 20852
rect 13748 20812 13749 20852
rect 13707 20803 13749 20812
rect 13612 20768 13652 20777
rect 13612 20189 13652 20728
rect 13611 20180 13653 20189
rect 13611 20140 13612 20180
rect 13652 20140 13653 20180
rect 13611 20131 13653 20140
rect 13324 19720 13460 19760
rect 13516 20012 13556 20021
rect 13324 19424 13364 19720
rect 13516 19517 13556 19972
rect 13611 20012 13653 20021
rect 13611 19972 13612 20012
rect 13652 19972 13653 20012
rect 13611 19963 13653 19972
rect 13612 19878 13652 19963
rect 13611 19676 13653 19685
rect 13611 19636 13612 19676
rect 13652 19636 13653 19676
rect 13611 19627 13653 19636
rect 13515 19508 13557 19517
rect 13515 19468 13516 19508
rect 13556 19468 13557 19508
rect 13515 19459 13557 19468
rect 13324 19384 13460 19424
rect 13324 19256 13364 19267
rect 13324 19181 13364 19216
rect 13323 19172 13365 19181
rect 13323 19132 13324 19172
rect 13364 19132 13365 19172
rect 13323 19123 13365 19132
rect 13036 18880 13268 18920
rect 13036 18584 13076 18880
rect 13323 18836 13365 18845
rect 13323 18796 13324 18836
rect 13364 18796 13365 18836
rect 13323 18787 13365 18796
rect 13227 18752 13269 18761
rect 13227 18712 13228 18752
rect 13268 18712 13269 18752
rect 13227 18703 13269 18712
rect 13228 18618 13268 18703
rect 13036 18257 13076 18544
rect 13035 18248 13077 18257
rect 13035 18208 13036 18248
rect 13076 18208 13077 18248
rect 13035 18199 13077 18208
rect 13227 18248 13269 18257
rect 13227 18208 13228 18248
rect 13268 18208 13269 18248
rect 13227 18199 13269 18208
rect 13131 18164 13173 18173
rect 13131 18124 13132 18164
rect 13172 18124 13173 18164
rect 13131 18115 13173 18124
rect 13132 17996 13172 18115
rect 13036 17744 13076 17755
rect 13036 17669 13076 17704
rect 13035 17660 13077 17669
rect 13035 17620 13036 17660
rect 13076 17620 13077 17660
rect 13132 17660 13172 17956
rect 13228 17921 13268 18199
rect 13324 17996 13364 18787
rect 13420 18752 13460 19384
rect 13420 18712 13556 18752
rect 13420 18584 13460 18593
rect 13420 18173 13460 18544
rect 13419 18164 13461 18173
rect 13419 18124 13420 18164
rect 13460 18124 13461 18164
rect 13419 18115 13461 18124
rect 13324 17947 13364 17956
rect 13419 17996 13461 18005
rect 13419 17956 13420 17996
rect 13460 17956 13461 17996
rect 13419 17947 13461 17956
rect 13227 17912 13269 17921
rect 13227 17872 13228 17912
rect 13268 17872 13269 17912
rect 13227 17863 13269 17872
rect 13323 17660 13365 17669
rect 13132 17620 13324 17660
rect 13364 17620 13365 17660
rect 13035 17611 13077 17620
rect 13323 17611 13365 17620
rect 12748 17368 12980 17408
rect 12651 17240 12693 17249
rect 12364 17200 12500 17240
rect 12363 16820 12405 16829
rect 12363 16780 12364 16820
rect 12404 16780 12405 16820
rect 12363 16771 12405 16780
rect 12267 16148 12309 16157
rect 12267 16108 12268 16148
rect 12308 16108 12309 16148
rect 12267 16099 12309 16108
rect 12171 15728 12213 15737
rect 12171 15688 12172 15728
rect 12212 15688 12213 15728
rect 12171 15679 12213 15688
rect 11980 15560 12020 15569
rect 11883 15476 11925 15485
rect 11883 15436 11884 15476
rect 11924 15436 11925 15476
rect 11883 15427 11925 15436
rect 11787 15308 11829 15317
rect 11787 15268 11788 15308
rect 11828 15268 11829 15308
rect 11787 15259 11829 15268
rect 11980 15149 12020 15520
rect 11979 15140 12021 15149
rect 11979 15100 11980 15140
rect 12020 15100 12021 15140
rect 11979 15091 12021 15100
rect 11595 14888 11637 14897
rect 11595 14848 11596 14888
rect 11636 14848 11637 14888
rect 11595 14839 11637 14848
rect 11307 14636 11349 14645
rect 11307 14596 11308 14636
rect 11348 14596 11349 14636
rect 11307 14587 11349 14596
rect 11308 14502 11348 14587
rect 11404 14309 11444 14680
rect 11596 14720 11636 14729
rect 11596 14477 11636 14680
rect 11595 14468 11637 14477
rect 11595 14428 11596 14468
rect 11636 14428 11637 14468
rect 11595 14419 11637 14428
rect 11403 14300 11445 14309
rect 11403 14260 11404 14300
rect 11444 14260 11445 14300
rect 11403 14251 11445 14260
rect 11212 14176 11348 14216
rect 11014 14092 11060 14132
rect 10868 14008 10964 14048
rect 10828 13999 10868 14008
rect 10731 13880 10773 13889
rect 10731 13840 10732 13880
rect 10772 13840 10773 13880
rect 10731 13831 10773 13840
rect 10444 13336 10676 13376
rect 10444 13292 10484 13336
rect 10444 13243 10484 13252
rect 10348 13208 10388 13217
rect 10252 13168 10348 13208
rect 10348 13159 10388 13168
rect 10539 13208 10581 13217
rect 10539 13168 10540 13208
rect 10580 13168 10581 13208
rect 10539 13159 10581 13168
rect 10636 13208 10676 13217
rect 10732 13208 10772 13831
rect 10828 13460 10868 13469
rect 11020 13460 11060 14092
rect 11115 14048 11157 14057
rect 11115 14008 11116 14048
rect 11156 14008 11157 14048
rect 11115 13999 11157 14008
rect 11212 14048 11252 14059
rect 11116 13805 11156 13999
rect 11212 13973 11252 14008
rect 11211 13964 11253 13973
rect 11211 13924 11212 13964
rect 11252 13924 11253 13964
rect 11211 13915 11253 13924
rect 11115 13796 11157 13805
rect 11115 13756 11116 13796
rect 11156 13756 11157 13796
rect 11115 13747 11157 13756
rect 10868 13420 11060 13460
rect 10828 13411 10868 13420
rect 10676 13168 10772 13208
rect 11116 13208 11156 13217
rect 10636 13159 10676 13168
rect 10155 12704 10197 12713
rect 10155 12664 10156 12704
rect 10196 12664 10197 12704
rect 10155 12655 10197 12664
rect 10251 12620 10293 12629
rect 10251 12580 10252 12620
rect 10292 12580 10293 12620
rect 10251 12571 10293 12580
rect 10156 12536 10196 12547
rect 10156 12461 10196 12496
rect 10252 12536 10292 12571
rect 10252 12485 10292 12496
rect 10155 12452 10197 12461
rect 10155 12412 10156 12452
rect 10196 12412 10197 12452
rect 10155 12403 10197 12412
rect 10251 12368 10293 12377
rect 10251 12328 10252 12368
rect 10292 12328 10293 12368
rect 10251 12319 10293 12328
rect 10252 11285 10292 12319
rect 10251 11276 10293 11285
rect 10251 11236 10252 11276
rect 10292 11236 10293 11276
rect 10251 11227 10293 11236
rect 10443 10940 10485 10949
rect 10443 10900 10444 10940
rect 10484 10900 10485 10940
rect 10443 10891 10485 10900
rect 10156 10312 10388 10352
rect 10156 10184 10196 10312
rect 10156 10135 10196 10144
rect 10252 10184 10292 10195
rect 10252 10109 10292 10144
rect 10251 10100 10293 10109
rect 10251 10060 10252 10100
rect 10292 10060 10293 10100
rect 10251 10051 10293 10060
rect 10059 10016 10101 10025
rect 10059 9976 10060 10016
rect 10100 9976 10101 10016
rect 10059 9967 10101 9976
rect 10155 9932 10197 9941
rect 10155 9892 10156 9932
rect 10196 9892 10197 9932
rect 10155 9883 10197 9892
rect 9964 9680 10004 9689
rect 9867 9596 9909 9605
rect 9867 9556 9868 9596
rect 9908 9556 9909 9596
rect 9867 9547 9909 9556
rect 9772 9512 9812 9521
rect 9676 9472 9772 9512
rect 9580 9378 9620 9463
rect 9579 9092 9621 9101
rect 9579 9052 9580 9092
rect 9620 9052 9621 9092
rect 9579 9043 9621 9052
rect 9483 8252 9525 8261
rect 9483 8212 9484 8252
rect 9524 8212 9525 8252
rect 9483 8203 9525 8212
rect 9292 7951 9332 7960
rect 9580 7916 9620 9043
rect 9676 8345 9716 9472
rect 9772 9463 9812 9472
rect 9868 9512 9908 9547
rect 9868 9462 9908 9472
rect 9867 9260 9909 9269
rect 9867 9220 9868 9260
rect 9908 9220 9909 9260
rect 9964 9260 10004 9640
rect 10059 9512 10101 9521
rect 10059 9472 10060 9512
rect 10100 9472 10101 9512
rect 10059 9463 10101 9472
rect 10156 9512 10196 9883
rect 10257 9512 10297 9521
rect 10060 9378 10100 9463
rect 9964 9220 10100 9260
rect 9867 9211 9909 9220
rect 9772 8672 9812 8683
rect 9772 8597 9812 8632
rect 9771 8588 9813 8597
rect 9771 8548 9772 8588
rect 9812 8548 9813 8588
rect 9771 8539 9813 8548
rect 9675 8336 9717 8345
rect 9675 8296 9676 8336
rect 9716 8296 9717 8336
rect 9675 8287 9717 8296
rect 9771 8252 9813 8261
rect 9771 8212 9772 8252
rect 9812 8212 9813 8252
rect 9771 8203 9813 8212
rect 9676 8093 9716 8137
rect 9675 8084 9717 8093
rect 9675 8044 9676 8084
rect 9716 8044 9717 8084
rect 9675 8042 9717 8044
rect 9675 8035 9676 8042
rect 9716 8035 9717 8042
rect 9676 7993 9716 8002
rect 9772 7916 9812 8203
rect 9580 7876 9716 7916
rect 9484 7832 9524 7841
rect 9196 7792 9484 7832
rect 9484 7783 9524 7792
rect 9579 7748 9621 7757
rect 9100 7708 9236 7748
rect 9099 7496 9141 7505
rect 9099 7456 9100 7496
rect 9140 7456 9141 7496
rect 9099 7447 9141 7456
rect 9003 7412 9045 7421
rect 9003 7372 9004 7412
rect 9044 7372 9045 7412
rect 9003 7363 9045 7372
rect 8907 7328 8949 7337
rect 8907 7288 8908 7328
rect 8948 7288 8949 7328
rect 8907 7279 8949 7288
rect 8908 7001 8948 7279
rect 9003 7160 9045 7169
rect 9003 7120 9004 7160
rect 9044 7120 9045 7160
rect 9003 7111 9045 7120
rect 9100 7160 9140 7447
rect 9100 7111 9140 7120
rect 9004 7026 9044 7111
rect 8716 6952 8852 6992
rect 8907 6992 8949 7001
rect 8907 6952 8908 6992
rect 8948 6952 8949 6992
rect 8619 6656 8661 6665
rect 8619 6616 8620 6656
rect 8660 6616 8661 6656
rect 8619 6607 8661 6616
rect 8620 6488 8660 6607
rect 8620 6439 8660 6448
rect 8620 6320 8660 6329
rect 8716 6320 8756 6952
rect 8907 6943 8949 6952
rect 8908 6572 8948 6943
rect 8908 6532 9044 6572
rect 8812 6488 8852 6499
rect 8812 6413 8852 6448
rect 8811 6404 8853 6413
rect 8811 6364 8812 6404
rect 8852 6364 8853 6404
rect 8811 6355 8853 6364
rect 8660 6280 8756 6320
rect 8620 6271 8660 6280
rect 8619 6068 8661 6077
rect 8619 6028 8620 6068
rect 8660 6028 8661 6068
rect 8619 6019 8661 6028
rect 8428 5597 8468 5608
rect 8523 5648 8565 5657
rect 8523 5608 8524 5648
rect 8564 5608 8565 5648
rect 8523 5599 8565 5608
rect 8332 5188 8468 5228
rect 8235 5144 8277 5153
rect 8235 5104 8236 5144
rect 8276 5104 8277 5144
rect 8235 5095 8277 5104
rect 8236 3632 8276 5095
rect 8332 5060 8372 5069
rect 8332 4901 8372 5020
rect 8331 4892 8373 4901
rect 8331 4852 8332 4892
rect 8372 4852 8373 4892
rect 8331 4843 8373 4852
rect 8428 3968 8468 5188
rect 8236 3583 8276 3592
rect 8332 3928 8468 3968
rect 8524 4962 8564 4971
rect 7948 2575 7988 2584
rect 8139 2624 8181 2633
rect 8139 2584 8140 2624
rect 8180 2584 8181 2624
rect 8139 2575 8181 2584
rect 8332 2540 8372 3928
rect 8427 3800 8469 3809
rect 8427 3760 8428 3800
rect 8468 3760 8469 3800
rect 8427 3751 8469 3760
rect 8428 3548 8468 3751
rect 8524 3716 8564 4922
rect 8620 3893 8660 6019
rect 8907 5984 8949 5993
rect 8907 5944 8908 5984
rect 8948 5944 8949 5984
rect 8907 5935 8949 5944
rect 8908 5732 8948 5935
rect 8908 5683 8948 5692
rect 9004 5732 9044 6532
rect 9196 6497 9236 7708
rect 9579 7708 9580 7748
rect 9620 7708 9621 7748
rect 9579 7699 9621 7708
rect 9387 7580 9429 7589
rect 9387 7540 9388 7580
rect 9428 7540 9429 7580
rect 9387 7531 9429 7540
rect 9195 6488 9237 6497
rect 9195 6448 9196 6488
rect 9236 6448 9237 6488
rect 9195 6439 9237 6448
rect 9004 5683 9044 5692
rect 9388 5648 9428 7531
rect 9483 7412 9525 7421
rect 9483 7372 9484 7412
rect 9524 7372 9525 7412
rect 9483 7363 9525 7372
rect 9484 7244 9524 7363
rect 9580 7337 9620 7699
rect 9579 7328 9621 7337
rect 9579 7288 9580 7328
rect 9620 7288 9621 7328
rect 9579 7279 9621 7288
rect 9484 7195 9524 7204
rect 9580 7244 9620 7279
rect 9580 7193 9620 7204
rect 9676 6665 9716 7876
rect 9772 7867 9812 7876
rect 9868 7832 9908 9211
rect 9963 8672 10005 8681
rect 9963 8632 9964 8672
rect 10004 8632 10005 8672
rect 9963 8623 10005 8632
rect 9964 8588 10004 8623
rect 9964 8537 10004 8548
rect 9963 8336 10005 8345
rect 9963 8296 9964 8336
rect 10004 8296 10005 8336
rect 9963 8287 10005 8296
rect 9964 7916 10004 8287
rect 10060 8000 10100 9220
rect 10156 9101 10196 9472
rect 10252 9472 10257 9512
rect 10252 9463 10297 9472
rect 10155 9092 10197 9101
rect 10155 9052 10156 9092
rect 10196 9052 10197 9092
rect 10155 9043 10197 9052
rect 10156 8924 10196 8933
rect 10252 8924 10292 9463
rect 10348 9269 10388 10312
rect 10347 9260 10389 9269
rect 10347 9220 10348 9260
rect 10388 9220 10389 9260
rect 10347 9211 10389 9220
rect 10347 9092 10389 9101
rect 10347 9052 10348 9092
rect 10388 9052 10389 9092
rect 10347 9043 10389 9052
rect 10348 8933 10388 9043
rect 10196 8884 10292 8924
rect 10347 8924 10389 8933
rect 10347 8884 10348 8924
rect 10388 8884 10389 8924
rect 10156 8875 10196 8884
rect 10347 8875 10389 8884
rect 10444 8672 10484 10891
rect 10540 10352 10580 13159
rect 10636 12704 10676 12713
rect 11116 12704 11156 13168
rect 10676 12664 11156 12704
rect 11212 13208 11252 13217
rect 11308 13208 11348 14176
rect 11252 13168 11348 13208
rect 10636 12655 10676 12664
rect 11212 12620 11252 13168
rect 11308 12982 11348 12991
rect 11308 12881 11348 12942
rect 11307 12872 11349 12881
rect 11307 12832 11308 12872
rect 11348 12832 11349 12872
rect 11307 12823 11349 12832
rect 11404 12704 11444 14251
rect 11883 14216 11925 14225
rect 11883 14176 11884 14216
rect 11924 14176 11925 14216
rect 11883 14167 11925 14176
rect 11787 14132 11829 14141
rect 11787 14092 11788 14132
rect 11828 14092 11829 14132
rect 11787 14083 11829 14092
rect 11499 14048 11541 14057
rect 11692 14048 11732 14057
rect 11499 14008 11500 14048
rect 11540 14008 11541 14048
rect 11499 13999 11541 14008
rect 11596 14008 11692 14048
rect 11500 13880 11540 13999
rect 11596 13889 11636 14008
rect 11692 13999 11732 14008
rect 11788 13998 11828 14083
rect 11884 14048 11924 14167
rect 11884 13999 11924 14008
rect 11979 14048 12021 14057
rect 11979 14008 11980 14048
rect 12020 14008 12021 14048
rect 11979 13999 12021 14008
rect 12172 14048 12212 15679
rect 12267 15308 12309 15317
rect 12267 15268 12268 15308
rect 12308 15268 12309 15308
rect 12267 15259 12309 15268
rect 12268 14216 12308 15259
rect 12364 14309 12404 16771
rect 12363 14300 12405 14309
rect 12363 14260 12364 14300
rect 12404 14260 12405 14300
rect 12363 14251 12405 14260
rect 12268 14167 12308 14176
rect 12172 13999 12212 14008
rect 12363 14048 12405 14057
rect 12363 14008 12364 14048
rect 12404 14008 12405 14048
rect 12363 13999 12405 14008
rect 11980 13914 12020 13999
rect 12364 13914 12404 13999
rect 11500 13831 11540 13840
rect 11595 13880 11637 13889
rect 11595 13840 11596 13880
rect 11636 13840 11637 13880
rect 11595 13831 11637 13840
rect 12460 13721 12500 17200
rect 12651 17200 12652 17240
rect 12692 17200 12693 17240
rect 12651 17191 12693 17200
rect 12652 17072 12692 17191
rect 12652 17023 12692 17032
rect 12555 16988 12597 16997
rect 12555 16948 12556 16988
rect 12596 16948 12597 16988
rect 12555 16939 12597 16948
rect 12556 14477 12596 16939
rect 12748 14729 12788 17368
rect 12844 17240 12884 17249
rect 13420 17240 13460 17947
rect 12884 17200 13460 17240
rect 12844 17191 12884 17200
rect 13420 17072 13460 17200
rect 13420 17023 13460 17032
rect 12939 16736 12981 16745
rect 12939 16696 12940 16736
rect 12980 16696 12981 16736
rect 12939 16687 12981 16696
rect 12843 16652 12885 16661
rect 12843 16612 12844 16652
rect 12884 16612 12885 16652
rect 12843 16603 12885 16612
rect 12844 16232 12884 16603
rect 12747 14720 12789 14729
rect 12747 14680 12748 14720
rect 12788 14680 12789 14720
rect 12747 14671 12789 14680
rect 12844 14720 12884 16192
rect 12844 14645 12884 14680
rect 12843 14636 12885 14645
rect 12843 14596 12844 14636
rect 12884 14596 12885 14636
rect 12843 14587 12885 14596
rect 12651 14552 12693 14561
rect 12651 14512 12652 14552
rect 12692 14512 12693 14552
rect 12651 14503 12693 14512
rect 12555 14468 12597 14477
rect 12555 14428 12556 14468
rect 12596 14428 12597 14468
rect 12555 14419 12597 14428
rect 12555 14300 12597 14309
rect 12555 14260 12556 14300
rect 12596 14260 12597 14300
rect 12555 14251 12597 14260
rect 12556 14048 12596 14251
rect 12556 13999 12596 14008
rect 12652 14048 12692 14503
rect 12843 14300 12885 14309
rect 12843 14260 12844 14300
rect 12884 14260 12885 14300
rect 12843 14251 12885 14260
rect 12844 14216 12884 14251
rect 12844 14165 12884 14176
rect 12940 14141 12980 16687
rect 13516 16400 13556 18712
rect 13612 18509 13652 19627
rect 13611 18500 13653 18509
rect 13611 18460 13612 18500
rect 13652 18460 13653 18500
rect 13611 18451 13653 18460
rect 13611 18332 13653 18341
rect 13611 18292 13612 18332
rect 13652 18292 13653 18332
rect 13611 18283 13653 18292
rect 13612 17660 13652 18283
rect 13708 18173 13748 20803
rect 13707 18164 13749 18173
rect 13707 18124 13708 18164
rect 13748 18124 13749 18164
rect 13707 18115 13749 18124
rect 13708 17744 13748 17755
rect 13708 17669 13748 17704
rect 13612 17501 13652 17620
rect 13707 17660 13749 17669
rect 13707 17620 13708 17660
rect 13748 17620 13749 17660
rect 13707 17611 13749 17620
rect 13611 17492 13653 17501
rect 13611 17452 13612 17492
rect 13652 17452 13653 17492
rect 13611 17443 13653 17452
rect 13804 17240 13844 21064
rect 13612 17200 13844 17240
rect 13612 16484 13652 17200
rect 13900 17165 13940 21400
rect 13995 21272 14037 21281
rect 13995 21232 13996 21272
rect 14036 21232 14037 21272
rect 13995 21223 14037 21232
rect 13996 20273 14036 21223
rect 14092 20768 14132 20777
rect 14092 20525 14132 20728
rect 14091 20516 14133 20525
rect 14091 20476 14092 20516
rect 14132 20476 14133 20516
rect 14091 20467 14133 20476
rect 13995 20264 14037 20273
rect 13995 20224 13996 20264
rect 14036 20224 14037 20264
rect 13995 20215 14037 20224
rect 14092 20096 14132 20467
rect 14092 20047 14132 20056
rect 13995 20012 14037 20021
rect 13995 19972 13996 20012
rect 14036 19972 14037 20012
rect 13995 19963 14037 19972
rect 13996 19349 14036 19963
rect 13995 19340 14037 19349
rect 13995 19300 13996 19340
rect 14036 19300 14037 19340
rect 13995 19291 14037 19300
rect 14188 19004 14228 22147
rect 14284 22146 14324 22231
rect 14283 21776 14325 21785
rect 14283 21736 14284 21776
rect 14324 21736 14325 21776
rect 14283 21727 14325 21736
rect 14284 21197 14324 21727
rect 14283 21188 14325 21197
rect 14283 21148 14284 21188
rect 14324 21148 14325 21188
rect 14283 21139 14325 21148
rect 14284 20861 14324 21139
rect 14283 20852 14325 20861
rect 14283 20812 14284 20852
rect 14324 20812 14325 20852
rect 14283 20803 14325 20812
rect 14380 20180 14420 22240
rect 14284 20140 14420 20180
rect 14284 19517 14324 20140
rect 14283 19508 14325 19517
rect 14283 19468 14284 19508
rect 14324 19468 14325 19508
rect 14283 19459 14325 19468
rect 14092 18964 14228 19004
rect 13995 18836 14037 18845
rect 13995 18796 13996 18836
rect 14036 18796 14037 18836
rect 13995 18787 14037 18796
rect 13996 18005 14036 18787
rect 13995 17996 14037 18005
rect 13995 17956 13996 17996
rect 14036 17956 14037 17996
rect 13995 17947 14037 17956
rect 13996 17744 14036 17947
rect 13996 17695 14036 17704
rect 13899 17156 13941 17165
rect 13899 17116 13900 17156
rect 13940 17116 13941 17156
rect 13899 17107 13941 17116
rect 13708 17072 13748 17081
rect 13708 16661 13748 17032
rect 13804 17072 13844 17081
rect 13707 16652 13749 16661
rect 13707 16612 13708 16652
rect 13748 16612 13749 16652
rect 13707 16603 13749 16612
rect 13804 16568 13844 17032
rect 13900 16913 13940 17107
rect 14092 17072 14132 18964
rect 14476 18920 14516 24088
rect 14572 23876 14612 23885
rect 14572 22793 14612 23836
rect 14571 22784 14613 22793
rect 14571 22744 14572 22784
rect 14612 22744 14613 22784
rect 14571 22735 14613 22744
rect 14668 21281 14708 24676
rect 14956 24666 14996 24751
rect 15147 24632 15189 24641
rect 15147 24592 15148 24632
rect 15188 24592 15189 24632
rect 15147 24583 15189 24592
rect 14764 24548 14804 24559
rect 14764 24473 14804 24508
rect 15148 24498 15188 24583
rect 14763 24464 14805 24473
rect 14763 24424 14764 24464
rect 14804 24424 14805 24464
rect 14763 24415 14805 24424
rect 14763 23960 14805 23969
rect 14763 23920 14764 23960
rect 14804 23920 14805 23960
rect 14763 23911 14805 23920
rect 14764 23826 14804 23911
rect 14859 23792 14901 23801
rect 14859 23752 14860 23792
rect 14900 23752 14901 23792
rect 14859 23743 14901 23752
rect 15052 23792 15092 23801
rect 14763 23456 14805 23465
rect 14763 23416 14764 23456
rect 14804 23416 14805 23456
rect 14763 23407 14805 23416
rect 14764 23120 14804 23407
rect 14764 21869 14804 23080
rect 14860 22280 14900 23743
rect 14956 23288 14996 23297
rect 15052 23288 15092 23752
rect 15148 23792 15188 23801
rect 15148 23549 15188 23752
rect 15147 23540 15189 23549
rect 15147 23500 15148 23540
rect 15188 23500 15189 23540
rect 15147 23491 15189 23500
rect 15244 23288 15284 25507
rect 15436 25472 15476 27196
rect 15531 27068 15573 27077
rect 15531 27028 15532 27068
rect 15572 27028 15573 27068
rect 15531 27019 15573 27028
rect 15532 26934 15572 27019
rect 14996 23248 15092 23288
rect 15148 23248 15284 23288
rect 15340 25432 15476 25472
rect 14956 23239 14996 23248
rect 15051 22532 15093 22541
rect 15051 22492 15052 22532
rect 15092 22492 15093 22532
rect 15051 22483 15093 22492
rect 14860 22231 14900 22240
rect 14763 21860 14805 21869
rect 14763 21820 14764 21860
rect 14804 21820 14805 21860
rect 14763 21811 14805 21820
rect 14764 21533 14804 21811
rect 14763 21524 14805 21533
rect 14763 21484 14764 21524
rect 14804 21484 14805 21524
rect 14763 21475 14805 21484
rect 14667 21272 14709 21281
rect 14667 21232 14668 21272
rect 14708 21232 14709 21272
rect 14667 21223 14709 21232
rect 14620 20777 14660 20786
rect 14660 20737 14900 20768
rect 14620 20728 14900 20737
rect 14763 20600 14805 20609
rect 14763 20560 14764 20600
rect 14804 20560 14805 20600
rect 14763 20551 14805 20560
rect 14764 20466 14804 20551
rect 14764 20189 14804 20274
rect 14763 20180 14805 20189
rect 14763 20140 14764 20180
rect 14804 20140 14805 20180
rect 14763 20131 14805 20140
rect 14620 20054 14660 20063
rect 14620 20012 14660 20014
rect 14620 19972 14708 20012
rect 14571 19256 14613 19265
rect 14571 19216 14572 19256
rect 14612 19216 14613 19256
rect 14571 19207 14613 19216
rect 14572 19122 14612 19207
rect 14668 19172 14708 19972
rect 14764 19508 14804 19517
rect 14860 19508 14900 20728
rect 15052 20273 15092 22483
rect 15148 21776 15188 23248
rect 15244 23120 15284 23131
rect 15244 23045 15284 23080
rect 15243 23036 15285 23045
rect 15243 22996 15244 23036
rect 15284 22996 15285 23036
rect 15243 22987 15285 22996
rect 15340 22616 15380 25432
rect 15532 25388 15572 25397
rect 15628 25388 15668 28867
rect 15724 28328 15764 31471
rect 15915 31352 15957 31361
rect 15915 31312 15916 31352
rect 15956 31312 15957 31352
rect 15915 31303 15957 31312
rect 15819 31268 15861 31277
rect 15819 31228 15820 31268
rect 15860 31228 15861 31268
rect 15819 31219 15861 31228
rect 15820 30773 15860 31219
rect 15819 30764 15861 30773
rect 15819 30724 15820 30764
rect 15860 30724 15861 30764
rect 15819 30715 15861 30724
rect 15820 30512 15860 30715
rect 15916 30675 15956 31303
rect 16012 30680 16052 32311
rect 16204 32192 16244 32201
rect 16300 32192 16340 32563
rect 16396 32537 16436 32824
rect 16588 32621 16628 35932
rect 16972 35888 17012 36091
rect 16876 35804 16916 35815
rect 16876 35729 16916 35764
rect 16875 35720 16917 35729
rect 16875 35680 16876 35720
rect 16916 35680 16917 35720
rect 16875 35671 16917 35680
rect 16972 35552 17012 35848
rect 17260 35888 17300 36511
rect 17260 35839 17300 35848
rect 16684 35512 17012 35552
rect 16684 35225 16724 35512
rect 17356 35468 17396 36604
rect 16780 35428 17396 35468
rect 16683 35216 16725 35225
rect 16683 35176 16684 35216
rect 16724 35176 16725 35216
rect 16683 35167 16725 35176
rect 16684 34376 16724 34387
rect 16684 34301 16724 34336
rect 16683 34292 16725 34301
rect 16683 34252 16684 34292
rect 16724 34252 16725 34292
rect 16683 34243 16725 34252
rect 16780 32873 16820 35428
rect 17452 35384 17492 36688
rect 17740 36644 17780 37276
rect 18028 37267 18068 37276
rect 18123 37316 18165 37325
rect 18123 37276 18124 37316
rect 18164 37276 18165 37316
rect 18123 37267 18165 37276
rect 18124 37148 18164 37267
rect 17932 37108 18164 37148
rect 17835 36980 17877 36989
rect 17835 36940 17836 36980
rect 17876 36940 17877 36980
rect 17835 36931 17877 36940
rect 17644 36604 17780 36644
rect 17836 36728 17876 36931
rect 17644 35729 17684 36604
rect 17836 36392 17876 36688
rect 17932 36728 17972 37108
rect 18219 37064 18261 37073
rect 18219 37024 18220 37064
rect 18260 37024 18261 37064
rect 18219 37015 18261 37024
rect 18124 36905 18164 36990
rect 18123 36896 18165 36905
rect 18123 36856 18124 36896
rect 18164 36856 18165 36896
rect 18123 36847 18165 36856
rect 18027 36812 18069 36821
rect 18027 36772 18028 36812
rect 18068 36772 18069 36812
rect 18027 36763 18069 36772
rect 17932 36679 17972 36688
rect 18028 36714 18068 36763
rect 18124 36728 18164 36737
rect 18028 36688 18124 36714
rect 18028 36674 18164 36688
rect 17836 36352 17972 36392
rect 17740 35888 17780 35897
rect 17643 35720 17685 35729
rect 17643 35680 17644 35720
rect 17684 35680 17685 35720
rect 17643 35671 17685 35680
rect 17356 35344 17492 35384
rect 17163 35300 17205 35309
rect 17163 35260 17164 35300
rect 17204 35260 17205 35300
rect 17163 35251 17205 35260
rect 16972 35216 17012 35225
rect 16972 34301 17012 35176
rect 17164 35166 17204 35251
rect 17067 34796 17109 34805
rect 17067 34756 17068 34796
rect 17108 34756 17109 34796
rect 17067 34747 17109 34756
rect 17068 34376 17108 34747
rect 17068 34327 17108 34336
rect 16971 34292 17013 34301
rect 16971 34252 16972 34292
rect 17012 34252 17013 34292
rect 16971 34243 17013 34252
rect 17163 34292 17205 34301
rect 17163 34252 17164 34292
rect 17204 34252 17205 34292
rect 17163 34243 17205 34252
rect 16875 34208 16917 34217
rect 16875 34168 16876 34208
rect 16916 34168 16917 34208
rect 16875 34159 16917 34168
rect 16876 34074 16916 34159
rect 16876 33704 16916 33713
rect 17164 33704 17204 34243
rect 16916 33664 17204 33704
rect 16876 33655 16916 33664
rect 17068 33452 17108 33461
rect 16972 33412 17068 33452
rect 16875 33032 16917 33041
rect 16875 32992 16876 33032
rect 16916 32992 16917 33032
rect 16875 32983 16917 32992
rect 16779 32864 16821 32873
rect 16779 32824 16780 32864
rect 16820 32824 16821 32864
rect 16779 32815 16821 32824
rect 16683 32780 16725 32789
rect 16683 32740 16684 32780
rect 16724 32740 16725 32780
rect 16683 32731 16725 32740
rect 16587 32612 16629 32621
rect 16587 32572 16588 32612
rect 16628 32572 16629 32612
rect 16587 32563 16629 32572
rect 16395 32528 16437 32537
rect 16395 32488 16396 32528
rect 16436 32488 16437 32528
rect 16395 32479 16437 32488
rect 16244 32152 16340 32192
rect 16204 32143 16244 32152
rect 16395 32108 16437 32117
rect 16300 32068 16396 32108
rect 16436 32068 16437 32108
rect 16300 31688 16340 32068
rect 16395 32059 16437 32068
rect 16684 31772 16724 32731
rect 16684 31732 16820 31772
rect 16204 31648 16340 31688
rect 16108 31352 16148 31363
rect 16108 31277 16148 31312
rect 16107 31268 16149 31277
rect 16107 31228 16108 31268
rect 16148 31228 16149 31268
rect 16107 31219 16149 31228
rect 16108 30848 16148 30857
rect 16204 30848 16244 31648
rect 16683 31604 16725 31613
rect 16683 31564 16684 31604
rect 16724 31564 16725 31604
rect 16683 31555 16725 31564
rect 16299 31520 16341 31529
rect 16299 31480 16300 31520
rect 16340 31480 16341 31520
rect 16299 31471 16341 31480
rect 16300 31386 16340 31471
rect 16684 31394 16724 31555
rect 16491 31352 16533 31361
rect 16491 31312 16492 31352
rect 16532 31312 16533 31352
rect 16491 31303 16533 31312
rect 16588 31352 16628 31361
rect 16780 31361 16820 31732
rect 16684 31345 16724 31354
rect 16779 31352 16821 31361
rect 16492 31218 16532 31303
rect 16148 30808 16244 30848
rect 16108 30799 16148 30808
rect 16300 30680 16340 30689
rect 16012 30640 16300 30680
rect 15916 30596 15956 30635
rect 15916 30556 16244 30596
rect 15820 30472 16052 30512
rect 15915 30092 15957 30101
rect 15915 30052 15916 30092
rect 15956 30052 15957 30092
rect 15915 30043 15957 30052
rect 15916 29597 15956 30043
rect 16012 29840 16052 30472
rect 16107 30428 16149 30437
rect 16107 30388 16108 30428
rect 16148 30388 16149 30428
rect 16107 30379 16149 30388
rect 15915 29588 15957 29597
rect 15915 29548 15916 29588
rect 15956 29548 15957 29588
rect 15915 29539 15957 29548
rect 15819 29252 15861 29261
rect 15819 29212 15820 29252
rect 15860 29212 15861 29252
rect 15819 29203 15861 29212
rect 15820 29168 15860 29203
rect 15820 29117 15860 29128
rect 15724 27077 15764 28288
rect 15820 28328 15860 28339
rect 15820 28253 15860 28288
rect 15819 28244 15861 28253
rect 15819 28204 15820 28244
rect 15860 28204 15861 28244
rect 15819 28195 15861 28204
rect 15723 27068 15765 27077
rect 15916 27068 15956 29539
rect 16012 29177 16052 29800
rect 16011 29168 16053 29177
rect 16011 29128 16012 29168
rect 16052 29128 16053 29168
rect 16011 29119 16053 29128
rect 16108 29000 16148 30379
rect 16204 30092 16244 30556
rect 16204 30043 16244 30052
rect 16300 29000 16340 30640
rect 16588 30512 16628 31312
rect 16779 31312 16780 31352
rect 16820 31312 16821 31352
rect 16876 31352 16916 32983
rect 16972 32864 17012 33412
rect 17068 33403 17108 33412
rect 17067 33116 17109 33125
rect 17067 33076 17068 33116
rect 17108 33076 17109 33116
rect 17067 33067 17109 33076
rect 16972 32815 17012 32824
rect 17068 32864 17108 33067
rect 17068 32815 17108 32824
rect 16971 32444 17013 32453
rect 16971 32404 16972 32444
rect 17012 32404 17013 32444
rect 16971 32395 17013 32404
rect 16972 31949 17012 32395
rect 17067 32192 17109 32201
rect 17067 32152 17068 32192
rect 17108 32152 17109 32192
rect 17067 32143 17109 32152
rect 17164 32192 17204 33664
rect 17356 33545 17396 35344
rect 17451 35216 17493 35225
rect 17451 35176 17452 35216
rect 17492 35176 17493 35216
rect 17451 35167 17493 35176
rect 17548 35216 17588 35225
rect 17452 35082 17492 35167
rect 17548 34385 17588 35176
rect 17547 34376 17589 34385
rect 17547 34336 17548 34376
rect 17588 34336 17589 34376
rect 17547 34327 17589 34336
rect 17547 34208 17589 34217
rect 17547 34168 17548 34208
rect 17588 34168 17589 34208
rect 17547 34159 17589 34168
rect 17548 33704 17588 34159
rect 17644 33965 17684 35671
rect 17643 33956 17685 33965
rect 17643 33916 17644 33956
rect 17684 33916 17685 33956
rect 17643 33907 17685 33916
rect 17548 33655 17588 33664
rect 17643 33704 17685 33713
rect 17643 33664 17644 33704
rect 17684 33664 17685 33704
rect 17643 33655 17685 33664
rect 17644 33570 17684 33655
rect 17355 33536 17397 33545
rect 17355 33496 17356 33536
rect 17396 33496 17397 33536
rect 17355 33487 17397 33496
rect 17547 33536 17589 33545
rect 17547 33496 17548 33536
rect 17588 33496 17589 33536
rect 17547 33487 17589 33496
rect 17452 32864 17492 32873
rect 17452 32621 17492 32824
rect 17548 32864 17588 33487
rect 17740 33293 17780 35848
rect 17932 35561 17972 36352
rect 17931 35552 17973 35561
rect 17931 35512 17932 35552
rect 17972 35512 17973 35552
rect 17931 35503 17973 35512
rect 17932 35132 17972 35141
rect 17932 34469 17972 35092
rect 18028 35132 18068 35141
rect 17931 34460 17973 34469
rect 17931 34420 17932 34460
rect 17972 34420 17973 34460
rect 17931 34411 17973 34420
rect 17932 33788 17972 34411
rect 18028 34133 18068 35092
rect 18027 34124 18069 34133
rect 18027 34084 18028 34124
rect 18068 34084 18069 34124
rect 18027 34075 18069 34084
rect 17932 33748 18164 33788
rect 18028 33620 18068 33631
rect 18028 33545 18068 33580
rect 18124 33620 18164 33748
rect 18027 33536 18069 33545
rect 18027 33496 18028 33536
rect 18068 33496 18069 33536
rect 18027 33487 18069 33496
rect 17739 33284 17781 33293
rect 17739 33244 17740 33284
rect 17780 33244 17781 33284
rect 17739 33235 17781 33244
rect 18124 33032 18164 33580
rect 17451 32612 17493 32621
rect 17451 32572 17452 32612
rect 17492 32572 17493 32612
rect 17451 32563 17493 32572
rect 17548 32453 17588 32824
rect 17740 32992 18164 33032
rect 17547 32444 17589 32453
rect 17547 32404 17548 32444
rect 17588 32404 17589 32444
rect 17547 32395 17589 32404
rect 17164 32171 17492 32192
rect 17164 32152 17452 32171
rect 16971 31940 17013 31949
rect 16971 31900 16972 31940
rect 17012 31900 17013 31940
rect 17068 31940 17108 32143
rect 17164 32024 17204 32152
rect 17452 32122 17492 32131
rect 17164 31984 17396 32024
rect 17068 31900 17300 31940
rect 16971 31891 17013 31900
rect 17067 31772 17109 31781
rect 17067 31732 17068 31772
rect 17108 31732 17109 31772
rect 17067 31723 17109 31732
rect 17068 31604 17108 31723
rect 17068 31555 17108 31564
rect 16972 31352 17012 31361
rect 16876 31312 16972 31352
rect 16779 31303 16821 31312
rect 16972 31303 17012 31312
rect 17164 31339 17204 31348
rect 16683 31268 16725 31277
rect 16683 31228 16684 31268
rect 16724 31228 16725 31268
rect 16683 31219 16725 31228
rect 16396 30472 16628 30512
rect 16396 30092 16436 30472
rect 16684 30260 16724 31219
rect 16780 31184 16820 31193
rect 16820 31144 17012 31184
rect 16780 31135 16820 31144
rect 16684 30220 16820 30260
rect 16396 30043 16436 30052
rect 16683 30092 16725 30101
rect 16683 30052 16684 30092
rect 16724 30052 16725 30092
rect 16683 30043 16725 30052
rect 16396 29840 16436 29849
rect 16396 29345 16436 29800
rect 16587 29840 16629 29849
rect 16587 29800 16588 29840
rect 16628 29800 16629 29840
rect 16587 29791 16629 29800
rect 16684 29840 16724 30043
rect 16684 29791 16724 29800
rect 16588 29706 16628 29791
rect 16780 29668 16820 30220
rect 16875 29924 16917 29933
rect 16875 29884 16876 29924
rect 16916 29884 16917 29924
rect 16875 29875 16917 29884
rect 16876 29840 16916 29875
rect 16972 29840 17012 31144
rect 17164 31025 17204 31299
rect 17163 31016 17205 31025
rect 17163 30976 17164 31016
rect 17204 30976 17205 31016
rect 17163 30967 17205 30976
rect 17068 30092 17108 30101
rect 17260 30092 17300 31900
rect 17356 30605 17396 31984
rect 17451 31940 17493 31949
rect 17620 31940 17684 32024
rect 17451 31900 17452 31940
rect 17492 31900 17493 31940
rect 17451 31891 17493 31900
rect 17548 31900 17644 31940
rect 17740 31940 17780 32992
rect 18220 32948 18260 37015
rect 18412 36905 18452 37855
rect 18508 37652 18548 37864
rect 19276 37829 19316 38116
rect 19372 38106 19412 38191
rect 19563 38156 19605 38165
rect 19563 38116 19564 38156
rect 19604 38116 19605 38156
rect 19563 38107 19605 38116
rect 19564 38022 19604 38107
rect 19756 37988 19796 37997
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 19275 37820 19317 37829
rect 19275 37780 19276 37820
rect 19316 37780 19317 37820
rect 19275 37771 19317 37780
rect 19756 37661 19796 37948
rect 18508 37603 18548 37612
rect 19755 37652 19797 37661
rect 19755 37612 19756 37652
rect 19796 37612 19797 37652
rect 19755 37603 19797 37612
rect 19179 37568 19221 37577
rect 19179 37528 19180 37568
rect 19220 37528 19221 37568
rect 19179 37519 19221 37528
rect 18892 37400 18932 37409
rect 18796 37316 18836 37325
rect 18411 36896 18453 36905
rect 18411 36856 18412 36896
rect 18452 36856 18453 36896
rect 18411 36847 18453 36856
rect 18796 36812 18836 37276
rect 18892 37241 18932 37360
rect 19180 37400 19220 37519
rect 19756 37484 19796 37493
rect 18891 37232 18933 37241
rect 18891 37192 18892 37232
rect 18932 37192 18933 37232
rect 18891 37183 18933 37192
rect 19083 37064 19125 37073
rect 19083 37024 19084 37064
rect 19124 37024 19125 37064
rect 19083 37015 19125 37024
rect 18604 36772 18836 36812
rect 18316 36728 18356 36737
rect 18316 36569 18356 36688
rect 18507 36728 18549 36737
rect 18507 36688 18508 36728
rect 18548 36688 18549 36728
rect 18507 36679 18549 36688
rect 18411 36644 18453 36653
rect 18411 36604 18412 36644
rect 18452 36604 18453 36644
rect 18411 36595 18453 36604
rect 18315 36560 18357 36569
rect 18315 36520 18316 36560
rect 18356 36520 18357 36560
rect 18315 36511 18357 36520
rect 18412 36510 18452 36595
rect 18508 36594 18548 36679
rect 18604 36317 18644 36772
rect 18700 36644 18740 36653
rect 18700 36485 18740 36604
rect 19084 36644 19124 37015
rect 19180 36821 19220 37360
rect 19467 37400 19509 37409
rect 19467 37360 19468 37400
rect 19508 37360 19509 37400
rect 19467 37351 19509 37360
rect 19659 37400 19701 37409
rect 19659 37360 19660 37400
rect 19700 37360 19701 37400
rect 19659 37351 19701 37360
rect 19468 37266 19508 37351
rect 19564 37232 19604 37241
rect 19275 36896 19317 36905
rect 19275 36856 19276 36896
rect 19316 36856 19317 36896
rect 19275 36847 19317 36856
rect 19179 36812 19221 36821
rect 19179 36772 19180 36812
rect 19220 36772 19221 36812
rect 19179 36763 19221 36772
rect 19276 36762 19316 36847
rect 19564 36737 19604 37192
rect 19660 37073 19700 37351
rect 19659 37064 19701 37073
rect 19659 37024 19660 37064
rect 19700 37024 19701 37064
rect 19659 37015 19701 37024
rect 19563 36728 19605 36737
rect 19563 36688 19564 36728
rect 19604 36688 19605 36728
rect 19563 36679 19605 36688
rect 19084 36595 19124 36604
rect 19467 36644 19509 36653
rect 19467 36604 19468 36644
rect 19508 36604 19509 36644
rect 19467 36595 19509 36604
rect 18891 36560 18933 36569
rect 18891 36520 18892 36560
rect 18932 36520 18933 36560
rect 18891 36511 18933 36520
rect 18699 36476 18741 36485
rect 18699 36436 18700 36476
rect 18740 36436 18741 36476
rect 18699 36427 18741 36436
rect 18892 36426 18932 36511
rect 19468 36510 19508 36595
rect 19660 36476 19700 36485
rect 18603 36308 18645 36317
rect 18603 36268 18604 36308
rect 18644 36268 18645 36308
rect 18603 36259 18645 36268
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 18699 36224 18741 36233
rect 18699 36184 18700 36224
rect 18740 36184 18741 36224
rect 18699 36175 18741 36184
rect 18603 35972 18645 35981
rect 18603 35932 18604 35972
rect 18644 35932 18645 35972
rect 18603 35923 18645 35932
rect 18411 35552 18453 35561
rect 18411 35512 18412 35552
rect 18452 35512 18453 35552
rect 18411 35503 18453 35512
rect 18315 35216 18357 35225
rect 18315 35176 18316 35216
rect 18356 35176 18357 35216
rect 18315 35167 18357 35176
rect 18412 35216 18452 35503
rect 18508 35216 18548 35225
rect 18412 35176 18508 35216
rect 18316 34376 18356 35167
rect 18412 34721 18452 35176
rect 18508 35167 18548 35176
rect 18411 34712 18453 34721
rect 18411 34672 18412 34712
rect 18452 34672 18453 34712
rect 18411 34663 18453 34672
rect 18316 34301 18356 34336
rect 18315 34292 18357 34301
rect 18315 34252 18316 34292
rect 18356 34252 18357 34292
rect 18315 34243 18357 34252
rect 18412 33125 18452 34663
rect 18508 34208 18548 34217
rect 18604 34208 18644 35923
rect 18700 34553 18740 36175
rect 19467 36140 19509 36149
rect 19276 36100 19468 36140
rect 19508 36100 19509 36140
rect 18987 36056 19029 36065
rect 18987 36016 18988 36056
rect 19028 36016 19029 36056
rect 18987 36007 19029 36016
rect 18988 35888 19028 36007
rect 18892 35848 18988 35888
rect 18892 35225 18932 35848
rect 18988 35839 19028 35848
rect 19180 35720 19220 35729
rect 19084 35680 19180 35720
rect 18891 35216 18933 35225
rect 19084 35216 19124 35680
rect 19180 35671 19220 35680
rect 19179 35300 19221 35309
rect 19179 35260 19180 35300
rect 19220 35260 19221 35300
rect 19179 35251 19221 35260
rect 18891 35176 18892 35216
rect 18932 35176 18933 35216
rect 18891 35167 18933 35176
rect 19036 35206 19124 35216
rect 19076 35176 19124 35206
rect 19180 35166 19220 35251
rect 19036 35157 19076 35166
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18699 34544 18741 34553
rect 18699 34504 18700 34544
rect 18740 34504 18741 34544
rect 18699 34495 18741 34504
rect 18700 34376 18740 34495
rect 18700 34327 18740 34336
rect 19083 34208 19125 34217
rect 18604 34168 18740 34208
rect 18411 33116 18453 33125
rect 18411 33076 18412 33116
rect 18452 33076 18453 33116
rect 18411 33067 18453 33076
rect 18220 32908 18452 32948
rect 18028 32864 18068 32873
rect 18068 32824 18356 32864
rect 18028 32815 18068 32824
rect 17931 32360 17973 32369
rect 17931 32320 17932 32360
rect 17972 32320 17973 32360
rect 17931 32311 17973 32320
rect 17835 32192 17877 32201
rect 17835 32152 17836 32192
rect 17876 32152 17877 32192
rect 17835 32143 17877 32152
rect 17836 32058 17876 32143
rect 17740 31900 17876 31940
rect 17355 30596 17397 30605
rect 17355 30556 17356 30596
rect 17396 30556 17397 30596
rect 17355 30547 17397 30556
rect 17452 30512 17492 31891
rect 17548 31352 17588 31900
rect 17644 31891 17684 31900
rect 17548 31303 17588 31312
rect 17644 31352 17684 31361
rect 17547 30764 17589 30773
rect 17547 30724 17548 30764
rect 17588 30724 17589 30764
rect 17547 30715 17589 30724
rect 17548 30680 17588 30715
rect 17548 30629 17588 30640
rect 17452 30472 17588 30512
rect 17355 30428 17397 30437
rect 17355 30388 17356 30428
rect 17396 30388 17397 30428
rect 17355 30379 17397 30388
rect 17108 30052 17300 30092
rect 17068 30043 17108 30052
rect 17163 29924 17205 29933
rect 17163 29884 17164 29924
rect 17204 29884 17205 29924
rect 17163 29875 17205 29884
rect 17068 29840 17108 29849
rect 16972 29800 17068 29840
rect 16876 29789 16916 29800
rect 17068 29791 17108 29800
rect 16780 29628 16916 29668
rect 16395 29336 16437 29345
rect 16395 29296 16396 29336
rect 16436 29296 16437 29336
rect 16395 29287 16437 29296
rect 16587 29168 16629 29177
rect 16587 29128 16588 29168
rect 16628 29128 16629 29168
rect 16587 29119 16629 29128
rect 16108 28960 16244 29000
rect 16300 28960 16436 29000
rect 16107 28580 16149 28589
rect 16107 28540 16108 28580
rect 16148 28540 16149 28580
rect 16107 28531 16149 28540
rect 16108 28253 16148 28531
rect 16107 28244 16149 28253
rect 16107 28204 16108 28244
rect 16148 28204 16149 28244
rect 16107 28195 16149 28204
rect 15723 27028 15724 27068
rect 15764 27028 15765 27068
rect 15723 27019 15765 27028
rect 15820 27028 15956 27068
rect 15724 26816 15764 26825
rect 15820 26816 15860 27028
rect 15915 26900 15957 26909
rect 15915 26860 15916 26900
rect 15956 26860 15957 26900
rect 15915 26851 15957 26860
rect 15764 26776 15860 26816
rect 15724 26767 15764 26776
rect 15723 26648 15765 26657
rect 15723 26608 15724 26648
rect 15764 26608 15765 26648
rect 15723 26599 15765 26608
rect 15572 25348 15668 25388
rect 15532 25339 15572 25348
rect 15436 25304 15476 25315
rect 15436 25229 15476 25264
rect 15435 25220 15477 25229
rect 15435 25180 15436 25220
rect 15476 25180 15477 25220
rect 15435 25171 15477 25180
rect 15436 22793 15476 25171
rect 15724 25136 15764 26599
rect 15532 25096 15764 25136
rect 15532 23876 15572 25096
rect 15627 24548 15669 24557
rect 15627 24508 15628 24548
rect 15668 24508 15669 24548
rect 15627 24499 15669 24508
rect 15532 23827 15572 23836
rect 15628 23792 15668 24499
rect 15723 23876 15765 23885
rect 15723 23836 15724 23876
rect 15764 23836 15765 23876
rect 15723 23827 15765 23836
rect 15628 23204 15668 23752
rect 15532 23164 15668 23204
rect 15435 22784 15477 22793
rect 15435 22744 15436 22784
rect 15476 22744 15477 22784
rect 15435 22735 15477 22744
rect 15532 22709 15572 23164
rect 15627 23036 15669 23045
rect 15627 22996 15628 23036
rect 15668 22996 15669 23036
rect 15627 22987 15669 22996
rect 15531 22700 15573 22709
rect 15531 22660 15532 22700
rect 15572 22660 15573 22700
rect 15531 22651 15573 22660
rect 15340 22576 15476 22616
rect 15340 22285 15380 22294
rect 15340 21776 15380 22245
rect 15148 21736 15284 21776
rect 15148 21608 15188 21619
rect 15148 21533 15188 21568
rect 15147 21524 15189 21533
rect 15147 21484 15148 21524
rect 15188 21484 15189 21524
rect 15147 21475 15189 21484
rect 15244 21020 15284 21736
rect 15340 21727 15380 21736
rect 15340 21020 15380 21029
rect 15244 20980 15340 21020
rect 15340 20971 15380 20980
rect 15148 20852 15188 20861
rect 15188 20812 15284 20852
rect 15148 20803 15188 20812
rect 15051 20264 15093 20273
rect 15051 20224 15052 20264
rect 15092 20224 15093 20264
rect 15051 20215 15093 20224
rect 15244 20189 15284 20812
rect 15436 20432 15476 22576
rect 15531 22196 15573 22205
rect 15531 22156 15532 22196
rect 15572 22156 15573 22196
rect 15531 22147 15573 22156
rect 15532 22062 15572 22147
rect 15531 21692 15573 21701
rect 15531 21652 15532 21692
rect 15572 21652 15573 21692
rect 15531 21643 15573 21652
rect 15532 21608 15572 21643
rect 15532 21557 15572 21568
rect 15531 20768 15573 20777
rect 15531 20728 15532 20768
rect 15572 20728 15573 20768
rect 15531 20719 15573 20728
rect 15532 20634 15572 20719
rect 15628 20609 15668 22987
rect 15724 21113 15764 23827
rect 15820 22373 15860 26776
rect 15916 23213 15956 26851
rect 16108 25724 16148 28195
rect 16204 26405 16244 28960
rect 16299 28328 16341 28337
rect 16299 28288 16300 28328
rect 16340 28288 16341 28328
rect 16299 28279 16341 28288
rect 16300 28194 16340 28279
rect 16299 27068 16341 27077
rect 16299 27028 16300 27068
rect 16340 27028 16341 27068
rect 16299 27019 16341 27028
rect 16203 26396 16245 26405
rect 16203 26356 16204 26396
rect 16244 26356 16245 26396
rect 16203 26347 16245 26356
rect 16204 26144 16244 26347
rect 16204 26095 16244 26104
rect 16108 25684 16244 25724
rect 16011 25640 16053 25649
rect 16011 25600 16012 25640
rect 16052 25600 16053 25640
rect 16011 25591 16053 25600
rect 16012 25304 16052 25591
rect 16012 25255 16052 25264
rect 16108 23792 16148 23801
rect 15915 23204 15957 23213
rect 15915 23164 15916 23204
rect 15956 23164 15957 23204
rect 15915 23155 15957 23164
rect 16108 22961 16148 23752
rect 16204 23717 16244 25684
rect 16203 23708 16245 23717
rect 16203 23668 16204 23708
rect 16244 23668 16245 23708
rect 16203 23659 16245 23668
rect 16107 22952 16149 22961
rect 16107 22912 16108 22952
rect 16148 22912 16149 22952
rect 16107 22903 16149 22912
rect 15915 22868 15957 22877
rect 15915 22828 15916 22868
rect 15956 22828 15957 22868
rect 15915 22819 15957 22828
rect 15819 22364 15861 22373
rect 15819 22324 15820 22364
rect 15860 22324 15861 22364
rect 15819 22315 15861 22324
rect 15916 22280 15956 22819
rect 15916 21953 15956 22240
rect 15915 21944 15957 21953
rect 15915 21904 15916 21944
rect 15956 21904 15957 21944
rect 15915 21895 15957 21904
rect 16204 21365 16244 23659
rect 16203 21356 16245 21365
rect 16203 21316 16204 21356
rect 16244 21316 16245 21356
rect 16203 21307 16245 21316
rect 15723 21104 15765 21113
rect 15723 21064 15724 21104
rect 15764 21064 15765 21104
rect 15723 21055 15765 21064
rect 15724 20936 15764 20945
rect 15764 20896 15860 20936
rect 15724 20887 15764 20896
rect 15724 20768 15764 20777
rect 15627 20600 15669 20609
rect 15627 20560 15628 20600
rect 15668 20560 15669 20600
rect 15627 20551 15669 20560
rect 15340 20392 15476 20432
rect 15243 20180 15285 20189
rect 15243 20140 15244 20180
rect 15284 20140 15285 20180
rect 15243 20131 15285 20140
rect 14956 20096 14996 20105
rect 15148 20096 15188 20105
rect 14996 20056 15092 20096
rect 14956 20047 14996 20056
rect 14804 19468 14900 19508
rect 14764 19459 14804 19468
rect 14956 19265 14996 19350
rect 14955 19256 14997 19265
rect 14955 19216 14956 19256
rect 14996 19216 14997 19256
rect 14955 19207 14997 19216
rect 14668 19132 14900 19172
rect 14763 19004 14805 19013
rect 14763 18964 14764 19004
rect 14804 18964 14805 19004
rect 14763 18955 14805 18964
rect 14188 18880 14516 18920
rect 14188 17996 14228 18880
rect 14764 18626 14804 18955
rect 14860 18752 14900 19132
rect 14955 19088 14997 19097
rect 14955 19048 14956 19088
rect 14996 19048 14997 19088
rect 14955 19039 14997 19048
rect 14860 18703 14900 18712
rect 14956 18626 14996 19039
rect 15052 18845 15092 20056
rect 15148 20012 15188 20056
rect 15148 19972 15284 20012
rect 15147 19844 15189 19853
rect 15147 19804 15148 19844
rect 15188 19804 15189 19844
rect 15147 19795 15189 19804
rect 15148 19710 15188 19795
rect 15147 19424 15189 19433
rect 15147 19384 15148 19424
rect 15188 19384 15189 19424
rect 15147 19375 15189 19384
rect 15051 18836 15093 18845
rect 15051 18796 15052 18836
rect 15092 18796 15093 18836
rect 15051 18787 15093 18796
rect 15052 18626 15092 18635
rect 14283 18584 14325 18593
rect 14283 18544 14284 18584
rect 14324 18544 14325 18584
rect 14283 18535 14325 18544
rect 14667 18584 14709 18593
rect 14764 18586 14900 18626
rect 14667 18544 14668 18584
rect 14708 18544 14709 18584
rect 14667 18535 14709 18544
rect 14178 17956 14228 17996
rect 14178 17660 14218 17956
rect 14284 17786 14324 18535
rect 14668 18450 14708 18535
rect 14475 18248 14517 18257
rect 14475 18208 14476 18248
rect 14516 18208 14517 18248
rect 14475 18199 14517 18208
rect 14476 17954 14516 18199
rect 14379 17912 14421 17921
rect 14379 17872 14380 17912
rect 14420 17872 14421 17912
rect 14763 17996 14805 18005
rect 14763 17956 14764 17996
rect 14804 17956 14805 17996
rect 14763 17947 14805 17956
rect 14476 17905 14516 17914
rect 14379 17870 14421 17872
rect 14379 17863 14380 17870
rect 14420 17863 14421 17870
rect 14572 17837 14612 17922
rect 14380 17777 14420 17830
rect 14571 17828 14613 17837
rect 14764 17828 14804 17947
rect 14571 17788 14572 17828
rect 14612 17788 14613 17828
rect 14571 17779 14613 17788
rect 14668 17788 14804 17828
rect 14668 17786 14708 17788
rect 14284 17737 14324 17746
rect 14668 17737 14708 17746
rect 14860 17744 14900 18586
rect 14956 18586 15052 18626
rect 14956 18509 14996 18586
rect 15052 18577 15092 18586
rect 14955 18500 14997 18509
rect 14955 18460 14956 18500
rect 14996 18460 14997 18500
rect 14955 18451 14997 18460
rect 15051 18332 15093 18341
rect 15051 18292 15052 18332
rect 15092 18292 15093 18332
rect 15051 18283 15093 18292
rect 14475 17660 14517 17669
rect 14178 17620 14228 17660
rect 13996 17032 14132 17072
rect 13899 16904 13941 16913
rect 13899 16864 13900 16904
rect 13940 16864 13941 16904
rect 13899 16855 13941 16864
rect 13804 16528 13940 16568
rect 13612 16444 13748 16484
rect 13420 16360 13556 16400
rect 13036 16064 13076 16073
rect 13036 15569 13076 16024
rect 13420 15821 13460 16360
rect 13515 16232 13557 16241
rect 13515 16192 13516 16232
rect 13556 16192 13557 16232
rect 13515 16183 13557 16192
rect 13516 16098 13556 16183
rect 13419 15812 13461 15821
rect 13419 15772 13420 15812
rect 13460 15772 13461 15812
rect 13419 15763 13461 15772
rect 13323 15728 13365 15737
rect 13708 15728 13748 16444
rect 13803 15812 13845 15821
rect 13803 15772 13804 15812
rect 13844 15772 13845 15812
rect 13803 15763 13845 15772
rect 13323 15688 13324 15728
rect 13364 15688 13365 15728
rect 13323 15679 13365 15688
rect 13516 15688 13748 15728
rect 13131 15644 13173 15653
rect 13131 15604 13132 15644
rect 13172 15604 13173 15644
rect 13131 15595 13173 15604
rect 13035 15560 13077 15569
rect 13035 15520 13036 15560
rect 13076 15520 13077 15560
rect 13035 15511 13077 15520
rect 13132 15233 13172 15595
rect 13228 15560 13268 15569
rect 13131 15224 13173 15233
rect 13131 15184 13132 15224
rect 13172 15184 13173 15224
rect 13131 15175 13173 15184
rect 13228 14888 13268 15520
rect 13324 14972 13364 15679
rect 13419 15644 13461 15653
rect 13419 15604 13420 15644
rect 13460 15604 13461 15644
rect 13419 15595 13461 15604
rect 13420 15510 13460 15595
rect 13324 14923 13364 14932
rect 13132 14848 13268 14888
rect 13132 14729 13172 14848
rect 13131 14720 13173 14729
rect 13131 14680 13132 14720
rect 13172 14680 13173 14720
rect 13131 14671 13173 14680
rect 13228 14720 13268 14729
rect 13035 14552 13077 14561
rect 13228 14552 13268 14680
rect 13035 14512 13036 14552
rect 13076 14512 13268 14552
rect 13035 14503 13077 14512
rect 13036 14418 13076 14503
rect 12939 14132 12981 14141
rect 12939 14092 12940 14132
rect 12980 14092 12981 14132
rect 12939 14083 12981 14092
rect 12652 13999 12692 14008
rect 12843 14048 12885 14057
rect 12843 14008 12844 14048
rect 12884 14008 12885 14048
rect 12843 13999 12885 14008
rect 13036 14048 13076 14057
rect 12844 13914 12884 13999
rect 12555 13880 12597 13889
rect 12555 13840 12556 13880
rect 12596 13840 12597 13880
rect 12555 13831 12597 13840
rect 12459 13712 12501 13721
rect 12459 13672 12460 13712
rect 12500 13672 12501 13712
rect 12459 13663 12501 13672
rect 11787 13460 11829 13469
rect 11787 13420 11788 13460
rect 11828 13420 11829 13460
rect 11787 13411 11829 13420
rect 10924 12580 11252 12620
rect 11308 12664 11444 12704
rect 11500 13208 11540 13217
rect 11500 12704 11540 13168
rect 11692 13208 11732 13217
rect 11595 13040 11637 13049
rect 11595 13000 11596 13040
rect 11636 13000 11637 13040
rect 11595 12991 11637 13000
rect 11596 12906 11636 12991
rect 11692 12788 11732 13168
rect 11788 13208 11828 13411
rect 11788 13159 11828 13168
rect 12076 13208 12116 13217
rect 11979 12872 12021 12881
rect 11979 12832 11980 12872
rect 12020 12832 12021 12872
rect 11979 12823 12021 12832
rect 11692 12748 11924 12788
rect 11500 12664 11828 12704
rect 10731 12536 10773 12545
rect 10731 12496 10732 12536
rect 10772 12496 10773 12536
rect 10731 12487 10773 12496
rect 10828 12536 10868 12547
rect 10732 12402 10772 12487
rect 10828 12461 10868 12496
rect 10924 12536 10964 12580
rect 11308 12536 11348 12664
rect 10924 12487 10964 12496
rect 11212 12491 11252 12500
rect 10827 12452 10869 12461
rect 10827 12412 10828 12452
rect 10868 12412 10869 12452
rect 10827 12403 10869 12412
rect 11019 12452 11061 12461
rect 11019 12412 11020 12452
rect 11060 12412 11061 12452
rect 11019 12403 11061 12412
rect 11211 12412 11212 12461
rect 11252 12412 11253 12461
rect 11211 12403 11253 12412
rect 10923 11780 10965 11789
rect 10923 11740 10924 11780
rect 10964 11740 10965 11780
rect 10923 11731 10965 11740
rect 10731 11696 10773 11705
rect 10731 11656 10732 11696
rect 10772 11656 10773 11696
rect 10731 11647 10773 11656
rect 10732 11024 10772 11647
rect 10732 10865 10772 10984
rect 10731 10856 10773 10865
rect 10731 10816 10732 10856
rect 10772 10816 10773 10856
rect 10731 10807 10773 10816
rect 10540 10312 10772 10352
rect 10539 10184 10581 10193
rect 10539 10144 10540 10184
rect 10580 10144 10581 10184
rect 10539 10135 10581 10144
rect 10540 8840 10580 10135
rect 10636 9605 10676 9636
rect 10635 9596 10677 9605
rect 10635 9556 10636 9596
rect 10676 9556 10677 9596
rect 10635 9547 10677 9556
rect 10636 9512 10676 9547
rect 10636 9101 10676 9472
rect 10635 9092 10677 9101
rect 10635 9052 10636 9092
rect 10676 9052 10677 9092
rect 10635 9043 10677 9052
rect 10540 8800 10676 8840
rect 10636 8681 10676 8800
rect 10444 8597 10484 8632
rect 10540 8672 10580 8681
rect 10155 8588 10197 8597
rect 10155 8548 10156 8588
rect 10196 8548 10197 8588
rect 10155 8539 10197 8548
rect 10443 8588 10485 8597
rect 10443 8548 10444 8588
rect 10484 8548 10485 8588
rect 10443 8539 10485 8548
rect 10156 8261 10196 8539
rect 10444 8508 10484 8539
rect 10540 8345 10580 8632
rect 10635 8672 10677 8681
rect 10635 8632 10636 8672
rect 10676 8632 10677 8672
rect 10635 8623 10677 8632
rect 10539 8336 10581 8345
rect 10539 8296 10540 8336
rect 10580 8296 10581 8336
rect 10539 8287 10581 8296
rect 10155 8252 10197 8261
rect 10155 8212 10156 8252
rect 10196 8212 10197 8252
rect 10155 8203 10197 8212
rect 10060 7951 10100 7960
rect 10443 8000 10485 8009
rect 10443 7960 10444 8000
rect 10484 7960 10485 8000
rect 10443 7951 10485 7960
rect 9964 7867 10004 7876
rect 10444 7866 10484 7951
rect 9868 7783 9908 7792
rect 10059 7664 10101 7673
rect 10059 7624 10060 7664
rect 10100 7624 10101 7664
rect 10059 7615 10101 7624
rect 10060 7160 10100 7615
rect 10155 7496 10197 7505
rect 10155 7456 10156 7496
rect 10196 7456 10197 7496
rect 10155 7447 10197 7456
rect 10060 6917 10100 7120
rect 10059 6908 10101 6917
rect 10059 6868 10060 6908
rect 10100 6868 10101 6908
rect 10059 6859 10101 6868
rect 10156 6833 10196 7447
rect 10540 7337 10580 8287
rect 10539 7328 10581 7337
rect 10539 7288 10540 7328
rect 10580 7288 10581 7328
rect 10539 7279 10581 7288
rect 10732 7244 10772 10312
rect 10924 10268 10964 11731
rect 11020 11117 11060 12403
rect 11212 12356 11252 12403
rect 11308 11957 11348 12496
rect 11404 12536 11444 12545
rect 11307 11948 11349 11957
rect 11307 11908 11308 11948
rect 11348 11908 11349 11948
rect 11307 11899 11349 11908
rect 11404 11948 11444 12496
rect 11500 12536 11540 12545
rect 11692 12536 11732 12545
rect 11540 12496 11692 12536
rect 11500 12487 11540 12496
rect 11692 12487 11732 12496
rect 11692 12284 11732 12293
rect 11595 12116 11637 12125
rect 11595 12076 11596 12116
rect 11636 12076 11637 12116
rect 11595 12067 11637 12076
rect 11499 12032 11541 12041
rect 11499 11992 11500 12032
rect 11540 11992 11541 12032
rect 11499 11983 11541 11992
rect 11404 11899 11444 11908
rect 11212 11696 11252 11707
rect 11212 11621 11252 11656
rect 11211 11612 11253 11621
rect 11211 11572 11212 11612
rect 11252 11572 11253 11612
rect 11211 11563 11253 11572
rect 11403 11528 11445 11537
rect 11403 11488 11404 11528
rect 11444 11488 11445 11528
rect 11403 11479 11445 11488
rect 11404 11394 11444 11479
rect 11211 11276 11253 11285
rect 11211 11236 11212 11276
rect 11252 11236 11253 11276
rect 11211 11227 11253 11236
rect 11019 11108 11061 11117
rect 11019 11068 11020 11108
rect 11060 11068 11061 11108
rect 11019 11059 11061 11068
rect 11020 11024 11060 11059
rect 11020 10974 11060 10984
rect 11116 11024 11156 11033
rect 11116 10856 11156 10984
rect 11020 10816 11156 10856
rect 11020 10361 11060 10816
rect 11212 10772 11252 11227
rect 11307 11192 11349 11201
rect 11307 11152 11308 11192
rect 11348 11152 11349 11192
rect 11307 11143 11349 11152
rect 11308 10781 11348 11143
rect 11500 10949 11540 11983
rect 11596 11705 11636 12067
rect 11595 11696 11637 11705
rect 11595 11656 11596 11696
rect 11636 11656 11637 11696
rect 11595 11647 11637 11656
rect 11596 11562 11636 11647
rect 11499 10940 11541 10949
rect 11499 10900 11500 10940
rect 11540 10900 11541 10940
rect 11499 10891 11541 10900
rect 11596 10940 11636 10951
rect 11500 10806 11540 10891
rect 11596 10865 11636 10900
rect 11595 10856 11637 10865
rect 11595 10816 11596 10856
rect 11636 10816 11637 10856
rect 11595 10807 11637 10816
rect 11116 10732 11252 10772
rect 11307 10772 11349 10781
rect 11307 10732 11308 10772
rect 11348 10732 11349 10772
rect 11019 10352 11061 10361
rect 11019 10312 11020 10352
rect 11060 10312 11061 10352
rect 11019 10303 11061 10312
rect 10924 10219 10964 10228
rect 10828 10184 10868 10193
rect 10828 9773 10868 10144
rect 11019 10184 11061 10193
rect 11019 10144 11020 10184
rect 11060 10144 11061 10184
rect 11019 10135 11061 10144
rect 10923 10100 10965 10109
rect 10923 10060 10924 10100
rect 10964 10060 10965 10100
rect 10923 10051 10965 10060
rect 10924 9932 10964 10051
rect 11020 10050 11060 10135
rect 11116 9932 11156 10732
rect 11307 10723 11349 10732
rect 11692 10697 11732 12244
rect 11788 11201 11828 12664
rect 11884 12536 11924 12748
rect 11884 12461 11924 12496
rect 11980 12536 12020 12823
rect 11883 12452 11925 12461
rect 11883 12412 11884 12452
rect 11924 12412 11925 12452
rect 11883 12403 11925 12412
rect 11980 12293 12020 12496
rect 11979 12284 12021 12293
rect 11979 12244 11980 12284
rect 12020 12244 12021 12284
rect 11979 12235 12021 12244
rect 11979 12032 12021 12041
rect 11979 11992 11980 12032
rect 12020 11992 12021 12032
rect 11979 11983 12021 11992
rect 11980 11621 12020 11983
rect 11979 11612 12021 11621
rect 11979 11572 11980 11612
rect 12020 11572 12021 11612
rect 11979 11563 12021 11572
rect 12076 11537 12116 13168
rect 12172 13208 12212 13217
rect 12172 13049 12212 13168
rect 12267 13208 12309 13217
rect 12267 13168 12268 13208
rect 12308 13168 12309 13208
rect 12267 13159 12309 13168
rect 12556 13208 12596 13831
rect 13036 13805 13076 14008
rect 13035 13796 13077 13805
rect 13035 13756 13036 13796
rect 13076 13756 13077 13796
rect 13035 13747 13077 13756
rect 12651 13712 12693 13721
rect 12651 13672 12652 13712
rect 12692 13672 12693 13712
rect 12651 13663 12693 13672
rect 12556 13159 12596 13168
rect 12268 13074 12308 13159
rect 12171 13040 12213 13049
rect 12171 13000 12172 13040
rect 12212 13000 12213 13040
rect 12171 12991 12213 13000
rect 12364 13040 12404 13049
rect 12652 13040 12692 13663
rect 12844 13208 12884 13217
rect 12171 12872 12213 12881
rect 12364 12872 12404 13000
rect 12171 12832 12172 12872
rect 12212 12832 12404 12872
rect 12556 13000 12692 13040
rect 12748 13124 12788 13133
rect 12171 12823 12213 12832
rect 12556 12704 12596 13000
rect 12364 12664 12596 12704
rect 12172 12629 12212 12660
rect 12171 12620 12213 12629
rect 12171 12580 12172 12620
rect 12212 12580 12213 12620
rect 12171 12571 12213 12580
rect 12172 12536 12212 12571
rect 12172 11621 12212 12496
rect 12171 11612 12213 11621
rect 12171 11572 12172 11612
rect 12212 11572 12213 11612
rect 12171 11563 12213 11572
rect 12075 11528 12117 11537
rect 12075 11488 12076 11528
rect 12116 11488 12117 11528
rect 12075 11479 12117 11488
rect 11787 11192 11829 11201
rect 11787 11152 11788 11192
rect 11828 11152 11829 11192
rect 11787 11143 11829 11152
rect 12075 11192 12117 11201
rect 12075 11152 12076 11192
rect 12116 11152 12117 11192
rect 12075 11143 12117 11152
rect 12076 11024 12116 11143
rect 12076 10975 12116 10984
rect 12364 10865 12404 12664
rect 12748 12545 12788 13084
rect 12844 13049 12884 13168
rect 13035 13208 13077 13217
rect 13035 13168 13036 13208
rect 13076 13168 13077 13208
rect 13035 13159 13077 13168
rect 13132 13208 13172 13217
rect 12843 13040 12885 13049
rect 12843 13000 12844 13040
rect 12884 13000 12885 13040
rect 12843 12991 12885 13000
rect 12939 12872 12981 12881
rect 12939 12832 12940 12872
rect 12980 12832 12981 12872
rect 12939 12823 12981 12832
rect 12747 12536 12789 12545
rect 12747 12496 12748 12536
rect 12788 12496 12789 12536
rect 12747 12487 12789 12496
rect 12651 11948 12693 11957
rect 12651 11908 12652 11948
rect 12692 11908 12693 11948
rect 12651 11899 12693 11908
rect 12843 11948 12885 11957
rect 12843 11908 12844 11948
rect 12884 11908 12885 11948
rect 12843 11899 12885 11908
rect 12555 11528 12597 11537
rect 12555 11488 12556 11528
rect 12596 11488 12597 11528
rect 12555 11479 12597 11488
rect 12556 11019 12596 11479
rect 12556 10970 12596 10979
rect 12363 10856 12405 10865
rect 12363 10816 12364 10856
rect 12404 10816 12405 10856
rect 12363 10807 12405 10816
rect 11691 10688 11733 10697
rect 11691 10648 11692 10688
rect 11732 10648 11733 10688
rect 11691 10639 11733 10648
rect 11307 10520 11349 10529
rect 11307 10480 11308 10520
rect 11348 10480 11349 10520
rect 11307 10471 11349 10480
rect 11979 10520 12021 10529
rect 11979 10480 11980 10520
rect 12020 10480 12021 10520
rect 11979 10471 12021 10480
rect 11308 10268 11348 10471
rect 11403 10352 11445 10361
rect 11403 10312 11404 10352
rect 11444 10312 11445 10352
rect 11403 10303 11445 10312
rect 11980 10352 12020 10471
rect 12363 10436 12405 10445
rect 12363 10396 12364 10436
rect 12404 10396 12405 10436
rect 12363 10387 12405 10396
rect 11980 10303 12020 10312
rect 11308 10219 11348 10228
rect 11404 10218 11444 10303
rect 11500 10268 11540 10277
rect 11212 10184 11252 10193
rect 11212 10100 11252 10144
rect 11212 10060 11444 10100
rect 10924 9892 11348 9932
rect 10827 9764 10869 9773
rect 10827 9724 10828 9764
rect 10868 9724 10869 9764
rect 10827 9715 10869 9724
rect 11019 9680 11061 9689
rect 11019 9640 11020 9680
rect 11060 9640 11061 9680
rect 11019 9631 11061 9640
rect 10827 8672 10869 8681
rect 10827 8632 10828 8672
rect 10868 8632 10869 8672
rect 10827 8623 10869 8632
rect 10828 8538 10868 8623
rect 11020 8177 11060 9631
rect 11115 8672 11157 8681
rect 11115 8632 11116 8672
rect 11156 8632 11157 8672
rect 11115 8623 11157 8632
rect 11212 8672 11252 8681
rect 11116 8538 11156 8623
rect 11019 8168 11061 8177
rect 11019 8128 11020 8168
rect 11060 8128 11061 8168
rect 11019 8119 11061 8128
rect 11020 7916 11060 8119
rect 11212 8093 11252 8632
rect 11211 8084 11253 8093
rect 11211 8044 11212 8084
rect 11252 8044 11253 8084
rect 11211 8035 11253 8044
rect 11020 7876 11252 7916
rect 11116 7244 11156 7253
rect 10732 7204 11116 7244
rect 11116 7195 11156 7204
rect 10540 7165 10580 7174
rect 10155 6824 10197 6833
rect 10155 6784 10156 6824
rect 10196 6784 10197 6824
rect 10155 6775 10197 6784
rect 9675 6656 9717 6665
rect 9675 6616 9676 6656
rect 9716 6616 9717 6656
rect 9675 6607 9717 6616
rect 10060 6488 10100 6497
rect 10156 6488 10196 6775
rect 10540 6740 10580 7125
rect 10635 7076 10677 7085
rect 10635 7036 10636 7076
rect 10676 7036 10677 7076
rect 10635 7027 10677 7036
rect 10252 6700 10580 6740
rect 10252 6656 10292 6700
rect 10252 6607 10292 6616
rect 10443 6488 10485 6497
rect 10156 6448 10444 6488
rect 10484 6448 10485 6488
rect 10060 6245 10100 6448
rect 10443 6439 10485 6448
rect 10444 6354 10484 6439
rect 10059 6236 10101 6245
rect 10059 6196 10060 6236
rect 10100 6196 10101 6236
rect 10059 6187 10101 6196
rect 10155 5984 10197 5993
rect 10347 5984 10389 5993
rect 10155 5944 10156 5984
rect 10196 5944 10348 5984
rect 10388 5944 10389 5984
rect 10155 5935 10197 5944
rect 10347 5935 10389 5944
rect 9867 5900 9909 5909
rect 9867 5860 9868 5900
rect 9908 5860 9909 5900
rect 9867 5851 9909 5860
rect 9868 5816 9908 5851
rect 9868 5765 9908 5776
rect 10060 5732 10100 5741
rect 10100 5692 10196 5732
rect 10060 5683 10100 5692
rect 9388 5599 9428 5608
rect 9484 5648 9524 5657
rect 9484 5321 9524 5608
rect 9772 5480 9812 5489
rect 9483 5312 9525 5321
rect 9483 5272 9484 5312
rect 9524 5272 9525 5312
rect 9483 5263 9525 5272
rect 9675 5228 9717 5237
rect 9675 5188 9676 5228
rect 9716 5188 9717 5228
rect 9675 5179 9717 5188
rect 9387 5144 9429 5153
rect 9387 5104 9388 5144
rect 9428 5104 9429 5144
rect 9387 5095 9429 5104
rect 9003 4976 9045 4985
rect 9003 4936 9004 4976
rect 9044 4936 9045 4976
rect 9003 4927 9045 4936
rect 9004 4842 9044 4927
rect 9195 4892 9237 4901
rect 9195 4852 9196 4892
rect 9236 4852 9237 4892
rect 9195 4843 9237 4852
rect 8907 4304 8949 4313
rect 9100 4304 9140 4313
rect 8907 4264 8908 4304
rect 8948 4264 8949 4304
rect 8907 4255 8949 4264
rect 9004 4264 9100 4304
rect 8908 4136 8948 4255
rect 9004 4145 9044 4264
rect 9100 4255 9140 4264
rect 8908 4087 8948 4096
rect 9003 4136 9045 4145
rect 9003 4096 9004 4136
rect 9044 4096 9045 4136
rect 9003 4087 9045 4096
rect 9196 4052 9236 4843
rect 9291 4640 9333 4649
rect 9291 4600 9292 4640
rect 9332 4600 9333 4640
rect 9291 4591 9333 4600
rect 9292 4304 9332 4591
rect 9292 4255 9332 4264
rect 9100 4012 9236 4052
rect 8619 3884 8661 3893
rect 8619 3844 8620 3884
rect 8660 3844 8661 3884
rect 8619 3835 8661 3844
rect 8524 3676 8660 3716
rect 8524 3548 8564 3557
rect 8428 3508 8524 3548
rect 8620 3548 8660 3676
rect 8620 3508 8852 3548
rect 8524 3499 8564 3508
rect 8668 3422 8708 3431
rect 8668 3380 8708 3382
rect 8524 3340 8708 3380
rect 8428 2717 8468 2733
rect 8427 2708 8469 2717
rect 8427 2668 8428 2708
rect 8468 2668 8469 2708
rect 8427 2659 8469 2668
rect 8428 2638 8468 2659
rect 8428 2589 8468 2598
rect 8524 2540 8564 3340
rect 8812 3296 8852 3508
rect 9003 3380 9045 3389
rect 9003 3340 9004 3380
rect 9044 3340 9045 3380
rect 9003 3331 9045 3340
rect 8716 3256 8852 3296
rect 8716 2708 8756 3256
rect 8800 2708 8852 2719
rect 8716 2668 8948 2708
rect 8620 2549 8660 2634
rect 8716 2598 8769 2668
rect 8236 2500 8372 2540
rect 8428 2500 8564 2540
rect 8619 2540 8661 2549
rect 8720 2540 8762 2549
rect 8619 2500 8620 2540
rect 8660 2500 8661 2540
rect 7851 2456 7893 2465
rect 7851 2416 7852 2456
rect 7892 2416 7893 2456
rect 7851 2407 7893 2416
rect 7659 2204 7701 2213
rect 7659 2164 7660 2204
rect 7700 2164 7701 2204
rect 7659 2155 7701 2164
rect 7852 1961 7892 2407
rect 8236 2120 8276 2500
rect 8332 2120 8372 2129
rect 8236 2080 8332 2120
rect 8332 2071 8372 2080
rect 8140 2036 8180 2045
rect 8044 1996 8140 2036
rect 7851 1952 7893 1961
rect 7851 1912 7852 1952
rect 7892 1912 7893 1952
rect 7851 1903 7893 1912
rect 7948 1938 7988 1947
rect 7755 1280 7797 1289
rect 7755 1240 7756 1280
rect 7796 1240 7797 1280
rect 7755 1231 7797 1240
rect 7660 1112 7700 1121
rect 7564 1072 7660 1112
rect 7276 1063 7316 1072
rect 7660 1063 7700 1072
rect 7371 944 7413 953
rect 7371 904 7372 944
rect 7412 904 7413 944
rect 7371 895 7413 904
rect 7563 944 7605 953
rect 7563 904 7564 944
rect 7604 904 7605 944
rect 7563 895 7605 904
rect 7372 80 7412 895
rect 7564 80 7604 895
rect 7756 80 7796 1231
rect 7948 1028 7988 1898
rect 8044 1037 8084 1996
rect 8140 1987 8180 1996
rect 8235 1364 8277 1373
rect 8235 1324 8236 1364
rect 8276 1324 8277 1364
rect 8235 1315 8277 1324
rect 8139 1280 8181 1289
rect 8139 1240 8140 1280
rect 8180 1240 8181 1280
rect 8139 1231 8181 1240
rect 7852 988 7988 1028
rect 8043 1028 8085 1037
rect 8043 988 8044 1028
rect 8084 988 8085 1028
rect 7852 617 7892 988
rect 8043 979 8085 988
rect 7947 860 7989 869
rect 7947 820 7948 860
rect 7988 820 7989 860
rect 7947 811 7989 820
rect 7851 608 7893 617
rect 7851 568 7852 608
rect 7892 568 7893 608
rect 7851 559 7893 568
rect 7948 80 7988 811
rect 8140 80 8180 1231
rect 8236 1037 8276 1315
rect 8331 1280 8373 1289
rect 8331 1240 8332 1280
rect 8372 1240 8373 1280
rect 8331 1231 8373 1240
rect 8235 1028 8277 1037
rect 8235 988 8236 1028
rect 8276 988 8277 1028
rect 8235 979 8277 988
rect 8332 80 8372 1231
rect 8428 1205 8468 2500
rect 8619 2491 8661 2500
rect 8716 2500 8721 2540
rect 8761 2500 8762 2540
rect 8716 2491 8762 2500
rect 8523 1952 8565 1961
rect 8523 1912 8524 1952
rect 8564 1912 8565 1952
rect 8523 1903 8565 1912
rect 8524 1818 8564 1903
rect 8523 1280 8565 1289
rect 8523 1240 8524 1280
rect 8564 1240 8565 1280
rect 8523 1231 8565 1240
rect 8427 1196 8469 1205
rect 8427 1156 8428 1196
rect 8468 1156 8469 1196
rect 8427 1147 8469 1156
rect 8524 80 8564 1231
rect 8716 80 8756 2491
rect 8812 2456 8852 2465
rect 8812 2213 8852 2416
rect 8811 2204 8853 2213
rect 8811 2164 8812 2204
rect 8852 2164 8853 2204
rect 8811 2155 8853 2164
rect 8811 1448 8853 1457
rect 8811 1408 8812 1448
rect 8852 1408 8853 1448
rect 8811 1399 8853 1408
rect 8812 701 8852 1399
rect 8908 1364 8948 2668
rect 9004 2624 9044 3331
rect 9004 2575 9044 2584
rect 9100 2624 9140 4012
rect 9195 3464 9237 3473
rect 9195 3424 9196 3464
rect 9236 3424 9237 3464
rect 9195 3415 9237 3424
rect 9196 3330 9236 3415
rect 9388 3212 9428 5095
rect 9484 4901 9524 4986
rect 9579 4976 9621 4985
rect 9579 4936 9580 4976
rect 9620 4936 9621 4976
rect 9579 4927 9621 4936
rect 9483 4892 9525 4901
rect 9483 4852 9484 4892
rect 9524 4852 9525 4892
rect 9483 4843 9525 4852
rect 9580 4842 9620 4927
rect 9676 4724 9716 5179
rect 9100 2575 9140 2584
rect 9196 3172 9428 3212
rect 9484 4684 9716 4724
rect 9100 1364 9140 1373
rect 8908 1324 9100 1364
rect 9100 1315 9140 1324
rect 8908 1112 8948 1123
rect 9196 1112 9236 3172
rect 9291 2792 9333 2801
rect 9291 2752 9292 2792
rect 9332 2752 9333 2792
rect 9291 2743 9333 2752
rect 9292 2658 9332 2743
rect 9484 1280 9524 4684
rect 9772 4649 9812 5440
rect 9963 4976 10005 4985
rect 9963 4936 9964 4976
rect 10004 4936 10005 4976
rect 9963 4927 10005 4936
rect 10060 4976 10100 4985
rect 9964 4842 10004 4927
rect 9771 4640 9813 4649
rect 9771 4600 9772 4640
rect 9812 4600 9813 4640
rect 9771 4591 9813 4600
rect 10060 4481 10100 4936
rect 10059 4472 10101 4481
rect 10059 4432 10060 4472
rect 10100 4432 10101 4472
rect 10059 4423 10101 4432
rect 9579 4304 9621 4313
rect 9579 4264 9580 4304
rect 9620 4264 9621 4304
rect 9579 4255 9621 4264
rect 9580 4231 9620 4255
rect 9580 4169 9620 4191
rect 9964 4220 10004 4229
rect 9772 3968 9812 3977
rect 9812 3928 9908 3968
rect 9772 3919 9812 3928
rect 9675 3884 9717 3893
rect 9675 3844 9676 3884
rect 9716 3844 9717 3884
rect 9675 3835 9717 3844
rect 9676 3464 9716 3835
rect 9676 3415 9716 3424
rect 9771 3380 9813 3389
rect 9771 3340 9772 3380
rect 9812 3340 9813 3380
rect 9771 3331 9813 3340
rect 9772 3246 9812 3331
rect 9771 2624 9813 2633
rect 9771 2584 9772 2624
rect 9812 2584 9813 2624
rect 9771 2575 9813 2584
rect 9772 2490 9812 2575
rect 9580 2456 9620 2465
rect 9580 2129 9620 2416
rect 9675 2204 9717 2213
rect 9675 2164 9676 2204
rect 9716 2164 9717 2204
rect 9675 2155 9717 2164
rect 9579 2120 9621 2129
rect 9579 2080 9580 2120
rect 9620 2080 9621 2120
rect 9579 2071 9621 2080
rect 9388 1240 9524 1280
rect 9291 1196 9333 1205
rect 9291 1156 9292 1196
rect 9332 1156 9333 1196
rect 9291 1147 9333 1156
rect 8908 1037 8948 1072
rect 9100 1072 9236 1112
rect 8907 1028 8949 1037
rect 8907 988 8908 1028
rect 8948 988 8949 1028
rect 8907 979 8949 988
rect 8811 692 8853 701
rect 8811 652 8812 692
rect 8852 652 8853 692
rect 8811 643 8853 652
rect 8907 356 8949 365
rect 8907 316 8908 356
rect 8948 316 8949 356
rect 8907 307 8949 316
rect 8908 80 8948 307
rect 9100 80 9140 1072
rect 9292 1062 9332 1147
rect 9388 776 9428 1240
rect 9676 1112 9716 2155
rect 9771 1952 9813 1961
rect 9771 1912 9772 1952
rect 9812 1912 9813 1952
rect 9771 1903 9813 1912
rect 9772 1793 9812 1903
rect 9771 1784 9813 1793
rect 9771 1744 9772 1784
rect 9812 1744 9813 1784
rect 9771 1735 9813 1744
rect 9771 1364 9813 1373
rect 9771 1324 9772 1364
rect 9812 1324 9813 1364
rect 9771 1315 9813 1324
rect 9676 1063 9716 1072
rect 9484 953 9524 1038
rect 9483 944 9525 953
rect 9483 904 9484 944
rect 9524 904 9525 944
rect 9483 895 9525 904
rect 9388 736 9524 776
rect 9291 692 9333 701
rect 9291 652 9292 692
rect 9332 652 9333 692
rect 9291 643 9333 652
rect 9292 80 9332 643
rect 9484 80 9524 736
rect 9772 692 9812 1315
rect 9676 652 9812 692
rect 9676 80 9716 652
rect 9868 608 9908 3928
rect 9964 2549 10004 4180
rect 10156 4145 10196 5692
rect 10443 5648 10485 5657
rect 10443 5608 10444 5648
rect 10484 5608 10485 5648
rect 10443 5599 10485 5608
rect 10444 5514 10484 5599
rect 10252 5480 10292 5489
rect 10155 4136 10197 4145
rect 10155 4096 10156 4136
rect 10196 4096 10197 4136
rect 10155 4087 10197 4096
rect 10156 3968 10196 3977
rect 10060 3928 10156 3968
rect 9963 2540 10005 2549
rect 9963 2500 9964 2540
rect 10004 2500 10005 2540
rect 9963 2491 10005 2500
rect 9963 2120 10005 2129
rect 9963 2080 9964 2120
rect 10004 2080 10005 2120
rect 9963 2071 10005 2080
rect 9964 1986 10004 2071
rect 9963 1112 10005 1121
rect 9963 1072 9964 1112
rect 10004 1072 10005 1112
rect 9963 1063 10005 1072
rect 9772 568 9908 608
rect 9772 197 9812 568
rect 9771 188 9813 197
rect 9964 188 10004 1063
rect 9771 148 9772 188
rect 9812 148 9813 188
rect 9771 139 9813 148
rect 9868 148 10004 188
rect 9868 80 9908 148
rect 10060 80 10100 3928
rect 10156 3919 10196 3928
rect 10252 3632 10292 5440
rect 10347 5396 10389 5405
rect 10347 5356 10348 5396
rect 10388 5356 10389 5396
rect 10347 5347 10389 5356
rect 10348 5060 10388 5347
rect 10443 5312 10485 5321
rect 10443 5272 10444 5312
rect 10484 5272 10485 5312
rect 10443 5263 10485 5272
rect 10348 5011 10388 5020
rect 10444 4220 10484 5263
rect 10539 5060 10581 5069
rect 10539 5020 10540 5060
rect 10580 5020 10581 5060
rect 10539 5011 10581 5020
rect 10444 4171 10484 4180
rect 10348 4136 10388 4145
rect 10348 3809 10388 4096
rect 10540 4136 10580 5011
rect 10636 4976 10676 7027
rect 10636 4927 10676 4936
rect 10732 6992 10772 7001
rect 10732 4388 10772 6952
rect 10924 6992 10964 7001
rect 10924 5153 10964 6952
rect 11212 6833 11252 7876
rect 11308 7589 11348 9892
rect 11404 9101 11444 10060
rect 11500 9689 11540 10228
rect 11884 10268 11924 10277
rect 11595 10184 11637 10193
rect 11595 10144 11596 10184
rect 11636 10144 11637 10184
rect 11595 10135 11637 10144
rect 11788 10184 11828 10195
rect 11596 10050 11636 10135
rect 11788 10109 11828 10144
rect 11787 10100 11829 10109
rect 11787 10060 11788 10100
rect 11828 10060 11829 10100
rect 11787 10051 11829 10060
rect 11499 9680 11541 9689
rect 11884 9680 11924 10228
rect 12076 10268 12116 10277
rect 11979 10016 12021 10025
rect 11979 9976 11980 10016
rect 12020 9976 12021 10016
rect 11979 9967 12021 9976
rect 11499 9640 11500 9680
rect 11540 9640 11541 9680
rect 11499 9631 11541 9640
rect 11596 9640 11924 9680
rect 11403 9092 11445 9101
rect 11403 9052 11404 9092
rect 11444 9052 11445 9092
rect 11403 9043 11445 9052
rect 11404 8924 11444 8933
rect 11596 8924 11636 9640
rect 11884 9512 11924 9521
rect 11444 8884 11636 8924
rect 11788 9472 11884 9512
rect 11404 8875 11444 8884
rect 11788 8840 11828 9472
rect 11884 9463 11924 9472
rect 11883 9260 11925 9269
rect 11883 9220 11884 9260
rect 11924 9220 11925 9260
rect 11883 9211 11925 9220
rect 11596 8800 11828 8840
rect 11499 8504 11541 8513
rect 11499 8464 11500 8504
rect 11540 8464 11541 8504
rect 11499 8455 11541 8464
rect 11403 8252 11445 8261
rect 11403 8212 11404 8252
rect 11444 8212 11445 8252
rect 11403 8203 11445 8212
rect 11404 7925 11444 8203
rect 11403 7916 11445 7925
rect 11403 7876 11404 7916
rect 11444 7876 11445 7916
rect 11403 7867 11445 7876
rect 11307 7580 11349 7589
rect 11307 7540 11308 7580
rect 11348 7540 11349 7580
rect 11307 7531 11349 7540
rect 11500 7244 11540 8455
rect 11596 8000 11636 8800
rect 11788 8672 11828 8681
rect 11785 8632 11788 8672
rect 11785 8623 11828 8632
rect 11691 8588 11733 8597
rect 11691 8548 11692 8588
rect 11732 8548 11733 8588
rect 11691 8539 11733 8548
rect 11692 8454 11732 8539
rect 11785 8513 11825 8623
rect 11884 8597 11924 9211
rect 11883 8588 11925 8597
rect 11883 8548 11884 8588
rect 11924 8548 11925 8588
rect 11883 8539 11925 8548
rect 11784 8504 11826 8513
rect 11784 8464 11785 8504
rect 11825 8464 11826 8504
rect 11784 8455 11826 8464
rect 11980 8345 12020 9967
rect 12076 9848 12116 10228
rect 12364 10226 12404 10387
rect 12652 10361 12692 11899
rect 12844 11696 12884 11899
rect 12748 11108 12788 11117
rect 12651 10352 12693 10361
rect 12651 10312 12652 10352
rect 12692 10312 12693 10352
rect 12651 10303 12693 10312
rect 12172 10184 12212 10193
rect 12556 10193 12596 10272
rect 12364 10177 12404 10186
rect 12459 10184 12501 10193
rect 12172 10100 12212 10144
rect 12459 10144 12460 10184
rect 12500 10144 12501 10184
rect 12459 10135 12501 10144
rect 12556 10184 12604 10193
rect 12603 10144 12604 10184
rect 12556 10135 12604 10144
rect 12652 10184 12692 10303
rect 12652 10135 12692 10144
rect 12172 10060 12305 10100
rect 12265 9932 12305 10060
rect 12364 10025 12404 10110
rect 12363 10016 12405 10025
rect 12363 9976 12364 10016
rect 12404 9976 12405 10016
rect 12460 10016 12500 10135
rect 12460 9976 12692 10016
rect 12363 9967 12405 9976
rect 12265 9892 12308 9932
rect 12268 9848 12308 9892
rect 12076 9808 12212 9848
rect 12268 9808 12500 9848
rect 12075 9680 12117 9689
rect 12075 9640 12076 9680
rect 12116 9640 12117 9680
rect 12075 9631 12117 9640
rect 12076 9546 12116 9631
rect 12172 9437 12212 9808
rect 12460 9764 12500 9808
rect 12460 9724 12603 9764
rect 12267 9680 12309 9689
rect 12267 9640 12268 9680
rect 12308 9640 12309 9680
rect 12267 9631 12309 9640
rect 12268 9512 12308 9631
rect 12563 9596 12603 9724
rect 12652 9680 12692 9976
rect 12748 9689 12788 11068
rect 12844 10361 12884 11656
rect 12940 10436 12980 12823
rect 13036 11948 13076 13159
rect 13132 13049 13172 13168
rect 13228 13208 13268 13217
rect 13131 13040 13173 13049
rect 13131 13000 13132 13040
rect 13172 13000 13173 13040
rect 13131 12991 13173 13000
rect 13132 12629 13172 12991
rect 13131 12620 13173 12629
rect 13131 12580 13132 12620
rect 13172 12580 13173 12620
rect 13131 12571 13173 12580
rect 13228 12491 13268 13168
rect 13516 12881 13556 15688
rect 13707 15560 13749 15569
rect 13707 15520 13708 15560
rect 13748 15520 13749 15560
rect 13707 15511 13749 15520
rect 13611 15392 13653 15401
rect 13611 15352 13612 15392
rect 13652 15352 13653 15392
rect 13611 15343 13653 15352
rect 13612 15258 13652 15343
rect 13612 14720 13652 14729
rect 13708 14720 13748 15511
rect 13652 14680 13748 14720
rect 13612 14057 13652 14680
rect 13611 14048 13653 14057
rect 13611 14008 13612 14048
rect 13652 14008 13653 14048
rect 13611 13999 13653 14008
rect 13611 13880 13653 13889
rect 13611 13840 13612 13880
rect 13652 13840 13653 13880
rect 13611 13831 13653 13840
rect 13612 13292 13652 13831
rect 13612 13243 13652 13252
rect 13708 13292 13748 13301
rect 13804 13292 13844 15763
rect 13900 15560 13940 16528
rect 13996 16073 14036 17032
rect 14091 16904 14133 16913
rect 14091 16864 14092 16904
rect 14132 16864 14133 16904
rect 14091 16855 14133 16864
rect 14092 16770 14132 16855
rect 14188 16652 14228 17620
rect 14475 17620 14476 17660
rect 14516 17620 14517 17660
rect 14475 17611 14517 17620
rect 14476 17240 14516 17611
rect 14860 17501 14900 17704
rect 14859 17492 14901 17501
rect 14859 17452 14860 17492
rect 14900 17452 14901 17492
rect 14859 17443 14901 17452
rect 15052 17333 15092 18283
rect 15051 17324 15093 17333
rect 15051 17284 15052 17324
rect 15092 17284 15093 17324
rect 15051 17275 15093 17284
rect 14380 17200 14516 17240
rect 14283 16652 14325 16661
rect 14188 16612 14284 16652
rect 14324 16612 14325 16652
rect 14283 16603 14325 16612
rect 13995 16064 14037 16073
rect 13995 16024 13996 16064
rect 14036 16024 14037 16064
rect 13995 16015 14037 16024
rect 13996 15728 14036 16015
rect 13996 15688 14228 15728
rect 13900 14888 13940 15520
rect 13996 15560 14036 15571
rect 13996 15485 14036 15520
rect 13995 15476 14037 15485
rect 13995 15436 13996 15476
rect 14036 15436 14037 15476
rect 13995 15427 14037 15436
rect 13900 14848 14132 14888
rect 13899 14720 13941 14729
rect 13899 14680 13900 14720
rect 13940 14680 13941 14720
rect 13899 14671 13941 14680
rect 13900 14586 13940 14671
rect 13995 14636 14037 14645
rect 13995 14596 13996 14636
rect 14036 14596 14037 14636
rect 13995 14587 14037 14596
rect 13996 14502 14036 14587
rect 13995 13964 14037 13973
rect 13995 13924 13996 13964
rect 14036 13924 14037 13964
rect 13995 13915 14037 13924
rect 13899 13880 13941 13889
rect 13899 13840 13900 13880
rect 13940 13840 13941 13880
rect 13899 13831 13941 13840
rect 13748 13252 13844 13292
rect 13515 12872 13557 12881
rect 13515 12832 13516 12872
rect 13556 12832 13557 12872
rect 13515 12823 13557 12832
rect 13323 12788 13365 12797
rect 13323 12748 13324 12788
rect 13364 12748 13365 12788
rect 13323 12739 13365 12748
rect 13036 11899 13076 11908
rect 13132 12451 13268 12491
rect 13324 12536 13364 12739
rect 13611 12620 13653 12629
rect 13611 12580 13612 12620
rect 13652 12580 13653 12620
rect 13611 12571 13653 12580
rect 13420 12536 13460 12545
rect 13324 12496 13420 12536
rect 13132 11780 13172 12451
rect 13324 11957 13364 12496
rect 13420 12487 13460 12496
rect 13612 12486 13652 12571
rect 13323 11948 13365 11957
rect 13323 11908 13324 11948
rect 13364 11908 13365 11948
rect 13323 11899 13365 11908
rect 13419 11864 13461 11873
rect 13419 11824 13420 11864
rect 13460 11824 13461 11864
rect 13419 11815 13461 11824
rect 13132 11740 13364 11780
rect 13036 11528 13076 11537
rect 13036 11360 13076 11488
rect 13228 11528 13268 11537
rect 13036 11320 13172 11360
rect 13035 11024 13077 11033
rect 13035 10984 13036 11024
rect 13076 10984 13077 11024
rect 13035 10975 13077 10984
rect 13036 10890 13076 10975
rect 12940 10396 13076 10436
rect 12843 10352 12885 10361
rect 12843 10312 12844 10352
rect 12884 10312 12885 10352
rect 12843 10303 12885 10312
rect 12844 10184 12884 10193
rect 12844 10109 12884 10144
rect 12843 10100 12885 10109
rect 12843 10060 12844 10100
rect 12884 10060 12885 10100
rect 12843 10051 12885 10060
rect 12844 10049 12884 10051
rect 12940 10016 12980 10027
rect 12940 9941 12980 9976
rect 12939 9932 12981 9941
rect 12939 9892 12940 9932
rect 12980 9892 12981 9932
rect 12939 9883 12981 9892
rect 12939 9764 12981 9773
rect 12939 9724 12940 9764
rect 12980 9724 12981 9764
rect 12939 9715 12981 9724
rect 12652 9631 12692 9640
rect 12747 9680 12789 9689
rect 12747 9640 12748 9680
rect 12788 9640 12789 9680
rect 12747 9631 12789 9640
rect 12556 9556 12603 9596
rect 12556 9512 12596 9556
rect 12268 9463 12308 9472
rect 12412 9489 12452 9498
rect 12171 9428 12213 9437
rect 12171 9388 12172 9428
rect 12212 9388 12213 9428
rect 12171 9379 12213 9388
rect 12412 9344 12452 9449
rect 12809 9497 12849 9506
rect 12412 9304 12500 9344
rect 12267 9260 12309 9269
rect 12267 9220 12268 9260
rect 12308 9220 12309 9260
rect 12267 9211 12309 9220
rect 12171 9092 12213 9101
rect 12171 9052 12172 9092
rect 12212 9052 12213 9092
rect 12171 9043 12213 9052
rect 12076 8672 12116 8681
rect 11691 8336 11733 8345
rect 11691 8296 11692 8336
rect 11732 8296 11733 8336
rect 11691 8287 11733 8296
rect 11979 8336 12021 8345
rect 11979 8296 11980 8336
rect 12020 8296 12021 8336
rect 11979 8287 12021 8296
rect 11692 8177 11732 8287
rect 11691 8168 11733 8177
rect 11691 8128 11692 8168
rect 11732 8128 11733 8168
rect 11691 8119 11733 8128
rect 11884 8084 11924 8095
rect 11884 8009 11924 8044
rect 11979 8084 12021 8093
rect 11979 8044 11980 8084
rect 12020 8044 12021 8084
rect 11979 8035 12021 8044
rect 11692 8000 11732 8009
rect 11596 7960 11692 8000
rect 11692 7841 11732 7960
rect 11883 8000 11925 8009
rect 11883 7960 11884 8000
rect 11924 7960 11925 8000
rect 11883 7951 11925 7960
rect 11691 7832 11733 7841
rect 11691 7792 11692 7832
rect 11732 7792 11733 7832
rect 11691 7783 11733 7792
rect 11500 7195 11540 7204
rect 11788 7160 11828 7169
rect 11595 7076 11637 7085
rect 11595 7036 11596 7076
rect 11636 7036 11637 7076
rect 11595 7027 11637 7036
rect 11308 6992 11348 7001
rect 11211 6824 11253 6833
rect 11211 6784 11212 6824
rect 11252 6784 11253 6824
rect 11211 6775 11253 6784
rect 11211 6488 11253 6497
rect 11211 6448 11212 6488
rect 11252 6448 11253 6488
rect 11211 6439 11253 6448
rect 10923 5144 10965 5153
rect 10923 5104 10924 5144
rect 10964 5104 10965 5144
rect 10923 5095 10965 5104
rect 11115 5060 11157 5069
rect 11115 5020 11116 5060
rect 11156 5020 11157 5060
rect 11115 5011 11157 5020
rect 10924 4976 10964 4985
rect 10540 4087 10580 4096
rect 10636 4348 10772 4388
rect 10828 4936 10924 4976
rect 10347 3800 10389 3809
rect 10347 3760 10348 3800
rect 10388 3760 10389 3800
rect 10347 3751 10389 3760
rect 10252 3592 10484 3632
rect 10155 3464 10197 3473
rect 10155 3424 10156 3464
rect 10196 3424 10197 3464
rect 10155 3415 10197 3424
rect 10252 3464 10292 3473
rect 10156 3330 10196 3415
rect 10252 2129 10292 3424
rect 10347 3464 10389 3473
rect 10347 3424 10348 3464
rect 10388 3424 10389 3464
rect 10347 3415 10389 3424
rect 10348 2381 10388 3415
rect 10347 2372 10389 2381
rect 10347 2332 10348 2372
rect 10388 2332 10389 2372
rect 10347 2323 10389 2332
rect 10251 2120 10293 2129
rect 10251 2080 10252 2120
rect 10292 2080 10293 2120
rect 10251 2071 10293 2080
rect 10156 1952 10196 1961
rect 10348 1952 10388 2323
rect 10196 1912 10388 1952
rect 10156 1037 10196 1912
rect 10251 1700 10293 1709
rect 10251 1660 10252 1700
rect 10292 1660 10293 1700
rect 10251 1651 10293 1660
rect 10155 1028 10197 1037
rect 10155 988 10156 1028
rect 10196 988 10197 1028
rect 10155 979 10197 988
rect 10252 80 10292 1651
rect 10444 80 10484 3592
rect 10636 2885 10676 4348
rect 10828 4313 10868 4936
rect 10924 4927 10964 4936
rect 11116 4926 11156 5011
rect 10924 4808 10964 4817
rect 10964 4768 11156 4808
rect 10924 4759 10964 4768
rect 10923 4556 10965 4565
rect 10923 4516 10924 4556
rect 10964 4516 10965 4556
rect 10923 4507 10965 4516
rect 10924 4388 10964 4507
rect 10924 4339 10964 4348
rect 10827 4304 10869 4313
rect 10827 4264 10828 4304
rect 10868 4264 10869 4304
rect 10827 4255 10869 4264
rect 10732 4136 10772 4145
rect 10732 3893 10772 4096
rect 10923 4136 10965 4145
rect 10923 4096 10924 4136
rect 10964 4096 10965 4136
rect 10923 4087 10965 4096
rect 11116 4136 11156 4768
rect 11212 4229 11252 6439
rect 11308 5237 11348 6952
rect 11499 6740 11541 6749
rect 11404 6700 11500 6740
rect 11540 6700 11541 6740
rect 11307 5228 11349 5237
rect 11307 5188 11308 5228
rect 11348 5188 11349 5228
rect 11307 5179 11349 5188
rect 11308 4962 11348 4987
rect 11308 4901 11348 4922
rect 11307 4892 11349 4901
rect 11307 4852 11308 4892
rect 11348 4852 11349 4892
rect 11307 4843 11349 4852
rect 11404 4565 11444 6700
rect 11499 6691 11541 6700
rect 11596 4976 11636 7027
rect 11692 6992 11732 7001
rect 11692 6749 11732 6952
rect 11691 6740 11733 6749
rect 11691 6700 11692 6740
rect 11732 6700 11733 6740
rect 11691 6691 11733 6700
rect 11692 6488 11732 6499
rect 11692 6413 11732 6448
rect 11691 6404 11733 6413
rect 11691 6364 11692 6404
rect 11732 6364 11733 6404
rect 11691 6355 11733 6364
rect 11692 5648 11732 5657
rect 11692 5489 11732 5608
rect 11691 5480 11733 5489
rect 11691 5440 11692 5480
rect 11732 5440 11733 5480
rect 11691 5431 11733 5440
rect 11788 5144 11828 7120
rect 11884 6656 11924 6665
rect 11980 6656 12020 8035
rect 12076 8009 12116 8632
rect 12075 8000 12117 8009
rect 12075 7960 12076 8000
rect 12116 7960 12117 8000
rect 12075 7951 12117 7960
rect 12076 7866 12116 7951
rect 12172 7832 12212 9043
rect 12268 8765 12308 9211
rect 12363 9092 12405 9101
rect 12363 9052 12364 9092
rect 12404 9052 12405 9092
rect 12363 9043 12405 9052
rect 12267 8756 12309 8765
rect 12267 8716 12268 8756
rect 12308 8716 12309 8756
rect 12267 8707 12309 8716
rect 12267 8084 12309 8093
rect 12267 8044 12268 8084
rect 12308 8044 12309 8084
rect 12267 8035 12309 8044
rect 12268 8000 12308 8035
rect 12268 7949 12308 7960
rect 12364 8000 12404 9043
rect 12460 8933 12500 9304
rect 12459 8924 12501 8933
rect 12459 8884 12460 8924
rect 12500 8884 12501 8924
rect 12459 8875 12501 8884
rect 12460 8672 12500 8681
rect 12460 8009 12500 8632
rect 12556 8177 12596 9472
rect 12652 9483 12692 9492
rect 12849 9457 12884 9497
rect 12809 9448 12884 9457
rect 12652 9437 12692 9443
rect 12651 9428 12693 9437
rect 12651 9388 12652 9428
rect 12692 9388 12693 9428
rect 12651 9379 12693 9388
rect 12652 9348 12692 9379
rect 12844 9176 12884 9448
rect 12940 9344 12980 9715
rect 13036 9512 13076 10396
rect 13036 9463 13076 9472
rect 13036 9344 13076 9353
rect 12940 9304 13036 9344
rect 13132 9344 13172 11320
rect 13228 10184 13268 11488
rect 13324 11285 13364 11740
rect 13420 11696 13460 11815
rect 13420 11647 13460 11656
rect 13708 11369 13748 13252
rect 13900 12620 13940 13831
rect 13996 12629 14036 13915
rect 14092 13721 14132 14848
rect 14091 13712 14133 13721
rect 14091 13672 14092 13712
rect 14132 13672 14133 13712
rect 14091 13663 14133 13672
rect 14188 13208 14228 15688
rect 14283 15560 14325 15569
rect 14283 15520 14284 15560
rect 14324 15520 14325 15560
rect 14283 15511 14325 15520
rect 14284 15426 14324 15511
rect 14275 15056 14317 15065
rect 14275 15016 14276 15056
rect 14316 15016 14324 15056
rect 14275 15007 14324 15016
rect 14284 14972 14324 15007
rect 14284 14923 14324 14932
rect 14380 14804 14420 17200
rect 14476 17072 14516 17083
rect 14476 16997 14516 17032
rect 14475 16988 14517 16997
rect 14475 16948 14476 16988
rect 14516 16948 14517 16988
rect 14475 16939 14517 16948
rect 14763 16232 14805 16241
rect 14763 16192 14764 16232
rect 14804 16192 14805 16232
rect 14763 16183 14805 16192
rect 14764 16098 14804 16183
rect 14955 16064 14997 16073
rect 14955 16024 14956 16064
rect 14996 16024 14997 16064
rect 14955 16015 14997 16024
rect 14956 15930 14996 16015
rect 15052 15821 15092 17275
rect 15148 16325 15188 19375
rect 15244 17753 15284 19972
rect 15243 17744 15285 17753
rect 15243 17704 15244 17744
rect 15284 17704 15285 17744
rect 15243 17695 15285 17704
rect 15340 16661 15380 20392
rect 15435 20096 15477 20105
rect 15435 20056 15436 20096
rect 15476 20056 15477 20096
rect 15435 20047 15477 20056
rect 15436 19962 15476 20047
rect 15532 20012 15572 20021
rect 15435 19340 15477 19349
rect 15435 19300 15436 19340
rect 15476 19300 15477 19340
rect 15435 19291 15477 19300
rect 15339 16652 15381 16661
rect 15339 16612 15340 16652
rect 15380 16612 15381 16652
rect 15339 16603 15381 16612
rect 15147 16316 15189 16325
rect 15147 16276 15148 16316
rect 15188 16276 15189 16316
rect 15147 16267 15189 16276
rect 15244 16232 15284 16241
rect 15244 15989 15284 16192
rect 15340 16232 15380 16241
rect 15436 16232 15476 19291
rect 15532 18929 15572 19972
rect 15724 20012 15764 20728
rect 15628 19928 15668 19937
rect 15531 18920 15573 18929
rect 15531 18880 15532 18920
rect 15572 18880 15573 18920
rect 15531 18871 15573 18880
rect 15628 17669 15668 19888
rect 15724 19349 15764 19972
rect 15820 20096 15860 20896
rect 15915 20852 15957 20861
rect 15915 20812 15916 20852
rect 15956 20812 15957 20852
rect 15915 20803 15957 20812
rect 15916 20768 15956 20803
rect 16204 20777 16244 20862
rect 15916 20717 15956 20728
rect 16012 20768 16052 20777
rect 16203 20768 16245 20777
rect 16052 20728 16148 20768
rect 16012 20719 16052 20728
rect 16011 20600 16053 20609
rect 16011 20560 16012 20600
rect 16052 20560 16053 20600
rect 16011 20551 16053 20560
rect 15723 19340 15765 19349
rect 15723 19300 15724 19340
rect 15764 19300 15765 19340
rect 15723 19291 15765 19300
rect 15820 19265 15860 20056
rect 16012 20096 16052 20551
rect 16012 20047 16052 20056
rect 15915 20012 15957 20021
rect 15915 19972 15916 20012
rect 15956 19972 15957 20012
rect 15915 19963 15957 19972
rect 15819 19256 15861 19265
rect 15819 19216 15820 19256
rect 15860 19216 15861 19256
rect 15819 19207 15861 19216
rect 15627 17660 15669 17669
rect 15627 17620 15628 17660
rect 15668 17620 15669 17660
rect 15627 17611 15669 17620
rect 15723 17156 15765 17165
rect 15723 17116 15724 17156
rect 15764 17116 15765 17156
rect 15723 17107 15765 17116
rect 15724 17072 15764 17107
rect 15724 17021 15764 17032
rect 15819 17072 15861 17081
rect 15819 17032 15820 17072
rect 15860 17032 15861 17072
rect 15819 17023 15861 17032
rect 15820 16904 15860 17023
rect 15916 16988 15956 19963
rect 16011 19844 16053 19853
rect 16011 19804 16012 19844
rect 16052 19804 16053 19844
rect 16011 19795 16053 19804
rect 16012 17072 16052 19795
rect 16108 18425 16148 20728
rect 16203 20728 16204 20768
rect 16244 20728 16245 20768
rect 16203 20719 16245 20728
rect 16204 20600 16244 20609
rect 16204 20357 16244 20560
rect 16203 20348 16245 20357
rect 16203 20308 16204 20348
rect 16244 20308 16245 20348
rect 16203 20299 16245 20308
rect 16203 19760 16245 19769
rect 16203 19720 16204 19760
rect 16244 19720 16245 19760
rect 16203 19711 16245 19720
rect 16204 19256 16244 19711
rect 16300 19433 16340 27019
rect 16396 26405 16436 28960
rect 16588 27656 16628 29119
rect 16780 28333 16820 28342
rect 16683 28160 16725 28169
rect 16683 28120 16684 28160
rect 16724 28120 16725 28160
rect 16683 28111 16725 28120
rect 16588 26825 16628 27616
rect 16587 26816 16629 26825
rect 16587 26776 16588 26816
rect 16628 26776 16629 26816
rect 16587 26767 16629 26776
rect 16491 26480 16533 26489
rect 16491 26440 16492 26480
rect 16532 26440 16533 26480
rect 16491 26431 16533 26440
rect 16395 26396 16437 26405
rect 16395 26356 16396 26396
rect 16436 26356 16437 26396
rect 16395 26347 16437 26356
rect 16396 26144 16436 26153
rect 16492 26144 16532 26431
rect 16588 26237 16628 26767
rect 16684 26480 16724 28111
rect 16780 27824 16820 28293
rect 16780 27775 16820 27784
rect 16684 26440 16820 26480
rect 16587 26228 16629 26237
rect 16587 26188 16588 26228
rect 16628 26188 16629 26228
rect 16587 26179 16629 26188
rect 16436 26104 16532 26144
rect 16396 26095 16436 26104
rect 16683 26060 16725 26069
rect 16683 26020 16684 26060
rect 16724 26020 16725 26060
rect 16683 26011 16725 26020
rect 16540 25313 16580 25322
rect 16580 25273 16628 25304
rect 16540 25264 16628 25273
rect 16588 24800 16628 25264
rect 16684 25220 16724 26011
rect 16684 25171 16724 25180
rect 16780 25052 16820 26440
rect 16588 24751 16628 24760
rect 16684 25012 16820 25052
rect 16396 24632 16436 24641
rect 16436 24592 16532 24632
rect 16396 24583 16436 24592
rect 16395 24296 16437 24305
rect 16395 24256 16396 24296
rect 16436 24256 16437 24296
rect 16395 24247 16437 24256
rect 16396 20693 16436 24247
rect 16492 23708 16532 24592
rect 16684 24305 16724 25012
rect 16876 24380 16916 29628
rect 17067 29168 17109 29177
rect 17067 29128 17068 29168
rect 17108 29128 17109 29168
rect 17067 29119 17109 29128
rect 17068 29034 17108 29119
rect 16972 28244 17012 28253
rect 17164 28244 17204 29875
rect 17356 29840 17396 30379
rect 17356 29791 17396 29800
rect 17452 29840 17492 29849
rect 17452 29420 17492 29800
rect 17356 29380 17492 29420
rect 17260 28916 17300 28925
rect 17260 28328 17300 28876
rect 17260 28279 17300 28288
rect 17356 28328 17396 29380
rect 17548 29336 17588 30472
rect 17644 30269 17684 31312
rect 17739 30428 17781 30437
rect 17739 30388 17740 30428
rect 17780 30388 17781 30428
rect 17739 30379 17781 30388
rect 17740 30294 17780 30379
rect 17643 30260 17685 30269
rect 17643 30220 17644 30260
rect 17684 30220 17685 30260
rect 17643 30211 17685 30220
rect 17644 29672 17684 30211
rect 17739 30092 17781 30101
rect 17739 30052 17740 30092
rect 17780 30052 17781 30092
rect 17836 30092 17876 31900
rect 17932 31436 17972 32311
rect 18220 32201 18260 32286
rect 18028 32192 18068 32201
rect 18219 32192 18261 32201
rect 18068 32152 18164 32192
rect 18028 32143 18068 32152
rect 18027 32024 18069 32033
rect 18027 31984 18028 32024
rect 18068 31984 18069 32024
rect 18124 32024 18164 32152
rect 18219 32152 18220 32192
rect 18260 32152 18261 32192
rect 18219 32143 18261 32152
rect 18220 32024 18260 32033
rect 18124 31984 18220 32024
rect 18027 31975 18069 31984
rect 18220 31975 18260 31984
rect 18028 31890 18068 31975
rect 18028 31436 18068 31445
rect 17932 31396 18028 31436
rect 17932 30773 17972 31396
rect 18028 31387 18068 31396
rect 18123 31436 18165 31445
rect 18123 31396 18124 31436
rect 18164 31396 18165 31436
rect 18123 31387 18165 31396
rect 18124 31302 18164 31387
rect 18123 31184 18165 31193
rect 18123 31144 18124 31184
rect 18164 31144 18165 31184
rect 18123 31135 18165 31144
rect 17931 30764 17973 30773
rect 17931 30724 17932 30764
rect 17972 30724 17973 30764
rect 17931 30715 17973 30724
rect 17836 30052 18068 30092
rect 17739 30043 17781 30052
rect 17740 29924 17780 30043
rect 17836 29924 17876 29933
rect 17740 29884 17836 29924
rect 17836 29875 17876 29884
rect 17932 29840 17972 29849
rect 17644 29632 17876 29672
rect 17548 29296 17684 29336
rect 17451 29252 17493 29261
rect 17451 29212 17452 29252
rect 17492 29212 17493 29252
rect 17451 29203 17493 29212
rect 17012 28204 17204 28244
rect 16972 28195 17012 28204
rect 17356 28160 17396 28288
rect 17164 28120 17396 28160
rect 17164 27749 17204 28120
rect 17452 27992 17492 29203
rect 17547 29168 17589 29177
rect 17547 29128 17548 29168
rect 17588 29128 17589 29168
rect 17547 29119 17589 29128
rect 17548 29034 17588 29119
rect 17644 29000 17684 29296
rect 17644 28960 17780 29000
rect 17547 28916 17589 28925
rect 17547 28876 17548 28916
rect 17588 28876 17589 28916
rect 17547 28867 17589 28876
rect 17260 27952 17492 27992
rect 17163 27740 17205 27749
rect 17163 27700 17164 27740
rect 17204 27700 17205 27740
rect 17163 27691 17205 27700
rect 17068 27572 17108 27581
rect 16971 26816 17013 26825
rect 16971 26776 16972 26816
rect 17012 26776 17013 26816
rect 16971 26767 17013 26776
rect 16972 26682 17012 26767
rect 16971 26396 17013 26405
rect 16971 26356 16972 26396
rect 17012 26356 17013 26396
rect 16971 26347 17013 26356
rect 16780 24340 16916 24380
rect 16972 24548 17012 26347
rect 17068 26321 17108 27532
rect 17260 27488 17300 27952
rect 17548 27833 17588 28867
rect 17643 28328 17685 28337
rect 17643 28288 17644 28328
rect 17684 28288 17685 28328
rect 17643 28279 17685 28288
rect 17740 28328 17780 28960
rect 17355 27824 17397 27833
rect 17355 27784 17356 27824
rect 17396 27784 17397 27824
rect 17355 27775 17397 27784
rect 17547 27824 17589 27833
rect 17547 27784 17548 27824
rect 17588 27784 17589 27824
rect 17547 27775 17589 27784
rect 17260 27439 17300 27448
rect 17163 26984 17205 26993
rect 17163 26944 17164 26984
rect 17204 26944 17205 26984
rect 17163 26935 17205 26944
rect 17164 26850 17204 26935
rect 17163 26396 17205 26405
rect 17163 26356 17164 26396
rect 17204 26356 17205 26396
rect 17163 26347 17205 26356
rect 17067 26312 17109 26321
rect 17067 26272 17068 26312
rect 17108 26272 17109 26312
rect 17067 26263 17109 26272
rect 17164 25145 17204 26347
rect 17259 25892 17301 25901
rect 17259 25852 17260 25892
rect 17300 25852 17301 25892
rect 17259 25843 17301 25852
rect 17260 25304 17300 25843
rect 17356 25817 17396 27775
rect 17452 27572 17492 27581
rect 17452 27413 17492 27532
rect 17644 27488 17684 28279
rect 17740 28169 17780 28288
rect 17836 28328 17876 29632
rect 17836 28253 17876 28288
rect 17835 28244 17877 28253
rect 17835 28204 17836 28244
rect 17876 28204 17877 28244
rect 17835 28195 17877 28204
rect 17739 28160 17781 28169
rect 17739 28120 17740 28160
rect 17780 28120 17781 28160
rect 17739 28111 17781 28120
rect 17836 27656 17876 27665
rect 17836 27497 17876 27616
rect 17644 27439 17684 27448
rect 17835 27488 17877 27497
rect 17835 27448 17836 27488
rect 17876 27448 17877 27488
rect 17835 27439 17877 27448
rect 17451 27404 17493 27413
rect 17451 27364 17452 27404
rect 17492 27364 17493 27404
rect 17451 27355 17493 27364
rect 17932 27245 17972 29800
rect 18028 29513 18068 30052
rect 18027 29504 18069 29513
rect 18027 29464 18028 29504
rect 18068 29464 18069 29504
rect 18027 29455 18069 29464
rect 17931 27236 17973 27245
rect 17931 27196 17932 27236
rect 17972 27196 17973 27236
rect 17931 27187 17973 27196
rect 17451 26984 17493 26993
rect 18028 26984 18068 29455
rect 17451 26944 17452 26984
rect 17492 26944 17493 26984
rect 17451 26935 17493 26944
rect 17932 26944 18068 26984
rect 17452 26816 17492 26935
rect 17452 26767 17492 26776
rect 17548 26816 17588 26856
rect 17548 26741 17588 26776
rect 17932 26816 17972 26944
rect 17547 26732 17589 26741
rect 17547 26692 17548 26732
rect 17588 26692 17589 26732
rect 17547 26683 17589 26692
rect 17355 25808 17397 25817
rect 17355 25768 17356 25808
rect 17396 25768 17397 25808
rect 17355 25759 17397 25768
rect 17260 25255 17300 25264
rect 17356 25304 17396 25313
rect 17548 25304 17588 26683
rect 17739 26396 17781 26405
rect 17739 26356 17740 26396
rect 17780 26356 17781 26396
rect 17739 26347 17781 26356
rect 17643 26228 17685 26237
rect 17643 26188 17644 26228
rect 17684 26188 17685 26228
rect 17643 26179 17685 26188
rect 17644 26144 17684 26179
rect 17644 26093 17684 26104
rect 17643 25808 17685 25817
rect 17643 25768 17644 25808
rect 17684 25768 17685 25808
rect 17643 25759 17685 25768
rect 17396 25264 17588 25304
rect 17356 25255 17396 25264
rect 17163 25136 17205 25145
rect 17163 25096 17164 25136
rect 17204 25096 17205 25136
rect 17163 25087 17205 25096
rect 17355 25136 17397 25145
rect 17355 25096 17356 25136
rect 17396 25096 17397 25136
rect 17355 25087 17397 25096
rect 17259 24800 17301 24809
rect 17259 24760 17260 24800
rect 17300 24760 17301 24800
rect 17259 24751 17301 24760
rect 17260 24666 17300 24751
rect 17068 24548 17108 24557
rect 16972 24508 17068 24548
rect 16683 24296 16725 24305
rect 16683 24256 16684 24296
rect 16724 24256 16725 24296
rect 16683 24247 16725 24256
rect 16636 23801 16676 23810
rect 16676 23761 16724 23792
rect 16636 23752 16724 23761
rect 16492 23668 16628 23708
rect 16491 23456 16533 23465
rect 16491 23416 16492 23456
rect 16532 23416 16533 23456
rect 16491 23407 16533 23416
rect 16492 23120 16532 23407
rect 16492 23071 16532 23080
rect 16588 22289 16628 23668
rect 16684 23288 16724 23752
rect 16780 23708 16820 24340
rect 16972 23708 17012 24508
rect 17068 24499 17108 24508
rect 17163 24548 17205 24557
rect 17163 24508 17164 24548
rect 17204 24508 17205 24548
rect 17163 24499 17205 24508
rect 16780 23659 16820 23668
rect 16876 23668 17012 23708
rect 16779 23372 16821 23381
rect 16779 23332 16780 23372
rect 16820 23332 16821 23372
rect 16779 23323 16821 23332
rect 16684 23239 16724 23248
rect 16780 22532 16820 23323
rect 16876 22709 16916 23668
rect 17068 23624 17108 23633
rect 16972 23584 17068 23624
rect 16972 23120 17012 23584
rect 17068 23575 17108 23584
rect 17068 23288 17108 23297
rect 17164 23288 17204 24499
rect 17260 23801 17300 23806
rect 17259 23797 17301 23801
rect 17259 23752 17260 23797
rect 17300 23752 17301 23797
rect 17259 23743 17301 23752
rect 17260 23662 17300 23743
rect 17356 23540 17396 25087
rect 17451 24716 17493 24725
rect 17451 24676 17452 24716
rect 17492 24676 17493 24716
rect 17451 24667 17493 24676
rect 17452 24548 17492 24667
rect 17644 24632 17684 25759
rect 17740 25649 17780 26347
rect 17835 25892 17877 25901
rect 17835 25852 17836 25892
rect 17876 25852 17877 25892
rect 17835 25843 17877 25852
rect 17836 25758 17876 25843
rect 17739 25640 17781 25649
rect 17739 25600 17740 25640
rect 17780 25600 17781 25640
rect 17739 25591 17781 25600
rect 17740 25397 17780 25428
rect 17739 25388 17781 25397
rect 17739 25348 17740 25388
rect 17780 25348 17781 25388
rect 17932 25388 17972 26776
rect 18027 26816 18069 26825
rect 18027 26776 18028 26816
rect 18068 26776 18069 26816
rect 18027 26767 18069 26776
rect 18028 25472 18068 26767
rect 18124 26144 18164 31135
rect 18219 30764 18261 30773
rect 18219 30724 18220 30764
rect 18260 30724 18261 30764
rect 18219 30715 18261 30724
rect 18220 30680 18260 30715
rect 18220 30521 18260 30640
rect 18219 30512 18261 30521
rect 18219 30472 18220 30512
rect 18260 30472 18261 30512
rect 18219 30463 18261 30472
rect 18219 28748 18261 28757
rect 18219 28708 18220 28748
rect 18260 28708 18261 28748
rect 18219 28699 18261 28708
rect 18220 28580 18260 28699
rect 18316 28664 18356 32824
rect 18412 32360 18452 32908
rect 18508 32878 18548 34168
rect 18604 33713 18644 33798
rect 18603 33704 18645 33713
rect 18603 33664 18604 33704
rect 18644 33664 18645 33704
rect 18603 33655 18645 33664
rect 18603 33536 18645 33545
rect 18603 33496 18604 33536
rect 18644 33496 18645 33536
rect 18603 33487 18645 33496
rect 18508 32829 18548 32838
rect 18604 32537 18644 33487
rect 18700 32780 18740 34168
rect 19083 34168 19084 34208
rect 19124 34168 19125 34208
rect 19083 34159 19125 34168
rect 19084 33699 19124 34159
rect 19276 33872 19316 36100
rect 19467 36091 19509 36100
rect 19371 35972 19413 35981
rect 19371 35932 19372 35972
rect 19412 35932 19413 35972
rect 19371 35923 19413 35932
rect 19372 35838 19412 35923
rect 19563 35720 19605 35729
rect 19563 35680 19564 35720
rect 19604 35680 19605 35720
rect 19563 35671 19605 35680
rect 19564 35586 19604 35671
rect 19660 35300 19700 36436
rect 19756 36149 19796 37444
rect 19852 36821 19892 38200
rect 19948 38156 19988 38165
rect 19948 37409 19988 38116
rect 20140 37988 20180 37997
rect 20180 37948 20660 37988
rect 20140 37939 20180 37948
rect 20235 37820 20277 37829
rect 20235 37780 20236 37820
rect 20276 37780 20277 37820
rect 20235 37771 20277 37780
rect 20236 37652 20276 37771
rect 20236 37603 20276 37612
rect 19947 37400 19989 37409
rect 19947 37360 19948 37400
rect 19988 37360 19989 37400
rect 19947 37351 19989 37360
rect 20127 37389 20167 37398
rect 20043 37316 20085 37325
rect 20127 37316 20167 37349
rect 20043 37276 20044 37316
rect 20084 37276 20167 37316
rect 20043 37267 20085 37276
rect 19947 37232 19989 37241
rect 19947 37192 19948 37232
rect 19988 37192 19989 37232
rect 19947 37183 19989 37192
rect 19948 37098 19988 37183
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19947 36980 19989 36989
rect 19947 36940 19948 36980
rect 19988 36940 19989 36980
rect 19947 36931 19989 36940
rect 19851 36812 19893 36821
rect 19851 36772 19852 36812
rect 19892 36772 19893 36812
rect 19851 36763 19893 36772
rect 19852 36644 19892 36653
rect 19948 36644 19988 36931
rect 19892 36604 19988 36644
rect 19852 36595 19892 36604
rect 20044 36560 20084 36569
rect 20084 36520 20564 36560
rect 20044 36511 20084 36520
rect 19755 36140 19797 36149
rect 19755 36100 19756 36140
rect 19796 36100 19797 36140
rect 19755 36091 19797 36100
rect 19564 35260 19700 35300
rect 19756 35972 19796 35981
rect 19467 35048 19509 35057
rect 19467 35008 19468 35048
rect 19508 35008 19509 35048
rect 19467 34999 19509 35008
rect 19468 34914 19508 34999
rect 19276 33823 19316 33832
rect 19371 33872 19413 33881
rect 19371 33832 19372 33872
rect 19412 33832 19413 33872
rect 19371 33823 19413 33832
rect 19084 33650 19124 33659
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 19084 33116 19124 33125
rect 19372 33116 19412 33823
rect 19467 33620 19509 33629
rect 19467 33580 19468 33620
rect 19508 33580 19509 33620
rect 19467 33571 19509 33580
rect 19468 33486 19508 33571
rect 19124 33076 19412 33116
rect 19084 33067 19124 33076
rect 18891 32948 18933 32957
rect 18891 32908 18892 32948
rect 18932 32908 18933 32948
rect 18891 32899 18933 32908
rect 19372 32948 19412 32957
rect 18892 32864 18932 32899
rect 18892 32813 18932 32824
rect 19083 32864 19125 32873
rect 19083 32824 19084 32864
rect 19124 32824 19125 32864
rect 19083 32815 19125 32824
rect 18700 32731 18740 32740
rect 19084 32730 19124 32815
rect 19372 32789 19412 32908
rect 19564 32864 19604 35260
rect 19660 35132 19700 35141
rect 19660 34889 19700 35092
rect 19659 34880 19701 34889
rect 19659 34840 19660 34880
rect 19700 34840 19701 34880
rect 19659 34831 19701 34840
rect 19756 33881 19796 35932
rect 20127 35888 20167 35897
rect 19852 35848 20127 35888
rect 19852 35561 19892 35848
rect 20127 35839 20167 35848
rect 20235 35804 20277 35813
rect 20235 35764 20236 35804
rect 20276 35764 20277 35804
rect 20235 35755 20277 35764
rect 19948 35720 19988 35729
rect 19851 35552 19893 35561
rect 19851 35512 19852 35552
rect 19892 35512 19893 35552
rect 19851 35503 19893 35512
rect 19851 35132 19893 35141
rect 19851 35092 19852 35132
rect 19892 35092 19893 35132
rect 19851 35083 19893 35092
rect 19852 34998 19892 35083
rect 19948 34553 19988 35680
rect 20236 35670 20276 35755
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 20044 34964 20084 34973
rect 19947 34544 19989 34553
rect 19947 34504 19948 34544
rect 19988 34504 19989 34544
rect 19947 34495 19989 34504
rect 19948 34397 19988 34406
rect 19851 34292 19893 34301
rect 19948 34292 19988 34357
rect 19851 34252 19852 34292
rect 19892 34252 19988 34292
rect 19851 34243 19893 34252
rect 20044 34208 20084 34924
rect 20140 34217 20180 34302
rect 19948 34168 20084 34208
rect 20139 34208 20181 34217
rect 20139 34168 20140 34208
rect 20180 34168 20181 34208
rect 19755 33872 19797 33881
rect 19755 33832 19756 33872
rect 19796 33832 19797 33872
rect 19755 33823 19797 33832
rect 19756 33620 19796 33629
rect 19948 33620 19988 34168
rect 20139 34159 20181 34168
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 19660 33580 19756 33620
rect 19660 33041 19700 33580
rect 19756 33571 19796 33580
rect 19852 33580 19988 33620
rect 19755 33200 19797 33209
rect 19755 33160 19756 33200
rect 19796 33160 19797 33200
rect 19755 33151 19797 33160
rect 19659 33032 19701 33041
rect 19659 32992 19660 33032
rect 19700 32992 19701 33032
rect 19659 32983 19701 32992
rect 19756 32948 19796 33151
rect 19756 32899 19796 32908
rect 19564 32824 19700 32864
rect 19371 32780 19413 32789
rect 19371 32740 19372 32780
rect 19412 32740 19413 32780
rect 19660 32780 19700 32824
rect 19660 32740 19796 32780
rect 19371 32731 19413 32740
rect 19564 32696 19604 32705
rect 19604 32656 19700 32696
rect 19564 32647 19604 32656
rect 18603 32528 18645 32537
rect 18603 32488 18604 32528
rect 18644 32488 18645 32528
rect 18603 32479 18645 32488
rect 18412 32320 18548 32360
rect 18412 32192 18452 32201
rect 18412 31613 18452 32152
rect 18411 31604 18453 31613
rect 18411 31564 18412 31604
rect 18452 31564 18453 31604
rect 18411 31555 18453 31564
rect 18411 31436 18453 31445
rect 18411 31396 18412 31436
rect 18452 31396 18453 31436
rect 18411 31387 18453 31396
rect 18412 29840 18452 31387
rect 18508 30773 18548 32320
rect 18604 32285 18644 32479
rect 19180 32360 19220 32369
rect 19220 32320 19508 32360
rect 19180 32311 19220 32320
rect 18603 32276 18645 32285
rect 18603 32236 18604 32276
rect 18644 32236 18645 32276
rect 18603 32227 18645 32236
rect 18604 32108 18644 32117
rect 18604 31865 18644 32068
rect 18988 32108 19028 32117
rect 19372 32108 19412 32119
rect 19028 32068 19316 32108
rect 18988 32059 19028 32068
rect 18796 31940 18836 31949
rect 18700 31900 18796 31940
rect 18603 31856 18645 31865
rect 18603 31816 18604 31856
rect 18644 31816 18645 31856
rect 18603 31807 18645 31816
rect 18700 31529 18740 31900
rect 18796 31891 18836 31900
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18795 31604 18837 31613
rect 18795 31564 18796 31604
rect 18836 31564 18837 31604
rect 18795 31555 18837 31564
rect 18699 31520 18741 31529
rect 18699 31480 18700 31520
rect 18740 31480 18741 31520
rect 18699 31471 18741 31480
rect 18604 31352 18644 31363
rect 18604 31277 18644 31312
rect 18603 31268 18645 31277
rect 18603 31228 18604 31268
rect 18644 31228 18645 31268
rect 18603 31219 18645 31228
rect 18796 31100 18836 31555
rect 18891 31436 18933 31445
rect 18891 31396 18892 31436
rect 18932 31396 18933 31436
rect 18891 31387 18933 31396
rect 18604 31060 18836 31100
rect 18507 30764 18549 30773
rect 18507 30724 18508 30764
rect 18548 30724 18549 30764
rect 18507 30715 18549 30724
rect 18412 29791 18452 29800
rect 18316 28624 18452 28664
rect 18220 28540 18261 28580
rect 18221 28496 18261 28540
rect 18221 28456 18278 28496
rect 18238 28412 18278 28456
rect 18412 28412 18452 28624
rect 18238 28372 18356 28412
rect 18412 28372 18463 28412
rect 18316 28328 18356 28372
rect 18423 28333 18463 28372
rect 18423 28293 18551 28333
rect 18316 28279 18356 28288
rect 18219 28244 18261 28253
rect 18511 28244 18551 28293
rect 18219 28204 18220 28244
rect 18260 28204 18261 28244
rect 18219 28195 18261 28204
rect 18508 28204 18551 28244
rect 18124 26095 18164 26104
rect 18220 25481 18260 28195
rect 18411 27236 18453 27245
rect 18411 27196 18412 27236
rect 18452 27196 18453 27236
rect 18411 27187 18453 27196
rect 18315 25724 18357 25733
rect 18315 25684 18316 25724
rect 18356 25684 18357 25724
rect 18315 25675 18357 25684
rect 18219 25472 18261 25481
rect 18028 25432 18164 25472
rect 17932 25348 18068 25388
rect 17739 25339 17781 25348
rect 17740 25304 17780 25339
rect 17740 25229 17780 25264
rect 17836 25304 17876 25313
rect 17739 25220 17781 25229
rect 17739 25180 17740 25220
rect 17780 25180 17781 25220
rect 17739 25171 17781 25180
rect 17836 25145 17876 25264
rect 17931 25220 17973 25229
rect 17931 25180 17932 25220
rect 17972 25180 17973 25220
rect 17931 25171 17973 25180
rect 17835 25136 17877 25145
rect 17835 25096 17836 25136
rect 17876 25096 17877 25136
rect 17835 25087 17877 25096
rect 17836 24632 17876 24641
rect 17644 24592 17836 24632
rect 17836 24583 17876 24592
rect 17452 24499 17492 24508
rect 17644 24464 17684 24473
rect 17932 24464 17972 25171
rect 17684 24424 17972 24464
rect 17644 24415 17684 24424
rect 17931 24296 17973 24305
rect 17931 24256 17932 24296
rect 17972 24256 17973 24296
rect 17931 24247 17973 24256
rect 17740 23792 17780 23803
rect 17740 23717 17780 23752
rect 17739 23708 17781 23717
rect 17739 23668 17740 23708
rect 17780 23668 17781 23708
rect 17739 23659 17781 23668
rect 17108 23248 17204 23288
rect 17260 23500 17396 23540
rect 17739 23540 17781 23549
rect 17739 23500 17740 23540
rect 17780 23500 17781 23540
rect 17068 23239 17108 23248
rect 16972 23071 17012 23080
rect 17164 23120 17204 23129
rect 16875 22700 16917 22709
rect 16875 22660 16876 22700
rect 16916 22660 16917 22700
rect 16875 22651 16917 22660
rect 17164 22541 17204 23080
rect 17163 22532 17205 22541
rect 16780 22492 17108 22532
rect 16587 22280 16629 22289
rect 16587 22240 16588 22280
rect 16628 22240 16629 22280
rect 16587 22231 16629 22240
rect 16779 22280 16821 22289
rect 16779 22240 16780 22280
rect 16820 22240 16821 22280
rect 16779 22231 16821 22240
rect 16780 21608 16820 22231
rect 16684 21568 16780 21608
rect 16491 20768 16533 20777
rect 16491 20728 16492 20768
rect 16532 20728 16533 20768
rect 16491 20719 16533 20728
rect 16588 20768 16628 20777
rect 16395 20684 16437 20693
rect 16395 20644 16396 20684
rect 16436 20644 16437 20684
rect 16395 20635 16437 20644
rect 16492 20634 16532 20719
rect 16395 20432 16437 20441
rect 16395 20392 16396 20432
rect 16436 20392 16437 20432
rect 16395 20383 16437 20392
rect 16396 19508 16436 20383
rect 16491 20348 16533 20357
rect 16491 20308 16492 20348
rect 16532 20308 16533 20348
rect 16491 20299 16533 20308
rect 16396 19459 16436 19468
rect 16299 19424 16341 19433
rect 16299 19384 16300 19424
rect 16340 19384 16341 19424
rect 16299 19375 16341 19384
rect 16204 18593 16244 19216
rect 16396 19088 16436 19097
rect 16300 19048 16396 19088
rect 16300 18761 16340 19048
rect 16396 19039 16436 19048
rect 16395 18920 16437 18929
rect 16395 18880 16396 18920
rect 16436 18880 16437 18920
rect 16395 18871 16437 18880
rect 16299 18752 16341 18761
rect 16299 18712 16300 18752
rect 16340 18712 16341 18752
rect 16299 18703 16341 18712
rect 16203 18584 16245 18593
rect 16300 18584 16340 18593
rect 16203 18544 16204 18584
rect 16244 18544 16300 18584
rect 16203 18535 16245 18544
rect 16300 18535 16340 18544
rect 16107 18416 16149 18425
rect 16107 18376 16108 18416
rect 16148 18376 16149 18416
rect 16107 18367 16149 18376
rect 16108 17744 16148 17753
rect 16204 17744 16244 18535
rect 16299 17996 16341 18005
rect 16299 17956 16300 17996
rect 16340 17956 16341 17996
rect 16396 17996 16436 18871
rect 16492 18668 16532 20299
rect 16588 19601 16628 20728
rect 16684 20273 16724 21568
rect 16780 21559 16820 21568
rect 16971 21524 17013 21533
rect 16971 21484 16972 21524
rect 17012 21484 17013 21524
rect 16971 21475 17013 21484
rect 16972 21356 17012 21475
rect 16876 21316 16972 21356
rect 16876 20777 16916 21316
rect 16972 21307 17012 21316
rect 16971 20936 17013 20945
rect 16971 20896 16972 20936
rect 17012 20896 17013 20936
rect 16971 20887 17013 20896
rect 16972 20852 17012 20887
rect 16972 20801 17012 20812
rect 17068 20852 17108 22492
rect 17163 22492 17164 22532
rect 17204 22492 17205 22532
rect 17163 22483 17205 22492
rect 17163 22280 17205 22289
rect 17163 22240 17164 22280
rect 17204 22240 17205 22280
rect 17163 22231 17205 22240
rect 17164 22146 17204 22231
rect 17163 21608 17205 21617
rect 17163 21568 17164 21608
rect 17204 21568 17205 21608
rect 17163 21559 17205 21568
rect 17164 21474 17204 21559
rect 17068 20803 17108 20812
rect 16875 20768 16917 20777
rect 16875 20728 16876 20768
rect 16916 20728 16917 20768
rect 16875 20719 16917 20728
rect 16779 20516 16821 20525
rect 16779 20476 16780 20516
rect 16820 20476 16821 20516
rect 16779 20467 16821 20476
rect 16683 20264 16725 20273
rect 16683 20224 16684 20264
rect 16724 20224 16725 20264
rect 16683 20215 16725 20224
rect 16587 19592 16629 19601
rect 16587 19552 16588 19592
rect 16628 19552 16629 19592
rect 16587 19543 16629 19552
rect 16588 19256 16628 19265
rect 16588 18845 16628 19216
rect 16684 19256 16724 19267
rect 16684 19181 16724 19216
rect 16683 19172 16725 19181
rect 16683 19132 16684 19172
rect 16724 19132 16725 19172
rect 16683 19123 16725 19132
rect 16587 18836 16629 18845
rect 16587 18796 16588 18836
rect 16628 18796 16629 18836
rect 16587 18787 16629 18796
rect 16780 18752 16820 20467
rect 16876 20105 16916 20719
rect 17260 20525 17300 23500
rect 17739 23491 17781 23500
rect 17355 23120 17397 23129
rect 17355 23080 17356 23120
rect 17396 23080 17397 23120
rect 17355 23071 17397 23080
rect 17356 22986 17396 23071
rect 17548 22280 17588 22289
rect 17355 22196 17397 22205
rect 17355 22156 17356 22196
rect 17396 22156 17397 22196
rect 17355 22147 17397 22156
rect 17356 22062 17396 22147
rect 17548 22121 17588 22240
rect 17547 22112 17589 22121
rect 17547 22072 17548 22112
rect 17588 22072 17589 22112
rect 17547 22063 17589 22072
rect 17644 22112 17684 22121
rect 17644 21785 17684 22072
rect 17643 21776 17685 21785
rect 17643 21736 17644 21776
rect 17684 21736 17685 21776
rect 17643 21727 17685 21736
rect 17355 21440 17397 21449
rect 17355 21400 17356 21440
rect 17396 21400 17397 21440
rect 17355 21391 17397 21400
rect 17259 20516 17301 20525
rect 17259 20476 17260 20516
rect 17300 20476 17301 20516
rect 17259 20467 17301 20476
rect 17259 20264 17301 20273
rect 17259 20224 17260 20264
rect 17300 20224 17301 20264
rect 17259 20215 17301 20224
rect 16875 20096 16917 20105
rect 16875 20056 16876 20096
rect 16916 20056 16917 20096
rect 16875 20047 16917 20056
rect 17260 20096 17300 20215
rect 17260 20047 17300 20056
rect 17259 19592 17301 19601
rect 17259 19552 17260 19592
rect 17300 19552 17301 19592
rect 17259 19543 17301 19552
rect 16971 19340 17013 19349
rect 16971 19300 16972 19340
rect 17012 19300 17013 19340
rect 16971 19291 17013 19300
rect 16875 19256 16917 19265
rect 16875 19216 16876 19256
rect 16916 19216 16917 19256
rect 16875 19207 16917 19216
rect 16972 19256 17012 19291
rect 16876 19122 16916 19207
rect 16972 19205 17012 19216
rect 17127 19256 17167 19265
rect 17167 19216 17204 19256
rect 17127 19207 17204 19216
rect 16972 19088 17012 19097
rect 16780 18712 16916 18752
rect 16492 18628 16628 18668
rect 16491 18416 16533 18425
rect 16491 18376 16492 18416
rect 16532 18376 16533 18416
rect 16491 18367 16533 18376
rect 16492 18282 16532 18367
rect 16492 17996 16532 18005
rect 16396 17956 16492 17996
rect 16299 17947 16341 17956
rect 16492 17947 16532 17956
rect 16300 17862 16340 17947
rect 16148 17704 16244 17744
rect 16299 17744 16341 17753
rect 16299 17704 16300 17744
rect 16340 17704 16341 17744
rect 16108 17695 16148 17704
rect 16299 17695 16341 17704
rect 16107 17576 16149 17585
rect 16107 17536 16108 17576
rect 16148 17536 16149 17576
rect 16107 17527 16149 17536
rect 16108 17324 16148 17527
rect 16108 17284 16244 17324
rect 16108 17072 16148 17081
rect 16012 17032 16108 17072
rect 16108 17023 16148 17032
rect 16204 16988 16244 17284
rect 15916 16948 16052 16988
rect 15724 16864 15860 16904
rect 15627 16484 15669 16493
rect 15627 16444 15628 16484
rect 15668 16444 15669 16484
rect 15627 16435 15669 16444
rect 15380 16192 15476 16232
rect 15340 16183 15380 16192
rect 15243 15980 15285 15989
rect 15243 15940 15244 15980
rect 15284 15940 15285 15980
rect 15243 15931 15285 15940
rect 15051 15812 15093 15821
rect 15051 15772 15052 15812
rect 15092 15772 15093 15812
rect 15051 15763 15093 15772
rect 14763 15728 14805 15737
rect 14763 15688 14764 15728
rect 14804 15688 14805 15728
rect 14763 15679 14805 15688
rect 14956 15728 14996 15737
rect 14764 15560 14804 15679
rect 14606 15545 14646 15554
rect 14764 15511 14804 15520
rect 14860 15560 14900 15569
rect 14606 15224 14646 15505
rect 14860 15317 14900 15520
rect 14859 15308 14901 15317
rect 14859 15268 14860 15308
rect 14900 15268 14901 15308
rect 14859 15259 14901 15268
rect 14572 15184 14646 15224
rect 14572 15065 14612 15184
rect 14763 15140 14805 15149
rect 14763 15100 14764 15140
rect 14804 15100 14805 15140
rect 14763 15091 14805 15100
rect 14571 15056 14613 15065
rect 14571 15016 14572 15056
rect 14612 15016 14613 15056
rect 14571 15007 14613 15016
rect 14667 14888 14709 14897
rect 14667 14848 14668 14888
rect 14708 14848 14709 14888
rect 14667 14839 14709 14848
rect 14091 12872 14133 12881
rect 14091 12832 14092 12872
rect 14132 12832 14133 12872
rect 14091 12823 14133 12832
rect 13900 12571 13940 12580
rect 13995 12620 14037 12629
rect 13995 12580 13996 12620
rect 14036 12580 14037 12620
rect 13995 12571 14037 12580
rect 13803 12536 13845 12545
rect 13803 12496 13804 12536
rect 13844 12496 13845 12536
rect 13803 12487 13845 12496
rect 13996 12536 14036 12571
rect 13804 12402 13844 12487
rect 13996 12486 14036 12496
rect 14092 12536 14132 12823
rect 13803 11444 13845 11453
rect 13803 11404 13804 11444
rect 13844 11404 13845 11444
rect 13803 11395 13845 11404
rect 13707 11360 13749 11369
rect 13707 11320 13708 11360
rect 13748 11320 13749 11360
rect 13707 11311 13749 11320
rect 13323 11276 13365 11285
rect 13323 11236 13324 11276
rect 13364 11236 13365 11276
rect 13323 11227 13365 11236
rect 13611 11192 13653 11201
rect 13611 11152 13612 11192
rect 13652 11152 13653 11192
rect 13611 11143 13653 11152
rect 13323 11108 13365 11117
rect 13323 11068 13324 11108
rect 13364 11068 13365 11108
rect 13323 11059 13365 11068
rect 13324 10193 13364 11059
rect 13228 9941 13268 10144
rect 13323 10184 13365 10193
rect 13323 10144 13324 10184
rect 13364 10144 13365 10184
rect 13323 10135 13365 10144
rect 13324 10050 13364 10135
rect 13227 9932 13269 9941
rect 13227 9892 13228 9932
rect 13268 9892 13269 9932
rect 13227 9883 13269 9892
rect 13227 9764 13269 9773
rect 13227 9724 13228 9764
rect 13268 9724 13269 9764
rect 13227 9715 13269 9724
rect 13228 9512 13268 9715
rect 13515 9596 13557 9605
rect 13515 9556 13516 9596
rect 13556 9556 13557 9596
rect 13515 9547 13557 9556
rect 13228 9463 13268 9472
rect 13516 9462 13556 9547
rect 13323 9428 13365 9437
rect 13323 9388 13324 9428
rect 13364 9388 13365 9428
rect 13323 9379 13365 9388
rect 13132 9304 13268 9344
rect 13036 9295 13076 9304
rect 12844 9136 13172 9176
rect 12651 9092 12693 9101
rect 12651 9052 12652 9092
rect 12692 9052 12693 9092
rect 12651 9043 12693 9052
rect 12555 8168 12597 8177
rect 12555 8128 12556 8168
rect 12596 8128 12597 8168
rect 12555 8119 12597 8128
rect 12364 7951 12404 7960
rect 12459 8000 12501 8009
rect 12459 7960 12460 8000
rect 12500 7960 12501 8000
rect 12459 7951 12501 7960
rect 12652 8000 12692 9043
rect 13132 8924 13172 9136
rect 13132 8875 13172 8884
rect 12747 8756 12789 8765
rect 13228 8756 13268 9304
rect 13324 8765 13364 9379
rect 13419 9008 13461 9017
rect 13419 8968 13420 9008
rect 13460 8968 13461 9008
rect 13419 8959 13461 8968
rect 12747 8716 12748 8756
rect 12788 8716 12789 8756
rect 12747 8707 12789 8716
rect 12940 8716 13268 8756
rect 13323 8756 13365 8765
rect 13323 8716 13324 8756
rect 13364 8716 13365 8756
rect 12748 8672 12788 8707
rect 12748 8621 12788 8632
rect 12844 8588 12884 8597
rect 12747 8504 12789 8513
rect 12747 8464 12748 8504
rect 12788 8464 12789 8504
rect 12747 8455 12789 8464
rect 12748 8168 12788 8455
rect 12844 8429 12884 8548
rect 12843 8420 12885 8429
rect 12843 8380 12844 8420
rect 12884 8380 12885 8420
rect 12843 8371 12885 8380
rect 12748 8119 12788 8128
rect 12652 7951 12692 7960
rect 12844 8000 12884 8009
rect 12940 8000 12980 8716
rect 13323 8707 13365 8716
rect 13420 8681 13460 8959
rect 13612 8840 13652 11143
rect 13707 10772 13749 10781
rect 13707 10732 13708 10772
rect 13748 10732 13749 10772
rect 13707 10723 13749 10732
rect 13708 10277 13748 10723
rect 13707 10268 13749 10277
rect 13707 10228 13708 10268
rect 13748 10228 13749 10268
rect 13707 10219 13749 10228
rect 13804 10268 13844 11395
rect 13899 11276 13941 11285
rect 13899 11236 13900 11276
rect 13940 11236 13941 11276
rect 13899 11227 13941 11236
rect 13804 10219 13844 10228
rect 13708 10134 13748 10219
rect 13803 10100 13845 10109
rect 13803 10060 13804 10100
rect 13844 10060 13845 10100
rect 13803 10051 13845 10060
rect 13707 9932 13749 9941
rect 13707 9892 13708 9932
rect 13748 9892 13749 9932
rect 13707 9883 13749 9892
rect 13708 9507 13748 9883
rect 13708 9458 13748 9467
rect 13516 8800 13652 8840
rect 13419 8672 13461 8681
rect 13419 8632 13420 8672
rect 13460 8632 13461 8672
rect 13419 8623 13461 8632
rect 13035 8588 13077 8597
rect 13035 8548 13036 8588
rect 13076 8548 13077 8588
rect 13035 8539 13077 8548
rect 12884 7960 12980 8000
rect 13036 8000 13076 8539
rect 13516 8504 13556 8800
rect 13611 8672 13653 8681
rect 13611 8632 13612 8672
rect 13652 8632 13653 8672
rect 13611 8623 13653 8632
rect 13612 8513 13652 8623
rect 12844 7951 12884 7960
rect 13036 7951 13076 7960
rect 13228 8464 13556 8504
rect 13611 8504 13653 8513
rect 13611 8464 13612 8504
rect 13652 8464 13653 8504
rect 12268 7832 12308 7841
rect 12172 7792 12268 7832
rect 12268 7783 12308 7792
rect 12267 7664 12309 7673
rect 12267 7624 12268 7664
rect 12308 7624 12309 7664
rect 12267 7615 12309 7624
rect 12075 7496 12117 7505
rect 12075 7456 12076 7496
rect 12116 7456 12117 7496
rect 12075 7447 12117 7456
rect 11924 6616 12020 6656
rect 12076 7160 12116 7447
rect 12268 7169 12308 7615
rect 12363 7580 12405 7589
rect 12363 7540 12364 7580
rect 12404 7540 12405 7580
rect 12363 7531 12405 7540
rect 11884 6607 11924 6616
rect 12076 6572 12116 7120
rect 12172 7160 12212 7169
rect 12172 7001 12212 7120
rect 12267 7160 12309 7169
rect 12267 7120 12268 7160
rect 12308 7120 12309 7160
rect 12267 7111 12309 7120
rect 12171 6992 12213 7001
rect 12171 6952 12172 6992
rect 12212 6952 12213 6992
rect 12171 6943 12213 6952
rect 11980 6532 12116 6572
rect 11884 5900 11924 5909
rect 11980 5900 12020 6532
rect 12076 6446 12116 6455
rect 12075 6406 12076 6413
rect 12116 6406 12117 6413
rect 12075 6404 12117 6406
rect 12075 6364 12076 6404
rect 12116 6364 12117 6404
rect 12075 6355 12117 6364
rect 12076 6311 12116 6355
rect 12172 6329 12212 6943
rect 12171 6320 12213 6329
rect 12171 6280 12172 6320
rect 12212 6280 12213 6320
rect 12171 6271 12213 6280
rect 11924 5860 12020 5900
rect 11884 5851 11924 5860
rect 11980 5657 12020 5860
rect 11979 5648 12021 5657
rect 11979 5608 11980 5648
rect 12020 5608 12021 5648
rect 11979 5599 12021 5608
rect 12172 5573 12212 5604
rect 12171 5564 12213 5573
rect 12171 5524 12172 5564
rect 12212 5524 12213 5564
rect 12171 5515 12213 5524
rect 12172 5480 12212 5515
rect 11788 5104 12020 5144
rect 11788 4976 11828 4985
rect 11596 4936 11788 4976
rect 11788 4927 11828 4936
rect 11883 4976 11925 4985
rect 11883 4936 11884 4976
rect 11924 4936 11925 4976
rect 11883 4927 11925 4936
rect 11499 4892 11541 4901
rect 11499 4852 11500 4892
rect 11540 4852 11541 4892
rect 11499 4843 11541 4852
rect 11403 4556 11445 4565
rect 11403 4516 11404 4556
rect 11444 4516 11445 4556
rect 11403 4507 11445 4516
rect 11307 4304 11349 4313
rect 11307 4264 11308 4304
rect 11348 4264 11349 4304
rect 11307 4255 11349 4264
rect 11211 4220 11253 4229
rect 11211 4180 11212 4220
rect 11252 4180 11253 4220
rect 11211 4171 11253 4180
rect 11116 4087 11156 4096
rect 11308 4136 11348 4255
rect 11308 4087 11348 4096
rect 11403 4136 11445 4145
rect 11403 4096 11404 4136
rect 11444 4096 11445 4136
rect 11403 4087 11445 4096
rect 10827 4052 10869 4061
rect 10827 4012 10828 4052
rect 10868 4012 10869 4052
rect 10827 4003 10869 4012
rect 10731 3884 10773 3893
rect 10731 3844 10732 3884
rect 10772 3844 10773 3884
rect 10731 3835 10773 3844
rect 10731 3380 10773 3389
rect 10731 3340 10732 3380
rect 10772 3340 10773 3380
rect 10731 3331 10773 3340
rect 10732 3246 10772 3331
rect 10635 2876 10677 2885
rect 10635 2836 10636 2876
rect 10676 2836 10677 2876
rect 10635 2827 10677 2836
rect 10731 2792 10773 2801
rect 10731 2752 10732 2792
rect 10772 2752 10773 2792
rect 10731 2743 10773 2752
rect 10539 1952 10581 1961
rect 10539 1912 10540 1952
rect 10580 1912 10581 1952
rect 10539 1903 10581 1912
rect 10540 1625 10580 1903
rect 10539 1616 10581 1625
rect 10539 1576 10540 1616
rect 10580 1576 10581 1616
rect 10539 1567 10581 1576
rect 10732 1205 10772 2743
rect 10828 2549 10868 4003
rect 10924 4002 10964 4087
rect 11404 4002 11444 4087
rect 11211 3968 11253 3977
rect 11211 3928 11212 3968
rect 11252 3928 11253 3968
rect 11211 3919 11253 3928
rect 11212 3834 11252 3919
rect 11500 3464 11540 4843
rect 11691 4556 11733 4565
rect 11691 4516 11692 4556
rect 11732 4516 11733 4556
rect 11691 4507 11733 4516
rect 11595 4220 11637 4229
rect 11595 4180 11596 4220
rect 11636 4180 11637 4220
rect 11595 4171 11637 4180
rect 11596 4086 11636 4171
rect 11692 4061 11732 4507
rect 11884 4145 11924 4927
rect 11980 4817 12020 5104
rect 11979 4808 12021 4817
rect 11979 4768 11980 4808
rect 12020 4768 12021 4808
rect 11979 4759 12021 4768
rect 12075 4724 12117 4733
rect 12075 4684 12076 4724
rect 12116 4684 12117 4724
rect 12075 4675 12117 4684
rect 12076 4145 12116 4675
rect 11883 4136 11925 4145
rect 12075 4136 12117 4145
rect 11883 4096 11884 4136
rect 11924 4096 12020 4136
rect 11883 4087 11925 4096
rect 11691 4052 11733 4061
rect 11691 4012 11692 4052
rect 11732 4012 11733 4052
rect 11691 4003 11733 4012
rect 11980 3977 12020 4096
rect 12075 4096 12076 4136
rect 12116 4096 12117 4136
rect 12075 4087 12117 4096
rect 12076 4002 12116 4087
rect 11595 3968 11637 3977
rect 11595 3928 11596 3968
rect 11636 3928 11637 3968
rect 11595 3919 11637 3928
rect 11788 3968 11828 3977
rect 11979 3968 12021 3977
rect 11828 3928 11924 3968
rect 11788 3919 11828 3928
rect 11116 3380 11156 3389
rect 10924 3212 10964 3221
rect 10827 2540 10869 2549
rect 10827 2500 10828 2540
rect 10868 2500 10869 2540
rect 10827 2491 10869 2500
rect 10924 1625 10964 3172
rect 11020 2624 11060 2633
rect 11020 2549 11060 2584
rect 11019 2540 11061 2549
rect 11019 2500 11020 2540
rect 11060 2500 11061 2540
rect 11019 2491 11061 2500
rect 11020 2213 11060 2491
rect 11019 2204 11061 2213
rect 11019 2164 11020 2204
rect 11060 2164 11061 2204
rect 11019 2155 11061 2164
rect 11116 1952 11156 3340
rect 11308 3212 11348 3221
rect 11212 2801 11252 2814
rect 11211 2792 11253 2801
rect 11211 2752 11212 2792
rect 11252 2752 11253 2792
rect 11211 2743 11253 2752
rect 11212 2719 11252 2743
rect 11212 2670 11252 2679
rect 11211 2540 11253 2549
rect 11211 2500 11212 2540
rect 11252 2500 11253 2540
rect 11211 2491 11253 2500
rect 11020 1912 11156 1952
rect 10923 1616 10965 1625
rect 10923 1576 10924 1616
rect 10964 1576 10965 1616
rect 10923 1567 10965 1576
rect 11020 1289 11060 1912
rect 11116 1364 11156 1373
rect 11212 1364 11252 2491
rect 11308 1457 11348 3172
rect 11500 2633 11540 3424
rect 11596 3464 11636 3919
rect 11691 3800 11733 3809
rect 11691 3760 11692 3800
rect 11732 3760 11733 3800
rect 11691 3751 11733 3760
rect 11596 3415 11636 3424
rect 11692 3464 11732 3751
rect 11692 3415 11732 3424
rect 11787 3464 11829 3473
rect 11787 3424 11788 3464
rect 11828 3424 11829 3464
rect 11787 3415 11829 3424
rect 11788 3330 11828 3415
rect 11787 3212 11829 3221
rect 11787 3172 11788 3212
rect 11828 3172 11829 3212
rect 11787 3163 11829 3172
rect 11595 2876 11637 2885
rect 11595 2836 11596 2876
rect 11636 2836 11637 2876
rect 11595 2827 11637 2836
rect 11499 2624 11541 2633
rect 11499 2584 11500 2624
rect 11540 2584 11541 2624
rect 11499 2575 11541 2584
rect 11404 2456 11444 2465
rect 11444 2416 11540 2456
rect 11404 2407 11444 2416
rect 11403 2120 11445 2129
rect 11403 2080 11404 2120
rect 11444 2080 11445 2120
rect 11403 2071 11445 2080
rect 11404 1952 11444 2071
rect 11404 1903 11444 1912
rect 11500 1793 11540 2416
rect 11596 1868 11636 2827
rect 11788 2708 11828 3163
rect 11884 2876 11924 3928
rect 11979 3928 11980 3968
rect 12020 3928 12021 3968
rect 11979 3919 12021 3928
rect 12075 3800 12117 3809
rect 12075 3760 12076 3800
rect 12116 3760 12117 3800
rect 12075 3751 12117 3760
rect 12076 3632 12116 3751
rect 12076 3583 12116 3592
rect 12075 3464 12117 3473
rect 12075 3424 12076 3464
rect 12116 3424 12117 3464
rect 12075 3415 12117 3424
rect 11884 2836 12020 2876
rect 11884 2708 11924 2717
rect 11788 2668 11884 2708
rect 11884 2659 11924 2668
rect 11980 2540 12020 2836
rect 12076 2637 12116 3415
rect 12172 3221 12212 5440
rect 12268 4976 12308 7111
rect 12364 6161 12404 7531
rect 12556 7160 12596 7171
rect 12556 7085 12596 7120
rect 12651 7160 12693 7169
rect 12651 7120 12652 7160
rect 12692 7120 12693 7160
rect 12651 7111 12693 7120
rect 13132 7160 13172 7169
rect 13228 7160 13268 8464
rect 13611 8455 13653 8464
rect 13804 8345 13844 10051
rect 13803 8336 13845 8345
rect 13803 8296 13804 8336
rect 13844 8296 13845 8336
rect 13803 8287 13845 8296
rect 13324 8000 13364 8009
rect 13516 8000 13556 8009
rect 13364 7960 13460 8000
rect 13324 7951 13364 7960
rect 13324 7748 13364 7757
rect 13324 7169 13364 7708
rect 13172 7120 13268 7160
rect 13323 7160 13365 7169
rect 13323 7120 13324 7160
rect 13364 7120 13365 7160
rect 13132 7111 13172 7120
rect 13323 7111 13365 7120
rect 12555 7076 12597 7085
rect 12555 7036 12556 7076
rect 12596 7036 12597 7076
rect 12555 7027 12597 7036
rect 12652 7026 12692 7111
rect 13420 7085 13460 7960
rect 13516 7505 13556 7960
rect 13612 8000 13652 8009
rect 13515 7496 13557 7505
rect 13515 7456 13516 7496
rect 13556 7456 13557 7496
rect 13515 7447 13557 7456
rect 13612 7421 13652 7960
rect 13708 8000 13748 8009
rect 13611 7412 13653 7421
rect 13611 7372 13612 7412
rect 13652 7372 13653 7412
rect 13611 7363 13653 7372
rect 13708 7337 13748 7960
rect 13804 8000 13844 8009
rect 13515 7328 13557 7337
rect 13515 7288 13516 7328
rect 13556 7288 13557 7328
rect 13515 7279 13557 7288
rect 13707 7328 13749 7337
rect 13707 7288 13708 7328
rect 13748 7288 13749 7328
rect 13707 7279 13749 7288
rect 13419 7076 13461 7085
rect 13419 7036 13420 7076
rect 13460 7036 13461 7076
rect 13419 7027 13461 7036
rect 12939 6656 12981 6665
rect 12939 6616 12940 6656
rect 12980 6616 12981 6656
rect 12939 6607 12981 6616
rect 13516 6656 13556 7279
rect 13612 7165 13652 7174
rect 13804 7160 13844 7960
rect 13900 7580 13940 11227
rect 14092 10940 14132 12496
rect 14188 11201 14228 13168
rect 14284 14764 14420 14804
rect 14571 14804 14613 14813
rect 14571 14764 14572 14804
rect 14612 14764 14613 14804
rect 14284 14048 14324 14764
rect 14571 14755 14613 14764
rect 14476 14720 14516 14729
rect 14476 14309 14516 14680
rect 14572 14670 14612 14755
rect 14668 14754 14708 14839
rect 14764 14804 14804 15091
rect 14764 14755 14804 14764
rect 14860 14720 14900 14729
rect 14956 14720 14996 15688
rect 15147 15644 15189 15653
rect 15147 15604 15148 15644
rect 15188 15604 15189 15644
rect 15147 15595 15189 15604
rect 15052 15560 15092 15571
rect 15052 15485 15092 15520
rect 15148 15560 15188 15595
rect 15051 15476 15093 15485
rect 15051 15436 15052 15476
rect 15092 15436 15093 15476
rect 15051 15427 15093 15436
rect 15148 15149 15188 15520
rect 15147 15140 15189 15149
rect 15147 15100 15148 15140
rect 15188 15100 15189 15140
rect 15147 15091 15189 15100
rect 15436 15065 15476 16192
rect 15435 15056 15477 15065
rect 15435 15016 15436 15056
rect 15476 15016 15477 15056
rect 15435 15007 15477 15016
rect 15628 14813 15668 16435
rect 15724 16316 15764 16864
rect 15916 16820 15956 16829
rect 15724 16267 15764 16276
rect 15819 16316 15861 16325
rect 15819 16276 15820 16316
rect 15860 16276 15861 16316
rect 15819 16267 15861 16276
rect 15820 16182 15860 16267
rect 15723 16064 15765 16073
rect 15723 16024 15724 16064
rect 15764 16024 15765 16064
rect 15723 16015 15765 16024
rect 15724 15560 15764 16015
rect 15916 15989 15956 16780
rect 15915 15980 15957 15989
rect 15915 15940 15916 15980
rect 15956 15940 15957 15980
rect 15915 15931 15957 15940
rect 15724 15511 15764 15520
rect 15819 15560 15861 15569
rect 15819 15520 15820 15560
rect 15860 15520 15861 15560
rect 15819 15511 15861 15520
rect 15820 15426 15860 15511
rect 15627 14804 15669 14813
rect 15627 14764 15628 14804
rect 15668 14764 15669 14804
rect 15627 14755 15669 14764
rect 14900 14680 14996 14720
rect 15340 14720 15380 14729
rect 14860 14671 14900 14680
rect 15051 14636 15093 14645
rect 15051 14596 15052 14636
rect 15092 14596 15093 14636
rect 15051 14587 15093 14596
rect 15052 14309 15092 14587
rect 14475 14300 14517 14309
rect 14475 14260 14476 14300
rect 14516 14260 14517 14300
rect 14475 14251 14517 14260
rect 15051 14300 15093 14309
rect 15051 14260 15052 14300
rect 15092 14260 15093 14300
rect 15340 14300 15380 14680
rect 15340 14260 15572 14300
rect 15051 14251 15093 14260
rect 14763 14216 14805 14225
rect 14763 14176 14764 14216
rect 14804 14176 14805 14216
rect 14763 14167 14805 14176
rect 14476 14132 14516 14143
rect 14476 14057 14516 14092
rect 14284 12797 14324 14008
rect 14475 14048 14517 14057
rect 14475 14008 14476 14048
rect 14516 14008 14517 14048
rect 14475 13999 14517 14008
rect 14668 14048 14708 14059
rect 14668 13973 14708 14008
rect 14764 14048 14804 14167
rect 14956 14132 14996 14141
rect 14996 14092 15092 14132
rect 14956 14083 14996 14092
rect 14764 13999 14804 14008
rect 14859 14048 14901 14057
rect 14859 14008 14860 14048
rect 14900 14008 14901 14048
rect 15052 14048 15092 14092
rect 15148 14048 15188 14057
rect 15052 14008 15148 14048
rect 14859 13999 14901 14008
rect 15148 13999 15188 14008
rect 15340 14048 15380 14057
rect 14667 13964 14709 13973
rect 14667 13924 14668 13964
rect 14708 13924 14709 13964
rect 14667 13915 14709 13924
rect 14475 13628 14517 13637
rect 14475 13588 14476 13628
rect 14516 13588 14517 13628
rect 14475 13579 14517 13588
rect 14283 12788 14325 12797
rect 14283 12748 14284 12788
rect 14324 12748 14325 12788
rect 14283 12739 14325 12748
rect 14476 12545 14516 13579
rect 14716 13217 14756 13226
rect 14860 13208 14900 13999
rect 15243 13964 15285 13973
rect 15340 13964 15380 14008
rect 15243 13924 15244 13964
rect 15284 13924 15380 13964
rect 15436 14048 15476 14057
rect 15243 13915 15285 13924
rect 15148 13796 15188 13805
rect 14756 13177 14900 13208
rect 14716 13168 14900 13177
rect 15052 13208 15092 13217
rect 15148 13208 15188 13756
rect 15243 13628 15285 13637
rect 15243 13588 15244 13628
rect 15284 13588 15285 13628
rect 15243 13579 15285 13588
rect 15092 13168 15188 13208
rect 15244 13208 15284 13579
rect 15436 13469 15476 14008
rect 15435 13460 15477 13469
rect 15435 13420 15436 13460
rect 15476 13420 15477 13460
rect 15435 13411 15477 13420
rect 15435 13292 15477 13301
rect 15532 13292 15572 14260
rect 16012 14216 16052 16948
rect 16204 16939 16244 16948
rect 16300 16904 16340 17695
rect 16491 17240 16533 17249
rect 16491 17200 16492 17240
rect 16532 17200 16533 17240
rect 16491 17191 16533 17200
rect 16492 17072 16532 17191
rect 16588 17072 16628 18628
rect 16779 18584 16821 18593
rect 16779 18544 16780 18584
rect 16820 18544 16821 18584
rect 16779 18535 16821 18544
rect 16780 18450 16820 18535
rect 16876 17912 16916 18712
rect 16972 18080 17012 19048
rect 17164 18845 17204 19207
rect 17163 18836 17205 18845
rect 17163 18796 17164 18836
rect 17204 18796 17205 18836
rect 17163 18787 17205 18796
rect 17068 18677 17108 18708
rect 17067 18668 17109 18677
rect 17067 18628 17068 18668
rect 17108 18628 17109 18668
rect 17067 18619 17109 18628
rect 17068 18584 17108 18619
rect 17164 18593 17204 18678
rect 17068 18509 17108 18544
rect 17163 18584 17205 18593
rect 17163 18544 17164 18584
rect 17204 18544 17205 18584
rect 17163 18535 17205 18544
rect 17067 18500 17109 18509
rect 17067 18460 17068 18500
rect 17108 18460 17109 18500
rect 17067 18451 17109 18460
rect 17163 18416 17205 18425
rect 17163 18376 17164 18416
rect 17204 18376 17205 18416
rect 17163 18367 17205 18376
rect 16972 18040 17108 18080
rect 16711 17872 16916 17912
rect 16971 17912 17013 17921
rect 16971 17872 16972 17912
rect 17012 17872 17013 17912
rect 16711 17828 16751 17872
rect 16971 17863 17013 17872
rect 16684 17788 16751 17828
rect 16684 17249 16724 17788
rect 16780 17744 16822 17753
rect 16780 17704 16781 17744
rect 16821 17704 16822 17744
rect 16780 17695 16822 17704
rect 16876 17744 16916 17755
rect 16780 17660 16820 17695
rect 16876 17669 16916 17704
rect 16780 17611 16820 17620
rect 16875 17660 16917 17669
rect 16875 17620 16876 17660
rect 16916 17620 16917 17660
rect 16875 17611 16917 17620
rect 16779 17492 16821 17501
rect 16779 17452 16780 17492
rect 16820 17452 16821 17492
rect 16779 17443 16821 17452
rect 16683 17240 16725 17249
rect 16683 17200 16684 17240
rect 16724 17200 16725 17240
rect 16683 17191 16725 17200
rect 16684 17072 16724 17081
rect 16588 17032 16684 17072
rect 16396 16988 16436 16999
rect 16396 16913 16436 16948
rect 16300 16855 16340 16864
rect 16395 16904 16437 16913
rect 16395 16864 16396 16904
rect 16436 16864 16437 16904
rect 16395 16855 16437 16864
rect 16299 16232 16341 16241
rect 16299 16192 16300 16232
rect 16340 16192 16341 16232
rect 16299 16183 16341 16192
rect 16300 16098 16340 16183
rect 16492 15728 16532 17032
rect 16684 17023 16724 17032
rect 16780 16988 16820 17443
rect 16780 16939 16820 16948
rect 16972 16988 17012 17863
rect 17068 17072 17108 18040
rect 17164 17744 17204 18367
rect 17164 17695 17204 17704
rect 17068 17023 17108 17032
rect 16972 16939 17012 16948
rect 16876 16904 16916 16913
rect 16876 16409 16916 16864
rect 17260 16409 17300 19543
rect 17356 19256 17396 21391
rect 17547 21356 17589 21365
rect 17547 21316 17548 21356
rect 17588 21316 17589 21356
rect 17547 21307 17589 21316
rect 17451 20768 17493 20777
rect 17451 20728 17452 20768
rect 17492 20728 17493 20768
rect 17451 20719 17493 20728
rect 17548 20768 17588 21307
rect 17643 21188 17685 21197
rect 17643 21148 17644 21188
rect 17684 21148 17685 21188
rect 17643 21139 17685 21148
rect 17452 20180 17492 20719
rect 17548 20189 17588 20728
rect 17452 20131 17492 20140
rect 17547 20180 17589 20189
rect 17547 20140 17548 20180
rect 17588 20140 17589 20180
rect 17547 20131 17589 20140
rect 17547 19592 17589 19601
rect 17547 19552 17548 19592
rect 17588 19552 17589 19592
rect 17547 19543 17589 19552
rect 17548 19508 17588 19543
rect 17548 19457 17588 19468
rect 17451 19340 17493 19349
rect 17451 19300 17452 19340
rect 17492 19300 17493 19340
rect 17451 19291 17493 19300
rect 17356 19207 17396 19216
rect 17452 19004 17492 19291
rect 17547 19256 17589 19265
rect 17547 19216 17548 19256
rect 17588 19216 17589 19256
rect 17547 19207 17589 19216
rect 17548 19122 17588 19207
rect 17452 18964 17588 19004
rect 17451 18836 17493 18845
rect 17451 18796 17452 18836
rect 17492 18796 17493 18836
rect 17451 18787 17493 18796
rect 17355 18500 17397 18509
rect 17355 18460 17356 18500
rect 17396 18460 17397 18500
rect 17355 18451 17397 18460
rect 17356 17249 17396 18451
rect 17452 18416 17492 18787
rect 17452 18367 17492 18376
rect 17451 18248 17493 18257
rect 17451 18208 17452 18248
rect 17492 18208 17493 18248
rect 17451 18199 17493 18208
rect 17452 17744 17492 18199
rect 17548 17996 17588 18964
rect 17548 17947 17588 17956
rect 17452 17695 17492 17704
rect 17355 17240 17397 17249
rect 17355 17200 17356 17240
rect 17396 17200 17397 17240
rect 17355 17191 17397 17200
rect 17356 17072 17396 17083
rect 17356 16997 17396 17032
rect 17355 16988 17397 16997
rect 17355 16948 17356 16988
rect 17396 16948 17397 16988
rect 17355 16939 17397 16948
rect 16875 16400 16917 16409
rect 16875 16360 16876 16400
rect 16916 16360 16917 16400
rect 16875 16351 16917 16360
rect 17259 16400 17301 16409
rect 17259 16360 17260 16400
rect 17300 16360 17301 16400
rect 17259 16351 17301 16360
rect 16780 16237 16820 16246
rect 16780 16073 16820 16197
rect 17260 16232 17300 16241
rect 17452 16232 17492 16241
rect 17300 16192 17396 16232
rect 17260 16183 17300 16192
rect 16779 16064 16821 16073
rect 16779 16024 16780 16064
rect 16820 16024 16821 16064
rect 16779 16015 16821 16024
rect 16972 16064 17012 16073
rect 16875 15896 16917 15905
rect 16875 15856 16876 15896
rect 16916 15856 16917 15896
rect 16875 15847 16917 15856
rect 16492 15688 16820 15728
rect 16203 15560 16245 15569
rect 16203 15520 16204 15560
rect 16244 15520 16245 15560
rect 16203 15511 16245 15520
rect 16780 15560 16820 15688
rect 16780 15511 16820 15520
rect 16204 15426 16244 15511
rect 16300 15476 16340 15485
rect 16300 15317 16340 15436
rect 16683 15476 16725 15485
rect 16683 15436 16684 15476
rect 16724 15436 16725 15476
rect 16683 15427 16725 15436
rect 16395 15392 16437 15401
rect 16395 15352 16396 15392
rect 16436 15352 16437 15392
rect 16395 15343 16437 15352
rect 16299 15308 16341 15317
rect 16299 15268 16300 15308
rect 16340 15268 16341 15308
rect 16299 15259 16341 15268
rect 16396 15233 16436 15343
rect 16395 15224 16437 15233
rect 16395 15184 16396 15224
rect 16436 15184 16437 15224
rect 16395 15175 16437 15184
rect 16299 15140 16341 15149
rect 16299 15100 16300 15140
rect 16340 15100 16341 15140
rect 16299 15091 16341 15100
rect 16300 14393 16340 15091
rect 16587 14972 16629 14981
rect 16587 14932 16588 14972
rect 16628 14932 16629 14972
rect 16587 14923 16629 14932
rect 16491 14720 16533 14729
rect 16491 14680 16492 14720
rect 16532 14680 16533 14720
rect 16491 14671 16533 14680
rect 16588 14720 16628 14923
rect 16588 14671 16628 14680
rect 16299 14384 16341 14393
rect 16299 14344 16300 14384
rect 16340 14344 16341 14384
rect 16299 14335 16341 14344
rect 16204 14216 16244 14225
rect 16012 14176 16204 14216
rect 16204 14167 16244 14176
rect 15627 14048 15669 14057
rect 15627 14008 15628 14048
rect 15668 14008 15669 14048
rect 15627 13999 15669 14008
rect 15724 14048 15764 14057
rect 15628 13914 15668 13999
rect 15724 13889 15764 14008
rect 15820 14048 15860 14057
rect 15723 13880 15765 13889
rect 15723 13840 15724 13880
rect 15764 13840 15765 13880
rect 15723 13831 15765 13840
rect 15627 13460 15669 13469
rect 15627 13420 15628 13460
rect 15668 13420 15669 13460
rect 15627 13411 15669 13420
rect 15435 13252 15436 13292
rect 15476 13252 15572 13292
rect 15435 13243 15477 13252
rect 15052 13159 15092 13168
rect 15244 13159 15284 13168
rect 15339 13208 15381 13217
rect 15339 13168 15340 13208
rect 15380 13168 15381 13208
rect 15339 13159 15381 13168
rect 15436 13208 15476 13243
rect 14859 13040 14901 13049
rect 14859 13000 14860 13040
rect 14900 13000 14901 13040
rect 14859 12991 14901 13000
rect 15148 13040 15188 13049
rect 15340 13040 15380 13159
rect 15436 13157 15476 13168
rect 15188 13000 15380 13040
rect 15148 12991 15188 13000
rect 14860 12906 14900 12991
rect 15243 12872 15285 12881
rect 15243 12832 15244 12872
rect 15284 12832 15285 12872
rect 15243 12823 15285 12832
rect 14571 12788 14613 12797
rect 14571 12748 14572 12788
rect 14612 12748 14613 12788
rect 14571 12739 14613 12748
rect 14284 12536 14324 12545
rect 14284 12041 14324 12496
rect 14475 12536 14517 12545
rect 14475 12496 14476 12536
rect 14516 12496 14517 12536
rect 14475 12487 14517 12496
rect 14283 12032 14325 12041
rect 14283 11992 14284 12032
rect 14324 11992 14325 12032
rect 14283 11983 14325 11992
rect 14283 11864 14325 11873
rect 14283 11824 14284 11864
rect 14324 11824 14325 11864
rect 14283 11815 14325 11824
rect 14187 11192 14229 11201
rect 14187 11152 14188 11192
rect 14228 11152 14229 11192
rect 14187 11143 14229 11152
rect 13996 10900 14132 10940
rect 14284 11024 14324 11815
rect 14476 11369 14516 12487
rect 14572 12461 14612 12739
rect 14571 12452 14613 12461
rect 14571 12412 14572 12452
rect 14612 12412 14613 12452
rect 14571 12403 14613 12412
rect 14571 12116 14613 12125
rect 14571 12076 14572 12116
rect 14612 12076 14613 12116
rect 14571 12067 14613 12076
rect 14572 11696 14612 12067
rect 15051 11948 15093 11957
rect 15051 11908 15052 11948
rect 15092 11908 15093 11948
rect 15051 11899 15093 11908
rect 14668 11696 14708 11724
rect 14572 11656 14668 11696
rect 14475 11360 14517 11369
rect 14475 11320 14476 11360
rect 14516 11320 14517 11360
rect 14475 11311 14517 11320
rect 13996 9260 14036 10900
rect 14284 10781 14324 10984
rect 14572 10940 14612 11656
rect 14668 11647 14708 11656
rect 15052 11696 15092 11899
rect 15052 11647 15092 11656
rect 15147 11696 15189 11705
rect 15147 11656 15148 11696
rect 15188 11656 15189 11696
rect 15147 11647 15189 11656
rect 14860 11528 14900 11537
rect 14860 11033 14900 11488
rect 15051 11360 15093 11369
rect 15051 11320 15052 11360
rect 15092 11320 15093 11360
rect 15051 11311 15093 11320
rect 14859 11024 14901 11033
rect 14859 10984 14860 11024
rect 14900 10984 14901 11024
rect 14859 10975 14901 10984
rect 15052 11024 15092 11311
rect 14380 10900 14612 10940
rect 14283 10772 14325 10781
rect 14283 10732 14284 10772
rect 14324 10732 14325 10772
rect 14283 10723 14325 10732
rect 14091 10268 14133 10277
rect 14091 10228 14092 10268
rect 14132 10228 14133 10268
rect 14091 10219 14133 10228
rect 14092 9344 14132 10219
rect 14284 10184 14324 10195
rect 14284 10109 14324 10144
rect 14283 10100 14325 10109
rect 14283 10060 14284 10100
rect 14324 10060 14325 10100
rect 14283 10051 14325 10060
rect 14187 9764 14229 9773
rect 14187 9724 14188 9764
rect 14228 9724 14229 9764
rect 14187 9715 14229 9724
rect 14188 9512 14228 9715
rect 14188 9463 14228 9472
rect 14092 9304 14324 9344
rect 13996 9220 14132 9260
rect 13995 8756 14037 8765
rect 13995 8716 13996 8756
rect 14036 8716 14037 8756
rect 13995 8707 14037 8716
rect 13996 8000 14036 8707
rect 14092 8345 14132 9220
rect 14091 8336 14133 8345
rect 14091 8296 14092 8336
rect 14132 8296 14133 8336
rect 14091 8287 14133 8296
rect 14091 8168 14133 8177
rect 14091 8128 14092 8168
rect 14132 8128 14133 8168
rect 14091 8119 14133 8128
rect 14092 8034 14132 8119
rect 13996 7951 14036 7960
rect 14187 8000 14229 8009
rect 14187 7960 14188 8000
rect 14228 7960 14229 8000
rect 14187 7951 14229 7960
rect 14188 7866 14228 7951
rect 13900 7540 14132 7580
rect 13995 7412 14037 7421
rect 13995 7372 13996 7412
rect 14036 7372 14037 7412
rect 13995 7363 14037 7372
rect 13996 7278 14036 7363
rect 13612 7085 13652 7125
rect 13708 7120 13844 7160
rect 13995 7160 14037 7169
rect 13995 7120 13996 7160
rect 14036 7120 14037 7160
rect 13611 7076 13653 7085
rect 13611 7036 13612 7076
rect 13652 7036 13653 7076
rect 13611 7027 13653 7036
rect 13708 6824 13748 7120
rect 13995 7111 14037 7120
rect 13899 7076 13941 7085
rect 13899 7036 13900 7076
rect 13940 7036 13941 7076
rect 13899 7027 13941 7036
rect 12843 6488 12885 6497
rect 12843 6448 12844 6488
rect 12884 6448 12885 6488
rect 12843 6439 12885 6448
rect 12363 6152 12405 6161
rect 12363 6112 12364 6152
rect 12404 6112 12405 6152
rect 12363 6103 12405 6112
rect 12459 5900 12501 5909
rect 12459 5860 12460 5900
rect 12500 5860 12501 5900
rect 12459 5851 12501 5860
rect 12364 5648 12404 5657
rect 12364 5237 12404 5608
rect 12460 5648 12500 5851
rect 12460 5405 12500 5608
rect 12556 5648 12596 5657
rect 12459 5396 12501 5405
rect 12459 5356 12460 5396
rect 12500 5356 12501 5396
rect 12459 5347 12501 5356
rect 12363 5228 12405 5237
rect 12363 5188 12364 5228
rect 12404 5188 12405 5228
rect 12363 5179 12405 5188
rect 12556 5060 12596 5608
rect 12844 5489 12884 6439
rect 12940 5648 12980 6607
rect 13516 6581 13556 6616
rect 13612 6784 13748 6824
rect 13804 6992 13844 7001
rect 13515 6572 13557 6581
rect 13515 6532 13516 6572
rect 13556 6532 13557 6572
rect 13515 6523 13557 6532
rect 13323 6488 13365 6497
rect 13516 6492 13556 6523
rect 13323 6448 13324 6488
rect 13364 6448 13365 6488
rect 13323 6439 13365 6448
rect 13227 6404 13269 6413
rect 13227 6364 13228 6404
rect 13268 6364 13269 6404
rect 13227 6355 13269 6364
rect 12940 5599 12980 5608
rect 13035 5648 13077 5657
rect 13035 5608 13036 5648
rect 13076 5608 13077 5648
rect 13035 5599 13077 5608
rect 13132 5648 13172 5657
rect 13036 5514 13076 5599
rect 12652 5480 12692 5489
rect 12843 5480 12885 5489
rect 12692 5440 12788 5480
rect 12652 5431 12692 5440
rect 12651 5228 12693 5237
rect 12651 5188 12652 5228
rect 12692 5188 12693 5228
rect 12748 5228 12788 5440
rect 12843 5440 12844 5480
rect 12884 5440 12885 5480
rect 12843 5431 12885 5440
rect 13132 5405 13172 5608
rect 13228 5648 13268 6355
rect 13324 6354 13364 6439
rect 13419 6236 13461 6245
rect 13419 6196 13420 6236
rect 13460 6196 13461 6236
rect 13419 6187 13461 6196
rect 13323 5900 13365 5909
rect 13323 5860 13324 5900
rect 13364 5860 13365 5900
rect 13323 5851 13365 5860
rect 13324 5741 13364 5851
rect 13323 5732 13365 5741
rect 13323 5692 13324 5732
rect 13364 5692 13365 5732
rect 13323 5683 13365 5692
rect 13131 5396 13173 5405
rect 13131 5356 13132 5396
rect 13172 5356 13173 5396
rect 13131 5347 13173 5356
rect 12748 5188 13172 5228
rect 12651 5179 12693 5188
rect 12460 5020 12596 5060
rect 12268 4927 12308 4936
rect 12363 4976 12405 4985
rect 12363 4936 12364 4976
rect 12404 4936 12405 4976
rect 12363 4927 12405 4936
rect 12364 4842 12404 4927
rect 12460 4901 12500 5020
rect 12652 4985 12692 5179
rect 12651 4976 12693 4985
rect 12651 4936 12652 4976
rect 12692 4936 12693 4976
rect 12651 4927 12693 4936
rect 12748 4976 12788 4985
rect 12748 4901 12788 4936
rect 12843 4976 12885 4985
rect 12843 4936 12844 4976
rect 12884 4936 12885 4976
rect 12843 4927 12885 4936
rect 13132 4976 13172 5188
rect 13132 4927 13172 4936
rect 12459 4892 12501 4901
rect 12459 4852 12460 4892
rect 12500 4852 12501 4892
rect 12459 4843 12501 4852
rect 12747 4892 12789 4901
rect 12747 4852 12748 4892
rect 12788 4852 12789 4892
rect 12747 4843 12789 4852
rect 12555 4808 12597 4817
rect 12555 4768 12556 4808
rect 12596 4768 12597 4808
rect 12555 4759 12597 4768
rect 12363 4724 12405 4733
rect 12363 4684 12364 4724
rect 12404 4684 12405 4724
rect 12363 4675 12405 4684
rect 12268 3464 12308 3475
rect 12268 3389 12308 3424
rect 12267 3380 12309 3389
rect 12267 3340 12268 3380
rect 12308 3340 12309 3380
rect 12267 3331 12309 3340
rect 12171 3212 12213 3221
rect 12171 3172 12172 3212
rect 12212 3172 12213 3212
rect 12171 3163 12213 3172
rect 12171 2708 12213 2717
rect 12171 2668 12172 2708
rect 12212 2668 12213 2708
rect 12171 2659 12213 2668
rect 12076 2588 12116 2597
rect 12172 2574 12212 2659
rect 12268 2624 12308 2633
rect 12364 2624 12404 4675
rect 12459 4556 12501 4565
rect 12459 4516 12460 4556
rect 12500 4516 12501 4556
rect 12459 4507 12501 4516
rect 12460 2717 12500 4507
rect 12459 2708 12501 2717
rect 12459 2668 12460 2708
rect 12500 2668 12501 2708
rect 12459 2659 12501 2668
rect 12308 2584 12404 2624
rect 12268 2575 12308 2584
rect 11980 2500 12116 2540
rect 11596 1819 11636 1828
rect 11692 2456 11732 2465
rect 11499 1784 11541 1793
rect 11499 1744 11500 1784
rect 11540 1744 11541 1784
rect 11499 1735 11541 1744
rect 11595 1616 11637 1625
rect 11595 1576 11596 1616
rect 11636 1576 11637 1616
rect 11595 1567 11637 1576
rect 11307 1448 11349 1457
rect 11307 1408 11308 1448
rect 11348 1408 11349 1448
rect 11307 1399 11349 1408
rect 11156 1324 11252 1364
rect 11116 1315 11156 1324
rect 11019 1280 11061 1289
rect 11019 1240 11020 1280
rect 11060 1240 11061 1280
rect 11019 1231 11061 1240
rect 10731 1196 10773 1205
rect 10731 1156 10732 1196
rect 10772 1156 10773 1196
rect 10731 1147 10773 1156
rect 10924 1112 10964 1121
rect 10924 365 10964 1072
rect 11308 1112 11348 1121
rect 11211 944 11253 953
rect 11211 904 11212 944
rect 11252 904 11253 944
rect 11211 895 11253 904
rect 11019 524 11061 533
rect 11019 484 11020 524
rect 11060 484 11061 524
rect 11019 475 11061 484
rect 10923 356 10965 365
rect 10923 316 10924 356
rect 10964 316 10965 356
rect 10923 307 10965 316
rect 10635 272 10677 281
rect 10635 232 10636 272
rect 10676 232 10677 272
rect 10635 223 10677 232
rect 10636 80 10676 223
rect 10827 104 10869 113
rect 10827 80 10828 104
rect 5108 64 5128 80
rect 5048 0 5128 64
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 0 8008 80
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 64 10828 80
rect 10868 80 10869 104
rect 11020 80 11060 475
rect 11212 80 11252 895
rect 11308 524 11348 1072
rect 11308 484 11540 524
rect 11500 281 11540 484
rect 11499 272 11541 281
rect 11499 232 11500 272
rect 11540 232 11541 272
rect 11499 223 11541 232
rect 11403 188 11445 197
rect 11403 148 11404 188
rect 11444 148 11445 188
rect 11403 139 11445 148
rect 11404 80 11444 139
rect 11596 80 11636 1567
rect 11692 1364 11732 2416
rect 11979 2288 12021 2297
rect 11979 2248 11980 2288
rect 12020 2248 12021 2288
rect 11979 2239 12021 2248
rect 11980 2120 12020 2239
rect 11980 2071 12020 2080
rect 11788 1700 11828 1709
rect 11788 1541 11828 1660
rect 11787 1532 11829 1541
rect 11787 1492 11788 1532
rect 11828 1492 11829 1532
rect 11787 1483 11829 1492
rect 11692 1324 11828 1364
rect 11788 80 11828 1324
rect 12076 1280 12116 2500
rect 12460 2456 12500 2465
rect 12171 2372 12213 2381
rect 12171 2332 12172 2372
rect 12212 2332 12213 2372
rect 12171 2323 12213 2332
rect 12172 2129 12212 2323
rect 12460 2213 12500 2416
rect 12556 2381 12596 4759
rect 12748 2969 12788 4843
rect 12844 4313 12884 4927
rect 13131 4724 13173 4733
rect 13131 4684 13132 4724
rect 13172 4684 13173 4724
rect 13131 4675 13173 4684
rect 13132 4590 13172 4675
rect 13131 4388 13173 4397
rect 13131 4348 13132 4388
rect 13172 4348 13173 4388
rect 13228 4388 13268 5608
rect 13420 5648 13460 6187
rect 13515 5732 13557 5741
rect 13515 5692 13516 5732
rect 13556 5692 13557 5732
rect 13515 5683 13557 5692
rect 13420 5599 13460 5608
rect 13516 5598 13556 5683
rect 13612 5648 13652 6784
rect 13707 6656 13749 6665
rect 13707 6616 13708 6656
rect 13748 6616 13749 6656
rect 13707 6607 13749 6616
rect 13708 6488 13748 6607
rect 13804 6497 13844 6952
rect 13708 6439 13748 6448
rect 13803 6488 13845 6497
rect 13803 6448 13804 6488
rect 13844 6448 13845 6488
rect 13803 6439 13845 6448
rect 13900 6488 13940 7027
rect 13996 7026 14036 7111
rect 13900 6413 13940 6448
rect 13996 6488 14036 6497
rect 13899 6404 13941 6413
rect 13899 6364 13900 6404
rect 13940 6364 13941 6404
rect 13899 6355 13941 6364
rect 13707 6236 13749 6245
rect 13707 6196 13708 6236
rect 13748 6196 13749 6236
rect 13707 6187 13749 6196
rect 13708 6102 13748 6187
rect 13899 5900 13941 5909
rect 13899 5860 13900 5900
rect 13940 5860 13941 5900
rect 13899 5851 13941 5860
rect 13612 5599 13652 5608
rect 13900 5648 13940 5851
rect 13900 5599 13940 5608
rect 13419 5480 13461 5489
rect 13419 5440 13420 5480
rect 13460 5440 13461 5480
rect 13419 5431 13461 5440
rect 13803 5480 13845 5489
rect 13996 5480 14036 6448
rect 14092 5825 14132 7540
rect 14188 7160 14228 7171
rect 14188 7085 14228 7120
rect 14284 7160 14324 9304
rect 14380 7505 14420 10900
rect 14860 10890 14900 10975
rect 14476 10772 14516 10781
rect 14764 10772 14804 10781
rect 14516 10732 14708 10772
rect 14476 10723 14516 10732
rect 14668 10268 14708 10732
rect 14764 10445 14804 10732
rect 14859 10772 14901 10781
rect 14859 10732 14860 10772
rect 14900 10732 14901 10772
rect 14859 10723 14901 10732
rect 14763 10436 14805 10445
rect 14763 10396 14764 10436
rect 14804 10396 14805 10436
rect 14763 10387 14805 10396
rect 14668 10228 14804 10268
rect 14571 10100 14613 10109
rect 14571 10060 14572 10100
rect 14612 10060 14613 10100
rect 14571 10051 14613 10060
rect 14475 9596 14517 9605
rect 14475 9556 14476 9596
rect 14516 9556 14517 9596
rect 14475 9547 14517 9556
rect 14476 8177 14516 9547
rect 14572 8588 14612 10051
rect 14668 9605 14708 10228
rect 14764 10198 14804 10228
rect 14764 10149 14804 10158
rect 14763 9932 14805 9941
rect 14763 9892 14764 9932
rect 14804 9892 14805 9932
rect 14763 9883 14805 9892
rect 14667 9596 14709 9605
rect 14667 9556 14668 9596
rect 14708 9556 14709 9596
rect 14667 9547 14709 9556
rect 14764 9512 14804 9883
rect 14764 9463 14804 9472
rect 14668 9428 14708 9437
rect 14668 9185 14708 9388
rect 14667 9176 14709 9185
rect 14667 9136 14668 9176
rect 14708 9136 14709 9176
rect 14667 9127 14709 9136
rect 14860 8840 14900 10723
rect 15052 10277 15092 10984
rect 15148 10352 15188 11647
rect 15244 10529 15284 12823
rect 15628 12704 15668 13411
rect 15436 12664 15668 12704
rect 15436 12293 15476 12664
rect 15724 12620 15764 12629
rect 15820 12620 15860 14008
rect 15916 14048 15956 14057
rect 15916 13637 15956 14008
rect 16108 14048 16148 14057
rect 16300 14048 16340 14057
rect 16011 13880 16053 13889
rect 16011 13840 16012 13880
rect 16052 13840 16053 13880
rect 16011 13831 16053 13840
rect 15915 13628 15957 13637
rect 15915 13588 15916 13628
rect 15956 13588 15957 13628
rect 15915 13579 15957 13588
rect 15764 12580 15956 12620
rect 15724 12571 15764 12580
rect 15532 12536 15572 12547
rect 15532 12461 15572 12496
rect 15916 12536 15956 12580
rect 15916 12487 15956 12496
rect 15531 12452 15573 12461
rect 15531 12412 15532 12452
rect 15572 12412 15573 12452
rect 15531 12403 15573 12412
rect 16012 12368 16052 13831
rect 16108 13217 16148 14008
rect 16204 14008 16300 14048
rect 16107 13208 16149 13217
rect 16107 13168 16108 13208
rect 16148 13168 16149 13208
rect 16107 13159 16149 13168
rect 16107 13040 16149 13049
rect 16107 13000 16108 13040
rect 16148 13000 16149 13040
rect 16107 12991 16149 13000
rect 16108 12536 16148 12991
rect 16108 12487 16148 12496
rect 15628 12328 16052 12368
rect 16108 12368 16148 12377
rect 16204 12368 16244 14008
rect 16300 13999 16340 14008
rect 16492 14048 16532 14671
rect 16588 14216 16628 14225
rect 16684 14216 16724 15427
rect 16779 14636 16821 14645
rect 16779 14596 16780 14636
rect 16820 14596 16821 14636
rect 16779 14587 16821 14596
rect 16780 14502 16820 14587
rect 16876 14552 16916 15847
rect 16972 15401 17012 16024
rect 17164 16064 17204 16073
rect 16971 15392 17013 15401
rect 16971 15352 16972 15392
rect 17012 15352 17013 15392
rect 16971 15343 17013 15352
rect 16971 15140 17013 15149
rect 16971 15100 16972 15140
rect 17012 15100 17013 15140
rect 16971 15091 17013 15100
rect 16972 14972 17012 15091
rect 17164 14981 17204 16024
rect 17259 15980 17301 15989
rect 17259 15940 17260 15980
rect 17300 15940 17301 15980
rect 17259 15931 17301 15940
rect 17260 15555 17300 15931
rect 17260 15506 17300 15515
rect 17259 15392 17301 15401
rect 17259 15352 17260 15392
rect 17300 15352 17301 15392
rect 17259 15343 17301 15352
rect 16972 14923 17012 14932
rect 17163 14972 17205 14981
rect 17163 14932 17164 14972
rect 17204 14932 17205 14972
rect 17163 14923 17205 14932
rect 17260 14888 17300 15343
rect 17356 14897 17396 16192
rect 17452 15821 17492 16192
rect 17451 15812 17493 15821
rect 17451 15772 17452 15812
rect 17492 15772 17493 15812
rect 17644 15812 17684 21139
rect 17740 19928 17780 23491
rect 17836 22280 17876 22289
rect 17836 22037 17876 22240
rect 17835 22028 17877 22037
rect 17835 21988 17836 22028
rect 17876 21988 17877 22028
rect 17835 21979 17877 21988
rect 17932 21197 17972 24247
rect 18028 23549 18068 25348
rect 18124 25304 18164 25432
rect 18219 25432 18220 25472
rect 18260 25432 18261 25472
rect 18219 25423 18261 25432
rect 18316 25304 18356 25675
rect 18124 25264 18260 25304
rect 18123 25136 18165 25145
rect 18123 25096 18124 25136
rect 18164 25096 18165 25136
rect 18123 25087 18165 25096
rect 18027 23540 18069 23549
rect 18027 23500 18028 23540
rect 18068 23500 18069 23540
rect 18027 23491 18069 23500
rect 18124 22625 18164 25087
rect 18220 23792 18260 25264
rect 18316 25255 18356 25264
rect 18412 24893 18452 27187
rect 18508 26816 18548 28204
rect 18508 26405 18548 26776
rect 18507 26396 18549 26405
rect 18507 26356 18508 26396
rect 18548 26356 18549 26396
rect 18507 26347 18549 26356
rect 18507 26228 18549 26237
rect 18507 26188 18508 26228
rect 18548 26188 18549 26228
rect 18507 26179 18549 26188
rect 18508 25481 18548 26179
rect 18507 25472 18549 25481
rect 18507 25432 18508 25472
rect 18548 25432 18549 25472
rect 18507 25423 18549 25432
rect 18604 25397 18644 31060
rect 18699 30680 18741 30689
rect 18699 30640 18700 30680
rect 18740 30640 18741 30680
rect 18699 30631 18741 30640
rect 18700 29168 18740 30631
rect 18892 30437 18932 31387
rect 19132 31361 19172 31370
rect 19172 31321 19220 31352
rect 19132 31312 19220 31321
rect 19180 30857 19220 31312
rect 19276 31268 19316 32068
rect 19372 32033 19412 32068
rect 19371 32024 19413 32033
rect 19371 31984 19372 32024
rect 19412 31984 19413 32024
rect 19371 31975 19413 31984
rect 19468 31604 19508 32320
rect 19276 31219 19316 31228
rect 19372 31564 19508 31604
rect 19564 31940 19604 31949
rect 19179 30848 19221 30857
rect 19179 30808 19180 30848
rect 19220 30808 19221 30848
rect 19179 30799 19221 30808
rect 19275 30764 19317 30773
rect 19275 30724 19276 30764
rect 19316 30724 19317 30764
rect 19275 30715 19317 30724
rect 18891 30428 18933 30437
rect 18891 30388 18892 30428
rect 18932 30388 18933 30428
rect 18891 30379 18933 30388
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 18940 29849 18980 29858
rect 18980 29809 19028 29840
rect 18940 29800 19028 29809
rect 18988 29336 19028 29800
rect 19084 29756 19124 29765
rect 19276 29756 19316 30715
rect 19372 30101 19412 31564
rect 19467 31436 19509 31445
rect 19467 31396 19468 31436
rect 19508 31396 19509 31436
rect 19467 31387 19509 31396
rect 19468 31302 19508 31387
rect 19564 31109 19604 31900
rect 19660 31445 19700 32656
rect 19756 32369 19796 32740
rect 19755 32360 19797 32369
rect 19755 32320 19756 32360
rect 19796 32320 19797 32360
rect 19755 32311 19797 32320
rect 19756 32108 19796 32117
rect 19756 31697 19796 32068
rect 19852 32033 19892 33580
rect 20139 33536 20181 33545
rect 20139 33496 20140 33536
rect 20180 33496 20181 33536
rect 20139 33487 20181 33496
rect 19947 33452 19989 33461
rect 19947 33412 19948 33452
rect 19988 33412 19989 33452
rect 19947 33403 19989 33412
rect 19948 33318 19988 33403
rect 20140 33402 20180 33487
rect 20139 33116 20181 33125
rect 20139 33076 20140 33116
rect 20180 33076 20181 33116
rect 20139 33067 20181 33076
rect 20140 33032 20180 33067
rect 20524 33041 20564 36520
rect 20620 33377 20660 37948
rect 20716 37157 20756 40384
rect 21195 40384 21196 40424
rect 21236 40384 21237 40424
rect 21195 40375 21237 40384
rect 20811 40088 20853 40097
rect 20811 40048 20812 40088
rect 20852 40048 20853 40088
rect 20811 40039 20853 40048
rect 20812 39593 20852 40039
rect 20811 39584 20853 39593
rect 20811 39544 20812 39584
rect 20852 39544 20853 39584
rect 20811 39535 20853 39544
rect 21003 37232 21045 37241
rect 21003 37192 21004 37232
rect 21044 37192 21045 37232
rect 21003 37183 21045 37192
rect 20715 37148 20757 37157
rect 20715 37108 20716 37148
rect 20756 37108 20757 37148
rect 20715 37099 20757 37108
rect 20715 36896 20757 36905
rect 20715 36856 20716 36896
rect 20756 36856 20757 36896
rect 20715 36847 20757 36856
rect 20716 33713 20756 36847
rect 20811 35972 20853 35981
rect 20811 35932 20812 35972
rect 20852 35932 20853 35972
rect 20811 35923 20853 35932
rect 20812 34049 20852 35923
rect 20811 34040 20853 34049
rect 20811 34000 20812 34040
rect 20852 34000 20853 34040
rect 20811 33991 20853 34000
rect 20715 33704 20757 33713
rect 20715 33664 20716 33704
rect 20756 33664 20757 33704
rect 20715 33655 20757 33664
rect 20619 33368 20661 33377
rect 20619 33328 20620 33368
rect 20660 33328 20661 33368
rect 20619 33319 20661 33328
rect 20140 32981 20180 32992
rect 20523 33032 20565 33041
rect 20523 32992 20524 33032
rect 20564 32992 20565 33032
rect 20523 32983 20565 32992
rect 19948 32696 19988 32705
rect 19948 32108 19988 32656
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 19948 32068 20084 32108
rect 19851 32024 19893 32033
rect 19851 31984 19852 32024
rect 19892 31984 19893 32024
rect 19851 31975 19893 31984
rect 19948 31940 19988 31949
rect 19755 31688 19797 31697
rect 19755 31648 19756 31688
rect 19796 31648 19797 31688
rect 19755 31639 19797 31648
rect 19948 31445 19988 31900
rect 19659 31436 19701 31445
rect 19659 31396 19660 31436
rect 19700 31396 19701 31436
rect 19659 31387 19701 31396
rect 19852 31436 19892 31445
rect 19755 31352 19797 31361
rect 19755 31312 19756 31352
rect 19796 31312 19797 31352
rect 19755 31303 19797 31312
rect 19659 31184 19701 31193
rect 19659 31144 19660 31184
rect 19700 31144 19701 31184
rect 19659 31135 19701 31144
rect 19563 31100 19605 31109
rect 19563 31060 19564 31100
rect 19604 31060 19605 31100
rect 19563 31051 19605 31060
rect 19660 31050 19700 31135
rect 19659 30848 19701 30857
rect 19659 30808 19660 30848
rect 19700 30808 19701 30848
rect 19659 30799 19701 30808
rect 19660 30714 19700 30799
rect 19468 30680 19508 30691
rect 19756 30689 19796 31303
rect 19852 30773 19892 31396
rect 19947 31436 19989 31445
rect 19947 31396 19948 31436
rect 19988 31396 19989 31436
rect 19947 31387 19989 31396
rect 20044 31361 20084 32068
rect 20043 31352 20085 31361
rect 20043 31312 20044 31352
rect 20084 31312 20085 31352
rect 20043 31303 20085 31312
rect 20044 31184 20084 31193
rect 19948 31144 20044 31184
rect 19851 30764 19893 30773
rect 19851 30724 19852 30764
rect 19892 30724 19893 30764
rect 19851 30715 19893 30724
rect 19468 30605 19508 30640
rect 19755 30680 19797 30689
rect 19755 30640 19756 30680
rect 19796 30640 19797 30680
rect 19755 30631 19797 30640
rect 19467 30596 19509 30605
rect 19467 30556 19468 30596
rect 19508 30556 19509 30596
rect 19467 30547 19509 30556
rect 19852 30596 19892 30605
rect 19371 30092 19413 30101
rect 19852 30092 19892 30556
rect 19371 30052 19372 30092
rect 19412 30052 19413 30092
rect 19371 30043 19413 30052
rect 19468 30052 19892 30092
rect 19371 29924 19413 29933
rect 19371 29884 19372 29924
rect 19412 29884 19413 29924
rect 19371 29875 19413 29884
rect 19372 29790 19412 29875
rect 19124 29716 19316 29756
rect 19084 29707 19124 29716
rect 19468 29672 19508 30052
rect 19755 29924 19797 29933
rect 19755 29884 19756 29924
rect 19796 29884 19797 29924
rect 19755 29875 19797 29884
rect 19756 29790 19796 29875
rect 19948 29849 19988 31144
rect 20044 31135 20084 31144
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 20044 30428 20084 30437
rect 19947 29840 19989 29849
rect 19947 29800 19948 29840
rect 19988 29800 19989 29840
rect 19947 29791 19989 29800
rect 20044 29681 20084 30388
rect 21004 30353 21044 37183
rect 21196 35645 21236 40375
rect 21195 35636 21237 35645
rect 21195 35596 21196 35636
rect 21236 35596 21237 35636
rect 21195 35587 21237 35596
rect 21195 33452 21237 33461
rect 21195 33412 21196 33452
rect 21236 33412 21237 33452
rect 21195 33403 21237 33412
rect 21196 32780 21236 33403
rect 21388 32780 21428 41383
rect 21100 32740 21236 32780
rect 21292 32740 21428 32780
rect 21003 30344 21045 30353
rect 21003 30304 21004 30344
rect 21044 30304 21045 30344
rect 21003 30295 21045 30304
rect 18988 29287 19028 29296
rect 19276 29632 19508 29672
rect 19564 29672 19604 29681
rect 19948 29672 19988 29681
rect 19604 29632 19892 29672
rect 18796 29168 18836 29196
rect 18700 29128 18796 29168
rect 18603 25388 18645 25397
rect 18603 25348 18604 25388
rect 18644 25348 18645 25388
rect 18603 25339 18645 25348
rect 18700 25136 18740 29128
rect 18796 29119 18836 29128
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18987 28496 19029 28505
rect 18987 28456 18988 28496
rect 19028 28456 19029 28496
rect 18987 28447 19029 28456
rect 18796 28333 18836 28342
rect 18796 27749 18836 28293
rect 18891 28244 18933 28253
rect 18891 28204 18892 28244
rect 18932 28204 18933 28244
rect 18891 28195 18933 28204
rect 18988 28244 19028 28447
rect 19276 28421 19316 29632
rect 19564 29623 19604 29632
rect 19372 29093 19412 29178
rect 19371 29084 19413 29093
rect 19756 29084 19796 29093
rect 19371 29044 19372 29084
rect 19412 29044 19413 29084
rect 19371 29035 19413 29044
rect 19468 29044 19756 29084
rect 19468 28505 19508 29044
rect 19756 29035 19796 29044
rect 19564 28916 19604 28925
rect 19604 28876 19700 28916
rect 19564 28867 19604 28876
rect 19467 28496 19509 28505
rect 19467 28456 19468 28496
rect 19508 28456 19509 28496
rect 19467 28447 19509 28456
rect 19275 28412 19317 28421
rect 19275 28372 19276 28412
rect 19316 28372 19317 28412
rect 19275 28363 19317 28372
rect 19372 28412 19412 28421
rect 18988 28195 19028 28204
rect 18795 27740 18837 27749
rect 18795 27700 18796 27740
rect 18836 27700 18837 27740
rect 18795 27691 18837 27700
rect 18892 27665 18932 28195
rect 19275 27740 19317 27749
rect 19275 27700 19276 27740
rect 19316 27700 19317 27740
rect 19275 27691 19317 27700
rect 18891 27656 18933 27665
rect 18891 27616 18892 27656
rect 18932 27616 18933 27656
rect 18891 27607 18933 27616
rect 19084 27656 19124 27665
rect 19084 27404 19124 27616
rect 19276 27606 19316 27691
rect 19084 27364 19316 27404
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 19276 27068 19316 27364
rect 19372 27077 19412 28372
rect 19564 28160 19604 28169
rect 19467 27572 19509 27581
rect 19467 27532 19468 27572
rect 19508 27532 19509 27572
rect 19467 27523 19509 27532
rect 19468 27438 19508 27523
rect 18892 27028 19316 27068
rect 19371 27068 19413 27077
rect 19371 27028 19372 27068
rect 19412 27028 19413 27068
rect 18892 26237 18932 27028
rect 19371 27019 19413 27028
rect 19564 26993 19604 28120
rect 19660 28085 19700 28876
rect 19756 28412 19796 28421
rect 19659 28076 19701 28085
rect 19659 28036 19660 28076
rect 19700 28036 19701 28076
rect 19659 28027 19701 28036
rect 19660 27413 19700 27498
rect 19659 27404 19701 27413
rect 19659 27364 19660 27404
rect 19700 27364 19701 27404
rect 19659 27355 19701 27364
rect 19756 27236 19796 28372
rect 19852 27749 19892 29632
rect 19948 29261 19988 29632
rect 20043 29672 20085 29681
rect 20043 29632 20044 29672
rect 20084 29632 20085 29672
rect 20043 29623 20085 29632
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 21100 29420 21140 32740
rect 21292 29420 21332 32740
rect 21387 30176 21429 30185
rect 21387 30136 21388 30176
rect 21428 30136 21429 30176
rect 21387 30127 21429 30136
rect 21004 29380 21140 29420
rect 21196 29380 21332 29420
rect 19947 29252 19989 29261
rect 19947 29212 19948 29252
rect 19988 29212 19989 29252
rect 19947 29203 19989 29212
rect 19947 29000 19989 29009
rect 19947 28960 19948 29000
rect 19988 28960 19989 29000
rect 19947 28951 19989 28960
rect 19948 28866 19988 28951
rect 19947 28160 19989 28169
rect 19947 28120 19948 28160
rect 19988 28120 19989 28160
rect 19947 28111 19989 28120
rect 20907 28160 20949 28169
rect 20907 28120 20908 28160
rect 20948 28120 20949 28160
rect 20907 28111 20949 28120
rect 19948 28026 19988 28111
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 19851 27740 19893 27749
rect 19851 27700 19852 27740
rect 19892 27700 19893 27740
rect 19851 27691 19893 27700
rect 19852 27572 19892 27581
rect 19892 27532 19988 27572
rect 19852 27523 19892 27532
rect 19851 27404 19893 27413
rect 19851 27364 19852 27404
rect 19892 27364 19893 27404
rect 19851 27355 19893 27364
rect 19660 27196 19796 27236
rect 19563 26984 19605 26993
rect 19563 26944 19564 26984
rect 19604 26944 19605 26984
rect 19563 26935 19605 26944
rect 19372 26900 19412 26909
rect 19036 26825 19076 26834
rect 19076 26785 19316 26816
rect 19036 26776 19316 26785
rect 19179 26648 19221 26657
rect 19179 26608 19180 26648
rect 19220 26608 19221 26648
rect 19179 26599 19221 26608
rect 19180 26514 19220 26599
rect 19276 26312 19316 26776
rect 19372 26489 19412 26860
rect 19660 26741 19700 27196
rect 19756 26900 19796 26909
rect 19659 26732 19701 26741
rect 19659 26692 19660 26732
rect 19700 26692 19701 26732
rect 19659 26683 19701 26692
rect 19563 26648 19605 26657
rect 19563 26608 19564 26648
rect 19604 26608 19605 26648
rect 19563 26599 19605 26608
rect 19564 26514 19604 26599
rect 19371 26480 19413 26489
rect 19371 26440 19372 26480
rect 19412 26440 19413 26480
rect 19371 26431 19413 26440
rect 19564 26312 19604 26321
rect 19276 26272 19564 26312
rect 19564 26263 19604 26272
rect 18891 26228 18933 26237
rect 19756 26228 19796 26860
rect 18891 26188 18892 26228
rect 18932 26188 18933 26228
rect 18891 26179 18933 26188
rect 19372 26153 19412 26228
rect 19660 26188 19796 26228
rect 19275 26144 19317 26153
rect 19275 26104 19276 26144
rect 19316 26104 19317 26144
rect 19275 26095 19317 26104
rect 19372 26144 19424 26153
rect 19660 26144 19700 26188
rect 19423 26104 19424 26144
rect 19372 26095 19424 26104
rect 19468 26104 19700 26144
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18891 25472 18933 25481
rect 18891 25432 18892 25472
rect 18932 25432 18933 25472
rect 18891 25423 18933 25432
rect 18508 25096 18740 25136
rect 18796 25309 18836 25318
rect 18411 24884 18453 24893
rect 18411 24844 18412 24884
rect 18452 24844 18453 24884
rect 18411 24835 18453 24844
rect 18315 24632 18357 24641
rect 18315 24592 18316 24632
rect 18356 24592 18357 24632
rect 18315 24583 18357 24592
rect 18220 23381 18260 23752
rect 18316 23792 18356 24583
rect 18219 23372 18261 23381
rect 18219 23332 18220 23372
rect 18260 23332 18261 23372
rect 18219 23323 18261 23332
rect 18123 22616 18165 22625
rect 18123 22576 18124 22616
rect 18164 22576 18165 22616
rect 18123 22567 18165 22576
rect 18124 21701 18164 22567
rect 18123 21692 18165 21701
rect 18123 21652 18124 21692
rect 18164 21652 18165 21692
rect 18123 21643 18165 21652
rect 18027 21608 18069 21617
rect 18027 21568 18028 21608
rect 18068 21568 18069 21608
rect 18027 21559 18069 21568
rect 17931 21188 17973 21197
rect 17931 21148 17932 21188
rect 17972 21148 17973 21188
rect 17931 21139 17973 21148
rect 17835 21104 17877 21113
rect 17835 21064 17836 21104
rect 17876 21064 17877 21104
rect 17835 21055 17877 21064
rect 17836 20861 17876 21055
rect 17835 20852 17877 20861
rect 17835 20812 17836 20852
rect 17876 20812 17877 20852
rect 17835 20803 17877 20812
rect 17836 20096 17876 20803
rect 18028 20782 18068 21559
rect 18316 21365 18356 23752
rect 18412 23129 18452 24835
rect 18411 23120 18453 23129
rect 18411 23080 18412 23120
rect 18452 23080 18453 23120
rect 18508 23120 18548 25096
rect 18796 24809 18836 25269
rect 18795 24800 18837 24809
rect 18795 24760 18796 24800
rect 18836 24760 18837 24800
rect 18795 24751 18837 24760
rect 18892 24632 18932 25423
rect 19276 25397 19316 26095
rect 19371 25976 19413 25985
rect 19371 25936 19372 25976
rect 19412 25936 19413 25976
rect 19371 25927 19413 25936
rect 19275 25388 19317 25397
rect 19275 25348 19276 25388
rect 19316 25348 19317 25388
rect 19275 25339 19317 25348
rect 19372 25388 19412 25927
rect 19372 25339 19412 25348
rect 18988 25220 19028 25229
rect 19468 25220 19508 26104
rect 19755 26060 19797 26069
rect 19755 26020 19756 26060
rect 19796 26020 19797 26060
rect 19852 26060 19892 27355
rect 19948 27077 19988 27532
rect 20044 27404 20084 27413
rect 19947 27068 19989 27077
rect 19947 27028 19948 27068
rect 19988 27028 19989 27068
rect 19947 27019 19989 27028
rect 19947 26816 19989 26825
rect 19947 26776 19948 26816
rect 19988 26776 19989 26816
rect 19947 26767 19989 26776
rect 19948 26648 19988 26767
rect 20044 26657 20084 27364
rect 19948 26599 19988 26608
rect 20043 26648 20085 26657
rect 20043 26608 20044 26648
rect 20084 26608 20085 26648
rect 20043 26599 20085 26608
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 20908 26321 20948 28111
rect 20907 26312 20949 26321
rect 20907 26272 20908 26312
rect 20948 26272 20949 26312
rect 20907 26263 20949 26272
rect 19852 26020 20084 26060
rect 19755 26011 19797 26020
rect 19756 25926 19796 26011
rect 19948 25892 19988 25901
rect 19852 25852 19948 25892
rect 19755 25388 19797 25397
rect 19755 25348 19756 25388
rect 19796 25348 19797 25388
rect 19755 25339 19797 25348
rect 19756 25254 19796 25339
rect 19028 25180 19508 25220
rect 18988 25171 19028 25180
rect 19564 25136 19604 25145
rect 19275 24800 19317 24809
rect 19275 24760 19276 24800
rect 19316 24760 19317 24800
rect 19275 24751 19317 24760
rect 19276 24666 19316 24751
rect 19084 24632 19124 24641
rect 18892 24592 19084 24632
rect 19084 24583 19124 24592
rect 19468 24548 19508 24559
rect 19468 24473 19508 24508
rect 19467 24464 19509 24473
rect 19467 24424 19468 24464
rect 19508 24424 19509 24464
rect 19467 24415 19509 24424
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 19564 24137 19604 25096
rect 19852 24809 19892 25852
rect 19948 25843 19988 25852
rect 20044 25145 20084 26020
rect 21004 25985 21044 29380
rect 21003 25976 21045 25985
rect 21003 25936 21004 25976
rect 21044 25936 21045 25976
rect 21003 25927 21045 25936
rect 21196 25229 21236 29380
rect 21291 29168 21333 29177
rect 21291 29128 21292 29168
rect 21332 29128 21333 29168
rect 21291 29119 21333 29128
rect 21195 25220 21237 25229
rect 21195 25180 21196 25220
rect 21236 25180 21237 25220
rect 21195 25171 21237 25180
rect 19948 25136 19988 25145
rect 19851 24800 19893 24809
rect 19851 24760 19852 24800
rect 19892 24760 19893 24800
rect 19851 24751 19893 24760
rect 19755 24632 19797 24641
rect 19755 24592 19756 24632
rect 19796 24592 19797 24632
rect 19755 24583 19797 24592
rect 19852 24632 19892 24641
rect 19660 24380 19700 24389
rect 19563 24128 19605 24137
rect 19563 24088 19564 24128
rect 19604 24088 19605 24128
rect 19563 24079 19605 24088
rect 19372 23960 19412 23969
rect 19412 23920 19604 23960
rect 19372 23911 19412 23920
rect 18700 23792 18740 23803
rect 18700 23717 18740 23752
rect 18796 23792 18836 23801
rect 18699 23708 18741 23717
rect 18699 23668 18700 23708
rect 18740 23668 18741 23708
rect 18699 23659 18741 23668
rect 18604 23120 18644 23129
rect 18796 23120 18836 23752
rect 19084 23792 19124 23801
rect 18508 23080 18604 23120
rect 18411 23071 18453 23080
rect 18604 22289 18644 23080
rect 18700 23080 18836 23120
rect 18987 23120 19029 23129
rect 18987 23080 18988 23120
rect 19028 23080 19029 23120
rect 18411 22280 18453 22289
rect 18411 22240 18412 22280
rect 18452 22240 18453 22280
rect 18411 22231 18453 22240
rect 18603 22280 18645 22289
rect 18603 22240 18604 22280
rect 18644 22240 18645 22280
rect 18603 22231 18645 22240
rect 18412 21608 18452 22231
rect 18700 22205 18740 23080
rect 18987 23071 19029 23080
rect 18988 22986 19028 23071
rect 18796 22877 18836 22962
rect 19084 22961 19124 23752
rect 19179 23792 19221 23801
rect 19179 23752 19180 23792
rect 19220 23752 19221 23792
rect 19179 23743 19221 23752
rect 19372 23792 19412 23801
rect 19180 23288 19220 23743
rect 19372 23288 19412 23752
rect 19564 23792 19604 23920
rect 19564 23743 19604 23752
rect 19660 23297 19700 24340
rect 19756 24044 19796 24583
rect 19852 24557 19892 24592
rect 19850 24548 19892 24557
rect 19850 24508 19851 24548
rect 19891 24508 19892 24548
rect 19850 24499 19892 24508
rect 19852 24380 19892 24389
rect 19852 24044 19892 24340
rect 19948 24305 19988 25096
rect 20043 25136 20085 25145
rect 20043 25096 20044 25136
rect 20084 25096 20085 25136
rect 20043 25087 20085 25096
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20043 24632 20085 24641
rect 20043 24592 20044 24632
rect 20084 24592 20085 24632
rect 20043 24583 20085 24592
rect 20044 24498 20084 24583
rect 19947 24296 19989 24305
rect 19947 24256 19948 24296
rect 19988 24256 19989 24296
rect 19947 24247 19989 24256
rect 19852 24004 20084 24044
rect 19756 23995 19796 24004
rect 19947 23876 19989 23885
rect 19947 23836 19948 23876
rect 19988 23836 19989 23876
rect 19947 23827 19989 23836
rect 19756 23792 19796 23801
rect 19796 23752 19892 23792
rect 19756 23743 19796 23752
rect 19468 23288 19508 23297
rect 19180 23248 19316 23288
rect 19372 23248 19468 23288
rect 19179 23120 19221 23129
rect 19179 23080 19180 23120
rect 19220 23080 19221 23120
rect 19179 23071 19221 23080
rect 19276 23120 19316 23248
rect 19468 23239 19508 23248
rect 19659 23288 19701 23297
rect 19659 23248 19660 23288
rect 19700 23248 19701 23288
rect 19659 23239 19701 23248
rect 19564 23120 19604 23129
rect 19180 22986 19220 23071
rect 19276 23045 19316 23080
rect 19468 23080 19564 23120
rect 19275 23036 19317 23045
rect 19275 22996 19276 23036
rect 19316 22996 19317 23036
rect 19275 22987 19317 22996
rect 19083 22952 19125 22961
rect 19083 22912 19084 22952
rect 19124 22912 19125 22952
rect 19083 22903 19125 22912
rect 19276 22877 19316 22987
rect 19371 22952 19413 22961
rect 19371 22912 19372 22952
rect 19412 22912 19413 22952
rect 19371 22903 19413 22912
rect 18795 22868 18837 22877
rect 18795 22828 18796 22868
rect 18836 22828 18837 22868
rect 18795 22819 18837 22828
rect 19275 22868 19317 22877
rect 19275 22828 19276 22868
rect 19316 22828 19317 22868
rect 19275 22819 19317 22828
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 19275 22532 19317 22541
rect 19275 22492 19276 22532
rect 19316 22492 19317 22532
rect 19275 22483 19317 22492
rect 19276 22398 19316 22483
rect 19083 22280 19125 22289
rect 19083 22240 19084 22280
rect 19124 22240 19125 22280
rect 19083 22231 19125 22240
rect 18699 22196 18741 22205
rect 18699 22156 18700 22196
rect 18740 22156 18741 22196
rect 18699 22147 18741 22156
rect 19084 22146 19124 22231
rect 19372 21785 19412 22903
rect 19468 22280 19508 23080
rect 19564 23071 19604 23080
rect 19660 23120 19700 23129
rect 19563 22868 19605 22877
rect 19563 22828 19564 22868
rect 19604 22828 19605 22868
rect 19563 22819 19605 22828
rect 19468 22205 19508 22240
rect 19564 22280 19604 22819
rect 19660 22709 19700 23080
rect 19756 23120 19796 23131
rect 19756 23045 19796 23080
rect 19755 23036 19797 23045
rect 19755 22996 19756 23036
rect 19796 22996 19797 23036
rect 19755 22987 19797 22996
rect 19659 22700 19701 22709
rect 19659 22660 19660 22700
rect 19700 22660 19701 22700
rect 19659 22651 19701 22660
rect 19659 22532 19701 22541
rect 19659 22492 19660 22532
rect 19700 22492 19701 22532
rect 19659 22483 19701 22492
rect 19564 22231 19604 22240
rect 19660 22280 19700 22483
rect 19660 22231 19700 22240
rect 19756 22280 19796 22289
rect 19852 22280 19892 23752
rect 19948 23742 19988 23827
rect 20044 23624 20084 24004
rect 19948 23584 20084 23624
rect 20140 23624 20180 23633
rect 20180 23584 20564 23624
rect 19948 23288 19988 23584
rect 20140 23575 20180 23584
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 19948 23248 20084 23288
rect 19948 23109 19988 23118
rect 19948 23045 19988 23069
rect 19947 23036 19989 23045
rect 19947 22996 19948 23036
rect 19988 22996 19989 23036
rect 19947 22987 19989 22996
rect 19948 22974 19988 22987
rect 19947 22868 19989 22877
rect 19947 22828 19948 22868
rect 19988 22828 19989 22868
rect 19947 22819 19989 22828
rect 19948 22734 19988 22819
rect 19948 22364 19988 22373
rect 20044 22364 20084 23248
rect 20140 23120 20180 23129
rect 20140 22961 20180 23080
rect 20236 23120 20276 23129
rect 20139 22952 20181 22961
rect 20139 22912 20140 22952
rect 20180 22912 20181 22952
rect 20139 22903 20181 22912
rect 20236 22793 20276 23080
rect 20235 22784 20277 22793
rect 20235 22744 20236 22784
rect 20276 22744 20277 22784
rect 20235 22735 20277 22744
rect 20524 22625 20564 23584
rect 20523 22616 20565 22625
rect 20523 22576 20524 22616
rect 20564 22576 20565 22616
rect 20523 22567 20565 22576
rect 19988 22324 20084 22364
rect 19948 22315 19988 22324
rect 19796 22240 19892 22280
rect 19756 22231 19796 22240
rect 19467 22196 19509 22205
rect 19467 22156 19468 22196
rect 19508 22156 19509 22196
rect 19467 22147 19509 22156
rect 20140 22121 20180 22206
rect 20139 22112 20181 22121
rect 20139 22072 20140 22112
rect 20180 22072 20181 22112
rect 20139 22063 20181 22072
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 19371 21776 19413 21785
rect 19371 21736 19372 21776
rect 19412 21736 19413 21776
rect 19371 21727 19413 21736
rect 20043 21776 20085 21785
rect 20043 21736 20044 21776
rect 20084 21736 20085 21776
rect 20043 21727 20085 21736
rect 18604 21692 18644 21703
rect 18604 21617 18644 21652
rect 18795 21692 18837 21701
rect 18795 21652 18796 21692
rect 18836 21652 18837 21692
rect 18795 21643 18837 21652
rect 19084 21652 19316 21692
rect 18412 21559 18452 21568
rect 18603 21608 18645 21617
rect 18796 21608 18836 21643
rect 18603 21568 18604 21608
rect 18644 21568 18740 21608
rect 18603 21559 18645 21568
rect 18315 21356 18357 21365
rect 18315 21316 18316 21356
rect 18356 21316 18357 21356
rect 18315 21307 18357 21316
rect 18028 20733 18068 20742
rect 18507 20768 18549 20777
rect 18507 20728 18508 20768
rect 18548 20728 18549 20768
rect 18507 20719 18549 20728
rect 18604 20768 18644 20777
rect 18219 20684 18261 20693
rect 18219 20644 18220 20684
rect 18260 20644 18261 20684
rect 18219 20635 18261 20644
rect 18220 20550 18260 20635
rect 18508 20634 18548 20719
rect 18412 20600 18452 20609
rect 18028 20273 18068 20358
rect 18027 20264 18069 20273
rect 18027 20224 18028 20264
rect 18068 20224 18069 20264
rect 18027 20215 18069 20224
rect 18412 20180 18452 20560
rect 18507 20348 18549 20357
rect 18507 20308 18508 20348
rect 18548 20308 18549 20348
rect 18507 20299 18549 20308
rect 18220 20140 18452 20180
rect 17836 20047 17876 20056
rect 17931 20096 17973 20105
rect 17931 20056 17932 20096
rect 17972 20056 17973 20096
rect 17931 20047 17973 20056
rect 18123 20096 18165 20105
rect 18123 20056 18124 20096
rect 18164 20056 18165 20096
rect 18123 20047 18165 20056
rect 17932 19962 17972 20047
rect 18027 20012 18069 20021
rect 18027 19972 18028 20012
rect 18068 19972 18069 20012
rect 18027 19963 18069 19972
rect 17740 19888 17876 19928
rect 17739 19760 17781 19769
rect 17739 19720 17740 19760
rect 17780 19720 17781 19760
rect 17739 19711 17781 19720
rect 17740 19256 17780 19711
rect 17740 19207 17780 19216
rect 17836 18677 17876 19888
rect 17835 18668 17877 18677
rect 17835 18628 17836 18668
rect 17876 18628 17877 18668
rect 17835 18619 17877 18628
rect 17740 18584 17780 18593
rect 17740 18173 17780 18544
rect 17931 18332 17973 18341
rect 17931 18292 17932 18332
rect 17972 18292 17973 18332
rect 17931 18283 17973 18292
rect 17739 18164 17781 18173
rect 17739 18124 17740 18164
rect 17780 18124 17781 18164
rect 17739 18115 17781 18124
rect 17740 17744 17780 17753
rect 17740 17165 17780 17704
rect 17739 17156 17781 17165
rect 17739 17116 17740 17156
rect 17780 17116 17781 17156
rect 17739 17107 17781 17116
rect 17644 15772 17780 15812
rect 17451 15763 17493 15772
rect 17452 15644 17492 15653
rect 17355 14888 17397 14897
rect 17260 14848 17302 14888
rect 17262 14804 17302 14848
rect 17355 14848 17356 14888
rect 17396 14848 17397 14888
rect 17355 14839 17397 14848
rect 17260 14764 17302 14804
rect 17260 14762 17300 14764
rect 17260 14713 17300 14722
rect 17356 14720 17396 14729
rect 17452 14720 17492 15604
rect 17644 15560 17684 15569
rect 17644 15401 17684 15520
rect 17643 15392 17685 15401
rect 17643 15352 17644 15392
rect 17684 15352 17685 15392
rect 17643 15343 17685 15352
rect 17547 14972 17589 14981
rect 17547 14932 17548 14972
rect 17588 14932 17589 14972
rect 17547 14923 17589 14932
rect 17396 14680 17492 14720
rect 17356 14671 17396 14680
rect 17355 14552 17397 14561
rect 16876 14512 17108 14552
rect 16779 14384 16821 14393
rect 16779 14344 16780 14384
rect 16820 14344 16821 14384
rect 16779 14335 16821 14344
rect 16628 14176 16724 14216
rect 16588 14167 16628 14176
rect 16492 13999 16532 14008
rect 16684 14048 16724 14057
rect 16780 14048 16820 14335
rect 17068 14216 17108 14512
rect 17355 14512 17356 14552
rect 17396 14512 17397 14552
rect 17355 14503 17397 14512
rect 17068 14167 17108 14176
rect 16875 14132 16917 14141
rect 16875 14092 16876 14132
rect 16916 14092 16917 14132
rect 16875 14083 16917 14092
rect 17163 14132 17205 14141
rect 17163 14092 17164 14132
rect 17204 14092 17205 14132
rect 17163 14083 17205 14092
rect 16724 14008 16820 14048
rect 16684 13999 16724 14008
rect 16876 13964 16916 14083
rect 16876 13915 16916 13924
rect 16491 13544 16533 13553
rect 16491 13504 16492 13544
rect 16532 13504 16533 13544
rect 16491 13495 16533 13504
rect 16148 12328 16244 12368
rect 16300 12536 16340 12545
rect 15435 12284 15477 12293
rect 15435 12244 15436 12284
rect 15476 12244 15477 12284
rect 15435 12235 15477 12244
rect 15436 10529 15476 12235
rect 15628 11360 15668 12328
rect 16108 12319 16148 12328
rect 16300 11948 16340 12496
rect 15820 11908 16340 11948
rect 16396 12452 16436 12461
rect 15628 11320 15764 11360
rect 15627 11024 15669 11033
rect 15627 10984 15628 11024
rect 15668 10984 15669 11024
rect 15627 10975 15669 10984
rect 15243 10520 15285 10529
rect 15243 10480 15244 10520
rect 15284 10480 15285 10520
rect 15243 10471 15285 10480
rect 15435 10520 15477 10529
rect 15435 10480 15436 10520
rect 15476 10480 15477 10520
rect 15435 10471 15477 10480
rect 15148 10312 15476 10352
rect 15051 10268 15093 10277
rect 15051 10228 15052 10268
rect 15092 10228 15093 10268
rect 15051 10219 15093 10228
rect 15244 10184 15284 10193
rect 14668 8800 14900 8840
rect 14956 10016 14996 10025
rect 14668 8714 14708 8800
rect 14668 8665 14708 8674
rect 14572 8548 14804 8588
rect 14571 8336 14613 8345
rect 14571 8296 14572 8336
rect 14612 8296 14613 8336
rect 14571 8287 14613 8296
rect 14475 8168 14517 8177
rect 14475 8128 14476 8168
rect 14516 8128 14517 8168
rect 14475 8119 14517 8128
rect 14572 8000 14612 8287
rect 14764 8009 14804 8548
rect 14860 8504 14900 8513
rect 14860 8345 14900 8464
rect 14859 8336 14901 8345
rect 14859 8296 14860 8336
rect 14900 8296 14901 8336
rect 14859 8287 14901 8296
rect 14859 8168 14901 8177
rect 14859 8128 14860 8168
rect 14900 8128 14901 8168
rect 14859 8119 14901 8128
rect 14572 7951 14612 7960
rect 14763 8000 14805 8009
rect 14763 7960 14764 8000
rect 14804 7960 14805 8000
rect 14763 7951 14805 7960
rect 14860 8000 14900 8119
rect 14956 8084 14996 9976
rect 15244 9932 15284 10144
rect 15052 9892 15284 9932
rect 15340 10016 15380 10025
rect 15052 9260 15092 9892
rect 15147 9764 15189 9773
rect 15147 9724 15148 9764
rect 15188 9724 15189 9764
rect 15147 9715 15189 9724
rect 15148 9521 15188 9715
rect 15243 9596 15285 9605
rect 15243 9556 15244 9596
rect 15284 9556 15285 9596
rect 15243 9547 15285 9556
rect 15147 9512 15189 9521
rect 15147 9472 15148 9512
rect 15188 9472 15189 9512
rect 15147 9463 15189 9472
rect 15244 9512 15284 9547
rect 15148 9378 15188 9463
rect 15244 9461 15284 9472
rect 15243 9344 15285 9353
rect 15243 9304 15244 9344
rect 15284 9304 15285 9344
rect 15243 9295 15285 9304
rect 15052 9220 15188 9260
rect 15148 8765 15188 9220
rect 15244 8924 15284 9295
rect 15340 9017 15380 9976
rect 15339 9008 15381 9017
rect 15339 8968 15340 9008
rect 15380 8968 15381 9008
rect 15339 8959 15381 8968
rect 15244 8884 15292 8924
rect 15252 8840 15292 8884
rect 15244 8800 15292 8840
rect 15147 8756 15189 8765
rect 15147 8716 15148 8756
rect 15188 8716 15189 8756
rect 15147 8707 15189 8716
rect 14956 8035 14996 8044
rect 15052 8672 15092 8681
rect 14860 7951 14900 7960
rect 14667 7580 14709 7589
rect 14667 7540 14668 7580
rect 14708 7540 14709 7580
rect 14667 7531 14709 7540
rect 14379 7496 14421 7505
rect 14379 7456 14380 7496
rect 14420 7456 14421 7496
rect 14379 7447 14421 7456
rect 14668 7412 14708 7531
rect 14668 7363 14708 7372
rect 14476 7160 14516 7169
rect 14284 7111 14324 7120
rect 14380 7120 14476 7160
rect 14187 7076 14229 7085
rect 14187 7036 14188 7076
rect 14228 7036 14229 7076
rect 14187 7027 14229 7036
rect 14380 6824 14420 7120
rect 14476 7111 14516 7120
rect 14668 7160 14708 7169
rect 14188 6784 14420 6824
rect 14091 5816 14133 5825
rect 14091 5776 14092 5816
rect 14132 5776 14133 5816
rect 14091 5767 14133 5776
rect 14092 5648 14132 5767
rect 14188 5741 14228 6784
rect 14380 6656 14420 6665
rect 14668 6656 14708 7120
rect 14420 6616 14708 6656
rect 14380 6607 14420 6616
rect 14283 6572 14325 6581
rect 14283 6532 14284 6572
rect 14324 6532 14325 6572
rect 14283 6523 14325 6532
rect 14284 6488 14324 6523
rect 14284 6437 14324 6448
rect 14475 6488 14517 6497
rect 14475 6448 14476 6488
rect 14516 6448 14517 6488
rect 14475 6439 14517 6448
rect 14667 6488 14709 6497
rect 14667 6448 14668 6488
rect 14708 6448 14709 6488
rect 14667 6439 14709 6448
rect 14476 6354 14516 6439
rect 14668 6354 14708 6439
rect 14379 6320 14421 6329
rect 14379 6280 14380 6320
rect 14420 6280 14421 6320
rect 14379 6271 14421 6280
rect 14283 6236 14325 6245
rect 14283 6196 14284 6236
rect 14324 6196 14325 6236
rect 14283 6187 14325 6196
rect 14187 5732 14229 5741
rect 14187 5692 14188 5732
rect 14228 5692 14229 5732
rect 14187 5683 14229 5692
rect 14092 5599 14132 5608
rect 13803 5440 13804 5480
rect 13844 5440 14036 5480
rect 13803 5431 13845 5440
rect 13323 4976 13365 4985
rect 13323 4936 13324 4976
rect 13364 4936 13365 4976
rect 13323 4927 13365 4936
rect 13420 4976 13460 5431
rect 13515 5396 13557 5405
rect 13707 5396 13749 5405
rect 13515 5356 13516 5396
rect 13556 5356 13557 5396
rect 13515 5347 13557 5356
rect 13612 5356 13708 5396
rect 13748 5356 13749 5396
rect 13420 4927 13460 4936
rect 13324 4842 13364 4927
rect 13516 4817 13556 5347
rect 13612 4901 13652 5356
rect 13707 5347 13749 5356
rect 13804 5346 13844 5431
rect 13899 5228 13941 5237
rect 13899 5188 13900 5228
rect 13940 5188 13941 5228
rect 13899 5179 13941 5188
rect 13708 4976 13748 4985
rect 13611 4892 13653 4901
rect 13611 4852 13612 4892
rect 13652 4852 13653 4892
rect 13611 4843 13653 4852
rect 13515 4808 13557 4817
rect 13515 4768 13516 4808
rect 13556 4768 13557 4808
rect 13515 4759 13557 4768
rect 13708 4556 13748 4936
rect 13804 4976 13844 4985
rect 13804 4733 13844 4936
rect 13900 4976 13940 5179
rect 14187 5060 14229 5069
rect 14187 5020 14188 5060
rect 14228 5020 14229 5060
rect 14187 5011 14229 5020
rect 13900 4927 13940 4936
rect 13995 4976 14037 4985
rect 13995 4936 13996 4976
rect 14036 4936 14037 4976
rect 13995 4927 14037 4936
rect 14188 4976 14228 5011
rect 13996 4842 14036 4927
rect 14188 4925 14228 4936
rect 13803 4724 13845 4733
rect 13803 4684 13804 4724
rect 13844 4684 13845 4724
rect 13803 4675 13845 4684
rect 13708 4516 13844 4556
rect 13516 4388 13556 4397
rect 13228 4348 13516 4388
rect 13131 4339 13173 4348
rect 13516 4339 13556 4348
rect 12843 4304 12885 4313
rect 12843 4264 12844 4304
rect 12884 4264 12885 4304
rect 12843 4255 12885 4264
rect 13132 3809 13172 4339
rect 13324 4136 13364 4145
rect 13228 4096 13324 4136
rect 13131 3800 13173 3809
rect 13131 3760 13132 3800
rect 13172 3760 13173 3800
rect 13131 3751 13173 3760
rect 13228 3389 13268 4096
rect 13324 4087 13364 4096
rect 13708 4136 13748 4145
rect 13323 3800 13365 3809
rect 13323 3760 13324 3800
rect 13364 3760 13365 3800
rect 13323 3751 13365 3760
rect 13227 3380 13269 3389
rect 13227 3340 13228 3380
rect 13268 3340 13269 3380
rect 13227 3331 13269 3340
rect 12747 2960 12789 2969
rect 12747 2920 12748 2960
rect 12788 2920 12789 2960
rect 12747 2911 12789 2920
rect 12651 2624 12693 2633
rect 12651 2584 12652 2624
rect 12692 2584 12693 2624
rect 12651 2575 12693 2584
rect 12652 2490 12692 2575
rect 12555 2372 12597 2381
rect 12555 2332 12556 2372
rect 12596 2332 12597 2372
rect 12555 2323 12597 2332
rect 12459 2204 12501 2213
rect 12459 2164 12460 2204
rect 12500 2164 12501 2204
rect 12459 2155 12501 2164
rect 13035 2204 13077 2213
rect 13035 2164 13036 2204
rect 13076 2164 13077 2204
rect 13035 2155 13077 2164
rect 12171 2120 12213 2129
rect 12171 2080 12172 2120
rect 12212 2080 12213 2120
rect 12171 2071 12213 2080
rect 12555 2120 12597 2129
rect 12555 2080 12556 2120
rect 12596 2080 12597 2120
rect 12555 2071 12597 2080
rect 12172 1952 12212 2071
rect 12172 1903 12212 1912
rect 12171 1784 12213 1793
rect 12171 1744 12172 1784
rect 12212 1744 12213 1784
rect 12171 1735 12213 1744
rect 11980 1240 12116 1280
rect 11980 80 12020 1240
rect 12172 80 12212 1735
rect 12363 1532 12405 1541
rect 12363 1492 12364 1532
rect 12404 1492 12405 1532
rect 12363 1483 12405 1492
rect 12364 80 12404 1483
rect 12556 1112 12596 2071
rect 12747 1784 12789 1793
rect 12747 1744 12748 1784
rect 12788 1744 12789 1784
rect 12747 1735 12789 1744
rect 12748 1364 12788 1735
rect 12748 1315 12788 1324
rect 12940 1289 12980 1374
rect 12939 1280 12981 1289
rect 12939 1240 12940 1280
rect 12980 1240 12981 1280
rect 12939 1231 12981 1240
rect 12460 1072 12556 1112
rect 12460 197 12500 1072
rect 12556 1063 12596 1072
rect 12940 1112 12980 1121
rect 13036 1112 13076 2155
rect 13131 2120 13173 2129
rect 13131 2080 13132 2120
rect 13172 2080 13173 2120
rect 13131 2071 13173 2080
rect 13132 1625 13172 2071
rect 13324 1625 13364 3751
rect 13611 3716 13653 3725
rect 13611 3676 13612 3716
rect 13652 3676 13653 3716
rect 13611 3667 13653 3676
rect 13515 3464 13557 3473
rect 13515 3424 13516 3464
rect 13556 3424 13557 3464
rect 13515 3415 13557 3424
rect 13516 3330 13556 3415
rect 13612 3212 13652 3667
rect 13708 3380 13748 4096
rect 13804 4136 13844 4516
rect 14091 4472 14133 4481
rect 14091 4432 14092 4472
rect 14132 4432 14133 4472
rect 14091 4423 14133 4432
rect 13995 4220 14037 4229
rect 13804 4087 13844 4096
rect 13900 4180 13996 4220
rect 14036 4180 14037 4220
rect 13900 4136 13940 4180
rect 13995 4171 14037 4180
rect 13900 4087 13940 4096
rect 13996 3968 14036 3977
rect 13899 3716 13941 3725
rect 13899 3676 13900 3716
rect 13940 3676 13941 3716
rect 13899 3667 13941 3676
rect 13900 3464 13940 3667
rect 13996 3473 14036 3928
rect 13900 3415 13940 3424
rect 13995 3464 14037 3473
rect 13995 3424 13996 3464
rect 14036 3424 14037 3464
rect 13995 3415 14037 3424
rect 13708 3340 13844 3380
rect 13708 3212 13748 3221
rect 13612 3172 13708 3212
rect 13708 3163 13748 3172
rect 13515 3044 13557 3053
rect 13515 3004 13516 3044
rect 13556 3004 13557 3044
rect 13515 2995 13557 3004
rect 13419 2456 13461 2465
rect 13419 2416 13420 2456
rect 13460 2416 13461 2456
rect 13419 2407 13461 2416
rect 13420 1952 13460 2407
rect 13420 1903 13460 1912
rect 13131 1616 13173 1625
rect 13131 1576 13132 1616
rect 13172 1576 13173 1616
rect 13131 1567 13173 1576
rect 13323 1616 13365 1625
rect 13323 1576 13324 1616
rect 13364 1576 13365 1616
rect 13323 1567 13365 1576
rect 13323 1280 13365 1289
rect 13323 1240 13324 1280
rect 13364 1240 13365 1280
rect 13323 1231 13365 1240
rect 12980 1072 13076 1112
rect 13131 1112 13173 1121
rect 13131 1072 13132 1112
rect 13172 1072 13173 1112
rect 12940 1063 12980 1072
rect 13131 1063 13173 1072
rect 13228 1112 13268 1123
rect 13132 978 13172 1063
rect 13228 1037 13268 1072
rect 13227 1028 13269 1037
rect 13227 988 13228 1028
rect 13268 988 13269 1028
rect 13227 979 13269 988
rect 12555 944 12597 953
rect 12555 904 12556 944
rect 12596 904 12597 944
rect 12555 895 12597 904
rect 12939 944 12981 953
rect 12939 904 12940 944
rect 12980 904 12981 944
rect 12939 895 12981 904
rect 12459 188 12501 197
rect 12459 148 12460 188
rect 12500 148 12501 188
rect 12459 139 12501 148
rect 12556 80 12596 895
rect 12747 524 12789 533
rect 12747 484 12748 524
rect 12788 484 12789 524
rect 12747 475 12789 484
rect 12748 80 12788 475
rect 12940 80 12980 895
rect 13131 860 13173 869
rect 13131 820 13132 860
rect 13172 820 13173 860
rect 13131 811 13173 820
rect 13132 80 13172 811
rect 13324 80 13364 1231
rect 13419 1112 13461 1121
rect 13419 1072 13420 1112
rect 13460 1072 13461 1112
rect 13419 1063 13461 1072
rect 13516 1112 13556 2995
rect 13707 2708 13749 2717
rect 13707 2668 13708 2708
rect 13748 2668 13749 2708
rect 13707 2659 13749 2668
rect 13611 2120 13653 2129
rect 13611 2080 13612 2120
rect 13652 2080 13653 2120
rect 13611 2071 13653 2080
rect 13612 1952 13652 2071
rect 13612 1903 13652 1912
rect 13708 1784 13748 2659
rect 13804 1793 13844 3340
rect 14092 2876 14132 4423
rect 14187 4220 14229 4229
rect 14187 4180 14188 4220
rect 14228 4180 14229 4220
rect 14187 4171 14229 4180
rect 14092 2827 14132 2836
rect 13899 2792 13941 2801
rect 13899 2752 13900 2792
rect 13940 2752 13941 2792
rect 13899 2743 13941 2752
rect 13900 2624 13940 2743
rect 13900 2575 13940 2584
rect 13516 1063 13556 1072
rect 13612 1744 13748 1784
rect 13803 1784 13845 1793
rect 13803 1744 13804 1784
rect 13844 1744 13845 1784
rect 13612 1112 13652 1744
rect 13803 1735 13845 1744
rect 14188 1709 14228 4171
rect 14284 4136 14324 6187
rect 14284 4087 14324 4096
rect 14283 2960 14325 2969
rect 14283 2920 14284 2960
rect 14324 2920 14325 2960
rect 14283 2911 14325 2920
rect 14284 2624 14324 2911
rect 14284 2575 14324 2584
rect 14187 1700 14229 1709
rect 14187 1660 14188 1700
rect 14228 1660 14229 1700
rect 14187 1651 14229 1660
rect 13707 1616 13749 1625
rect 13707 1576 13708 1616
rect 13748 1576 13749 1616
rect 13707 1567 13749 1576
rect 13612 1063 13652 1072
rect 13708 1112 13748 1567
rect 14380 1448 14420 6271
rect 14764 5909 14804 7951
rect 15052 7832 15092 8632
rect 15148 8504 15188 8513
rect 15244 8504 15284 8800
rect 15339 8672 15381 8681
rect 15339 8632 15340 8672
rect 15380 8632 15381 8672
rect 15339 8623 15381 8632
rect 15340 8538 15380 8623
rect 15188 8464 15284 8504
rect 15148 8455 15188 8464
rect 15147 8336 15189 8345
rect 15147 8296 15148 8336
rect 15188 8296 15189 8336
rect 15147 8287 15189 8296
rect 14956 7792 15092 7832
rect 14859 7664 14901 7673
rect 14859 7624 14860 7664
rect 14900 7624 14901 7664
rect 14859 7615 14901 7624
rect 14763 5900 14805 5909
rect 14763 5860 14764 5900
rect 14804 5860 14805 5900
rect 14763 5851 14805 5860
rect 14860 5069 14900 7615
rect 14956 7160 14996 7792
rect 15052 7337 15092 7422
rect 15051 7328 15093 7337
rect 15051 7288 15052 7328
rect 15092 7288 15093 7328
rect 15051 7279 15093 7288
rect 14956 6917 14996 7120
rect 15052 7160 15092 7169
rect 14955 6908 14997 6917
rect 14955 6868 14956 6908
rect 14996 6868 14997 6908
rect 14955 6859 14997 6868
rect 15052 5909 15092 7120
rect 15148 6824 15188 8287
rect 15244 7916 15284 8464
rect 15436 8345 15476 10312
rect 15532 10184 15572 10195
rect 15532 10109 15572 10144
rect 15628 10184 15668 10975
rect 15628 10135 15668 10144
rect 15531 10100 15573 10109
rect 15531 10060 15532 10100
rect 15572 10060 15573 10100
rect 15531 10051 15573 10060
rect 15724 9680 15764 11320
rect 15820 10436 15860 11908
rect 16300 11696 16340 11707
rect 16300 11621 16340 11656
rect 16299 11612 16341 11621
rect 16299 11572 16300 11612
rect 16340 11572 16341 11612
rect 16299 11563 16341 11572
rect 16107 11360 16149 11369
rect 16396 11360 16436 12412
rect 16492 12368 16532 13495
rect 16876 13460 16916 13469
rect 16492 12319 16532 12328
rect 16588 13420 16876 13460
rect 16588 12452 16628 13420
rect 16876 13411 16916 13420
rect 16971 13376 17013 13385
rect 16971 13336 16972 13376
rect 17012 13336 17013 13376
rect 16971 13327 17013 13336
rect 16683 13208 16725 13217
rect 16683 13168 16684 13208
rect 16724 13168 16820 13208
rect 16683 13159 16725 13168
rect 16684 13074 16724 13159
rect 16588 12116 16628 12412
rect 16492 12076 16628 12116
rect 16684 12536 16724 12545
rect 16492 11696 16532 12076
rect 16588 11948 16628 11957
rect 16684 11948 16724 12496
rect 16780 11957 16820 13168
rect 16876 12452 16916 12461
rect 16972 12452 17012 13327
rect 17068 13208 17108 13217
rect 17068 12713 17108 13168
rect 17067 12704 17109 12713
rect 17067 12664 17068 12704
rect 17108 12664 17109 12704
rect 17067 12655 17109 12664
rect 16916 12412 17012 12452
rect 16876 12403 16916 12412
rect 17068 12368 17108 12377
rect 17164 12368 17204 14083
rect 17259 14048 17301 14057
rect 17259 14008 17260 14048
rect 17300 14008 17301 14048
rect 17259 13999 17301 14008
rect 17260 13914 17300 13999
rect 17259 12536 17301 12545
rect 17259 12496 17260 12536
rect 17300 12496 17301 12536
rect 17259 12487 17301 12496
rect 17260 12402 17300 12487
rect 17108 12328 17204 12368
rect 17068 12319 17108 12328
rect 16628 11908 16724 11948
rect 16779 11948 16821 11957
rect 16779 11908 16780 11948
rect 16820 11908 16821 11948
rect 16588 11899 16628 11908
rect 16779 11899 16821 11908
rect 16588 11696 16628 11705
rect 16492 11656 16588 11696
rect 16588 11647 16628 11656
rect 16684 11696 16724 11705
rect 16491 11528 16533 11537
rect 16491 11488 16492 11528
rect 16532 11488 16533 11528
rect 16491 11479 16533 11488
rect 15820 10387 15860 10396
rect 15916 11320 16108 11360
rect 16148 11320 16149 11360
rect 15819 10184 15861 10193
rect 15819 10144 15820 10184
rect 15860 10144 15861 10184
rect 15819 10135 15861 10144
rect 15820 10050 15860 10135
rect 15916 10016 15956 11320
rect 16107 11311 16149 11320
rect 16204 11320 16436 11360
rect 16011 10688 16053 10697
rect 16011 10648 16012 10688
rect 16052 10648 16053 10688
rect 16011 10639 16053 10648
rect 16012 10184 16052 10639
rect 16107 10352 16149 10361
rect 16107 10312 16108 10352
rect 16148 10312 16149 10352
rect 16107 10303 16149 10312
rect 16204 10352 16244 11320
rect 16492 11276 16532 11479
rect 16300 11236 16532 11276
rect 16300 11024 16340 11236
rect 16300 10975 16340 10984
rect 16684 10949 16724 11656
rect 16780 11537 16820 11899
rect 16876 11696 16916 11705
rect 16779 11528 16821 11537
rect 16779 11488 16780 11528
rect 16820 11488 16821 11528
rect 16779 11479 16821 11488
rect 16779 11024 16821 11033
rect 16779 10984 16780 11024
rect 16820 10984 16821 11024
rect 16779 10975 16821 10984
rect 16683 10940 16725 10949
rect 16683 10900 16684 10940
rect 16724 10900 16725 10940
rect 16683 10891 16725 10900
rect 16395 10772 16437 10781
rect 16395 10732 16396 10772
rect 16436 10732 16437 10772
rect 16395 10723 16437 10732
rect 16492 10772 16532 10781
rect 16780 10772 16820 10975
rect 16876 10781 16916 11656
rect 16972 11696 17012 11705
rect 16972 10949 17012 11656
rect 17127 11696 17167 11705
rect 17127 11360 17167 11656
rect 17356 11537 17396 14503
rect 17451 14468 17493 14477
rect 17451 14428 17452 14468
rect 17492 14428 17493 14468
rect 17451 14419 17493 14428
rect 17452 12629 17492 14419
rect 17451 12620 17493 12629
rect 17451 12580 17452 12620
rect 17492 12580 17493 12620
rect 17451 12571 17493 12580
rect 17451 11780 17493 11789
rect 17451 11740 17452 11780
rect 17492 11740 17493 11780
rect 17451 11731 17493 11740
rect 17452 11646 17492 11731
rect 17548 11705 17588 14923
rect 17644 14720 17684 14731
rect 17644 14645 17684 14680
rect 17643 14636 17685 14645
rect 17643 14596 17644 14636
rect 17684 14596 17685 14636
rect 17643 14587 17685 14596
rect 17643 14300 17685 14309
rect 17643 14260 17644 14300
rect 17684 14260 17685 14300
rect 17643 14251 17685 14260
rect 17644 12965 17684 14251
rect 17643 12956 17685 12965
rect 17643 12916 17644 12956
rect 17684 12916 17685 12956
rect 17643 12907 17685 12916
rect 17643 12704 17685 12713
rect 17643 12664 17644 12704
rect 17684 12664 17685 12704
rect 17643 12655 17685 12664
rect 17644 11948 17684 12655
rect 17644 11899 17684 11908
rect 17547 11696 17589 11705
rect 17547 11656 17548 11696
rect 17588 11656 17589 11696
rect 17547 11647 17589 11656
rect 17355 11528 17397 11537
rect 17355 11488 17356 11528
rect 17396 11488 17397 11528
rect 17355 11479 17397 11488
rect 17740 11360 17780 15772
rect 17932 15401 17972 18283
rect 17931 15392 17973 15401
rect 17931 15352 17932 15392
rect 17972 15352 17973 15392
rect 17931 15343 17973 15352
rect 17835 13124 17877 13133
rect 17835 13084 17836 13124
rect 17876 13084 17877 13124
rect 17835 13075 17877 13084
rect 17836 11948 17876 13075
rect 18028 12713 18068 19963
rect 18124 19962 18164 20047
rect 18220 19265 18260 20140
rect 18316 20054 18356 20063
rect 18508 20054 18548 20299
rect 18604 20273 18644 20728
rect 18700 20768 18740 21568
rect 18796 21557 18836 21568
rect 19084 21615 19124 21652
rect 19084 21566 19124 21575
rect 19276 21608 19316 21652
rect 19276 21533 19316 21568
rect 19372 21608 19412 21617
rect 19275 21524 19317 21533
rect 19275 21484 19276 21524
rect 19316 21484 19317 21524
rect 19275 21475 19317 21484
rect 19372 21365 19412 21568
rect 19467 21608 19509 21617
rect 19467 21568 19468 21608
rect 19508 21568 19509 21608
rect 19467 21559 19509 21568
rect 19564 21608 19604 21617
rect 19756 21608 19796 21617
rect 19604 21568 19756 21608
rect 19564 21559 19604 21568
rect 19756 21559 19796 21568
rect 19948 21608 19988 21619
rect 19468 21474 19508 21559
rect 19948 21533 19988 21568
rect 20044 21608 20084 21727
rect 20044 21559 20084 21568
rect 19947 21524 19989 21533
rect 19947 21484 19948 21524
rect 19988 21484 19989 21524
rect 19947 21475 19989 21484
rect 19755 21440 19797 21449
rect 19755 21400 19756 21440
rect 19796 21400 19797 21440
rect 19755 21391 19797 21400
rect 19084 21356 19124 21365
rect 19371 21356 19413 21365
rect 19124 21316 19316 21356
rect 19084 21307 19124 21316
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 19276 21104 19316 21316
rect 19371 21316 19372 21356
rect 19412 21316 19413 21356
rect 19371 21307 19413 21316
rect 19207 21064 19316 21104
rect 19207 21020 19247 21064
rect 19372 21029 19412 21307
rect 19756 21306 19796 21391
rect 18700 20719 18740 20728
rect 18988 20980 19247 21020
rect 19371 21020 19413 21029
rect 19371 20980 19372 21020
rect 19412 20980 19413 21020
rect 18603 20264 18645 20273
rect 18603 20224 18604 20264
rect 18644 20224 18645 20264
rect 18603 20215 18645 20224
rect 18988 20105 19028 20980
rect 19371 20971 19413 20980
rect 19563 21020 19605 21029
rect 19563 20980 19564 21020
rect 19604 20980 19605 21020
rect 19563 20971 19605 20980
rect 19276 20936 19316 20945
rect 19083 20852 19125 20861
rect 19083 20812 19084 20852
rect 19124 20812 19125 20852
rect 19083 20803 19125 20812
rect 19180 20852 19220 20861
rect 19084 20768 19124 20803
rect 19084 20717 19124 20728
rect 19180 20516 19220 20812
rect 19084 20476 19220 20516
rect 18316 19853 18356 20014
rect 18412 20014 18548 20054
rect 18700 20096 18740 20105
rect 18412 20012 18452 20014
rect 18412 19963 18452 19972
rect 18604 20012 18644 20021
rect 18508 19886 18548 19895
rect 18315 19844 18357 19853
rect 18315 19804 18316 19844
rect 18356 19804 18357 19844
rect 18315 19795 18357 19804
rect 18508 19685 18548 19846
rect 18507 19676 18549 19685
rect 18507 19636 18508 19676
rect 18548 19636 18549 19676
rect 18507 19627 18549 19636
rect 18219 19256 18261 19265
rect 18219 19216 18220 19256
rect 18260 19216 18261 19256
rect 18219 19207 18261 19216
rect 18604 18761 18644 19972
rect 18700 18929 18740 20056
rect 18987 20096 19029 20105
rect 18987 20056 18988 20096
rect 19028 20056 19029 20096
rect 18987 20047 19029 20056
rect 18892 19928 18932 19937
rect 19084 19928 19124 20476
rect 19276 20357 19316 20896
rect 19372 20852 19412 20861
rect 19275 20348 19317 20357
rect 19275 20308 19276 20348
rect 19316 20308 19317 20348
rect 19275 20299 19317 20308
rect 19275 20180 19317 20189
rect 19275 20140 19276 20180
rect 19316 20140 19317 20180
rect 19275 20131 19317 20140
rect 18932 19888 19124 19928
rect 19180 20096 19220 20105
rect 18892 19879 18932 19888
rect 19180 19844 19220 20056
rect 19276 20096 19316 20131
rect 19276 20045 19316 20056
rect 19180 19804 19316 19844
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 18988 19256 19028 19265
rect 18699 18920 18741 18929
rect 18699 18880 18700 18920
rect 18740 18880 18741 18920
rect 18699 18871 18741 18880
rect 18603 18752 18645 18761
rect 18603 18712 18604 18752
rect 18644 18712 18645 18752
rect 18603 18703 18645 18712
rect 18411 18668 18453 18677
rect 18411 18628 18412 18668
rect 18452 18628 18453 18668
rect 18411 18619 18453 18628
rect 18219 18416 18261 18425
rect 18219 18376 18220 18416
rect 18260 18376 18261 18416
rect 18219 18367 18261 18376
rect 18123 18080 18165 18089
rect 18123 18040 18124 18080
rect 18164 18040 18165 18080
rect 18123 18031 18165 18040
rect 18124 14804 18164 18031
rect 18124 14755 18164 14764
rect 18220 13040 18260 18367
rect 18315 16736 18357 16745
rect 18315 16696 18316 16736
rect 18356 16696 18357 16736
rect 18315 16687 18357 16696
rect 18316 14972 18356 16687
rect 18412 15317 18452 18619
rect 18988 18584 19028 19216
rect 19179 19256 19221 19265
rect 19179 19216 19180 19256
rect 19220 19216 19221 19256
rect 19179 19207 19221 19216
rect 19180 19172 19220 19207
rect 19180 19121 19220 19132
rect 19276 18845 19316 19804
rect 19372 19013 19412 20812
rect 19468 20768 19508 20777
rect 19468 19433 19508 20728
rect 19564 20441 19604 20971
rect 20044 20936 20084 20945
rect 19852 20896 20044 20936
rect 19660 20768 19700 20777
rect 19563 20432 19605 20441
rect 19563 20392 19564 20432
rect 19604 20392 19605 20432
rect 19563 20383 19605 20392
rect 19564 20096 19604 20105
rect 19467 19424 19509 19433
rect 19467 19384 19468 19424
rect 19508 19384 19509 19424
rect 19467 19375 19509 19384
rect 19467 19256 19509 19265
rect 19564 19256 19604 20056
rect 19660 19601 19700 20728
rect 19852 20768 19892 20896
rect 20044 20887 20084 20896
rect 19852 20719 19892 20728
rect 20044 20768 20084 20779
rect 20044 20693 20084 20728
rect 20235 20768 20277 20777
rect 20235 20728 20236 20768
rect 20276 20728 20277 20768
rect 20235 20719 20277 20728
rect 20043 20684 20085 20693
rect 20043 20644 20044 20684
rect 20084 20644 20085 20684
rect 20043 20635 20085 20644
rect 20236 20634 20276 20719
rect 19755 20600 19797 20609
rect 19755 20560 19756 20600
rect 19796 20560 19797 20600
rect 19755 20551 19797 20560
rect 19756 20466 19796 20551
rect 19851 20432 19893 20441
rect 19851 20392 19852 20432
rect 19892 20392 19893 20432
rect 19851 20383 19893 20392
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 19852 20096 19892 20383
rect 19852 20047 19892 20056
rect 19948 20096 19988 20107
rect 19948 20021 19988 20056
rect 20140 20054 20180 20063
rect 19947 20012 19989 20021
rect 19947 19972 19948 20012
rect 19988 19972 19989 20012
rect 19947 19963 19989 19972
rect 19947 19844 19989 19853
rect 19947 19804 19948 19844
rect 19988 19804 19989 19844
rect 19947 19795 19989 19804
rect 19948 19710 19988 19795
rect 20140 19676 20180 20014
rect 20811 19928 20853 19937
rect 20811 19888 20812 19928
rect 20852 19888 20853 19928
rect 20811 19879 20853 19888
rect 20140 19636 20276 19676
rect 19659 19592 19701 19601
rect 19659 19552 19660 19592
rect 19700 19552 19701 19592
rect 19659 19543 19701 19552
rect 19659 19424 19701 19433
rect 19659 19384 19660 19424
rect 19700 19384 19701 19424
rect 19659 19375 19701 19384
rect 19467 19216 19468 19256
rect 19508 19216 19604 19256
rect 19467 19207 19509 19216
rect 19468 19122 19508 19207
rect 19371 19004 19413 19013
rect 19371 18964 19372 19004
rect 19412 18964 19413 19004
rect 19371 18955 19413 18964
rect 19563 18920 19605 18929
rect 19563 18880 19564 18920
rect 19604 18880 19605 18920
rect 19563 18871 19605 18880
rect 19275 18836 19317 18845
rect 19275 18796 19276 18836
rect 19316 18796 19317 18836
rect 19275 18787 19317 18796
rect 19179 18752 19221 18761
rect 19179 18712 19180 18752
rect 19220 18712 19221 18752
rect 19179 18703 19221 18712
rect 19371 18752 19413 18761
rect 19371 18712 19372 18752
rect 19412 18712 19413 18752
rect 19371 18703 19413 18712
rect 19564 18752 19604 18871
rect 19564 18703 19604 18712
rect 19180 18618 19220 18703
rect 18700 18544 18988 18584
rect 18700 17996 18740 18544
rect 18988 18535 19028 18544
rect 19372 18584 19412 18703
rect 19660 18593 19700 19375
rect 19756 19256 19796 19267
rect 20236 19265 20276 19636
rect 19756 19181 19796 19216
rect 20235 19256 20277 19265
rect 20235 19216 20236 19256
rect 20276 19216 20277 19256
rect 20235 19207 20277 19216
rect 19755 19172 19797 19181
rect 19755 19132 19756 19172
rect 19796 19132 19797 19172
rect 19755 19123 19797 19132
rect 19852 19172 19892 19183
rect 19852 19097 19892 19132
rect 20140 19097 20180 19141
rect 19851 19088 19893 19097
rect 19851 19048 19852 19088
rect 19892 19048 19893 19088
rect 19851 19039 19893 19048
rect 20139 19088 20181 19097
rect 20139 19048 20140 19088
rect 20180 19048 20181 19088
rect 20139 19046 20181 19048
rect 20139 19039 20140 19046
rect 19755 19004 19797 19013
rect 19755 18964 19756 19004
rect 19796 18964 19797 19004
rect 19755 18955 19797 18964
rect 19372 18535 19412 18544
rect 19468 18584 19508 18593
rect 19468 18341 19508 18544
rect 19659 18584 19701 18593
rect 19659 18544 19660 18584
rect 19700 18544 19701 18584
rect 19659 18535 19701 18544
rect 19756 18584 19796 18955
rect 19852 18761 19892 19039
rect 20180 19039 20181 19046
rect 20140 18997 20180 19006
rect 19947 18920 19989 18929
rect 19947 18880 19948 18920
rect 19988 18880 19989 18920
rect 19947 18871 19989 18880
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 19851 18752 19893 18761
rect 19851 18712 19852 18752
rect 19892 18712 19893 18752
rect 19851 18703 19893 18712
rect 19948 18593 19988 18871
rect 20331 18752 20373 18761
rect 20331 18712 20332 18752
rect 20372 18712 20373 18752
rect 20331 18703 20373 18712
rect 19660 18450 19700 18535
rect 19756 18341 19796 18544
rect 19911 18584 19988 18593
rect 19951 18544 19988 18584
rect 20140 18584 20180 18593
rect 19911 18535 19951 18544
rect 19467 18332 19509 18341
rect 19467 18292 19468 18332
rect 19508 18292 19509 18332
rect 19467 18283 19509 18292
rect 19755 18332 19797 18341
rect 19755 18292 19756 18332
rect 19796 18292 19797 18332
rect 19755 18283 19797 18292
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 20140 18089 20180 18544
rect 20235 18332 20277 18341
rect 20235 18292 20236 18332
rect 20276 18292 20277 18332
rect 20235 18283 20277 18292
rect 20139 18080 20181 18089
rect 20139 18040 20140 18080
rect 20180 18040 20181 18080
rect 20139 18031 20181 18040
rect 19179 17996 19221 18005
rect 18700 17956 19028 17996
rect 18988 17744 19028 17956
rect 19179 17956 19180 17996
rect 19220 17956 19221 17996
rect 19179 17947 19221 17956
rect 19947 17996 19989 18005
rect 19947 17956 19948 17996
rect 19988 17956 19989 17996
rect 19947 17947 19989 17956
rect 19180 17862 19220 17947
rect 19948 17862 19988 17947
rect 19371 17828 19413 17837
rect 19371 17788 19372 17828
rect 19412 17788 19413 17828
rect 19371 17779 19413 17788
rect 19755 17828 19797 17837
rect 19755 17788 19756 17828
rect 19796 17788 19797 17828
rect 19755 17779 19797 17788
rect 18988 17333 19028 17704
rect 19372 17694 19412 17779
rect 19756 17694 19796 17779
rect 19947 17660 19989 17669
rect 19947 17620 19948 17660
rect 19988 17620 19989 17660
rect 19947 17611 19989 17620
rect 19564 17576 19604 17585
rect 19468 17536 19564 17576
rect 19179 17408 19221 17417
rect 19179 17368 19180 17408
rect 19220 17368 19221 17408
rect 19179 17359 19221 17368
rect 18603 17324 18645 17333
rect 18603 17284 18604 17324
rect 18644 17284 18645 17324
rect 18603 17275 18645 17284
rect 18987 17324 19029 17333
rect 18987 17284 18988 17324
rect 19028 17284 19029 17324
rect 18987 17275 19029 17284
rect 18604 17072 18644 17275
rect 18795 17156 18837 17165
rect 18795 17116 18796 17156
rect 18836 17116 18837 17156
rect 18795 17107 18837 17116
rect 18507 16232 18549 16241
rect 18507 16192 18508 16232
rect 18548 16192 18549 16232
rect 18507 16183 18549 16192
rect 18604 16232 18644 17032
rect 18796 17022 18836 17107
rect 18988 17072 19028 17081
rect 18988 16829 19028 17032
rect 19084 16988 19124 16999
rect 19084 16913 19124 16948
rect 19083 16904 19125 16913
rect 19083 16864 19084 16904
rect 19124 16864 19125 16904
rect 19083 16855 19125 16864
rect 19180 16904 19220 17359
rect 19372 17072 19412 17081
rect 19180 16855 19220 16864
rect 19276 16988 19316 16997
rect 18987 16820 19029 16829
rect 18987 16780 18988 16820
rect 19028 16780 19029 16820
rect 18987 16771 19029 16780
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 18892 16400 18932 16409
rect 19276 16400 19316 16948
rect 18932 16360 19316 16400
rect 18892 16351 18932 16360
rect 18700 16232 18740 16241
rect 19180 16232 19220 16360
rect 18604 16192 18700 16232
rect 18740 16192 18932 16232
rect 18508 16073 18548 16183
rect 18507 16064 18549 16073
rect 18507 16024 18508 16064
rect 18548 16024 18549 16064
rect 18507 16015 18549 16024
rect 18411 15308 18453 15317
rect 18411 15268 18412 15308
rect 18452 15268 18453 15308
rect 18411 15259 18453 15268
rect 18411 15140 18453 15149
rect 18411 15100 18412 15140
rect 18452 15100 18453 15140
rect 18411 15091 18453 15100
rect 18316 14923 18356 14932
rect 18412 14048 18452 15091
rect 18508 14720 18548 16015
rect 18604 15149 18644 16192
rect 18700 16183 18740 16192
rect 18892 15560 18932 16192
rect 19180 16183 19220 16192
rect 19276 16232 19316 16241
rect 19276 15569 19316 16192
rect 19372 16064 19412 17032
rect 19468 16577 19508 17536
rect 19564 17527 19604 17536
rect 19948 17081 19988 17611
rect 20236 17576 20276 18283
rect 20332 17753 20372 18703
rect 20619 18584 20661 18593
rect 20619 18544 20620 18584
rect 20660 18544 20661 18584
rect 20619 18535 20661 18544
rect 20331 17744 20373 17753
rect 20331 17704 20332 17744
rect 20372 17704 20373 17744
rect 20331 17695 20373 17704
rect 20236 17536 20564 17576
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20126 17156 20168 17165
rect 20126 17116 20127 17156
rect 20167 17116 20168 17156
rect 20126 17107 20168 17116
rect 20127 17083 20167 17107
rect 19564 17072 19604 17081
rect 19467 16568 19509 16577
rect 19467 16528 19468 16568
rect 19508 16528 19509 16568
rect 19467 16519 19509 16528
rect 19564 16400 19604 17032
rect 19947 17072 19989 17081
rect 19947 17032 19948 17072
rect 19988 17032 19989 17072
rect 19947 17023 19989 17032
rect 19659 16988 19701 16997
rect 19659 16948 19660 16988
rect 19700 16948 19701 16988
rect 19659 16939 19701 16948
rect 19852 16988 19892 16997
rect 19660 16493 19700 16939
rect 19755 16904 19797 16913
rect 19755 16864 19756 16904
rect 19796 16864 19797 16904
rect 19755 16855 19797 16864
rect 19756 16770 19796 16855
rect 19659 16484 19701 16493
rect 19659 16444 19660 16484
rect 19700 16444 19701 16484
rect 19659 16435 19701 16444
rect 19372 16015 19412 16024
rect 19468 16360 19604 16400
rect 19468 16232 19508 16360
rect 19371 15896 19413 15905
rect 19371 15856 19372 15896
rect 19412 15856 19413 15896
rect 19371 15847 19413 15856
rect 18892 15511 18932 15520
rect 19275 15560 19317 15569
rect 19275 15520 19276 15560
rect 19316 15520 19317 15560
rect 19275 15511 19317 15520
rect 19372 15560 19412 15847
rect 19084 15308 19124 15317
rect 19372 15308 19412 15520
rect 19468 15485 19508 16192
rect 19563 16232 19605 16241
rect 19563 16192 19564 16232
rect 19604 16192 19605 16232
rect 19563 16183 19605 16192
rect 19721 16239 19761 16248
rect 19761 16199 19796 16239
rect 19721 16190 19796 16199
rect 19467 15476 19509 15485
rect 19467 15436 19468 15476
rect 19508 15436 19509 15476
rect 19467 15427 19509 15436
rect 19124 15268 19412 15308
rect 19084 15259 19124 15268
rect 18603 15140 18645 15149
rect 18603 15100 18604 15140
rect 18644 15100 18645 15140
rect 18603 15091 18645 15100
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 18603 14888 18645 14897
rect 18603 14848 18604 14888
rect 18644 14848 18645 14888
rect 18603 14839 18645 14848
rect 18508 14671 18548 14680
rect 18604 14720 18644 14839
rect 19083 14804 19125 14813
rect 19083 14764 19084 14804
rect 19124 14764 19125 14804
rect 19083 14755 19125 14764
rect 18796 14720 18836 14729
rect 18508 14048 18548 14057
rect 18316 14008 18508 14048
rect 18316 13217 18356 14008
rect 18508 13999 18548 14008
rect 18411 13544 18453 13553
rect 18411 13504 18412 13544
rect 18452 13504 18453 13544
rect 18411 13495 18453 13504
rect 18315 13208 18357 13217
rect 18315 13168 18316 13208
rect 18356 13168 18357 13208
rect 18315 13159 18357 13168
rect 18220 13000 18356 13040
rect 18027 12704 18069 12713
rect 18027 12664 18028 12704
rect 18068 12664 18069 12704
rect 18027 12655 18069 12664
rect 18027 12536 18069 12545
rect 18027 12496 18028 12536
rect 18068 12496 18069 12536
rect 18027 12487 18069 12496
rect 17836 11899 17876 11908
rect 17835 11696 17877 11705
rect 17835 11656 17836 11696
rect 17876 11656 17877 11696
rect 17835 11647 17877 11656
rect 18028 11696 18068 12487
rect 18028 11647 18068 11656
rect 18220 11696 18260 11707
rect 17836 11562 17876 11647
rect 18220 11621 18260 11656
rect 18219 11612 18261 11621
rect 18219 11572 18220 11612
rect 18260 11572 18261 11612
rect 18219 11563 18261 11572
rect 17127 11320 17492 11360
rect 17740 11320 17972 11360
rect 17068 11024 17108 11033
rect 16971 10940 17013 10949
rect 16971 10900 16972 10940
rect 17012 10900 17013 10940
rect 16971 10891 17013 10900
rect 16532 10732 16820 10772
rect 16875 10772 16917 10781
rect 16875 10732 16876 10772
rect 16916 10732 16917 10772
rect 16299 10436 16341 10445
rect 16299 10396 16300 10436
rect 16340 10396 16341 10436
rect 16299 10387 16341 10396
rect 16204 10303 16244 10312
rect 16108 10268 16148 10303
rect 16108 10217 16148 10228
rect 16300 10268 16340 10387
rect 16300 10219 16340 10228
rect 16012 10135 16052 10144
rect 16396 10184 16436 10723
rect 16492 10193 16532 10732
rect 16875 10723 16917 10732
rect 16683 10604 16725 10613
rect 16683 10564 16684 10604
rect 16724 10564 16725 10604
rect 16683 10555 16725 10564
rect 16587 10352 16629 10361
rect 16587 10312 16588 10352
rect 16628 10312 16629 10352
rect 16587 10303 16629 10312
rect 16588 10218 16628 10303
rect 16396 10135 16436 10144
rect 16491 10184 16533 10193
rect 16491 10144 16492 10184
rect 16532 10144 16533 10184
rect 16491 10135 16533 10144
rect 16299 10016 16341 10025
rect 15916 9976 16148 10016
rect 16011 9764 16053 9773
rect 16011 9724 16012 9764
rect 16052 9724 16053 9764
rect 16011 9715 16053 9724
rect 15532 9640 15764 9680
rect 15435 8336 15477 8345
rect 15435 8296 15436 8336
rect 15476 8296 15477 8336
rect 15435 8287 15477 8296
rect 15435 8084 15477 8093
rect 15435 8044 15436 8084
rect 15476 8044 15477 8084
rect 15435 8035 15477 8044
rect 15436 8000 15476 8035
rect 15244 7876 15380 7916
rect 15244 7748 15284 7757
rect 15244 7421 15284 7708
rect 15243 7412 15285 7421
rect 15243 7372 15244 7412
rect 15284 7372 15285 7412
rect 15243 7363 15285 7372
rect 15340 7337 15380 7876
rect 15436 7673 15476 7960
rect 15435 7664 15477 7673
rect 15435 7624 15436 7664
rect 15476 7624 15477 7664
rect 15532 7664 15572 9640
rect 15915 9596 15957 9605
rect 15915 9556 15916 9596
rect 15956 9556 15957 9596
rect 15915 9547 15957 9556
rect 15628 9512 15668 9521
rect 15628 9185 15668 9472
rect 15819 9512 15861 9521
rect 15819 9472 15820 9512
rect 15860 9472 15861 9512
rect 15819 9463 15861 9472
rect 15724 9428 15764 9437
rect 15724 9269 15764 9388
rect 15820 9344 15860 9463
rect 15916 9428 15956 9547
rect 16012 9512 16052 9715
rect 16012 9463 16052 9472
rect 15916 9379 15956 9388
rect 15820 9295 15860 9304
rect 15723 9260 15765 9269
rect 15723 9220 15724 9260
rect 15764 9220 15765 9260
rect 15723 9211 15765 9220
rect 15627 9176 15669 9185
rect 15627 9136 15628 9176
rect 15668 9136 15669 9176
rect 16108 9176 16148 9976
rect 16299 9976 16300 10016
rect 16340 9976 16341 10016
rect 16299 9967 16341 9976
rect 16300 9689 16340 9967
rect 16299 9680 16341 9689
rect 16299 9640 16300 9680
rect 16340 9640 16341 9680
rect 16299 9631 16341 9640
rect 16587 9680 16629 9689
rect 16587 9640 16588 9680
rect 16628 9640 16629 9680
rect 16587 9631 16629 9640
rect 16204 9512 16244 9523
rect 16204 9437 16244 9472
rect 16299 9512 16341 9521
rect 16299 9472 16300 9512
rect 16340 9472 16341 9512
rect 16299 9463 16341 9472
rect 16491 9512 16533 9521
rect 16491 9472 16492 9512
rect 16532 9472 16533 9512
rect 16491 9463 16533 9472
rect 16588 9512 16628 9631
rect 16588 9463 16628 9472
rect 16203 9428 16245 9437
rect 16203 9388 16204 9428
rect 16244 9388 16245 9428
rect 16203 9379 16245 9388
rect 16300 9428 16340 9463
rect 16300 9377 16340 9388
rect 16492 9428 16532 9463
rect 16492 9377 16532 9388
rect 16395 9344 16437 9353
rect 16395 9304 16396 9344
rect 16436 9304 16437 9344
rect 16395 9295 16437 9304
rect 16396 9210 16436 9295
rect 16108 9136 16340 9176
rect 15627 9127 15669 9136
rect 16203 9008 16245 9017
rect 16203 8968 16204 9008
rect 16244 8968 16245 9008
rect 16203 8959 16245 8968
rect 15627 7664 15669 7673
rect 15532 7624 15628 7664
rect 15668 7624 15669 7664
rect 15435 7615 15477 7624
rect 15627 7615 15669 7624
rect 15339 7328 15381 7337
rect 15339 7288 15340 7328
rect 15380 7288 15381 7328
rect 15339 7279 15381 7288
rect 15627 7328 15669 7337
rect 15627 7288 15628 7328
rect 15668 7288 15669 7328
rect 15627 7279 15669 7288
rect 15435 7244 15477 7253
rect 15435 7204 15436 7244
rect 15476 7204 15477 7244
rect 15435 7195 15477 7204
rect 15532 7244 15572 7253
rect 15244 7160 15284 7169
rect 15436 7160 15476 7195
rect 15284 7120 15380 7160
rect 15244 7111 15284 7120
rect 15340 6992 15380 7120
rect 15436 7109 15476 7120
rect 15532 7001 15572 7204
rect 15628 7194 15668 7279
rect 15731 7253 16148 7286
rect 15724 7246 16148 7253
rect 15724 7244 15771 7246
rect 15764 7204 15771 7244
rect 15724 7195 15764 7204
rect 15820 7160 15860 7169
rect 15531 6992 15573 7001
rect 15340 6952 15476 6992
rect 15148 6784 15284 6824
rect 15147 6656 15189 6665
rect 15147 6616 15148 6656
rect 15188 6616 15189 6656
rect 15147 6607 15189 6616
rect 15051 5900 15093 5909
rect 15051 5860 15052 5900
rect 15092 5860 15093 5900
rect 15051 5851 15093 5860
rect 14859 5060 14901 5069
rect 14859 5020 14860 5060
rect 14900 5020 14901 5060
rect 14859 5011 14901 5020
rect 14475 4976 14517 4985
rect 14475 4936 14476 4976
rect 14516 4936 14517 4976
rect 14475 4927 14517 4936
rect 14476 3809 14516 4927
rect 14475 3800 14517 3809
rect 15148 3800 15188 6607
rect 14475 3760 14476 3800
rect 14516 3760 14517 3800
rect 14475 3751 14517 3760
rect 15052 3760 15188 3800
rect 15052 3389 15092 3760
rect 15147 3632 15189 3641
rect 15147 3592 15148 3632
rect 15188 3592 15189 3632
rect 15147 3583 15189 3592
rect 15148 3464 15188 3583
rect 15148 3415 15188 3424
rect 15051 3380 15093 3389
rect 15051 3340 15052 3380
rect 15092 3340 15093 3380
rect 15051 3331 15093 3340
rect 15147 3296 15189 3305
rect 15147 3256 15148 3296
rect 15188 3256 15189 3296
rect 15147 3247 15189 3256
rect 15148 2801 15188 3247
rect 14955 2792 14997 2801
rect 14955 2752 14956 2792
rect 14996 2752 14997 2792
rect 14955 2743 14997 2752
rect 15147 2792 15189 2801
rect 15147 2752 15148 2792
rect 15188 2752 15189 2792
rect 15147 2743 15189 2752
rect 14092 1408 14420 1448
rect 14860 1952 14900 1961
rect 13899 1196 13941 1205
rect 13899 1156 13900 1196
rect 13940 1156 13941 1196
rect 13899 1147 13941 1156
rect 13708 1063 13748 1072
rect 13420 978 13460 1063
rect 13900 1062 13940 1147
rect 13515 944 13557 953
rect 13515 904 13516 944
rect 13556 904 13557 944
rect 13515 895 13557 904
rect 13707 944 13749 953
rect 13707 904 13708 944
rect 13748 904 13749 944
rect 13707 895 13749 904
rect 13516 80 13556 895
rect 13708 80 13748 895
rect 13899 692 13941 701
rect 13899 652 13900 692
rect 13940 652 13941 692
rect 13899 643 13941 652
rect 13900 80 13940 643
rect 14092 80 14132 1408
rect 14283 1280 14325 1289
rect 14283 1240 14284 1280
rect 14324 1240 14325 1280
rect 14283 1231 14325 1240
rect 14475 1280 14517 1289
rect 14475 1240 14476 1280
rect 14516 1240 14517 1280
rect 14188 944 14228 953
rect 14188 617 14228 904
rect 14187 608 14229 617
rect 14187 568 14188 608
rect 14228 568 14229 608
rect 14187 559 14229 568
rect 14284 80 14324 1231
rect 14380 1205 14420 1236
rect 14475 1231 14517 1240
rect 14667 1280 14709 1289
rect 14667 1240 14668 1280
rect 14708 1240 14709 1280
rect 14667 1231 14709 1240
rect 14379 1196 14421 1205
rect 14379 1156 14380 1196
rect 14420 1156 14421 1196
rect 14379 1147 14421 1156
rect 14380 1112 14420 1147
rect 14380 197 14420 1072
rect 14379 188 14421 197
rect 14379 148 14380 188
rect 14420 148 14421 188
rect 14379 139 14421 148
rect 14476 80 14516 1231
rect 14668 80 14708 1231
rect 14860 1205 14900 1912
rect 14859 1196 14901 1205
rect 14859 1156 14860 1196
rect 14900 1156 14901 1196
rect 14859 1147 14901 1156
rect 14956 1121 14996 2743
rect 15148 2288 15188 2743
rect 15244 2624 15284 6784
rect 15340 5648 15380 5657
rect 15340 4976 15380 5608
rect 15436 5573 15476 6952
rect 15531 6952 15532 6992
rect 15572 6952 15573 6992
rect 15531 6943 15573 6952
rect 15820 6329 15860 7120
rect 16011 7160 16053 7169
rect 16011 7120 16012 7160
rect 16052 7120 16053 7160
rect 16011 7111 16053 7120
rect 15915 7076 15957 7085
rect 15915 7036 15916 7076
rect 15956 7036 15957 7076
rect 15915 7027 15957 7036
rect 15916 6488 15956 7027
rect 16012 7026 16052 7111
rect 16108 6749 16148 7246
rect 16107 6740 16149 6749
rect 16107 6700 16108 6740
rect 16148 6700 16149 6740
rect 16107 6691 16149 6700
rect 16108 6656 16148 6691
rect 16108 6606 16148 6616
rect 15819 6320 15861 6329
rect 15819 6280 15820 6320
rect 15860 6280 15861 6320
rect 15819 6271 15861 6280
rect 15916 6245 15956 6448
rect 15915 6236 15957 6245
rect 15915 6196 15916 6236
rect 15956 6196 15957 6236
rect 15915 6187 15957 6196
rect 15531 5900 15573 5909
rect 15531 5860 15532 5900
rect 15572 5860 15573 5900
rect 16204 5900 16244 8959
rect 16300 8093 16340 9136
rect 16684 9092 16724 10555
rect 16779 10520 16821 10529
rect 16779 10480 16780 10520
rect 16820 10480 16821 10520
rect 16779 10471 16821 10480
rect 16780 9857 16820 10471
rect 16972 10445 17012 10891
rect 17068 10529 17108 10984
rect 17164 11024 17204 11033
rect 17204 10984 17396 11024
rect 17164 10975 17204 10984
rect 17163 10856 17205 10865
rect 17163 10816 17164 10856
rect 17204 10816 17205 10856
rect 17163 10807 17205 10816
rect 17067 10520 17109 10529
rect 17067 10480 17068 10520
rect 17108 10480 17109 10520
rect 17067 10471 17109 10480
rect 16971 10436 17013 10445
rect 16971 10396 16972 10436
rect 17012 10396 17013 10436
rect 16971 10387 17013 10396
rect 16875 10352 16917 10361
rect 16875 10312 16876 10352
rect 16916 10312 16917 10352
rect 16875 10303 16917 10312
rect 16876 10184 16916 10303
rect 16876 10135 16916 10144
rect 16972 10184 17012 10193
rect 16779 9848 16821 9857
rect 16779 9808 16780 9848
rect 16820 9808 16821 9848
rect 16779 9799 16821 9808
rect 16875 9512 16917 9521
rect 16875 9472 16876 9512
rect 16916 9472 16917 9512
rect 16875 9463 16917 9472
rect 16779 9260 16821 9269
rect 16779 9220 16780 9260
rect 16820 9220 16821 9260
rect 16779 9211 16821 9220
rect 16780 9126 16820 9211
rect 16396 9052 16724 9092
rect 16299 8084 16341 8093
rect 16299 8044 16300 8084
rect 16340 8044 16341 8084
rect 16299 8035 16341 8044
rect 16300 7841 16340 8035
rect 16299 7832 16341 7841
rect 16299 7792 16300 7832
rect 16340 7792 16341 7832
rect 16299 7783 16341 7792
rect 16396 6833 16436 9052
rect 16780 8924 16820 8933
rect 16876 8924 16916 9463
rect 16972 9428 17012 10144
rect 17164 9941 17204 10807
rect 17259 10184 17301 10193
rect 17259 10144 17260 10184
rect 17300 10144 17301 10184
rect 17259 10135 17301 10144
rect 17260 10050 17300 10135
rect 17163 9932 17205 9941
rect 17163 9892 17164 9932
rect 17204 9892 17205 9932
rect 17163 9883 17205 9892
rect 17164 9680 17204 9883
rect 17068 9640 17204 9680
rect 17068 9596 17108 9640
rect 17356 9596 17396 10984
rect 17452 10856 17492 11320
rect 17644 11024 17684 11035
rect 17644 10949 17684 10984
rect 17835 11024 17877 11033
rect 17835 10984 17836 11024
rect 17876 10984 17877 11024
rect 17835 10975 17877 10984
rect 17643 10940 17685 10949
rect 17643 10900 17644 10940
rect 17684 10900 17685 10940
rect 17643 10891 17685 10900
rect 17836 10890 17876 10975
rect 17452 10807 17492 10816
rect 17643 10772 17685 10781
rect 17643 10732 17644 10772
rect 17684 10732 17685 10772
rect 17643 10723 17685 10732
rect 17644 10638 17684 10723
rect 17739 10688 17781 10697
rect 17739 10648 17740 10688
rect 17780 10648 17781 10688
rect 17739 10639 17781 10648
rect 17643 10520 17685 10529
rect 17548 10480 17644 10520
rect 17684 10480 17685 10520
rect 17451 10352 17493 10361
rect 17451 10312 17452 10352
rect 17492 10312 17493 10352
rect 17451 10303 17493 10312
rect 17452 9848 17492 10303
rect 17548 10025 17588 10480
rect 17643 10471 17685 10480
rect 17643 10352 17685 10361
rect 17643 10312 17644 10352
rect 17684 10312 17685 10352
rect 17643 10303 17685 10312
rect 17740 10352 17780 10639
rect 17932 10604 17972 11320
rect 18124 11201 18164 11286
rect 18123 11192 18165 11201
rect 18123 11152 18124 11192
rect 18164 11152 18165 11192
rect 18123 11143 18165 11152
rect 18028 11024 18068 11033
rect 18219 11024 18261 11033
rect 18068 10984 18164 11024
rect 18028 10975 18068 10984
rect 17932 10564 18068 10604
rect 17740 10303 17780 10312
rect 17644 10184 17684 10303
rect 17740 10184 17780 10193
rect 17644 10144 17740 10184
rect 17740 10135 17780 10144
rect 17835 10100 17877 10109
rect 17835 10060 17836 10100
rect 17876 10060 17877 10100
rect 17835 10051 17877 10060
rect 17547 10016 17589 10025
rect 17547 9976 17548 10016
rect 17588 9976 17589 10016
rect 17547 9967 17589 9976
rect 17452 9808 17588 9848
rect 17068 9547 17108 9556
rect 17164 9556 17396 9596
rect 17164 9512 17204 9556
rect 17452 9512 17492 9521
rect 16972 9388 17108 9428
rect 16971 9260 17013 9269
rect 16971 9220 16972 9260
rect 17012 9220 17013 9260
rect 16971 9211 17013 9220
rect 16820 8884 16916 8924
rect 16780 8875 16820 8884
rect 16588 8672 16628 8681
rect 16779 8672 16821 8681
rect 16628 8632 16724 8672
rect 16588 8623 16628 8632
rect 16587 8420 16629 8429
rect 16587 8380 16588 8420
rect 16628 8380 16629 8420
rect 16587 8371 16629 8380
rect 16588 7085 16628 8371
rect 16684 8252 16724 8632
rect 16779 8632 16780 8672
rect 16820 8632 16821 8672
rect 16779 8623 16821 8632
rect 16780 8429 16820 8623
rect 16779 8420 16821 8429
rect 16779 8380 16780 8420
rect 16820 8380 16821 8420
rect 16779 8371 16821 8380
rect 16684 8212 16820 8252
rect 16684 8093 16724 8124
rect 16683 8084 16725 8093
rect 16683 8044 16684 8084
rect 16724 8044 16725 8084
rect 16683 8035 16725 8044
rect 16684 8000 16724 8035
rect 16684 7169 16724 7960
rect 16780 7841 16820 8212
rect 16875 8084 16917 8093
rect 16875 8044 16876 8084
rect 16916 8044 16917 8084
rect 16875 8035 16917 8044
rect 16876 7950 16916 8035
rect 16779 7832 16821 7841
rect 16779 7792 16780 7832
rect 16820 7792 16821 7832
rect 16972 7832 17012 9211
rect 17068 8681 17108 9388
rect 17164 9017 17204 9472
rect 17260 9472 17452 9512
rect 17163 9008 17205 9017
rect 17163 8968 17164 9008
rect 17204 8968 17205 9008
rect 17163 8959 17205 8968
rect 17067 8672 17109 8681
rect 17067 8632 17068 8672
rect 17108 8632 17109 8672
rect 17067 8623 17109 8632
rect 17164 8672 17204 8681
rect 17260 8672 17300 9472
rect 17452 9463 17492 9472
rect 17451 8672 17493 8681
rect 17204 8632 17396 8672
rect 17164 8623 17204 8632
rect 17259 8420 17301 8429
rect 17259 8380 17260 8420
rect 17300 8380 17301 8420
rect 17259 8371 17301 8380
rect 17068 8009 17108 8094
rect 17163 8084 17205 8093
rect 17163 8044 17164 8084
rect 17204 8044 17205 8084
rect 17163 8035 17205 8044
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17164 8000 17204 8035
rect 17164 7949 17204 7960
rect 17164 7832 17204 7841
rect 16972 7792 17164 7832
rect 16779 7783 16821 7792
rect 17164 7783 17204 7792
rect 17260 7664 17300 8371
rect 17356 8000 17396 8632
rect 17451 8632 17452 8672
rect 17492 8632 17493 8672
rect 17451 8623 17493 8632
rect 17452 8538 17492 8623
rect 17548 8588 17588 9808
rect 17643 9764 17685 9773
rect 17643 9724 17644 9764
rect 17684 9724 17685 9764
rect 17643 9715 17685 9724
rect 17548 8261 17588 8548
rect 17547 8252 17589 8261
rect 17547 8212 17548 8252
rect 17588 8212 17589 8252
rect 17547 8203 17589 8212
rect 17644 8168 17684 9715
rect 17739 9512 17781 9521
rect 17739 9472 17740 9512
rect 17780 9472 17781 9512
rect 17739 9463 17781 9472
rect 17836 9512 17876 10051
rect 17931 10016 17973 10025
rect 17931 9976 17932 10016
rect 17972 9976 17973 10016
rect 17931 9967 17973 9976
rect 17932 9882 17972 9967
rect 18028 9941 18068 10564
rect 18124 10352 18164 10984
rect 18219 10984 18220 11024
rect 18260 10984 18261 11024
rect 18219 10975 18261 10984
rect 18220 10890 18260 10975
rect 18124 10312 18260 10352
rect 18123 10184 18165 10193
rect 18123 10144 18124 10184
rect 18164 10144 18165 10184
rect 18123 10135 18165 10144
rect 18124 10050 18164 10135
rect 18027 9932 18069 9941
rect 18027 9892 18028 9932
rect 18068 9892 18069 9932
rect 18027 9883 18069 9892
rect 18027 9764 18069 9773
rect 18027 9724 18028 9764
rect 18068 9724 18069 9764
rect 18027 9715 18069 9724
rect 17931 9680 17973 9689
rect 17931 9640 17932 9680
rect 17972 9640 17973 9680
rect 17931 9631 17973 9640
rect 17932 9546 17972 9631
rect 17836 9463 17876 9472
rect 18028 9512 18068 9715
rect 18220 9689 18260 10312
rect 18219 9680 18261 9689
rect 18219 9640 18220 9680
rect 18260 9640 18261 9680
rect 18219 9631 18261 9640
rect 18123 9596 18165 9605
rect 18123 9556 18124 9596
rect 18164 9556 18165 9596
rect 18123 9547 18165 9556
rect 18028 9463 18068 9472
rect 18124 9512 18164 9547
rect 17740 9378 17780 9463
rect 17931 9428 17973 9437
rect 17931 9388 17932 9428
rect 17972 9388 17973 9428
rect 17931 9379 17973 9388
rect 17836 8924 17876 8933
rect 17932 8924 17972 9379
rect 17876 8884 17972 8924
rect 17836 8875 17876 8884
rect 18124 8840 18164 9472
rect 18225 9512 18265 9523
rect 18225 9437 18265 9472
rect 18224 9428 18266 9437
rect 18224 9388 18225 9428
rect 18265 9388 18266 9428
rect 18224 9379 18266 9388
rect 18219 9260 18261 9269
rect 18219 9220 18220 9260
rect 18260 9220 18261 9260
rect 18219 9211 18261 9220
rect 17932 8800 18164 8840
rect 17932 8756 17972 8800
rect 17644 8119 17684 8128
rect 17740 8716 17972 8756
rect 18124 8756 18164 8800
rect 17548 8000 17588 8009
rect 17396 7960 17548 8000
rect 17356 7951 17396 7960
rect 17355 7832 17397 7841
rect 17355 7792 17356 7832
rect 17396 7792 17397 7832
rect 17355 7783 17397 7792
rect 17164 7624 17300 7664
rect 16683 7160 16725 7169
rect 16683 7120 16684 7160
rect 16724 7120 16725 7160
rect 16683 7111 16725 7120
rect 16587 7076 16629 7085
rect 16587 7036 16588 7076
rect 16628 7036 16629 7076
rect 16587 7027 16629 7036
rect 16395 6824 16437 6833
rect 16395 6784 16396 6824
rect 16436 6784 16437 6824
rect 16395 6775 16437 6784
rect 16299 6740 16341 6749
rect 16299 6700 16300 6740
rect 16340 6700 16341 6740
rect 16299 6691 16341 6700
rect 16491 6740 16533 6749
rect 16491 6700 16492 6740
rect 16532 6700 16533 6740
rect 16491 6691 16533 6700
rect 16300 6488 16340 6691
rect 16300 6439 16340 6448
rect 16396 6488 16436 6497
rect 16492 6487 16532 6691
rect 16436 6448 16532 6487
rect 16396 6447 16532 6448
rect 16588 6616 17012 6656
rect 16588 6488 16628 6616
rect 16396 6439 16436 6447
rect 16588 6439 16628 6448
rect 16684 6488 16724 6497
rect 16300 6320 16342 6329
rect 16300 6280 16301 6320
rect 16341 6280 16342 6320
rect 16300 6271 16342 6280
rect 16587 6320 16629 6329
rect 16587 6280 16588 6320
rect 16628 6280 16629 6320
rect 16587 6271 16629 6280
rect 16300 6236 16340 6271
rect 16300 6187 16340 6196
rect 16204 5860 16340 5900
rect 15531 5851 15573 5860
rect 15532 5766 15572 5851
rect 15724 5657 15764 5742
rect 16204 5741 16244 5772
rect 16203 5732 16245 5741
rect 16203 5692 16204 5732
rect 16244 5692 16245 5732
rect 16203 5683 16245 5692
rect 15723 5648 15765 5657
rect 15723 5608 15724 5648
rect 15764 5608 15765 5648
rect 15723 5599 15765 5608
rect 15916 5648 15956 5657
rect 15435 5564 15477 5573
rect 15435 5524 15436 5564
rect 15476 5524 15477 5564
rect 15435 5515 15477 5524
rect 15436 5144 15476 5515
rect 15532 5480 15572 5489
rect 15819 5480 15861 5489
rect 15572 5440 15764 5480
rect 15532 5431 15572 5440
rect 15628 5144 15668 5153
rect 15436 5104 15628 5144
rect 15628 5095 15668 5104
rect 15436 4976 15476 4985
rect 15340 4936 15436 4976
rect 15724 4976 15764 5440
rect 15819 5440 15820 5480
rect 15860 5440 15861 5480
rect 15819 5431 15861 5440
rect 15820 5346 15860 5431
rect 15916 5321 15956 5608
rect 16011 5648 16053 5657
rect 16011 5608 16012 5648
rect 16052 5608 16053 5648
rect 16011 5599 16053 5608
rect 16204 5648 16244 5683
rect 15915 5312 15957 5321
rect 15915 5272 15916 5312
rect 15956 5272 15957 5312
rect 15915 5263 15957 5272
rect 15916 5144 15956 5153
rect 16012 5144 16052 5599
rect 16204 5573 16244 5608
rect 16203 5564 16245 5573
rect 16203 5524 16204 5564
rect 16244 5524 16245 5564
rect 16203 5515 16245 5524
rect 15956 5104 16052 5144
rect 15916 5095 15956 5104
rect 15820 4976 15860 4985
rect 15724 4936 15820 4976
rect 15340 2969 15380 4936
rect 15436 4927 15476 4936
rect 15820 4927 15860 4936
rect 16107 4976 16149 4985
rect 16107 4936 16108 4976
rect 16148 4936 16149 4976
rect 16107 4927 16149 4936
rect 16204 4976 16244 5515
rect 16300 5069 16340 5860
rect 16492 5648 16532 5657
rect 16492 5153 16532 5608
rect 16588 5648 16628 6271
rect 16684 5657 16724 6448
rect 16828 6487 16868 6496
rect 16972 6488 17012 6616
rect 17164 6581 17204 7624
rect 17260 7160 17300 7169
rect 17356 7160 17396 7783
rect 17452 7412 17492 7960
rect 17548 7951 17588 7960
rect 17740 8000 17780 8716
rect 18124 8707 18164 8716
rect 18028 8672 18068 8681
rect 17835 8504 17877 8513
rect 17835 8464 17836 8504
rect 17876 8464 17877 8504
rect 17835 8455 17877 8464
rect 17740 7951 17780 7960
rect 17547 7832 17589 7841
rect 17547 7792 17548 7832
rect 17588 7792 17589 7832
rect 17547 7783 17589 7792
rect 17452 7363 17492 7372
rect 17300 7120 17396 7160
rect 17260 7111 17300 7120
rect 17259 6992 17301 7001
rect 17259 6952 17260 6992
rect 17300 6952 17301 6992
rect 17259 6943 17301 6952
rect 17260 6614 17300 6943
rect 17163 6572 17205 6581
rect 17163 6532 17164 6572
rect 17204 6532 17205 6572
rect 17356 6581 17396 7120
rect 17260 6565 17300 6574
rect 17355 6572 17397 6581
rect 17163 6523 17205 6532
rect 17355 6532 17356 6572
rect 17396 6532 17397 6572
rect 17355 6523 17397 6532
rect 17068 6488 17108 6497
rect 16868 6447 16876 6487
rect 16972 6448 17068 6488
rect 16828 6438 16876 6447
rect 16836 6152 16876 6438
rect 17068 6152 17108 6448
rect 17451 6488 17493 6497
rect 17548 6488 17588 7783
rect 17739 7496 17781 7505
rect 17739 7456 17740 7496
rect 17780 7456 17781 7496
rect 17739 7447 17781 7456
rect 17643 6572 17685 6581
rect 17643 6532 17644 6572
rect 17684 6532 17685 6572
rect 17643 6523 17685 6532
rect 17451 6448 17452 6488
rect 17492 6448 17588 6488
rect 17451 6439 17493 6448
rect 17164 6404 17204 6413
rect 17164 6236 17204 6364
rect 17356 6404 17396 6413
rect 17164 6196 17300 6236
rect 16836 6112 16916 6152
rect 17068 6112 17204 6152
rect 16876 5900 16916 6112
rect 16876 5851 16916 5860
rect 17067 5732 17109 5741
rect 17067 5692 17068 5732
rect 17108 5692 17109 5732
rect 17067 5683 17109 5692
rect 17164 5732 17204 6112
rect 17164 5683 17204 5692
rect 16588 5396 16628 5608
rect 16683 5648 16725 5657
rect 16683 5608 16684 5648
rect 16724 5608 16725 5648
rect 16683 5599 16725 5608
rect 17068 5648 17108 5683
rect 17260 5657 17300 6196
rect 17068 5597 17108 5608
rect 17259 5648 17301 5657
rect 17259 5608 17260 5648
rect 17300 5608 17301 5648
rect 17259 5599 17301 5608
rect 17356 5480 17396 6364
rect 17452 6354 17492 6439
rect 17644 6404 17684 6523
rect 17740 6488 17780 7447
rect 17836 7160 17876 8455
rect 18028 8093 18068 8632
rect 18123 8588 18165 8597
rect 18123 8548 18124 8588
rect 18164 8548 18165 8588
rect 18123 8539 18165 8548
rect 18027 8084 18069 8093
rect 18027 8044 18028 8084
rect 18068 8044 18069 8084
rect 18027 8035 18069 8044
rect 18028 7916 18068 7925
rect 18028 7589 18068 7876
rect 18027 7580 18069 7589
rect 18027 7540 18028 7580
rect 18068 7540 18069 7580
rect 18027 7531 18069 7540
rect 17836 7111 17876 7120
rect 17740 6439 17780 6448
rect 17548 6364 17684 6404
rect 17451 6236 17493 6245
rect 17451 6196 17452 6236
rect 17492 6196 17493 6236
rect 17451 6187 17493 6196
rect 17452 5648 17492 6187
rect 17452 5599 17492 5608
rect 16876 5440 17396 5480
rect 16588 5356 16724 5396
rect 16587 5228 16629 5237
rect 16587 5188 16588 5228
rect 16628 5188 16629 5228
rect 16587 5179 16629 5188
rect 16491 5144 16533 5153
rect 16491 5104 16492 5144
rect 16532 5104 16533 5144
rect 16491 5095 16533 5104
rect 16299 5060 16341 5069
rect 16299 5020 16300 5060
rect 16340 5020 16341 5060
rect 16299 5011 16341 5020
rect 16588 5060 16628 5179
rect 16204 4927 16244 4936
rect 16491 4976 16533 4985
rect 16491 4936 16492 4976
rect 16532 4936 16533 4976
rect 16491 4927 16533 4936
rect 15915 4472 15957 4481
rect 15915 4432 15916 4472
rect 15956 4432 15957 4472
rect 15915 4423 15957 4432
rect 15819 4304 15861 4313
rect 15819 4264 15820 4304
rect 15860 4264 15861 4304
rect 15819 4255 15861 4264
rect 15532 4136 15572 4145
rect 15532 3641 15572 4096
rect 15723 4136 15765 4145
rect 15723 4096 15724 4136
rect 15764 4096 15765 4136
rect 15723 4087 15765 4096
rect 15724 4052 15764 4087
rect 15724 4001 15764 4012
rect 15627 3968 15669 3977
rect 15627 3928 15628 3968
rect 15668 3928 15669 3968
rect 15627 3919 15669 3928
rect 15531 3632 15573 3641
rect 15531 3592 15532 3632
rect 15572 3592 15573 3632
rect 15531 3583 15573 3592
rect 15628 3557 15668 3919
rect 15820 3884 15860 4255
rect 15724 3844 15860 3884
rect 15627 3548 15669 3557
rect 15627 3508 15628 3548
rect 15668 3508 15669 3548
rect 15627 3499 15669 3508
rect 15436 3464 15476 3473
rect 15436 3305 15476 3424
rect 15724 3464 15764 3844
rect 15819 3548 15861 3557
rect 15819 3508 15820 3548
rect 15860 3508 15861 3548
rect 15819 3499 15861 3508
rect 15724 3415 15764 3424
rect 15820 3414 15860 3499
rect 15435 3296 15477 3305
rect 15916 3296 15956 4423
rect 16011 4136 16053 4145
rect 16011 4096 16012 4136
rect 16052 4096 16053 4136
rect 16011 4087 16053 4096
rect 16108 4136 16148 4927
rect 16492 4842 16532 4927
rect 16588 4220 16628 5020
rect 16588 4171 16628 4180
rect 16108 4087 16148 4096
rect 16492 4136 16532 4145
rect 16012 4002 16052 4087
rect 16492 4052 16532 4096
rect 16684 4052 16724 5356
rect 16876 4808 16916 5440
rect 17356 5144 17396 5153
rect 17068 4976 17108 4985
rect 16876 4759 16916 4768
rect 16972 4936 17068 4976
rect 16779 4136 16821 4145
rect 16972 4136 17012 4936
rect 17068 4927 17108 4936
rect 17164 4976 17204 4985
rect 17204 4936 17300 4976
rect 17164 4927 17204 4936
rect 17163 4724 17205 4733
rect 17163 4684 17164 4724
rect 17204 4684 17205 4724
rect 17163 4675 17205 4684
rect 17067 4304 17109 4313
rect 17067 4264 17068 4304
rect 17108 4264 17109 4304
rect 17067 4255 17109 4264
rect 16779 4096 16780 4136
rect 16820 4096 17012 4136
rect 17068 4136 17108 4255
rect 16779 4087 16821 4096
rect 17068 4087 17108 4096
rect 16492 4012 16724 4052
rect 16491 3800 16533 3809
rect 16491 3760 16492 3800
rect 16532 3760 16533 3800
rect 16491 3751 16533 3760
rect 16395 3716 16437 3725
rect 16395 3676 16396 3716
rect 16436 3676 16437 3716
rect 16395 3667 16437 3676
rect 16203 3632 16245 3641
rect 16203 3592 16204 3632
rect 16244 3592 16245 3632
rect 16203 3583 16245 3592
rect 15435 3256 15436 3296
rect 15476 3256 15477 3296
rect 15435 3247 15477 3256
rect 15820 3256 15956 3296
rect 15723 3212 15765 3221
rect 15723 3172 15724 3212
rect 15764 3172 15765 3212
rect 15723 3163 15765 3172
rect 15339 2960 15381 2969
rect 15339 2920 15340 2960
rect 15380 2920 15381 2960
rect 15339 2911 15381 2920
rect 15532 2624 15572 2633
rect 15244 2584 15532 2624
rect 15532 2575 15572 2584
rect 15724 2624 15764 3163
rect 15724 2575 15764 2584
rect 15243 2288 15285 2297
rect 15820 2288 15860 3256
rect 16108 3212 16148 3221
rect 15915 2960 15957 2969
rect 15915 2920 15916 2960
rect 15956 2920 15957 2960
rect 15915 2911 15957 2920
rect 15148 2248 15244 2288
rect 15284 2248 15285 2288
rect 15243 2239 15285 2248
rect 15340 2248 15860 2288
rect 15244 1952 15284 2239
rect 15244 1903 15284 1912
rect 15340 1952 15380 2248
rect 15916 2120 15956 2911
rect 16011 2624 16053 2633
rect 16011 2584 16012 2624
rect 16052 2584 16053 2624
rect 16011 2575 16053 2584
rect 15820 2080 15956 2120
rect 15531 2036 15573 2045
rect 15531 1996 15532 2036
rect 15572 1996 15573 2036
rect 15531 1987 15573 1996
rect 15340 1903 15380 1912
rect 15436 1952 15476 1961
rect 15436 1793 15476 1912
rect 15532 1902 15572 1987
rect 15435 1784 15477 1793
rect 15435 1744 15436 1784
rect 15476 1744 15477 1784
rect 15435 1735 15477 1744
rect 15051 1700 15093 1709
rect 15051 1660 15052 1700
rect 15092 1660 15093 1700
rect 15051 1651 15093 1660
rect 15052 1566 15092 1651
rect 15435 1448 15477 1457
rect 15435 1408 15436 1448
rect 15476 1408 15477 1448
rect 15435 1399 15477 1408
rect 14955 1112 14997 1121
rect 14955 1072 14956 1112
rect 14996 1072 14997 1112
rect 14955 1063 14997 1072
rect 15243 860 15285 869
rect 15243 820 15244 860
rect 15284 820 15285 860
rect 15243 811 15285 820
rect 14859 524 14901 533
rect 14859 484 14860 524
rect 14900 484 14901 524
rect 14859 475 14901 484
rect 14860 80 14900 475
rect 15051 440 15093 449
rect 15051 400 15052 440
rect 15092 400 15093 440
rect 15051 391 15093 400
rect 15052 80 15092 391
rect 15244 80 15284 811
rect 15436 80 15476 1399
rect 15627 1112 15669 1121
rect 15627 1072 15628 1112
rect 15668 1072 15669 1112
rect 15820 1112 15860 2080
rect 15915 1952 15957 1961
rect 15915 1912 15916 1952
rect 15956 1912 15957 1952
rect 15915 1903 15957 1912
rect 15916 1818 15956 1903
rect 16012 1112 16052 2575
rect 16108 2549 16148 3172
rect 16107 2540 16149 2549
rect 16107 2500 16108 2540
rect 16148 2500 16149 2540
rect 16107 2491 16149 2500
rect 16204 1793 16244 3583
rect 16300 3296 16340 3305
rect 16300 2885 16340 3256
rect 16299 2876 16341 2885
rect 16299 2836 16300 2876
rect 16340 2836 16341 2876
rect 16299 2827 16341 2836
rect 16299 2540 16341 2549
rect 16299 2500 16300 2540
rect 16340 2500 16341 2540
rect 16396 2540 16436 3667
rect 16492 3305 16532 3751
rect 16587 3632 16629 3641
rect 16587 3592 16588 3632
rect 16628 3592 16629 3632
rect 16587 3583 16629 3592
rect 16491 3296 16533 3305
rect 16491 3256 16492 3296
rect 16532 3256 16533 3296
rect 16491 3247 16533 3256
rect 16396 2500 16532 2540
rect 16299 2491 16341 2500
rect 16203 1784 16245 1793
rect 16203 1744 16204 1784
rect 16244 1744 16245 1784
rect 16203 1735 16245 1744
rect 15820 1072 15956 1112
rect 15627 1063 15669 1072
rect 15628 978 15668 1063
rect 15820 944 15860 953
rect 15820 785 15860 904
rect 15819 776 15861 785
rect 15819 736 15820 776
rect 15860 736 15861 776
rect 15819 727 15861 736
rect 15819 440 15861 449
rect 15819 400 15820 440
rect 15860 400 15861 440
rect 15819 391 15861 400
rect 15627 272 15669 281
rect 15627 232 15628 272
rect 15668 232 15669 272
rect 15627 223 15669 232
rect 15628 80 15668 223
rect 15820 80 15860 391
rect 15916 356 15956 1072
rect 16052 1072 16148 1112
rect 16012 1063 16052 1072
rect 16108 449 16148 1072
rect 16107 440 16149 449
rect 16107 400 16108 440
rect 16148 400 16149 440
rect 16107 391 16149 400
rect 15916 316 16052 356
rect 16012 80 16052 316
rect 16204 80 16244 1735
rect 16300 1121 16340 2491
rect 16395 1448 16437 1457
rect 16395 1408 16396 1448
rect 16436 1408 16437 1448
rect 16395 1399 16437 1408
rect 16299 1112 16341 1121
rect 16299 1072 16300 1112
rect 16340 1072 16341 1112
rect 16299 1063 16341 1072
rect 16396 80 16436 1399
rect 16492 1205 16532 2500
rect 16491 1196 16533 1205
rect 16491 1156 16492 1196
rect 16532 1156 16533 1196
rect 16491 1147 16533 1156
rect 16588 80 16628 3583
rect 16683 3548 16725 3557
rect 16683 3508 16684 3548
rect 16724 3508 16725 3548
rect 16683 3499 16725 3508
rect 16684 3464 16724 3499
rect 16684 3413 16724 3424
rect 16780 3464 16820 4087
rect 17067 3800 17109 3809
rect 17067 3760 17068 3800
rect 17108 3760 17109 3800
rect 17067 3751 17109 3760
rect 17068 3632 17108 3751
rect 17068 3583 17108 3592
rect 16971 3548 17013 3557
rect 16971 3508 16972 3548
rect 17012 3508 17013 3548
rect 16971 3499 17013 3508
rect 16780 3415 16820 3424
rect 16876 3464 16916 3473
rect 16876 3296 16916 3424
rect 16972 3380 17012 3499
rect 16972 3340 17108 3380
rect 16780 3256 16916 3296
rect 16780 2717 16820 3256
rect 16875 3128 16917 3137
rect 16875 3088 16876 3128
rect 16916 3088 16917 3128
rect 16875 3079 16917 3088
rect 16779 2708 16821 2717
rect 16779 2668 16780 2708
rect 16820 2668 16821 2708
rect 16779 2659 16821 2668
rect 16876 1784 16916 3079
rect 16972 2624 17012 2633
rect 16972 1952 17012 2584
rect 17068 2204 17108 3340
rect 17164 2876 17204 4675
rect 17260 3641 17300 4936
rect 17356 4145 17396 5104
rect 17451 5060 17493 5069
rect 17451 5020 17452 5060
rect 17492 5020 17493 5060
rect 17451 5011 17493 5020
rect 17355 4136 17397 4145
rect 17355 4096 17356 4136
rect 17396 4096 17397 4136
rect 17355 4087 17397 4096
rect 17452 3968 17492 5011
rect 17548 4565 17588 6364
rect 18124 5228 18164 8539
rect 18220 8093 18260 9211
rect 18316 8177 18356 13000
rect 18412 12368 18452 13495
rect 18508 13460 18548 13469
rect 18604 13460 18644 14680
rect 18700 14680 18796 14720
rect 18700 13889 18740 14680
rect 18796 14671 18836 14680
rect 18796 14552 18836 14561
rect 18796 14048 18836 14512
rect 18892 14048 18932 14057
rect 18796 14008 18892 14048
rect 18892 13999 18932 14008
rect 18988 13964 19028 13975
rect 18988 13889 19028 13924
rect 18699 13880 18741 13889
rect 18699 13840 18700 13880
rect 18740 13840 18741 13880
rect 18699 13831 18741 13840
rect 18987 13880 19029 13889
rect 18987 13840 18988 13880
rect 19028 13840 19029 13880
rect 18987 13831 19029 13840
rect 19084 13880 19124 14755
rect 19179 14720 19221 14729
rect 19276 14720 19316 15268
rect 19564 15224 19604 16183
rect 19756 15737 19796 16190
rect 19755 15728 19797 15737
rect 19755 15688 19756 15728
rect 19796 15688 19797 15728
rect 19755 15679 19797 15688
rect 19659 15644 19701 15653
rect 19659 15604 19660 15644
rect 19700 15604 19701 15644
rect 19659 15595 19701 15604
rect 19660 15560 19700 15595
rect 19660 15509 19700 15520
rect 19756 15560 19796 15569
rect 19756 15401 19796 15520
rect 19755 15392 19797 15401
rect 19755 15352 19756 15392
rect 19796 15352 19797 15392
rect 19755 15343 19797 15352
rect 19659 15308 19701 15317
rect 19659 15268 19660 15308
rect 19700 15268 19701 15308
rect 19659 15259 19701 15268
rect 19179 14680 19180 14720
rect 19220 14680 19316 14720
rect 19372 15184 19604 15224
rect 19179 14671 19221 14680
rect 19180 14586 19220 14671
rect 19372 14393 19412 15184
rect 19467 14720 19509 14729
rect 19467 14680 19468 14720
rect 19508 14680 19509 14720
rect 19467 14671 19509 14680
rect 19468 14586 19508 14671
rect 19563 14636 19605 14645
rect 19563 14596 19564 14636
rect 19604 14596 19605 14636
rect 19563 14587 19605 14596
rect 19564 14502 19604 14587
rect 19371 14384 19413 14393
rect 19660 14384 19700 15259
rect 19755 14972 19797 14981
rect 19755 14932 19756 14972
rect 19796 14932 19797 14972
rect 19755 14923 19797 14932
rect 19852 14972 19892 16948
rect 19948 16938 19988 17023
rect 19947 16820 19989 16829
rect 19947 16780 19948 16820
rect 19988 16780 19989 16820
rect 20127 16820 20167 17043
rect 20235 16988 20277 16997
rect 20235 16948 20236 16988
rect 20276 16948 20277 16988
rect 20235 16939 20277 16948
rect 20236 16854 20276 16939
rect 20127 16780 20180 16820
rect 19947 16771 19989 16780
rect 19948 16484 19988 16771
rect 19948 16435 19988 16444
rect 20140 16274 20180 16780
rect 19948 16232 19988 16241
rect 20140 16225 20180 16234
rect 20236 16232 20276 16241
rect 19948 15905 19988 16192
rect 20236 16073 20276 16192
rect 20235 16064 20277 16073
rect 20235 16024 20236 16064
rect 20276 16024 20277 16064
rect 20235 16015 20277 16024
rect 19947 15896 19989 15905
rect 19947 15856 19948 15896
rect 19988 15856 19989 15896
rect 19947 15847 19989 15856
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20043 15728 20085 15737
rect 20043 15688 20044 15728
rect 20084 15688 20085 15728
rect 20043 15679 20085 15688
rect 19947 15644 19989 15653
rect 19947 15604 19948 15644
rect 19988 15604 19989 15644
rect 19947 15595 19989 15604
rect 19852 14923 19892 14932
rect 19371 14344 19372 14384
rect 19412 14344 19413 14384
rect 19371 14335 19413 14344
rect 19468 14344 19700 14384
rect 19276 14048 19316 14057
rect 19084 13831 19124 13840
rect 19180 13964 19220 13973
rect 19180 13805 19220 13924
rect 19179 13796 19221 13805
rect 19179 13756 19180 13796
rect 19220 13756 19221 13796
rect 19179 13747 19221 13756
rect 18699 13628 18741 13637
rect 18699 13588 18700 13628
rect 18740 13588 18741 13628
rect 18699 13579 18741 13588
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18548 13420 18644 13460
rect 18508 13411 18548 13420
rect 18700 13217 18740 13579
rect 18795 13376 18837 13385
rect 18795 13336 18796 13376
rect 18836 13336 18837 13376
rect 18795 13327 18837 13336
rect 19083 13376 19125 13385
rect 19083 13336 19084 13376
rect 19124 13336 19125 13376
rect 19083 13327 19125 13336
rect 18507 13208 18549 13217
rect 18507 13168 18508 13208
rect 18548 13168 18549 13208
rect 18507 13159 18549 13168
rect 18699 13208 18741 13217
rect 18699 13168 18700 13208
rect 18740 13168 18741 13208
rect 18699 13159 18741 13168
rect 18796 13208 18836 13327
rect 18508 12536 18548 13159
rect 18700 12704 18740 13159
rect 18700 12655 18740 12664
rect 18603 12620 18645 12629
rect 18603 12580 18604 12620
rect 18644 12580 18645 12620
rect 18603 12571 18645 12580
rect 18508 12487 18548 12496
rect 18412 12328 18548 12368
rect 18411 12032 18453 12041
rect 18411 11992 18412 12032
rect 18452 11992 18453 12032
rect 18411 11983 18453 11992
rect 18412 11024 18452 11983
rect 18412 10975 18452 10984
rect 18508 10109 18548 12328
rect 18604 10529 18644 12571
rect 18796 12545 18836 13168
rect 19084 13208 19124 13327
rect 19276 13292 19316 14008
rect 19468 14048 19508 14344
rect 19468 13999 19508 14008
rect 19756 14216 19796 14923
rect 19948 14720 19988 15595
rect 20044 15392 20084 15679
rect 20044 15343 20084 15352
rect 20235 14972 20277 14981
rect 20235 14932 20236 14972
rect 20276 14932 20277 14972
rect 20235 14923 20277 14932
rect 20236 14838 20276 14923
rect 20044 14720 20084 14729
rect 19948 14680 20044 14720
rect 20044 14671 20084 14680
rect 20236 14720 20276 14729
rect 20524 14720 20564 17536
rect 20620 14981 20660 18535
rect 20715 17240 20757 17249
rect 20715 17200 20716 17240
rect 20756 17200 20757 17240
rect 20715 17191 20757 17200
rect 20619 14972 20661 14981
rect 20619 14932 20620 14972
rect 20660 14932 20661 14972
rect 20619 14923 20661 14932
rect 20276 14680 20564 14720
rect 20236 14671 20276 14680
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 20236 14216 20276 14227
rect 19756 14176 19988 14216
rect 19564 13964 19604 13973
rect 19468 13460 19508 13469
rect 19564 13460 19604 13924
rect 19756 13964 19796 14176
rect 19756 13915 19796 13924
rect 19852 14048 19892 14057
rect 19659 13880 19701 13889
rect 19659 13840 19660 13880
rect 19700 13840 19701 13880
rect 19659 13831 19701 13840
rect 19660 13746 19700 13831
rect 19755 13796 19797 13805
rect 19755 13756 19756 13796
rect 19796 13756 19797 13796
rect 19755 13747 19797 13756
rect 19508 13420 19604 13460
rect 19660 13460 19700 13469
rect 19468 13411 19508 13420
rect 19660 13376 19700 13420
rect 19564 13336 19700 13376
rect 19564 13292 19604 13336
rect 19276 13252 19604 13292
rect 19084 13159 19124 13168
rect 19180 13208 19220 13217
rect 19659 13208 19701 13217
rect 19220 13168 19412 13208
rect 19180 13159 19220 13168
rect 19372 13049 19412 13168
rect 19659 13168 19660 13208
rect 19700 13168 19701 13208
rect 19659 13159 19701 13168
rect 19756 13208 19796 13747
rect 19852 13208 19892 14008
rect 19948 13712 19988 14176
rect 20236 14141 20276 14176
rect 20235 14132 20277 14141
rect 20235 14092 20236 14132
rect 20276 14092 20277 14132
rect 20235 14083 20277 14092
rect 20043 13964 20085 13973
rect 20043 13924 20044 13964
rect 20084 13924 20085 13964
rect 20043 13915 20085 13924
rect 20044 13830 20084 13915
rect 19948 13672 20084 13712
rect 19948 13217 19988 13302
rect 19947 13208 19989 13217
rect 19852 13168 19948 13208
rect 19988 13168 19989 13208
rect 19756 13159 19796 13168
rect 19947 13159 19989 13168
rect 20044 13208 20084 13672
rect 20044 13159 20084 13168
rect 20145 13208 20185 13217
rect 19660 13074 19700 13159
rect 19371 13040 19413 13049
rect 20145 13040 20185 13168
rect 19371 13000 19372 13040
rect 19412 13000 19413 13040
rect 19371 12991 19413 13000
rect 19948 13000 20185 13040
rect 18795 12536 18837 12545
rect 18795 12496 18796 12536
rect 18836 12496 18837 12536
rect 18795 12487 18837 12496
rect 19179 12536 19221 12545
rect 19179 12496 19180 12536
rect 19220 12496 19221 12536
rect 19179 12487 19221 12496
rect 19180 12402 19220 12487
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 19372 11957 19412 12991
rect 19755 12956 19797 12965
rect 19755 12916 19756 12956
rect 19796 12916 19797 12956
rect 19755 12907 19797 12916
rect 19563 12872 19605 12881
rect 19563 12832 19564 12872
rect 19604 12832 19605 12872
rect 19563 12823 19605 12832
rect 19468 12536 19508 12547
rect 19468 12461 19508 12496
rect 19564 12536 19604 12823
rect 19467 12452 19509 12461
rect 19467 12412 19468 12452
rect 19508 12412 19509 12452
rect 19467 12403 19509 12412
rect 19564 12041 19604 12496
rect 19563 12032 19605 12041
rect 19563 11992 19564 12032
rect 19604 11992 19605 12032
rect 19563 11983 19605 11992
rect 19371 11948 19413 11957
rect 19371 11908 19372 11948
rect 19412 11908 19413 11948
rect 19371 11899 19413 11908
rect 19756 11780 19796 12907
rect 19948 12788 19988 13000
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 19852 12748 19988 12788
rect 19852 12368 19892 12748
rect 20043 12704 20085 12713
rect 20043 12664 20044 12704
rect 20084 12664 20085 12704
rect 20043 12655 20085 12664
rect 19947 12620 19989 12629
rect 19947 12580 19948 12620
rect 19988 12580 19989 12620
rect 19947 12571 19989 12580
rect 19852 12319 19892 12328
rect 19948 11948 19988 12571
rect 20044 12452 20084 12655
rect 20716 12461 20756 17191
rect 20812 14141 20852 19879
rect 21292 19265 21332 29119
rect 21388 29009 21428 30127
rect 21387 29000 21429 29009
rect 21387 28960 21388 29000
rect 21428 28960 21429 29000
rect 21387 28951 21429 28960
rect 21291 19256 21333 19265
rect 21291 19216 21292 19256
rect 21332 19216 21333 19256
rect 21291 19207 21333 19216
rect 20907 18920 20949 18929
rect 20907 18880 20908 18920
rect 20948 18880 20949 18920
rect 20907 18871 20949 18880
rect 20811 14132 20853 14141
rect 20811 14092 20812 14132
rect 20852 14092 20853 14132
rect 20811 14083 20853 14092
rect 20044 12403 20084 12412
rect 20235 12452 20277 12461
rect 20235 12412 20236 12452
rect 20276 12412 20277 12452
rect 20235 12403 20277 12412
rect 20715 12452 20757 12461
rect 20715 12412 20716 12452
rect 20756 12412 20757 12452
rect 20715 12403 20757 12412
rect 20236 12368 20276 12403
rect 20236 12317 20276 12328
rect 20908 12125 20948 18871
rect 21003 17744 21045 17753
rect 21003 17704 21004 17744
rect 21044 17704 21045 17744
rect 21003 17695 21045 17704
rect 20523 12116 20565 12125
rect 20523 12076 20524 12116
rect 20564 12076 20565 12116
rect 20523 12067 20565 12076
rect 20907 12116 20949 12125
rect 20907 12076 20908 12116
rect 20948 12076 20949 12116
rect 20907 12067 20949 12076
rect 20044 11948 20084 11957
rect 19948 11908 20044 11948
rect 20044 11899 20084 11908
rect 19852 11780 19892 11789
rect 19756 11740 19852 11780
rect 19852 11731 19892 11740
rect 19468 11696 19508 11705
rect 19468 11360 19508 11656
rect 19372 11320 19508 11360
rect 19660 11528 19700 11537
rect 19660 11360 19700 11488
rect 20048 11360 20416 11369
rect 19660 11320 19796 11360
rect 19275 11024 19317 11033
rect 19275 10984 19276 11024
rect 19316 10984 19317 11024
rect 19275 10975 19317 10984
rect 19372 11024 19412 11320
rect 19660 11024 19700 11033
rect 19372 10984 19660 11024
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18603 10520 18645 10529
rect 18603 10480 18604 10520
rect 18644 10480 18645 10520
rect 18603 10471 18645 10480
rect 18699 10268 18741 10277
rect 18699 10228 18700 10268
rect 18740 10228 18741 10268
rect 18699 10219 18741 10228
rect 18507 10100 18549 10109
rect 18507 10060 18508 10100
rect 18548 10060 18549 10100
rect 18507 10051 18549 10060
rect 18603 10016 18645 10025
rect 18603 9976 18604 10016
rect 18644 9976 18645 10016
rect 18603 9967 18645 9976
rect 18507 9176 18549 9185
rect 18507 9136 18508 9176
rect 18548 9136 18549 9176
rect 18507 9127 18549 9136
rect 18508 8849 18548 9127
rect 18507 8840 18549 8849
rect 18507 8800 18508 8840
rect 18548 8800 18549 8840
rect 18507 8791 18549 8800
rect 18409 8765 18449 8783
rect 18408 8756 18450 8765
rect 18408 8716 18409 8756
rect 18449 8716 18452 8756
rect 18408 8707 18452 8716
rect 18412 8691 18452 8707
rect 18412 8642 18452 8651
rect 18508 8691 18548 8700
rect 18411 8588 18453 8597
rect 18411 8548 18412 8588
rect 18452 8548 18453 8588
rect 18411 8539 18453 8548
rect 18315 8168 18357 8177
rect 18315 8128 18316 8168
rect 18356 8128 18357 8168
rect 18315 8119 18357 8128
rect 18412 8168 18452 8539
rect 18508 8429 18548 8651
rect 18604 8513 18644 9967
rect 18700 8597 18740 10219
rect 18796 9512 18836 9523
rect 18796 9437 18836 9472
rect 19084 9512 19124 9521
rect 18795 9428 18837 9437
rect 18795 9388 18796 9428
rect 18836 9388 18837 9428
rect 18795 9379 18837 9388
rect 19084 9269 19124 9472
rect 19179 9512 19221 9521
rect 19179 9472 19180 9512
rect 19220 9472 19221 9512
rect 19179 9463 19221 9472
rect 19180 9378 19220 9463
rect 19276 9353 19316 10975
rect 19372 10445 19412 10984
rect 19660 10975 19700 10984
rect 19467 10688 19509 10697
rect 19467 10648 19468 10688
rect 19508 10648 19509 10688
rect 19467 10639 19509 10648
rect 19371 10436 19413 10445
rect 19371 10396 19372 10436
rect 19412 10396 19413 10436
rect 19371 10387 19413 10396
rect 19372 10184 19412 10387
rect 19372 10135 19412 10144
rect 19468 9605 19508 10639
rect 19756 10520 19796 11320
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 19947 11276 19989 11285
rect 19947 11236 19948 11276
rect 19988 11236 19989 11276
rect 19947 11227 19989 11236
rect 19948 10940 19988 11227
rect 20236 11192 20276 11201
rect 20524 11192 20564 12067
rect 20619 12032 20661 12041
rect 20619 11992 20620 12032
rect 20660 11992 20661 12032
rect 20619 11983 20661 11992
rect 20276 11152 20564 11192
rect 20236 11143 20276 11152
rect 20044 10940 20084 10949
rect 19948 10900 20044 10940
rect 20044 10891 20084 10900
rect 19852 10772 19892 10783
rect 19852 10697 19892 10732
rect 19851 10688 19893 10697
rect 19851 10648 19852 10688
rect 19892 10648 19893 10688
rect 19851 10639 19893 10648
rect 19756 10480 19988 10520
rect 19852 10277 19892 10321
rect 19851 10268 19893 10277
rect 19851 10228 19852 10268
rect 19892 10228 19893 10268
rect 19851 10226 19893 10228
rect 19851 10219 19852 10226
rect 19756 10184 19796 10193
rect 19892 10219 19893 10226
rect 19852 10177 19892 10186
rect 19948 10184 19988 10480
rect 19564 10016 19604 10025
rect 19756 10016 19796 10144
rect 19948 10100 19988 10144
rect 19604 9976 19796 10016
rect 19564 9967 19604 9976
rect 19467 9596 19509 9605
rect 19467 9556 19468 9596
rect 19508 9556 19509 9596
rect 19467 9547 19509 9556
rect 19660 9512 19700 9521
rect 19275 9344 19317 9353
rect 19275 9304 19276 9344
rect 19316 9304 19317 9344
rect 19275 9295 19317 9304
rect 19468 9344 19508 9353
rect 19660 9344 19700 9472
rect 19508 9304 19700 9344
rect 19756 9512 19796 9976
rect 19468 9295 19508 9304
rect 19083 9260 19125 9269
rect 19083 9220 19084 9260
rect 19124 9220 19125 9260
rect 19083 9211 19125 9220
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18795 8840 18837 8849
rect 18795 8800 18796 8840
rect 18836 8800 18837 8840
rect 18795 8791 18837 8800
rect 18699 8588 18741 8597
rect 18699 8548 18700 8588
rect 18740 8548 18741 8588
rect 18699 8539 18741 8548
rect 18603 8504 18645 8513
rect 18603 8464 18604 8504
rect 18644 8464 18645 8504
rect 18603 8455 18645 8464
rect 18507 8420 18549 8429
rect 18507 8380 18508 8420
rect 18548 8380 18549 8420
rect 18507 8371 18549 8380
rect 18412 8119 18452 8128
rect 18219 8084 18261 8093
rect 18796 8084 18836 8791
rect 19756 8681 19796 9472
rect 19852 10060 19988 10100
rect 18892 8672 18932 8681
rect 18892 8177 18932 8632
rect 18988 8672 19028 8681
rect 18988 8345 19028 8632
rect 19468 8672 19508 8681
rect 18987 8336 19029 8345
rect 18987 8296 18988 8336
rect 19028 8296 19029 8336
rect 18987 8287 19029 8296
rect 18891 8168 18933 8177
rect 18891 8128 18892 8168
rect 18932 8128 18933 8168
rect 18891 8119 18933 8128
rect 18219 8044 18220 8084
rect 18260 8044 18261 8084
rect 18219 8035 18261 8044
rect 18700 8044 18836 8084
rect 18508 8000 18548 8009
rect 18220 7748 18260 7759
rect 18220 7673 18260 7708
rect 18508 7673 18548 7960
rect 18604 8000 18644 8011
rect 18604 7925 18644 7960
rect 18700 8000 18740 8044
rect 18892 8000 18932 8009
rect 18700 7951 18740 7960
rect 18796 7960 18892 8000
rect 18603 7916 18645 7925
rect 18603 7876 18604 7916
rect 18644 7876 18645 7916
rect 18603 7867 18645 7876
rect 18796 7748 18836 7960
rect 18892 7951 18932 7960
rect 19083 8000 19125 8009
rect 19083 7960 19084 8000
rect 19124 7960 19125 8000
rect 19083 7951 19125 7960
rect 19276 8000 19316 8009
rect 19468 8000 19508 8632
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 19852 8588 19892 10060
rect 20044 10016 20084 10025
rect 19948 9976 20044 10016
rect 19948 9512 19988 9976
rect 20044 9967 20084 9976
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 20523 9680 20565 9689
rect 20523 9640 20524 9680
rect 20564 9640 20565 9680
rect 20523 9631 20565 9640
rect 20126 9596 20168 9605
rect 20126 9556 20127 9596
rect 20167 9556 20168 9596
rect 20126 9547 20168 9556
rect 19948 9463 19988 9472
rect 20127 9523 20167 9547
rect 19947 9344 19989 9353
rect 19947 9304 19948 9344
rect 19988 9304 19989 9344
rect 19947 9295 19989 9304
rect 19948 9210 19988 9295
rect 20127 9176 20167 9483
rect 20235 9428 20277 9437
rect 20235 9388 20236 9428
rect 20276 9388 20277 9428
rect 20235 9379 20277 9388
rect 20236 9294 20276 9379
rect 20044 9136 20167 9176
rect 20044 8840 20084 9136
rect 19948 8800 20084 8840
rect 19948 8686 19988 8800
rect 19948 8637 19988 8646
rect 19852 8548 19988 8588
rect 19316 7960 19412 8000
rect 19276 7951 19316 7960
rect 18988 7916 19028 7927
rect 18988 7841 19028 7876
rect 18987 7832 19029 7841
rect 18987 7792 18988 7832
rect 19028 7792 19029 7832
rect 18987 7783 19029 7792
rect 19084 7832 19124 7951
rect 19084 7783 19124 7792
rect 19180 7916 19220 7925
rect 18604 7708 18836 7748
rect 19180 7748 19220 7876
rect 19180 7708 19316 7748
rect 18219 7664 18261 7673
rect 18219 7624 18220 7664
rect 18260 7624 18261 7664
rect 18219 7615 18261 7624
rect 18507 7664 18549 7673
rect 18507 7624 18508 7664
rect 18548 7624 18549 7664
rect 18507 7615 18549 7624
rect 18507 7160 18549 7169
rect 18507 7120 18508 7160
rect 18548 7120 18549 7160
rect 18507 7111 18549 7120
rect 18508 5657 18548 7111
rect 18507 5648 18549 5657
rect 18507 5608 18508 5648
rect 18548 5608 18549 5648
rect 18507 5599 18549 5608
rect 18124 5188 18260 5228
rect 17740 5144 17780 5153
rect 17780 5104 18164 5144
rect 17740 5095 17780 5104
rect 17836 4976 17876 4985
rect 17547 4556 17589 4565
rect 17547 4516 17548 4556
rect 17588 4516 17589 4556
rect 17547 4507 17589 4516
rect 17643 4304 17685 4313
rect 17643 4264 17644 4304
rect 17684 4264 17685 4304
rect 17643 4255 17685 4264
rect 17356 3928 17492 3968
rect 17548 4141 17588 4150
rect 17259 3632 17301 3641
rect 17259 3592 17260 3632
rect 17300 3592 17301 3632
rect 17259 3583 17301 3592
rect 17260 3464 17300 3473
rect 17260 3305 17300 3424
rect 17356 3464 17396 3928
rect 17548 3641 17588 4101
rect 17644 4061 17684 4255
rect 17643 4052 17685 4061
rect 17643 4012 17644 4052
rect 17684 4012 17685 4052
rect 17643 4003 17685 4012
rect 17740 3968 17780 3977
rect 17740 3641 17780 3928
rect 17836 3809 17876 4936
rect 18028 4724 18068 4733
rect 17931 4136 17973 4145
rect 17931 4096 17932 4136
rect 17972 4096 17973 4136
rect 17931 4087 17973 4096
rect 18028 4136 18068 4684
rect 18028 4087 18068 4096
rect 17932 4002 17972 4087
rect 17835 3800 17877 3809
rect 17835 3760 17836 3800
rect 17876 3760 17877 3800
rect 17835 3751 17877 3760
rect 17547 3632 17589 3641
rect 17547 3592 17548 3632
rect 17588 3592 17589 3632
rect 17547 3583 17589 3592
rect 17739 3632 17781 3641
rect 17739 3592 17740 3632
rect 17780 3592 17781 3632
rect 17739 3583 17781 3592
rect 17548 3464 17588 3473
rect 17740 3464 17780 3473
rect 17356 3415 17396 3424
rect 17452 3424 17548 3464
rect 17259 3296 17301 3305
rect 17259 3256 17260 3296
rect 17300 3256 17301 3296
rect 17259 3247 17301 3256
rect 17356 2876 17396 2885
rect 17164 2836 17356 2876
rect 17356 2827 17396 2836
rect 17164 2549 17204 2634
rect 17163 2540 17205 2549
rect 17163 2500 17164 2540
rect 17204 2500 17205 2540
rect 17163 2491 17205 2500
rect 17068 2164 17396 2204
rect 17356 2120 17396 2164
rect 17356 2071 17396 2080
rect 17164 1952 17204 1961
rect 16972 1912 17164 1952
rect 17164 1793 17204 1912
rect 17452 1877 17492 3424
rect 17548 3415 17588 3424
rect 17644 3424 17740 3464
rect 17548 3212 17588 3221
rect 17548 3053 17588 3172
rect 17547 3044 17589 3053
rect 17547 3004 17548 3044
rect 17588 3004 17589 3044
rect 17547 2995 17589 3004
rect 17548 2801 17588 2886
rect 17547 2792 17589 2801
rect 17547 2752 17548 2792
rect 17588 2752 17589 2792
rect 17547 2743 17589 2752
rect 17548 2624 17588 2635
rect 17548 2549 17588 2584
rect 17547 2540 17589 2549
rect 17547 2500 17548 2540
rect 17588 2500 17589 2540
rect 17644 2540 17684 3424
rect 17740 3415 17780 3424
rect 17932 3464 17972 3473
rect 17739 3296 17781 3305
rect 17739 3256 17740 3296
rect 17780 3256 17781 3296
rect 17739 3247 17781 3256
rect 17740 3162 17780 3247
rect 17932 2801 17972 3424
rect 18028 3464 18068 3475
rect 18028 3389 18068 3424
rect 18027 3380 18069 3389
rect 18027 3340 18028 3380
rect 18068 3340 18069 3380
rect 18027 3331 18069 3340
rect 18028 2969 18068 3331
rect 18124 3221 18164 5104
rect 18220 4565 18260 5188
rect 18508 4985 18548 5070
rect 18315 4976 18357 4985
rect 18315 4936 18316 4976
rect 18356 4936 18357 4976
rect 18315 4927 18357 4936
rect 18412 4976 18452 4985
rect 18219 4556 18261 4565
rect 18219 4516 18220 4556
rect 18260 4516 18261 4556
rect 18219 4507 18261 4516
rect 18219 4388 18261 4397
rect 18219 4348 18220 4388
rect 18260 4348 18261 4388
rect 18219 4339 18261 4348
rect 18220 4254 18260 4339
rect 18220 4136 18260 4145
rect 18220 3809 18260 4096
rect 18219 3800 18261 3809
rect 18219 3760 18220 3800
rect 18260 3760 18261 3800
rect 18219 3751 18261 3760
rect 18219 3464 18261 3473
rect 18219 3424 18220 3464
rect 18260 3424 18261 3464
rect 18219 3415 18261 3424
rect 18220 3330 18260 3415
rect 18123 3212 18165 3221
rect 18123 3172 18124 3212
rect 18164 3172 18165 3212
rect 18123 3163 18165 3172
rect 18220 3212 18260 3221
rect 18027 2960 18069 2969
rect 18027 2920 18028 2960
rect 18068 2920 18069 2960
rect 18027 2911 18069 2920
rect 17931 2792 17973 2801
rect 17931 2752 17932 2792
rect 17972 2752 17973 2792
rect 17931 2743 17973 2752
rect 18028 2633 18068 2718
rect 18027 2624 18069 2633
rect 18027 2584 18028 2624
rect 18068 2584 18069 2624
rect 18027 2575 18069 2584
rect 18124 2549 18164 3163
rect 18123 2540 18165 2549
rect 17644 2500 17780 2540
rect 17547 2491 17589 2500
rect 17740 2045 17780 2500
rect 18123 2500 18124 2540
rect 18164 2500 18165 2540
rect 18123 2491 18165 2500
rect 18220 2213 18260 3172
rect 18316 2540 18356 4927
rect 18412 4817 18452 4936
rect 18507 4976 18549 4985
rect 18507 4936 18508 4976
rect 18548 4936 18549 4976
rect 18507 4927 18549 4936
rect 18411 4808 18453 4817
rect 18411 4768 18412 4808
rect 18452 4768 18453 4808
rect 18411 4759 18453 4768
rect 18508 4808 18548 4817
rect 18604 4808 18644 7708
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 19276 7412 19316 7708
rect 19372 7589 19412 7960
rect 19468 7757 19508 7960
rect 19852 8000 19892 8009
rect 19948 8000 19988 8548
rect 20140 8513 20180 8598
rect 20139 8504 20181 8513
rect 20139 8464 20140 8504
rect 20180 8464 20181 8504
rect 20139 8455 20181 8464
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 20043 8168 20085 8177
rect 20043 8128 20044 8168
rect 20084 8128 20276 8168
rect 20043 8119 20085 8128
rect 20044 8000 20084 8009
rect 19948 7960 20044 8000
rect 19564 7916 19604 7925
rect 19467 7748 19509 7757
rect 19467 7708 19468 7748
rect 19508 7708 19509 7748
rect 19467 7699 19509 7708
rect 19371 7580 19413 7589
rect 19371 7540 19372 7580
rect 19412 7540 19413 7580
rect 19371 7531 19413 7540
rect 19564 7412 19604 7876
rect 19756 7916 19796 7925
rect 19659 7832 19701 7841
rect 19659 7792 19660 7832
rect 19700 7792 19701 7832
rect 19659 7783 19701 7792
rect 19660 7698 19700 7783
rect 19659 7580 19701 7589
rect 19659 7540 19660 7580
rect 19700 7540 19701 7580
rect 19659 7531 19701 7540
rect 19276 7253 19316 7372
rect 19372 7372 19604 7412
rect 19275 7244 19317 7253
rect 19275 7204 19276 7244
rect 19316 7204 19317 7244
rect 19275 7195 19317 7204
rect 18987 7160 19029 7169
rect 19084 7160 19124 7188
rect 18987 7120 18988 7160
rect 19028 7120 19084 7160
rect 18987 7111 19029 7120
rect 19084 7111 19124 7120
rect 18988 6488 19028 7111
rect 18988 6439 19028 6448
rect 19372 6320 19412 7372
rect 19467 7244 19509 7253
rect 19467 7204 19468 7244
rect 19508 7204 19509 7244
rect 19467 7195 19509 7204
rect 19468 7160 19508 7195
rect 19468 7109 19508 7120
rect 19563 7160 19605 7169
rect 19563 7120 19564 7160
rect 19604 7120 19605 7160
rect 19563 7111 19605 7120
rect 19564 7026 19604 7111
rect 19660 6992 19700 7531
rect 19756 7328 19796 7876
rect 19852 7505 19892 7960
rect 20044 7951 20084 7960
rect 20236 8000 20276 8128
rect 20524 8000 20564 9631
rect 20620 8513 20660 11983
rect 20811 11948 20853 11957
rect 20811 11908 20812 11948
rect 20852 11908 20853 11948
rect 20811 11899 20853 11908
rect 20812 11201 20852 11899
rect 20811 11192 20853 11201
rect 20811 11152 20812 11192
rect 20852 11152 20853 11192
rect 20811 11143 20853 11152
rect 20715 11108 20757 11117
rect 20715 11068 20716 11108
rect 20756 11068 20757 11108
rect 20715 11059 20757 11068
rect 20619 8504 20661 8513
rect 20619 8464 20620 8504
rect 20660 8464 20661 8504
rect 20619 8455 20661 8464
rect 20716 8084 20756 11059
rect 21004 10193 21044 17695
rect 21099 14216 21141 14225
rect 21099 14176 21100 14216
rect 21140 14176 21141 14216
rect 21099 14167 21141 14176
rect 21003 10184 21045 10193
rect 21003 10144 21004 10184
rect 21044 10144 21045 10184
rect 21003 10135 21045 10144
rect 21003 9176 21045 9185
rect 21003 9136 21004 9176
rect 21044 9136 21045 9176
rect 21003 9127 21045 9136
rect 20236 7951 20276 7960
rect 20332 7960 20564 8000
rect 20620 8044 20756 8084
rect 20236 7832 20276 7841
rect 20332 7832 20372 7960
rect 20276 7792 20372 7832
rect 20236 7783 20276 7792
rect 19851 7496 19893 7505
rect 19851 7456 19852 7496
rect 19892 7456 19893 7496
rect 19851 7447 19893 7456
rect 19756 7288 19892 7328
rect 19755 7160 19797 7169
rect 19755 7120 19756 7160
rect 19796 7120 19797 7160
rect 19755 7111 19797 7120
rect 19852 7160 19892 7288
rect 19953 7160 19993 7169
rect 19660 6943 19700 6952
rect 19756 6749 19796 7111
rect 19755 6740 19797 6749
rect 19755 6700 19756 6740
rect 19796 6700 19797 6740
rect 19755 6691 19797 6700
rect 19852 6665 19892 7120
rect 19948 7120 19953 7160
rect 19948 7111 19993 7120
rect 19851 6656 19893 6665
rect 19851 6616 19852 6656
rect 19892 6616 19893 6656
rect 19851 6607 19893 6616
rect 19659 6488 19701 6497
rect 19659 6448 19660 6488
rect 19700 6448 19701 6488
rect 19659 6439 19701 6448
rect 19756 6488 19796 6499
rect 19372 6271 19412 6280
rect 19563 6320 19605 6329
rect 19563 6280 19564 6320
rect 19604 6280 19605 6320
rect 19563 6271 19605 6280
rect 19180 6236 19220 6245
rect 19220 6196 19316 6236
rect 19180 6187 19220 6196
rect 18699 6068 18741 6077
rect 18699 6028 18700 6068
rect 18740 6028 18741 6068
rect 18699 6019 18741 6028
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18700 5900 18740 6019
rect 18700 5860 19028 5900
rect 18699 5648 18741 5657
rect 18699 5608 18700 5648
rect 18740 5608 18741 5648
rect 18699 5599 18741 5608
rect 18700 5514 18740 5599
rect 18892 5480 18932 5489
rect 18796 5440 18892 5480
rect 18796 5069 18836 5440
rect 18892 5431 18932 5440
rect 18795 5060 18837 5069
rect 18795 5020 18796 5060
rect 18836 5020 18837 5060
rect 18795 5011 18837 5020
rect 18699 4976 18741 4985
rect 18699 4936 18700 4976
rect 18740 4936 18741 4976
rect 18699 4927 18741 4936
rect 18700 4842 18740 4927
rect 18548 4768 18644 4808
rect 18988 4808 19028 5860
rect 19180 5648 19220 5657
rect 19276 5648 19316 6196
rect 19467 5984 19509 5993
rect 19467 5944 19468 5984
rect 19508 5944 19509 5984
rect 19467 5935 19509 5944
rect 19468 5648 19508 5935
rect 19084 5608 19180 5648
rect 19220 5608 19316 5648
rect 19372 5608 19468 5648
rect 19084 4985 19124 5608
rect 19180 5599 19220 5608
rect 19179 5312 19221 5321
rect 19179 5272 19180 5312
rect 19220 5272 19221 5312
rect 19179 5263 19221 5272
rect 19180 5060 19220 5263
rect 19180 5011 19220 5020
rect 19275 5060 19317 5069
rect 19275 5020 19276 5060
rect 19316 5020 19317 5060
rect 19275 5011 19317 5020
rect 19083 4976 19125 4985
rect 19083 4936 19084 4976
rect 19124 4936 19125 4976
rect 19083 4927 19125 4936
rect 19276 4976 19316 5011
rect 19276 4925 19316 4936
rect 18988 4768 19316 4808
rect 18508 4759 18548 4768
rect 18892 4724 18932 4733
rect 18700 4684 18892 4724
rect 18411 4640 18453 4649
rect 18411 4600 18412 4640
rect 18452 4600 18453 4640
rect 18411 4591 18453 4600
rect 18412 4136 18452 4591
rect 18507 4304 18549 4313
rect 18507 4264 18508 4304
rect 18548 4264 18549 4304
rect 18507 4255 18549 4264
rect 18604 4304 18644 4313
rect 18508 4220 18548 4255
rect 18508 4169 18548 4180
rect 18412 3809 18452 4096
rect 18411 3800 18453 3809
rect 18411 3760 18412 3800
rect 18452 3760 18453 3800
rect 18604 3800 18644 4264
rect 18700 4220 18740 4684
rect 18892 4675 18932 4684
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18795 4388 18837 4397
rect 18795 4348 18796 4388
rect 18836 4348 18837 4388
rect 18795 4339 18837 4348
rect 19083 4388 19125 4397
rect 19083 4348 19084 4388
rect 19124 4348 19125 4388
rect 19083 4339 19125 4348
rect 18700 4171 18740 4180
rect 18796 4136 18836 4339
rect 18796 4087 18836 4096
rect 19084 4136 19124 4339
rect 19084 3893 19124 4096
rect 19276 4061 19316 4768
rect 19372 4136 19412 5608
rect 19468 5599 19508 5608
rect 19564 5648 19604 6271
rect 19564 5480 19604 5608
rect 19275 4052 19317 4061
rect 19275 4012 19276 4052
rect 19316 4012 19317 4052
rect 19275 4003 19317 4012
rect 19372 3977 19412 4096
rect 19468 5440 19604 5480
rect 19468 4136 19508 5440
rect 19660 5321 19700 6439
rect 19756 6413 19796 6448
rect 19755 6404 19797 6413
rect 19755 6364 19756 6404
rect 19796 6364 19797 6404
rect 19755 6355 19797 6364
rect 19659 5312 19701 5321
rect 19659 5272 19660 5312
rect 19700 5272 19701 5312
rect 19659 5263 19701 5272
rect 19756 5069 19796 6355
rect 19852 5900 19892 5909
rect 19948 5900 19988 7111
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20331 6656 20373 6665
rect 20331 6616 20332 6656
rect 20372 6616 20373 6656
rect 20331 6607 20373 6616
rect 20235 6572 20277 6581
rect 20235 6532 20236 6572
rect 20276 6532 20277 6572
rect 20235 6523 20277 6532
rect 19892 5860 19988 5900
rect 20044 6488 20084 6497
rect 19852 5851 19892 5860
rect 20044 5648 20084 6448
rect 20236 5900 20276 6523
rect 20236 5851 20276 5860
rect 19948 5608 20044 5648
rect 19851 5480 19893 5489
rect 19851 5440 19852 5480
rect 19892 5440 19893 5480
rect 19851 5431 19893 5440
rect 19755 5060 19797 5069
rect 19755 5020 19756 5060
rect 19796 5020 19797 5060
rect 19755 5011 19797 5020
rect 19564 4976 19604 4985
rect 19564 4481 19604 4936
rect 19852 4892 19892 5431
rect 19948 4985 19988 5608
rect 20044 5599 20084 5608
rect 20236 5648 20276 5657
rect 20332 5648 20372 6607
rect 20276 5608 20564 5648
rect 20236 5599 20276 5608
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19947 4976 19989 4985
rect 19947 4936 19948 4976
rect 19988 4936 19989 4976
rect 19947 4927 19989 4936
rect 19852 4843 19892 4852
rect 20043 4808 20085 4817
rect 20043 4768 20044 4808
rect 20084 4768 20085 4808
rect 20043 4759 20085 4768
rect 20044 4674 20084 4759
rect 19563 4472 19605 4481
rect 19563 4432 19564 4472
rect 19604 4432 19605 4472
rect 19563 4423 19605 4432
rect 19563 4304 19605 4313
rect 19563 4264 19564 4304
rect 19604 4264 19605 4304
rect 19563 4255 19605 4264
rect 19756 4304 19796 4313
rect 19468 4087 19508 4096
rect 19371 3968 19413 3977
rect 19371 3928 19372 3968
rect 19412 3928 19413 3968
rect 19371 3919 19413 3928
rect 19083 3884 19125 3893
rect 19083 3844 19084 3884
rect 19124 3844 19125 3884
rect 19083 3835 19125 3844
rect 19467 3800 19509 3809
rect 18604 3760 18740 3800
rect 18411 3751 18453 3760
rect 18412 3464 18452 3473
rect 18412 3305 18452 3424
rect 18604 3464 18644 3473
rect 18411 3296 18453 3305
rect 18411 3256 18412 3296
rect 18452 3256 18453 3296
rect 18411 3247 18453 3256
rect 18316 2500 18548 2540
rect 18219 2204 18261 2213
rect 18219 2164 18220 2204
rect 18260 2164 18261 2204
rect 18219 2155 18261 2164
rect 18027 2120 18069 2129
rect 18027 2080 18028 2120
rect 18068 2080 18069 2120
rect 18027 2071 18069 2080
rect 17739 2036 17781 2045
rect 17739 1996 17740 2036
rect 17780 1996 17781 2036
rect 17739 1987 17781 1996
rect 17931 1952 17973 1961
rect 17931 1912 17932 1952
rect 17972 1912 17973 1952
rect 17931 1903 17973 1912
rect 17451 1868 17493 1877
rect 17739 1868 17781 1877
rect 17451 1828 17452 1868
rect 17492 1828 17684 1868
rect 17451 1819 17493 1828
rect 17163 1784 17205 1793
rect 16876 1744 17108 1784
rect 16875 1532 16917 1541
rect 16875 1492 16876 1532
rect 16916 1492 16917 1532
rect 16875 1483 16917 1492
rect 16876 449 16916 1483
rect 16971 1280 17013 1289
rect 16971 1240 16972 1280
rect 17012 1240 17013 1280
rect 16971 1231 17013 1240
rect 16875 440 16917 449
rect 16875 400 16876 440
rect 16916 400 16917 440
rect 16875 391 16917 400
rect 16779 356 16821 365
rect 16779 316 16780 356
rect 16820 316 16821 356
rect 16779 307 16821 316
rect 16780 80 16820 307
rect 16972 80 17012 1231
rect 17068 1112 17108 1744
rect 17163 1744 17164 1784
rect 17204 1744 17205 1784
rect 17163 1735 17205 1744
rect 17451 1700 17493 1709
rect 17451 1660 17452 1700
rect 17492 1660 17493 1700
rect 17451 1651 17493 1660
rect 17548 1700 17588 1709
rect 17355 1196 17397 1205
rect 17355 1156 17356 1196
rect 17396 1156 17397 1196
rect 17355 1147 17397 1156
rect 17260 1112 17300 1121
rect 17068 1072 17260 1112
rect 17260 1063 17300 1072
rect 17163 188 17205 197
rect 17163 148 17164 188
rect 17204 148 17205 188
rect 17163 139 17205 148
rect 17164 80 17204 139
rect 17356 80 17396 1147
rect 17452 1112 17492 1651
rect 17548 1373 17588 1660
rect 17547 1364 17589 1373
rect 17547 1324 17548 1364
rect 17588 1324 17589 1364
rect 17547 1315 17589 1324
rect 17452 1063 17492 1072
rect 17644 1112 17684 1828
rect 17739 1828 17740 1868
rect 17780 1828 17781 1868
rect 17739 1819 17781 1828
rect 17740 1734 17780 1819
rect 17932 1818 17972 1903
rect 17931 1280 17973 1289
rect 17931 1240 17932 1280
rect 17972 1240 17973 1280
rect 17931 1231 17973 1240
rect 17740 1121 17780 1206
rect 17644 1063 17684 1072
rect 17739 1112 17781 1121
rect 17739 1072 17740 1112
rect 17780 1072 17781 1112
rect 17739 1063 17781 1072
rect 17547 1028 17589 1037
rect 17547 988 17548 1028
rect 17588 988 17589 1028
rect 17547 979 17589 988
rect 17548 894 17588 979
rect 17739 944 17781 953
rect 17739 904 17740 944
rect 17780 904 17781 944
rect 17739 895 17781 904
rect 17547 440 17589 449
rect 17547 400 17548 440
rect 17588 400 17589 440
rect 17547 391 17589 400
rect 17548 80 17588 391
rect 17740 80 17780 895
rect 17932 80 17972 1231
rect 18028 1112 18068 2071
rect 18508 1961 18548 2500
rect 18604 2129 18644 3424
rect 18700 3380 18740 3760
rect 19467 3760 19468 3800
rect 19508 3760 19509 3800
rect 19467 3751 19509 3760
rect 18700 3331 18740 3340
rect 18892 3592 19412 3632
rect 18892 3380 18932 3592
rect 18892 3331 18932 3340
rect 18988 3464 19028 3473
rect 18795 3296 18837 3305
rect 18795 3256 18796 3296
rect 18836 3256 18837 3296
rect 18795 3247 18837 3256
rect 18796 3162 18836 3247
rect 18988 3212 19028 3424
rect 19180 3464 19220 3592
rect 19180 3415 19220 3424
rect 19275 3464 19317 3473
rect 19275 3424 19276 3464
rect 19316 3424 19317 3464
rect 19275 3415 19317 3424
rect 19276 3330 19316 3415
rect 19180 3212 19220 3221
rect 18988 3172 19180 3212
rect 19180 3163 19220 3172
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 19372 2876 19412 3592
rect 19468 3464 19508 3751
rect 19468 3415 19508 3424
rect 19564 3464 19604 4255
rect 19756 3800 19796 4264
rect 19948 4145 19988 4230
rect 20121 4220 20163 4229
rect 20121 4180 20122 4220
rect 20162 4180 20163 4220
rect 20121 4171 20163 4180
rect 19947 4136 19989 4145
rect 19947 4096 19948 4136
rect 19988 4096 19989 4136
rect 19947 4087 19989 4096
rect 20122 4141 20162 4171
rect 20122 4085 20162 4101
rect 20044 3968 20084 3977
rect 19716 3760 19796 3800
rect 19852 3928 20044 3968
rect 19716 3473 19756 3760
rect 19564 3415 19604 3424
rect 19708 3464 19756 3473
rect 19748 3424 19756 3464
rect 19708 3415 19748 3424
rect 19563 3296 19605 3305
rect 19563 3256 19564 3296
rect 19604 3256 19605 3296
rect 19563 3247 19605 3256
rect 19755 3296 19797 3305
rect 19755 3256 19756 3296
rect 19796 3256 19797 3296
rect 19755 3247 19797 3256
rect 19468 2876 19508 2885
rect 19372 2836 19468 2876
rect 19468 2827 19508 2836
rect 19276 2624 19316 2633
rect 19276 2381 19316 2584
rect 19275 2372 19317 2381
rect 19275 2332 19276 2372
rect 19316 2332 19317 2372
rect 19275 2323 19317 2332
rect 18603 2120 18645 2129
rect 18603 2080 18604 2120
rect 18644 2080 18645 2120
rect 18603 2071 18645 2080
rect 18507 1952 18549 1961
rect 18507 1912 18508 1952
rect 18548 1912 18549 1952
rect 18507 1903 18549 1912
rect 19180 1952 19220 1961
rect 19276 1952 19316 2323
rect 19371 2288 19413 2297
rect 19371 2248 19372 2288
rect 19412 2248 19413 2288
rect 19371 2239 19413 2248
rect 19372 2120 19412 2239
rect 19372 2071 19412 2080
rect 19220 1912 19316 1952
rect 19180 1903 19220 1912
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 19276 1457 19316 1912
rect 19564 1952 19604 3247
rect 19659 2960 19701 2969
rect 19659 2920 19660 2960
rect 19700 2920 19701 2960
rect 19659 2911 19701 2920
rect 19660 2624 19700 2911
rect 19660 2575 19700 2584
rect 19756 2624 19796 3247
rect 19852 3044 19892 3928
rect 20044 3919 20084 3928
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 19947 3632 19989 3641
rect 19947 3592 19948 3632
rect 19988 3592 19989 3632
rect 19947 3583 19989 3592
rect 19948 3464 19988 3583
rect 20043 3548 20085 3557
rect 20043 3508 20044 3548
rect 20084 3508 20085 3548
rect 20043 3499 20085 3508
rect 19948 3415 19988 3424
rect 20044 3414 20084 3499
rect 20129 3451 20169 3460
rect 20129 3221 20169 3411
rect 20128 3212 20170 3221
rect 20128 3172 20129 3212
rect 20169 3172 20170 3212
rect 20128 3163 20170 3172
rect 19852 3004 19988 3044
rect 19851 2876 19893 2885
rect 19851 2836 19852 2876
rect 19892 2836 19893 2876
rect 19851 2827 19893 2836
rect 19756 2575 19796 2584
rect 19852 2540 19892 2827
rect 19948 2624 19988 3004
rect 19948 2575 19988 2584
rect 20140 2549 20180 2634
rect 19852 2491 19892 2500
rect 20139 2540 20181 2549
rect 20139 2500 20140 2540
rect 20180 2500 20181 2540
rect 20139 2491 20181 2500
rect 19947 2456 19989 2465
rect 19947 2416 19948 2456
rect 19988 2416 19989 2456
rect 19947 2407 19989 2416
rect 19851 2288 19893 2297
rect 19851 2248 19852 2288
rect 19892 2248 19893 2288
rect 19851 2239 19893 2248
rect 19660 2129 19700 2214
rect 19659 2120 19701 2129
rect 19659 2080 19660 2120
rect 19700 2080 19701 2120
rect 19659 2071 19701 2080
rect 19660 1952 19700 1961
rect 19564 1912 19660 1952
rect 19275 1448 19317 1457
rect 19275 1408 19276 1448
rect 19316 1408 19317 1448
rect 19275 1399 19317 1408
rect 18507 1280 18549 1289
rect 18507 1240 18508 1280
rect 18548 1240 18549 1280
rect 18507 1231 18549 1240
rect 18699 1280 18741 1289
rect 18699 1240 18700 1280
rect 18740 1240 18741 1280
rect 18699 1231 18741 1240
rect 18028 1063 18068 1072
rect 18315 692 18357 701
rect 18315 652 18316 692
rect 18356 652 18357 692
rect 18315 643 18357 652
rect 18123 104 18165 113
rect 18123 80 18124 104
rect 10868 64 10888 80
rect 10808 0 10888 64
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 0 17032 80
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 64 18124 80
rect 18164 80 18165 104
rect 18316 80 18356 643
rect 18508 80 18548 1231
rect 18700 80 18740 1231
rect 19276 1112 19316 1399
rect 19468 1364 19508 1373
rect 19564 1364 19604 1912
rect 19660 1903 19700 1912
rect 19852 1952 19892 2239
rect 19852 1903 19892 1912
rect 19948 1952 19988 2407
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 20236 2120 20276 2129
rect 20524 2120 20564 5608
rect 20276 2080 20564 2120
rect 20236 2071 20276 2080
rect 19948 1903 19988 1912
rect 20126 1952 20168 1961
rect 20126 1912 20127 1952
rect 20167 1912 20168 1952
rect 20126 1903 20168 1912
rect 20127 1818 20167 1903
rect 19851 1784 19893 1793
rect 19851 1744 19852 1784
rect 19892 1744 19893 1784
rect 19851 1735 19893 1744
rect 19508 1324 19604 1364
rect 19468 1315 19508 1324
rect 19852 1196 19892 1735
rect 19852 1147 19892 1156
rect 20236 1196 20276 1205
rect 20620 1196 20660 8044
rect 21004 5237 21044 9127
rect 21100 7169 21140 14167
rect 21195 10016 21237 10025
rect 21195 9976 21196 10016
rect 21236 9976 21237 10016
rect 21195 9967 21237 9976
rect 21099 7160 21141 7169
rect 21099 7120 21100 7160
rect 21140 7120 21141 7160
rect 21099 7111 21141 7120
rect 21003 5228 21045 5237
rect 21003 5188 21004 5228
rect 21044 5188 21045 5228
rect 21003 5179 21045 5188
rect 20715 4892 20757 4901
rect 20715 4852 20716 4892
rect 20756 4852 20757 4892
rect 20715 4843 20757 4852
rect 20716 3809 20756 4843
rect 20811 3968 20853 3977
rect 20811 3928 20812 3968
rect 20852 3928 20853 3968
rect 20811 3919 20853 3928
rect 20715 3800 20757 3809
rect 20715 3760 20716 3800
rect 20756 3760 20757 3800
rect 20715 3751 20757 3760
rect 20812 2465 20852 3919
rect 20811 2456 20853 2465
rect 20811 2416 20812 2456
rect 20852 2416 20853 2456
rect 20811 2407 20853 2416
rect 20276 1156 20660 1196
rect 20236 1147 20276 1156
rect 19276 1063 19316 1072
rect 20044 953 20084 1038
rect 19083 944 19125 953
rect 19083 904 19084 944
rect 19124 904 19125 944
rect 19083 895 19125 904
rect 19660 944 19700 953
rect 18891 440 18933 449
rect 18891 400 18892 440
rect 18932 400 18933 440
rect 18891 391 18933 400
rect 18892 80 18932 391
rect 19084 80 19124 895
rect 19467 776 19509 785
rect 19467 736 19468 776
rect 19508 736 19509 776
rect 19467 727 19509 736
rect 19275 608 19317 617
rect 19275 568 19276 608
rect 19316 568 19317 608
rect 19275 559 19317 568
rect 19276 80 19316 559
rect 19468 80 19508 727
rect 19660 533 19700 904
rect 20043 944 20085 953
rect 20043 904 20044 944
rect 20084 904 20085 944
rect 20043 895 20085 904
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 19659 524 19701 533
rect 19659 484 19660 524
rect 19700 484 19701 524
rect 19659 475 19701 484
rect 21196 113 21236 9967
rect 21195 104 21237 113
rect 18164 64 18184 80
rect 18104 0 18184 64
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
rect 21195 64 21196 104
rect 21236 64 21237 104
rect 21195 55 21237 64
<< via2 >>
rect 1228 42904 1268 42944
rect 1132 41560 1172 41600
rect 1036 40300 1076 40340
rect 76 39376 116 39416
rect 76 39040 116 39080
rect 940 37192 980 37232
rect 172 35344 212 35384
rect 76 33244 116 33284
rect 76 32992 116 33032
rect 76 32488 116 32528
rect 76 32320 116 32360
rect 556 34000 596 34040
rect 364 31480 404 31520
rect 364 31312 404 31352
rect 748 33664 788 33704
rect 652 31480 692 31520
rect 556 30388 596 30428
rect 172 25180 212 25220
rect 268 21820 308 21860
rect 76 20896 116 20936
rect 76 20224 116 20264
rect 76 17368 116 17408
rect 172 17284 212 17324
rect 76 16612 116 16652
rect 76 10144 116 10184
rect 76 8800 116 8840
rect 556 23920 596 23960
rect 556 19468 596 19508
rect 460 19216 500 19256
rect 460 18544 500 18584
rect 364 12076 404 12116
rect 940 30556 980 30596
rect 940 30388 980 30428
rect 844 30136 884 30176
rect 748 26020 788 26060
rect 748 25852 788 25892
rect 844 25516 884 25556
rect 748 16948 788 16988
rect 652 15772 692 15812
rect 460 11824 500 11864
rect 556 8968 596 9008
rect 556 7288 596 7328
rect 364 6280 404 6320
rect 1612 40888 1652 40928
rect 1420 40720 1460 40760
rect 1324 40384 1364 40424
rect 1324 39712 1364 39752
rect 1420 39376 1460 39416
rect 1324 38956 1364 38996
rect 1324 38116 1364 38156
rect 1516 38704 1556 38744
rect 1516 38368 1556 38408
rect 1420 37612 1460 37652
rect 1900 42064 1940 42104
rect 1804 40468 1844 40508
rect 1708 39040 1748 39080
rect 2284 42148 2324 42188
rect 1996 40300 2036 40340
rect 1996 40132 2036 40172
rect 1900 38200 1940 38240
rect 1708 38116 1748 38156
rect 1804 37948 1844 37988
rect 1612 37192 1652 37232
rect 1516 36940 1556 36980
rect 1228 35764 1268 35804
rect 1420 35932 1460 35972
rect 1612 35932 1652 35972
rect 1804 35932 1844 35972
rect 1324 35176 1364 35216
rect 1516 35092 1556 35132
rect 1420 35008 1460 35048
rect 1324 34924 1364 34964
rect 2572 41896 2612 41936
rect 2380 41560 2420 41600
rect 2380 41056 2420 41096
rect 2860 41224 2900 41264
rect 3340 42148 3380 42188
rect 3148 41560 3188 41600
rect 3340 41560 3380 41600
rect 3052 41056 3092 41096
rect 2956 40552 2996 40592
rect 2956 40384 2996 40424
rect 2860 40300 2900 40340
rect 2476 39040 2516 39080
rect 2572 38872 2612 38912
rect 2380 38368 2420 38408
rect 2284 38200 2324 38240
rect 2188 38116 2228 38156
rect 2188 36268 2228 36308
rect 2092 35932 2132 35972
rect 1996 35680 2036 35720
rect 1804 35176 1844 35216
rect 1324 34672 1364 34712
rect 1516 34588 1556 34628
rect 1708 33832 1748 33872
rect 1324 33496 1364 33536
rect 1228 32824 1268 32864
rect 1612 33664 1652 33704
rect 1612 33412 1652 33452
rect 2092 35176 2132 35216
rect 1900 34840 1940 34880
rect 1900 33580 1940 33620
rect 1996 33496 2036 33536
rect 2092 33412 2132 33452
rect 1804 32992 1844 33032
rect 1804 32824 1844 32864
rect 1612 32404 1652 32444
rect 1900 32404 1940 32444
rect 2188 32908 2228 32948
rect 2860 39544 2900 39584
rect 2956 38872 2996 38912
rect 2476 36688 2516 36728
rect 2572 36436 2612 36476
rect 2572 35764 2612 35804
rect 2380 35344 2420 35384
rect 2476 35176 2516 35216
rect 2380 33076 2420 33116
rect 2188 32656 2228 32696
rect 1324 32236 1364 32276
rect 1324 32068 1364 32108
rect 1228 31312 1268 31352
rect 1708 32068 1748 32108
rect 2092 32068 2132 32108
rect 1612 31984 1652 32024
rect 1228 30556 1268 30596
rect 1132 30136 1172 30176
rect 1420 29968 1460 30008
rect 1612 29968 1652 30008
rect 1324 29800 1364 29840
rect 1132 29044 1172 29084
rect 1324 28876 1364 28916
rect 1516 29632 1556 29672
rect 1900 31312 1940 31352
rect 1804 30640 1844 30680
rect 1708 29548 1748 29588
rect 1708 29212 1748 29252
rect 1516 28960 1556 29000
rect 1420 28372 1460 28412
rect 1516 28204 1556 28244
rect 1324 27448 1364 27488
rect 1228 27028 1268 27068
rect 1420 26860 1460 26900
rect 1132 26188 1172 26228
rect 1612 27616 1652 27656
rect 1612 26776 1652 26816
rect 1324 26440 1364 26480
rect 1420 26272 1460 26312
rect 1324 26104 1364 26144
rect 1516 26104 1556 26144
rect 1804 28456 1844 28496
rect 1804 27700 1844 27740
rect 2284 32320 2324 32360
rect 2188 30808 2228 30848
rect 1996 28120 2036 28160
rect 1905 26944 1945 26984
rect 2092 27700 2132 27740
rect 1996 26188 2036 26228
rect 1228 25936 1268 25976
rect 1324 25600 1364 25640
rect 1324 25432 1364 25472
rect 1036 23248 1076 23288
rect 1900 25012 1940 25052
rect 1324 24928 1364 24968
rect 1324 24424 1364 24464
rect 2092 25432 2132 25472
rect 1996 24172 2036 24212
rect 1516 23920 1556 23960
rect 2092 23920 2132 23960
rect 1420 23752 1460 23792
rect 1324 23584 1364 23624
rect 1324 23332 1364 23372
rect 1516 23248 1556 23288
rect 1708 23584 1748 23624
rect 1708 23080 1748 23120
rect 1900 23584 1940 23624
rect 2284 28876 2324 28916
rect 2572 35092 2612 35132
rect 2860 37108 2900 37148
rect 3148 40384 3188 40424
rect 3148 39712 3188 39752
rect 3916 42400 3956 42440
rect 3340 39880 3380 39920
rect 3340 39376 3380 39416
rect 3244 38956 3284 38996
rect 3340 38284 3380 38324
rect 3148 37780 3188 37820
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 3628 39124 3668 39164
rect 3532 39040 3572 39080
rect 3532 38704 3572 38744
rect 3916 38872 3956 38912
rect 3820 38704 3860 38744
rect 3052 36856 3092 36896
rect 2764 35932 2804 35972
rect 2764 34756 2804 34796
rect 2764 32992 2804 33032
rect 2764 32824 2804 32864
rect 2764 32572 2804 32612
rect 2476 32320 2516 32360
rect 3052 36688 3092 36728
rect 3244 37192 3284 37232
rect 3820 38200 3860 38240
rect 4204 39376 4244 39416
rect 4204 39040 4244 39080
rect 4204 38536 4244 38576
rect 4684 42064 4724 42104
rect 5260 42484 5300 42524
rect 5068 41728 5108 41768
rect 4492 41560 4532 41600
rect 4492 41224 4532 41264
rect 4684 40972 4724 41012
rect 4492 40804 4532 40844
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 5068 41392 5108 41432
rect 4972 41224 5012 41264
rect 5260 41224 5300 41264
rect 5740 42484 5780 42524
rect 5644 41476 5684 41516
rect 5356 40972 5396 41012
rect 5260 40552 5300 40592
rect 4780 40468 4820 40508
rect 4876 40384 4916 40424
rect 4396 39376 4436 39416
rect 4396 39124 4436 39164
rect 4396 38536 4436 38576
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3724 37612 3764 37652
rect 3628 37444 3668 37484
rect 3628 37192 3668 37232
rect 3244 36856 3284 36896
rect 3340 36688 3380 36728
rect 3532 36772 3572 36812
rect 2956 36436 2996 36476
rect 3436 36520 3476 36560
rect 3820 37192 3860 37232
rect 3916 36772 3956 36812
rect 4012 36604 4052 36644
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 3916 36100 3956 36140
rect 4012 35764 4052 35804
rect 3340 35428 3380 35468
rect 3340 34924 3380 34964
rect 2956 34336 2996 34376
rect 4012 35344 4052 35384
rect 3820 35092 3860 35132
rect 3532 35008 3572 35048
rect 4396 38200 4436 38240
rect 4204 36940 4244 36980
rect 4204 36604 4244 36644
rect 4204 36100 4244 36140
rect 4204 35176 4244 35216
rect 4108 35008 4148 35048
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 4204 34756 4244 34796
rect 3244 34336 3284 34376
rect 3148 34168 3188 34208
rect 2956 33580 2996 33620
rect 3148 33412 3188 33452
rect 2956 33328 2996 33368
rect 2764 31984 2804 32024
rect 2476 31480 2516 31520
rect 2668 31312 2708 31352
rect 2476 30556 2516 30596
rect 3532 34252 3572 34292
rect 4204 34168 4244 34208
rect 3532 34000 3572 34040
rect 3820 33832 3860 33872
rect 3436 33580 3476 33620
rect 3244 32992 3284 33032
rect 3148 32908 3188 32948
rect 3244 32824 3284 32864
rect 3052 32656 3092 32696
rect 3340 32572 3380 32612
rect 3244 32320 3284 32360
rect 4108 33664 4148 33704
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 3532 32992 3572 33032
rect 2956 31144 2996 31184
rect 2860 30556 2900 30596
rect 2668 29212 2708 29252
rect 2380 28540 2420 28580
rect 2284 26692 2324 26732
rect 2380 26608 2420 26648
rect 2092 23584 2132 23624
rect 1996 23248 2036 23288
rect 1804 22912 1844 22952
rect 1612 22744 1652 22784
rect 1708 22576 1748 22616
rect 1516 22492 1556 22532
rect 1516 21736 1556 21776
rect 1324 21652 1364 21692
rect 1036 21568 1076 21608
rect 940 17536 980 17576
rect 940 15688 980 15728
rect 940 10984 980 11024
rect 940 6280 980 6320
rect 844 4852 884 4892
rect 748 4768 788 4808
rect 268 4264 308 4304
rect 940 3928 980 3968
rect 172 3256 212 3296
rect 1420 21484 1460 21524
rect 1132 21400 1172 21440
rect 1324 20812 1364 20852
rect 1516 20980 1556 21020
rect 1420 19804 1460 19844
rect 1516 19720 1556 19760
rect 1324 19300 1364 19340
rect 1132 18208 1172 18248
rect 1516 19216 1556 19256
rect 1708 20560 1748 20600
rect 1708 19468 1748 19508
rect 1900 21736 1940 21776
rect 1804 18964 1844 19004
rect 1612 18796 1652 18836
rect 2476 25600 2516 25640
rect 2476 25264 2516 25304
rect 2860 29128 2900 29168
rect 2764 28792 2804 28832
rect 3436 31312 3476 31352
rect 3148 30052 3188 30092
rect 3244 29800 3284 29840
rect 3052 28960 3092 29000
rect 2764 28456 2804 28496
rect 2956 28204 2996 28244
rect 3724 32824 3764 32864
rect 3916 32320 3956 32360
rect 4204 32656 4244 32696
rect 4108 32068 4148 32108
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 4204 31144 4244 31184
rect 4108 30388 4148 30428
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 3628 30052 3668 30092
rect 3340 29464 3380 29504
rect 3244 29380 3284 29420
rect 3244 29212 3284 29252
rect 3244 28960 3284 29000
rect 3148 28456 3188 28496
rect 3148 28288 3188 28328
rect 3532 29380 3572 29420
rect 3052 27868 3092 27908
rect 2860 26692 2900 26732
rect 2764 26608 2804 26648
rect 2956 26272 2996 26312
rect 3244 28036 3284 28076
rect 3148 26272 3188 26312
rect 3052 25768 3092 25808
rect 2860 25516 2900 25556
rect 2668 25432 2708 25472
rect 2380 23584 2420 23624
rect 2476 23164 2516 23204
rect 2380 22324 2420 22364
rect 2188 22156 2228 22196
rect 2284 21988 2324 22028
rect 2092 21484 2132 21524
rect 1516 18376 1556 18416
rect 1612 17620 1652 17660
rect 1420 17116 1460 17156
rect 1324 17032 1364 17072
rect 1324 16444 1364 16484
rect 1612 17032 1652 17072
rect 1804 18460 1844 18500
rect 1804 17704 1844 17744
rect 3436 27448 3476 27488
rect 3340 27028 3380 27068
rect 3916 29800 3956 29840
rect 4588 38704 4628 38744
rect 4588 38116 4628 38156
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 4876 39796 4916 39836
rect 5452 39796 5492 39836
rect 5068 39628 5108 39668
rect 4972 39460 5012 39500
rect 5068 39124 5108 39164
rect 4972 39040 5012 39080
rect 5356 39628 5396 39668
rect 5452 39544 5492 39584
rect 5644 40804 5684 40844
rect 5644 40048 5684 40088
rect 5548 39040 5588 39080
rect 5260 38872 5300 38912
rect 5644 38872 5684 38912
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 5548 38620 5588 38660
rect 5068 38284 5108 38324
rect 4780 38200 4820 38240
rect 4876 37612 4916 37652
rect 4780 37528 4820 37568
rect 4972 37444 5012 37484
rect 4492 37192 4532 37232
rect 4684 37024 4724 37064
rect 4588 36772 4628 36812
rect 4492 36520 4532 36560
rect 4396 35848 4436 35888
rect 4588 35764 4628 35804
rect 4492 35680 4532 35720
rect 4588 35512 4628 35552
rect 4492 35176 4532 35216
rect 4396 34588 4436 34628
rect 4396 32740 4436 32780
rect 4492 32572 4532 32612
rect 4492 32068 4532 32108
rect 4396 31816 4436 31856
rect 5836 41644 5876 41684
rect 6028 40468 6068 40508
rect 5932 40132 5972 40172
rect 6796 41980 6836 42020
rect 6604 41560 6644 41600
rect 6796 41560 6836 41600
rect 6412 41308 6452 41348
rect 6412 41056 6452 41096
rect 6028 40048 6068 40088
rect 5836 39124 5876 39164
rect 5740 37696 5780 37736
rect 5644 37360 5684 37400
rect 5164 37192 5204 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 5164 36772 5204 36812
rect 5644 36772 5684 36812
rect 5548 36604 5588 36644
rect 5548 36352 5588 36392
rect 5356 36184 5396 36224
rect 5068 35848 5108 35888
rect 5260 35848 5300 35888
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4780 35260 4820 35300
rect 5164 35092 5204 35132
rect 4684 34588 4724 34628
rect 4780 34336 4820 34376
rect 5260 34504 5300 34544
rect 4684 33832 4724 33872
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4780 33664 4820 33704
rect 4684 32992 4724 33032
rect 4396 30892 4436 30932
rect 4588 31564 4628 31604
rect 4876 33580 4916 33620
rect 4876 32656 4916 32696
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 5548 35596 5588 35636
rect 5452 35176 5492 35216
rect 5452 34840 5492 34880
rect 5452 34588 5492 34628
rect 5452 34084 5492 34124
rect 6028 38284 6068 38324
rect 6028 36436 6068 36476
rect 6028 35596 6068 35636
rect 5836 35428 5876 35468
rect 6700 40636 6740 40676
rect 6508 40468 6548 40508
rect 6316 39040 6356 39080
rect 6316 38116 6356 38156
rect 6220 38032 6260 38072
rect 6220 35848 6260 35888
rect 6124 35344 6164 35384
rect 5644 35260 5684 35300
rect 5836 35260 5876 35300
rect 6028 35260 6068 35300
rect 5932 35176 5972 35216
rect 5740 35092 5780 35132
rect 5836 35008 5876 35048
rect 6124 35008 6164 35048
rect 5740 34084 5780 34124
rect 5644 34000 5684 34040
rect 5548 33160 5588 33200
rect 5452 32236 5492 32276
rect 4972 32152 5012 32192
rect 5260 32152 5300 32192
rect 5356 31900 5396 31940
rect 4876 31732 4916 31772
rect 4684 31480 4724 31520
rect 4972 31312 5012 31352
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4684 30640 4724 30680
rect 4492 30220 4532 30260
rect 4588 29800 4628 29840
rect 4300 29632 4340 29672
rect 4492 29632 4532 29672
rect 5068 30304 5108 30344
rect 4492 29464 4532 29504
rect 4492 29128 4532 29168
rect 3628 28876 3668 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3724 28540 3764 28580
rect 3628 28372 3668 28412
rect 3820 28456 3860 28496
rect 4012 28372 4052 28412
rect 3724 28036 3764 28076
rect 4204 28540 4244 28580
rect 4492 28708 4532 28748
rect 4300 27532 4340 27572
rect 4684 28876 4724 28916
rect 4588 28288 4628 28328
rect 4492 27700 4532 27740
rect 3916 27448 3956 27488
rect 4108 27364 4148 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 4012 27028 4052 27068
rect 3628 26944 3668 26984
rect 3532 26692 3572 26732
rect 3340 26608 3380 26648
rect 4300 27280 4340 27320
rect 3628 26608 3668 26648
rect 4204 26776 4244 26816
rect 4108 26524 4148 26564
rect 3820 26440 3860 26480
rect 4396 26440 4436 26480
rect 4204 26020 4244 26060
rect 3820 25852 3860 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 4108 25516 4148 25556
rect 3244 25264 3284 25304
rect 3628 25269 3668 25304
rect 3628 25264 3668 25269
rect 3436 25180 3476 25220
rect 3148 25012 3188 25052
rect 3052 24760 3092 24800
rect 3052 24508 3092 24548
rect 2860 23752 2900 23792
rect 3052 23500 3092 23540
rect 2956 23164 2996 23204
rect 2860 23080 2900 23120
rect 2764 21652 2804 21692
rect 2668 21568 2708 21608
rect 2284 20980 2324 21020
rect 3532 24592 3572 24632
rect 3340 23752 3380 23792
rect 3724 24340 3764 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3148 23080 3188 23120
rect 3148 22828 3188 22868
rect 3148 21988 3188 22028
rect 3148 21820 3188 21860
rect 3052 21568 3092 21608
rect 3436 21484 3476 21524
rect 2956 21064 2996 21104
rect 2476 20728 2516 20768
rect 2380 20476 2420 20516
rect 2284 18460 2324 18500
rect 2284 17620 2324 17660
rect 2188 17368 2228 17408
rect 2092 17284 2132 17324
rect 2284 17284 2324 17324
rect 2572 19720 2612 19760
rect 2764 19720 2804 19760
rect 2956 20812 2996 20852
rect 3340 20812 3380 20852
rect 3244 20392 3284 20432
rect 3148 20308 3188 20348
rect 2956 20140 2996 20180
rect 2956 19888 2996 19928
rect 3148 19888 3188 19928
rect 2572 19132 2612 19172
rect 2860 19216 2900 19256
rect 2956 18712 2996 18752
rect 2476 17788 2516 17828
rect 1996 17200 2036 17240
rect 1708 16528 1748 16568
rect 1900 16696 1940 16736
rect 2188 17032 2228 17072
rect 2092 16948 2132 16988
rect 1996 16528 2036 16568
rect 1516 16360 1556 16400
rect 2092 16360 2132 16400
rect 1132 15940 1172 15980
rect 1324 16192 1364 16232
rect 1228 15688 1268 15728
rect 1228 15436 1268 15476
rect 1516 16024 1556 16064
rect 1516 14848 1556 14888
rect 1708 16192 1748 16232
rect 1900 16108 1940 16148
rect 1516 14596 1556 14636
rect 1132 14344 1172 14384
rect 1324 14260 1364 14300
rect 1324 13756 1364 13796
rect 1324 13168 1364 13208
rect 1516 12748 1556 12788
rect 1324 12496 1364 12536
rect 1996 15268 2036 15308
rect 1996 15016 2036 15056
rect 1900 14680 1940 14720
rect 1804 14596 1844 14636
rect 1804 14344 1844 14384
rect 1996 14344 2036 14384
rect 1708 11824 1748 11864
rect 1324 11656 1364 11696
rect 1708 11656 1748 11696
rect 1612 10648 1652 10688
rect 1228 9976 1268 10016
rect 1420 9976 1460 10016
rect 1516 9472 1556 9512
rect 1900 14260 1940 14300
rect 1804 9724 1844 9764
rect 1804 9556 1844 9596
rect 1420 9388 1460 9428
rect 1228 8632 1268 8672
rect 1324 7960 1364 8000
rect 1996 14176 2036 14216
rect 2380 16276 2420 16316
rect 2188 14176 2228 14216
rect 2284 13840 2324 13880
rect 2284 13672 2324 13712
rect 2188 13420 2228 13460
rect 2092 12748 2132 12788
rect 1996 12160 2036 12200
rect 1996 9472 2036 9512
rect 1996 9136 2036 9176
rect 1900 7708 1940 7748
rect 1612 7624 1652 7664
rect 1804 7624 1844 7664
rect 1516 7540 1556 7580
rect 1612 7456 1652 7496
rect 1516 7288 1556 7328
rect 1324 7036 1364 7076
rect 1420 6700 1460 6740
rect 1900 7540 1940 7580
rect 1996 7372 2036 7412
rect 2188 12160 2228 12200
rect 2188 8884 2228 8924
rect 2188 8632 2228 8672
rect 2188 7960 2228 8000
rect 2092 7036 2132 7076
rect 1708 6952 1748 6992
rect 1708 6784 1748 6824
rect 1420 6196 1460 6236
rect 1612 6028 1652 6068
rect 1516 5776 1556 5816
rect 2092 6700 2132 6740
rect 1900 6532 1940 6572
rect 1804 6448 1844 6488
rect 1900 6112 1940 6152
rect 1324 5608 1364 5648
rect 1228 5356 1268 5396
rect 1420 5104 1460 5144
rect 1228 4768 1268 4808
rect 1228 4180 1268 4220
rect 1132 4012 1172 4052
rect 1228 3928 1268 3968
rect 2764 18544 2804 18584
rect 2860 18460 2900 18500
rect 2668 17956 2708 17996
rect 2956 18376 2996 18416
rect 2860 17704 2900 17744
rect 2956 17452 2996 17492
rect 2860 17368 2900 17408
rect 2860 16864 2900 16904
rect 2860 16444 2900 16484
rect 3436 20308 3476 20348
rect 3340 18880 3380 18920
rect 3148 18460 3188 18500
rect 3244 18376 3284 18416
rect 3148 16528 3188 16568
rect 3052 16276 3092 16316
rect 2476 14848 2516 14888
rect 3052 16024 3092 16064
rect 2764 14344 2804 14384
rect 2860 13924 2900 13964
rect 2572 13840 2612 13880
rect 3628 23248 3668 23288
rect 5068 29632 5108 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 4876 29128 4916 29168
rect 5356 28876 5396 28916
rect 4780 28204 4820 28244
rect 5260 28204 5300 28244
rect 4876 28120 4916 28160
rect 4780 27952 4820 27992
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4684 27616 4724 27656
rect 4684 27028 4724 27068
rect 4876 27616 4916 27656
rect 5356 26776 5396 26816
rect 4780 26524 4820 26564
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 4684 26188 4724 26228
rect 5164 26272 5204 26312
rect 4684 25684 4724 25724
rect 4300 24592 4340 24632
rect 4684 25348 4724 25388
rect 5068 25264 5108 25304
rect 5260 25600 5300 25640
rect 4492 25180 4532 25220
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4684 24424 4724 24464
rect 4492 24340 4532 24380
rect 4204 23416 4244 23456
rect 4012 23332 4052 23372
rect 3724 23080 3764 23120
rect 4108 23080 4148 23120
rect 4300 22996 4340 23036
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4684 23332 4724 23372
rect 5164 23080 5204 23120
rect 4588 22996 4628 23036
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3724 22492 3764 22532
rect 3628 22240 3668 22280
rect 4204 22828 4244 22868
rect 4396 22828 4436 22868
rect 4972 22828 5012 22868
rect 4108 21652 4148 21692
rect 3820 21568 3860 21608
rect 4492 22492 4532 22532
rect 4684 22408 4724 22448
rect 4300 22324 4340 22364
rect 4300 21736 4340 21776
rect 3628 21400 3668 21440
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 4204 21064 4244 21104
rect 4108 20644 4148 20684
rect 3820 20560 3860 20600
rect 3820 19804 3860 19844
rect 3532 19720 3572 19760
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3532 19216 3572 19256
rect 3628 19132 3668 19172
rect 3532 18460 3572 18500
rect 4492 20896 4532 20936
rect 4300 20812 4340 20852
rect 4588 19888 4628 19928
rect 4396 19720 4436 19760
rect 3820 19048 3860 19088
rect 4204 19048 4244 19088
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 4876 21652 4916 21692
rect 5260 21400 5300 21440
rect 5164 21316 5204 21356
rect 5356 21232 5396 21272
rect 4972 20644 5012 20684
rect 5356 20812 5396 20852
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 5164 20056 5204 20096
rect 4876 19972 4916 20012
rect 4780 19300 4820 19340
rect 5260 19132 5300 19172
rect 4396 18880 4436 18920
rect 4396 18628 4436 18668
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 5068 18628 5108 18668
rect 3436 18292 3476 18332
rect 3724 18292 3764 18332
rect 3436 16948 3476 16988
rect 3340 16780 3380 16820
rect 3244 16444 3284 16484
rect 3340 15940 3380 15980
rect 3340 15604 3380 15644
rect 3244 15520 3284 15560
rect 3244 15268 3284 15308
rect 3148 15184 3188 15224
rect 3148 14848 3188 14888
rect 3052 13252 3092 13292
rect 2572 12832 2612 12872
rect 2476 11656 2516 11696
rect 2476 8716 2516 8756
rect 2956 12328 2996 12368
rect 3340 14932 3380 14972
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 4204 18040 4244 18080
rect 4780 18292 4820 18332
rect 4684 18040 4724 18080
rect 4396 17788 4436 17828
rect 4588 17788 4628 17828
rect 4108 17704 4148 17744
rect 4300 17704 4340 17744
rect 3916 17116 3956 17156
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 4300 16528 4340 16568
rect 3820 16360 3860 16400
rect 3532 16276 3572 16316
rect 3532 16108 3572 16148
rect 3820 15688 3860 15728
rect 4012 15604 4052 15644
rect 4300 16192 4340 16232
rect 4204 16108 4244 16148
rect 4492 17704 4532 17744
rect 4588 16192 4628 16232
rect 4396 15688 4436 15728
rect 4108 15520 4148 15560
rect 4588 15520 4628 15560
rect 4204 15436 4244 15476
rect 3628 15268 3668 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 4204 15268 4244 15308
rect 4300 15184 4340 15224
rect 4108 14932 4148 14972
rect 3724 14848 3764 14888
rect 4108 14764 4148 14804
rect 3340 12832 3380 12872
rect 4300 14680 4340 14720
rect 3532 13924 3572 13964
rect 4492 13840 4532 13880
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3916 13336 3956 13376
rect 4300 13336 4340 13376
rect 3628 13168 3668 13208
rect 3532 12832 3572 12872
rect 2956 12076 2996 12116
rect 2956 11908 2996 11948
rect 2956 11572 2996 11612
rect 3148 11992 3188 12032
rect 3148 11404 3188 11444
rect 3052 11152 3092 11192
rect 2668 10648 2708 10688
rect 2380 8380 2420 8420
rect 2380 8128 2420 8168
rect 2572 8632 2612 8672
rect 2668 8212 2708 8252
rect 2668 7960 2708 8000
rect 2668 6868 2708 6908
rect 2380 6784 2420 6824
rect 2380 6616 2420 6656
rect 2476 6532 2516 6572
rect 2860 10816 2900 10856
rect 2860 9892 2900 9932
rect 3436 11404 3476 11444
rect 3436 11152 3476 11192
rect 4300 13000 4340 13040
rect 4492 13000 4532 13040
rect 4204 12832 4244 12872
rect 3628 12244 3668 12284
rect 3916 12244 3956 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 4684 14932 4724 14972
rect 5356 18040 5396 18080
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 5932 34840 5972 34880
rect 5740 33748 5780 33788
rect 5836 33664 5876 33704
rect 5644 29128 5684 29168
rect 6892 40300 6932 40340
rect 6892 39628 6932 39668
rect 6508 39376 6548 39416
rect 6796 39376 6836 39416
rect 6604 39040 6644 39080
rect 6892 39040 6932 39080
rect 6508 38872 6548 38912
rect 6892 38788 6932 38828
rect 6508 38032 6548 38072
rect 6412 35260 6452 35300
rect 6700 38200 6740 38240
rect 6892 38032 6932 38072
rect 7276 42400 7316 42440
rect 7180 41560 7220 41600
rect 7084 40216 7124 40256
rect 7564 41812 7604 41852
rect 7660 41728 7700 41768
rect 7372 41560 7412 41600
rect 7468 41476 7508 41516
rect 8140 42736 8180 42776
rect 8524 41812 8564 41852
rect 8332 41644 8372 41684
rect 7948 41560 7988 41600
rect 7084 39628 7124 39668
rect 7276 39544 7316 39584
rect 7084 39376 7124 39416
rect 6988 37864 7028 37904
rect 7276 39124 7316 39164
rect 6700 37780 6740 37820
rect 7468 39040 7508 39080
rect 7660 38368 7700 38408
rect 7852 39628 7892 39668
rect 8140 40972 8180 41012
rect 8044 39208 8084 39248
rect 8908 41728 8948 41768
rect 8332 40972 8372 41012
rect 8332 40216 8372 40256
rect 8524 40216 8564 40256
rect 8428 39628 8468 39668
rect 8140 38872 8180 38912
rect 7276 37696 7316 37736
rect 7468 37612 7508 37652
rect 6796 36016 6836 36056
rect 6412 35092 6452 35132
rect 6508 35008 6548 35048
rect 6508 34672 6548 34712
rect 6604 34588 6644 34628
rect 6508 33664 6548 33704
rect 6220 33580 6260 33620
rect 6124 32404 6164 32444
rect 6028 32236 6068 32276
rect 5932 31984 5972 32024
rect 6604 33580 6644 33620
rect 6316 33412 6356 33452
rect 6988 35764 7028 35804
rect 6988 35512 7028 35552
rect 7372 36436 7412 36476
rect 7372 36184 7412 36224
rect 7564 36184 7604 36224
rect 7276 36016 7316 36056
rect 8332 37612 8372 37652
rect 8140 36688 8180 36728
rect 7948 36268 7988 36308
rect 7564 35848 7604 35888
rect 7372 35596 7412 35636
rect 7852 35848 7892 35888
rect 8140 36436 8180 36476
rect 7660 35428 7700 35468
rect 7756 35344 7796 35384
rect 7660 35176 7700 35216
rect 7372 35008 7412 35048
rect 7084 34840 7124 34880
rect 6988 34336 7028 34376
rect 6700 33076 6740 33116
rect 6796 32740 6836 32780
rect 6508 32488 6548 32528
rect 6700 32236 6740 32276
rect 6508 31984 6548 32024
rect 6220 31564 6260 31604
rect 6220 31396 6260 31436
rect 6508 31228 6548 31268
rect 6604 31060 6644 31100
rect 6508 30808 6548 30848
rect 5548 28792 5588 28832
rect 6508 30388 6548 30428
rect 6316 30220 6356 30260
rect 6316 29716 6356 29756
rect 6700 29968 6740 30008
rect 6700 29632 6740 29672
rect 6124 29380 6164 29420
rect 6508 29296 6548 29336
rect 5740 28792 5780 28832
rect 5548 27196 5588 27236
rect 5548 27028 5588 27068
rect 6316 28876 6356 28916
rect 5932 28708 5972 28748
rect 6124 28708 6164 28748
rect 6508 28708 6548 28748
rect 6220 28540 6260 28580
rect 6124 28372 6164 28412
rect 6316 28372 6356 28412
rect 6220 28036 6260 28076
rect 6124 27952 6164 27992
rect 5836 25852 5876 25892
rect 6124 27028 6164 27068
rect 6220 26776 6260 26816
rect 6700 28372 6740 28412
rect 6700 28120 6740 28160
rect 7852 35092 7892 35132
rect 7660 35008 7700 35048
rect 7372 34168 7412 34208
rect 7084 33748 7124 33788
rect 7276 33748 7316 33788
rect 7372 33664 7412 33704
rect 7276 33580 7316 33620
rect 6988 32152 7028 32192
rect 7180 32404 7220 32444
rect 7084 31984 7124 32024
rect 6988 31900 7028 31940
rect 6892 31648 6932 31688
rect 6892 31480 6932 31520
rect 6892 28708 6932 28748
rect 6892 28372 6932 28412
rect 6892 27952 6932 27992
rect 6700 27616 6740 27656
rect 6604 27448 6644 27488
rect 6412 27364 6452 27404
rect 6700 27364 6740 27404
rect 6508 26776 6548 26816
rect 6028 25348 6068 25388
rect 5644 24844 5684 24884
rect 5548 24592 5588 24632
rect 6220 25516 6260 25556
rect 6124 24844 6164 24884
rect 5932 24592 5972 24632
rect 6508 26524 6548 26564
rect 6796 27112 6836 27152
rect 6700 26524 6740 26564
rect 6604 26440 6644 26480
rect 6892 26104 6932 26144
rect 7564 33748 7604 33788
rect 7564 33076 7604 33116
rect 8044 35008 8084 35048
rect 7756 34252 7796 34292
rect 7660 32992 7700 33032
rect 7756 32824 7796 32864
rect 7468 32572 7508 32612
rect 7564 32404 7604 32444
rect 7468 32152 7508 32192
rect 7372 31480 7412 31520
rect 7372 30724 7412 30764
rect 7276 28708 7316 28748
rect 7084 28120 7124 28160
rect 7276 27532 7316 27572
rect 7180 27112 7220 27152
rect 7276 26776 7316 26816
rect 7180 26608 7220 26648
rect 7180 26440 7220 26480
rect 7084 26272 7124 26312
rect 7276 26188 7316 26228
rect 7180 25180 7220 25220
rect 6988 24928 7028 24968
rect 7180 24928 7220 24968
rect 6412 24760 6452 24800
rect 6700 24760 6740 24800
rect 6988 24760 7028 24800
rect 5836 24508 5876 24548
rect 6028 24340 6068 24380
rect 6124 23920 6164 23960
rect 6604 24592 6644 24632
rect 6796 24592 6836 24632
rect 7180 24592 7220 24632
rect 6988 24340 7028 24380
rect 6700 23836 6740 23876
rect 5836 22912 5876 22952
rect 5548 21148 5588 21188
rect 5548 18712 5588 18752
rect 5548 17200 5588 17240
rect 5548 16192 5588 16232
rect 5452 15688 5492 15728
rect 5068 15520 5108 15560
rect 5260 15436 5300 15476
rect 5548 15520 5588 15560
rect 5452 15268 5492 15308
rect 5452 14932 5492 14972
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4780 14260 4820 14300
rect 4876 14176 4916 14216
rect 4876 13840 4916 13880
rect 5548 14344 5588 14384
rect 5740 19972 5780 20012
rect 5740 19300 5780 19340
rect 5740 19048 5780 19088
rect 5740 17452 5780 17492
rect 5740 16864 5780 16904
rect 5644 14176 5684 14216
rect 6028 22996 6068 23036
rect 6220 22828 6260 22868
rect 5932 22156 5972 22196
rect 6220 22240 6260 22280
rect 6028 21652 6068 21692
rect 6124 21568 6164 21608
rect 6604 23584 6644 23624
rect 6604 23248 6644 23288
rect 6412 22996 6452 23036
rect 7084 23752 7124 23792
rect 7276 24340 7316 24380
rect 7564 31984 7604 32024
rect 7468 29716 7508 29756
rect 7660 31312 7700 31352
rect 7564 29044 7604 29084
rect 7468 27952 7508 27992
rect 8236 36268 8276 36308
rect 8236 35848 8276 35888
rect 8332 35512 8372 35552
rect 8044 34336 8084 34376
rect 8140 34252 8180 34292
rect 8044 33076 8084 33116
rect 7948 32908 7988 32948
rect 8716 40888 8756 40928
rect 8716 40384 8756 40424
rect 8908 39880 8948 39920
rect 9388 41896 9428 41936
rect 9292 41560 9332 41600
rect 8908 38872 8948 38912
rect 8716 38368 8756 38408
rect 8716 38200 8756 38240
rect 8620 37276 8660 37316
rect 8908 38032 8948 38072
rect 8812 37360 8852 37400
rect 8812 36940 8852 36980
rect 8524 36436 8564 36476
rect 8524 36184 8564 36224
rect 8524 35932 8564 35972
rect 8236 33664 8276 33704
rect 8236 33412 8276 33452
rect 8236 32656 8276 32696
rect 8140 32488 8180 32528
rect 8140 31900 8180 31940
rect 7852 31480 7892 31520
rect 7852 31228 7892 31268
rect 7756 30640 7796 30680
rect 7756 29884 7796 29924
rect 8428 34420 8468 34460
rect 8524 33916 8564 33956
rect 8524 33664 8564 33704
rect 8428 33160 8468 33200
rect 8332 31984 8372 32024
rect 8812 36604 8852 36644
rect 9292 38704 9332 38744
rect 9196 38116 9236 38156
rect 9004 37612 9044 37652
rect 9100 37444 9140 37484
rect 9004 36772 9044 36812
rect 8908 36520 8948 36560
rect 8716 36436 8756 36476
rect 8812 35764 8852 35804
rect 8716 35512 8756 35552
rect 8812 35176 8852 35216
rect 9004 35176 9044 35216
rect 8812 35008 8852 35048
rect 9388 37612 9428 37652
rect 9388 37444 9428 37484
rect 9388 37108 9428 37148
rect 9292 36520 9332 36560
rect 9196 36100 9236 36140
rect 9100 34672 9140 34712
rect 8620 32824 8660 32864
rect 8812 34168 8852 34208
rect 8908 33328 8948 33368
rect 8812 32824 8852 32864
rect 8524 32488 8564 32528
rect 8620 32236 8660 32276
rect 8524 32152 8564 32192
rect 8428 31648 8468 31688
rect 8044 30388 8084 30428
rect 7948 29884 7988 29924
rect 7852 29380 7892 29420
rect 7852 29044 7892 29084
rect 7756 28792 7796 28832
rect 7756 28288 7796 28328
rect 7660 27532 7700 27572
rect 7564 26608 7604 26648
rect 7468 26440 7508 26480
rect 7468 26104 7508 26144
rect 7756 26944 7796 26984
rect 7756 26776 7796 26816
rect 7948 28876 7988 28916
rect 7948 28288 7988 28328
rect 7852 26524 7892 26564
rect 7660 25852 7700 25892
rect 7564 25684 7604 25724
rect 7468 24760 7508 24800
rect 7468 24592 7508 24632
rect 7468 24172 7508 24212
rect 7372 24004 7412 24044
rect 7180 23584 7220 23624
rect 6700 22408 6740 22448
rect 6988 22408 7028 22448
rect 6412 22072 6452 22112
rect 6508 21904 6548 21944
rect 6412 21820 6452 21860
rect 6316 21316 6356 21356
rect 6028 20812 6068 20852
rect 6220 20812 6260 20852
rect 6124 20644 6164 20684
rect 6028 20392 6068 20432
rect 5932 17620 5972 17660
rect 6124 19384 6164 19424
rect 6124 18880 6164 18920
rect 6316 17956 6356 17996
rect 6028 17368 6068 17408
rect 6124 17032 6164 17072
rect 6316 17116 6356 17156
rect 5836 16360 5876 16400
rect 5836 16192 5876 16232
rect 6028 16192 6068 16232
rect 5932 15688 5972 15728
rect 5836 14680 5876 14720
rect 6892 22240 6932 22280
rect 6796 21820 6836 21860
rect 6604 21568 6644 21608
rect 6700 21484 6740 21524
rect 6604 21148 6644 21188
rect 6508 16612 6548 16652
rect 6988 21484 7028 21524
rect 8620 31312 8660 31352
rect 8620 30388 8660 30428
rect 8524 30304 8564 30344
rect 8332 30052 8372 30092
rect 8236 29968 8276 30008
rect 8812 31480 8852 31520
rect 8812 30640 8852 30680
rect 8812 30220 8852 30260
rect 8812 29968 8852 30008
rect 9004 32572 9044 32612
rect 9388 35512 9428 35552
rect 9676 42568 9716 42608
rect 9868 41560 9908 41600
rect 9964 40888 10004 40928
rect 10636 41980 10676 42020
rect 10444 41644 10484 41684
rect 10252 41560 10292 41600
rect 10156 40888 10196 40928
rect 10060 40300 10100 40340
rect 10540 40552 10580 40592
rect 10444 40216 10484 40256
rect 10732 40888 10772 40928
rect 10732 40384 10772 40424
rect 10348 39292 10388 39332
rect 9772 38872 9812 38912
rect 10348 38788 10388 38828
rect 9676 38536 9716 38576
rect 10348 38536 10388 38576
rect 9964 37864 10004 37904
rect 9580 37612 9620 37652
rect 10060 37696 10100 37736
rect 9676 37192 9716 37232
rect 9580 36604 9620 36644
rect 9772 36940 9812 36980
rect 10636 39796 10676 39836
rect 10636 39124 10676 39164
rect 10540 39040 10580 39080
rect 10540 38200 10580 38240
rect 10540 37612 10580 37652
rect 10348 37528 10388 37568
rect 10252 37360 10292 37400
rect 10156 36688 10196 36728
rect 9772 36520 9812 36560
rect 10252 36268 10292 36308
rect 9676 36100 9716 36140
rect 9676 35932 9716 35972
rect 9580 35344 9620 35384
rect 9772 35848 9812 35888
rect 9292 33832 9332 33872
rect 9292 33664 9332 33704
rect 9196 32824 9236 32864
rect 9100 32152 9140 32192
rect 9100 31312 9140 31352
rect 9292 32152 9332 32192
rect 10060 35848 10100 35888
rect 10444 36688 10484 36728
rect 10732 37780 10772 37820
rect 10732 37444 10772 37484
rect 10732 36940 10772 36980
rect 10540 36436 10580 36476
rect 10540 36016 10580 36056
rect 10156 35596 10196 35636
rect 10348 35848 10388 35888
rect 10924 41980 10964 42020
rect 11116 42148 11156 42188
rect 11020 41560 11060 41600
rect 10924 39628 10964 39668
rect 10924 37948 10964 37988
rect 10924 36100 10964 36140
rect 9964 35260 10004 35300
rect 10252 35260 10292 35300
rect 10828 35260 10868 35300
rect 9580 33832 9620 33872
rect 9388 31144 9428 31184
rect 10924 34756 10964 34796
rect 10060 34588 10100 34628
rect 11116 37276 11156 37316
rect 11116 36184 11156 36224
rect 11404 41644 11444 41684
rect 11980 42484 12020 42524
rect 11596 41560 11636 41600
rect 12556 42148 12596 42188
rect 11788 41560 11828 41600
rect 12364 41560 12404 41600
rect 11308 39880 11348 39920
rect 11212 36100 11252 36140
rect 11116 36016 11156 36056
rect 11308 36016 11348 36056
rect 11212 35344 11252 35384
rect 11116 34756 11156 34796
rect 10060 34420 10100 34460
rect 9772 33580 9812 33620
rect 9868 32908 9908 32948
rect 10060 34168 10100 34208
rect 10348 34168 10388 34208
rect 10924 34336 10964 34376
rect 11020 34252 11060 34292
rect 10540 34000 10580 34040
rect 10156 33832 10196 33872
rect 10444 33832 10484 33872
rect 10636 33832 10676 33872
rect 10156 33580 10196 33620
rect 10348 33412 10388 33452
rect 10540 33664 10580 33704
rect 9964 32320 10004 32360
rect 10444 32656 10484 32696
rect 10636 32824 10676 32864
rect 10060 32068 10100 32108
rect 9676 31480 9716 31520
rect 9004 30388 9044 30428
rect 8908 29884 8948 29924
rect 8908 29716 8948 29756
rect 8812 29632 8852 29672
rect 8140 29212 8180 29252
rect 8428 29380 8468 29420
rect 8428 29212 8468 29252
rect 8236 28876 8276 28916
rect 8332 27028 8372 27068
rect 8140 26776 8180 26816
rect 8044 26020 8084 26060
rect 8044 25852 8084 25892
rect 7660 23920 7700 23960
rect 7948 23920 7988 23960
rect 7564 23584 7604 23624
rect 7468 23080 7508 23120
rect 8140 24424 8180 24464
rect 9580 30304 9620 30344
rect 8620 28708 8660 28748
rect 8524 28288 8564 28328
rect 9004 28288 9044 28328
rect 8812 27280 8852 27320
rect 9004 27784 9044 27824
rect 9580 30052 9620 30092
rect 9196 29380 9236 29420
rect 9196 28540 9236 28580
rect 9196 28372 9236 28412
rect 9004 27616 9044 27656
rect 9100 27532 9140 27572
rect 9388 29968 9428 30008
rect 9580 29884 9620 29924
rect 9388 29212 9428 29252
rect 9964 30472 10004 30512
rect 10252 31396 10292 31436
rect 10156 31228 10196 31268
rect 10060 29968 10100 30008
rect 9868 29716 9908 29756
rect 9868 29380 9908 29420
rect 9484 27616 9524 27656
rect 9196 27028 9236 27068
rect 9100 26860 9140 26900
rect 9388 26860 9428 26900
rect 9676 27028 9716 27068
rect 9772 26944 9812 26984
rect 9676 26860 9716 26900
rect 9772 26776 9812 26816
rect 8428 26608 8468 26648
rect 9292 26524 9332 26564
rect 8620 26440 8660 26480
rect 8812 26440 8852 26480
rect 9100 26440 9140 26480
rect 8716 26104 8756 26144
rect 8716 25768 8756 25808
rect 8716 25432 8756 25472
rect 8620 23752 8660 23792
rect 8332 23332 8372 23372
rect 7852 22744 7892 22784
rect 7276 22660 7316 22700
rect 7756 22660 7796 22700
rect 7372 22492 7412 22532
rect 7276 22408 7316 22448
rect 7180 21568 7220 21608
rect 7276 21484 7316 21524
rect 7084 21316 7124 21356
rect 6892 21148 6932 21188
rect 6700 19888 6740 19928
rect 7660 22072 7700 22112
rect 7756 21568 7796 21608
rect 7468 21484 7508 21524
rect 6892 20056 6932 20096
rect 6892 19888 6932 19928
rect 6796 18376 6836 18416
rect 6796 17956 6836 17996
rect 7084 19552 7124 19592
rect 7372 19216 7412 19256
rect 6988 19132 7028 19172
rect 6988 18712 7028 18752
rect 7084 18544 7124 18584
rect 6892 17284 6932 17324
rect 6700 17116 6740 17156
rect 6700 16948 6740 16988
rect 6796 16780 6836 16820
rect 6604 16528 6644 16568
rect 6412 16360 6452 16400
rect 6311 16192 6351 16232
rect 6412 16192 6452 16232
rect 6700 15520 6740 15560
rect 6604 15436 6644 15476
rect 6700 15268 6740 15308
rect 6508 15100 6548 15140
rect 6028 14680 6068 14720
rect 5260 13168 5300 13208
rect 5164 13000 5204 13040
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4780 11740 4820 11780
rect 5260 11740 5300 11780
rect 4396 11656 4436 11696
rect 4588 11656 4628 11696
rect 4876 11656 4916 11696
rect 4780 11572 4820 11612
rect 4588 11488 4628 11528
rect 4492 11404 4532 11444
rect 3724 11236 3764 11276
rect 3532 11068 3572 11108
rect 3148 10984 3188 11024
rect 3244 10900 3284 10940
rect 4396 10900 4436 10940
rect 3436 10816 3476 10856
rect 3724 10816 3764 10856
rect 4108 10816 4148 10856
rect 3340 10480 3380 10520
rect 3244 10144 3284 10184
rect 3052 9976 3092 10016
rect 2956 9724 2996 9764
rect 3244 9808 3284 9848
rect 3148 9640 3188 9680
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3532 10312 3572 10352
rect 4012 10312 4052 10352
rect 3532 10060 3572 10100
rect 4204 10648 4244 10688
rect 4204 10312 4244 10352
rect 3532 9556 3572 9596
rect 3724 9556 3764 9596
rect 3052 9472 3092 9512
rect 3436 9472 3476 9512
rect 3340 9220 3380 9260
rect 3244 8884 3284 8924
rect 2956 8548 2996 8588
rect 2188 6196 2228 6236
rect 2668 6196 2708 6236
rect 2092 6028 2132 6068
rect 1900 5440 1940 5480
rect 1612 4600 1652 4640
rect 1804 4432 1844 4472
rect 1708 4348 1748 4388
rect 1516 3760 1556 3800
rect 2284 5776 2324 5816
rect 2380 5608 2420 5648
rect 2188 5524 2228 5564
rect 2092 5188 2132 5228
rect 1996 5020 2036 5060
rect 1996 3928 2036 3968
rect 1708 3760 1748 3800
rect 1420 3592 1460 3632
rect 1324 2752 1364 2792
rect 1612 3676 1652 3716
rect 1516 2836 1556 2876
rect 1612 2752 1652 2792
rect 1708 2248 1748 2288
rect 1420 1408 1460 1448
rect 1708 1324 1748 1364
rect 1516 1156 1556 1196
rect 844 904 884 944
rect 1708 484 1748 524
rect 1900 3592 1940 3632
rect 2284 4180 2324 4220
rect 2188 4096 2228 4136
rect 2188 3844 2228 3884
rect 2092 3172 2132 3212
rect 2188 2584 2228 2624
rect 1996 1996 2036 2036
rect 2188 1576 2228 1616
rect 2092 1072 2132 1112
rect 1996 904 2036 944
rect 2284 1240 2324 1280
rect 2572 5608 2612 5648
rect 2476 3088 2516 3128
rect 2476 1240 2516 1280
rect 2572 1156 2612 1196
rect 2956 7792 2996 7832
rect 3244 6868 3284 6908
rect 3052 6196 3092 6236
rect 2956 6112 2996 6152
rect 3244 6112 3284 6152
rect 3148 4936 3188 4976
rect 2860 4684 2900 4724
rect 3244 4684 3284 4724
rect 3052 3256 3092 3296
rect 3820 9472 3860 9512
rect 4300 9472 4340 9512
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3532 8632 3572 8672
rect 3724 8296 3764 8336
rect 3724 8044 3764 8084
rect 5068 11488 5108 11528
rect 4780 11320 4820 11360
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 5068 11152 5108 11192
rect 4972 11068 5012 11108
rect 4780 10228 4820 10268
rect 5164 10900 5204 10940
rect 4684 10060 4724 10100
rect 4588 9976 4628 10016
rect 4492 9808 4532 9848
rect 4492 9640 4532 9680
rect 5068 10060 5108 10100
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 5548 13168 5588 13208
rect 5452 12748 5492 12788
rect 5740 13000 5780 13040
rect 5644 12580 5684 12620
rect 5548 10984 5588 11024
rect 5836 12664 5876 12704
rect 6220 14512 6260 14552
rect 6124 13420 6164 13460
rect 6124 13168 6164 13208
rect 6028 12748 6068 12788
rect 5836 12412 5876 12452
rect 4876 9640 4916 9680
rect 4300 8884 4340 8924
rect 4972 9052 5012 9092
rect 4684 8884 4724 8924
rect 4204 8632 4244 8672
rect 4108 7876 4148 7916
rect 4204 7792 4244 7832
rect 3628 7708 3668 7748
rect 3820 7708 3860 7748
rect 4396 8380 4436 8420
rect 4396 7876 4436 7916
rect 3532 7624 3572 7664
rect 4300 7624 4340 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3820 7372 3860 7412
rect 3436 7288 3476 7328
rect 4108 7288 4148 7328
rect 4012 7204 4052 7244
rect 3916 6952 3956 6992
rect 3724 6448 3764 6488
rect 4972 8716 5012 8756
rect 4876 8632 4916 8672
rect 4780 8548 4820 8588
rect 5356 8632 5396 8672
rect 5548 10144 5588 10184
rect 5740 10312 5780 10352
rect 5740 10060 5780 10100
rect 4588 7540 4628 7580
rect 4492 7372 4532 7412
rect 4204 7120 4244 7160
rect 3436 6196 3476 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 4204 5944 4244 5984
rect 3532 5776 3572 5816
rect 3436 4432 3476 4472
rect 4204 5440 4244 5480
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3628 3760 3668 3800
rect 3340 3592 3380 3632
rect 3532 3592 3572 3632
rect 4300 4096 4340 4136
rect 3820 4012 3860 4052
rect 4588 6700 4628 6740
rect 4684 6532 4724 6572
rect 4492 6112 4532 6152
rect 4492 4936 4532 4976
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4972 8128 5012 8168
rect 5068 7960 5108 8000
rect 5164 7792 5204 7832
rect 5452 8464 5492 8504
rect 5457 8212 5497 8252
rect 5260 7456 5300 7496
rect 5644 9472 5684 9512
rect 6316 13336 6356 13376
rect 6316 13000 6356 13040
rect 6508 13672 6548 13712
rect 7372 18376 7412 18416
rect 7180 17704 7220 17744
rect 7084 16948 7124 16988
rect 7180 16276 7220 16316
rect 6892 16108 6932 16148
rect 7084 16024 7124 16064
rect 7372 16612 7412 16652
rect 7276 15940 7316 15980
rect 6892 15604 6932 15644
rect 6988 15436 7028 15476
rect 7180 15604 7220 15644
rect 7276 15520 7316 15560
rect 7084 14680 7124 14720
rect 6604 13504 6644 13544
rect 6412 12496 6452 12536
rect 6700 13168 6740 13208
rect 6604 13000 6644 13040
rect 6028 12244 6068 12284
rect 6220 12244 6260 12284
rect 5932 11320 5972 11360
rect 6604 11740 6644 11780
rect 6892 14512 6932 14552
rect 6892 13588 6932 13628
rect 7180 14260 7220 14300
rect 6988 13252 7028 13292
rect 7180 13252 7220 13292
rect 6892 12328 6932 12368
rect 7084 12244 7124 12284
rect 6988 11824 7028 11864
rect 6988 11656 7028 11696
rect 6220 11068 6260 11108
rect 6412 11068 6452 11108
rect 6028 10984 6068 11024
rect 6028 10228 6068 10268
rect 6220 10060 6260 10100
rect 6124 9472 6164 9512
rect 6892 11320 6932 11360
rect 6604 11236 6644 11276
rect 6604 11068 6644 11108
rect 5740 8884 5780 8924
rect 6028 8800 6068 8840
rect 5740 8212 5780 8252
rect 5644 7372 5684 7412
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 5644 7036 5684 7076
rect 5548 6196 5588 6236
rect 4780 6028 4820 6068
rect 5356 5944 5396 5984
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4396 3844 4436 3884
rect 3724 3592 3764 3632
rect 3436 3340 3476 3380
rect 3340 3172 3380 3212
rect 3244 2920 3284 2960
rect 3148 2416 3188 2456
rect 2956 2248 2996 2288
rect 2860 1660 2900 1700
rect 2764 1240 2804 1280
rect 3436 2920 3476 2960
rect 3724 3424 3764 3464
rect 4588 4348 4628 4388
rect 4588 4096 4628 4136
rect 4492 3592 4532 3632
rect 4108 3508 4148 3548
rect 4012 3340 4052 3380
rect 4972 4852 5012 4892
rect 4876 4684 4916 4724
rect 4780 4348 4820 4388
rect 4780 4180 4820 4220
rect 5356 4516 5396 4556
rect 5356 4096 5396 4136
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 5452 3676 5492 3716
rect 4492 3340 4532 3380
rect 4204 3088 4244 3128
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 3532 2668 3572 2708
rect 3436 2416 3476 2456
rect 3052 1324 3092 1364
rect 3340 1240 3380 1280
rect 3628 2584 3668 2624
rect 4108 2248 4148 2288
rect 4012 2164 4052 2204
rect 4012 1912 4052 1952
rect 4684 3172 4724 3212
rect 4972 3592 5012 3632
rect 4972 3172 5012 3212
rect 4972 2836 5012 2876
rect 5068 2752 5108 2792
rect 4780 2668 4820 2708
rect 4588 2416 4628 2456
rect 4492 2332 4532 2372
rect 4204 2164 4244 2204
rect 4396 2164 4436 2204
rect 3628 1744 3668 1784
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 3148 1072 3188 1112
rect 3532 904 3572 944
rect 3436 820 3476 860
rect 4012 1324 4052 1364
rect 3916 1240 3956 1280
rect 4300 1492 4340 1532
rect 4204 1240 4244 1280
rect 4108 1072 4148 1112
rect 5260 2500 5300 2540
rect 5164 2416 5204 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 5068 2080 5108 2120
rect 4780 1240 4820 1280
rect 4684 1072 4724 1112
rect 5260 1156 5300 1196
rect 6316 9052 6356 9092
rect 6220 8800 6260 8840
rect 6220 8296 6260 8336
rect 6028 6616 6068 6656
rect 5932 5860 5972 5900
rect 6124 5776 6164 5816
rect 5740 5692 5780 5732
rect 5644 4852 5684 4892
rect 5836 5104 5876 5144
rect 5740 3424 5780 3464
rect 5644 2752 5684 2792
rect 6028 5524 6068 5564
rect 5932 4936 5972 4976
rect 5932 4264 5972 4304
rect 5932 3760 5972 3800
rect 5548 2584 5588 2624
rect 6124 4936 6164 4976
rect 6700 9052 6740 9092
rect 6700 8380 6740 8420
rect 6700 8212 6740 8252
rect 6508 7624 6548 7664
rect 6508 7372 6548 7412
rect 6796 7204 6836 7244
rect 6700 7036 6740 7076
rect 6508 6616 6548 6656
rect 6412 6280 6452 6320
rect 6604 6280 6644 6320
rect 6316 5272 6356 5312
rect 6988 9556 7028 9596
rect 7756 21148 7796 21188
rect 7564 19216 7604 19256
rect 7564 18544 7604 18584
rect 7852 19804 7892 19844
rect 7756 18124 7796 18164
rect 8140 22156 8180 22196
rect 8428 22072 8468 22112
rect 8044 19300 8084 19340
rect 8044 18544 8084 18584
rect 7948 18124 7988 18164
rect 7756 17620 7796 17660
rect 7660 16360 7700 16400
rect 7756 15436 7796 15476
rect 7660 15184 7700 15224
rect 7564 15016 7604 15056
rect 7564 14596 7604 14636
rect 7468 14008 7508 14048
rect 7468 13756 7508 13796
rect 7660 13504 7700 13544
rect 7468 13168 7508 13208
rect 7948 17620 7988 17660
rect 7948 17452 7988 17492
rect 8332 19972 8372 20012
rect 8236 19720 8276 19760
rect 8140 17788 8180 17828
rect 8524 21484 8564 21524
rect 8908 25852 8948 25892
rect 9004 23752 9044 23792
rect 8908 23164 8948 23204
rect 8812 20896 8852 20936
rect 9196 26188 9236 26228
rect 9388 26104 9428 26144
rect 9196 25348 9236 25388
rect 9580 26440 9620 26480
rect 9484 25348 9524 25388
rect 9388 25264 9428 25304
rect 9388 23752 9428 23792
rect 9484 23668 9524 23708
rect 9196 22576 9236 22616
rect 9292 21988 9332 22028
rect 9100 21568 9140 21608
rect 9004 21232 9044 21272
rect 9004 20896 9044 20936
rect 8620 19216 8660 19256
rect 8524 18544 8564 18584
rect 8812 19216 8852 19256
rect 8908 18712 8948 18752
rect 8524 17536 8564 17576
rect 8716 17620 8756 17660
rect 8620 17452 8660 17492
rect 8236 17032 8276 17072
rect 8236 16780 8276 16820
rect 8140 16192 8180 16232
rect 8428 16528 8468 16568
rect 8332 14848 8372 14888
rect 8332 14512 8372 14552
rect 7948 14344 7988 14384
rect 7852 13252 7892 13292
rect 7564 12580 7604 12620
rect 7372 12244 7412 12284
rect 7372 11656 7412 11696
rect 7276 11488 7316 11528
rect 7276 11236 7316 11276
rect 7180 11152 7220 11192
rect 7180 10060 7220 10100
rect 7564 11572 7604 11612
rect 7468 11320 7508 11360
rect 7468 10564 7508 10604
rect 7276 9724 7316 9764
rect 7084 8800 7124 8840
rect 7084 8548 7124 8588
rect 7180 8464 7220 8504
rect 7084 8296 7124 8336
rect 7084 8128 7124 8168
rect 7084 7792 7124 7832
rect 7660 11236 7700 11276
rect 7660 10648 7700 10688
rect 7948 11824 7988 11864
rect 7948 11656 7988 11696
rect 7948 11236 7988 11276
rect 8140 12328 8180 12368
rect 8332 13084 8372 13124
rect 8716 17116 8756 17156
rect 9388 21568 9428 21608
rect 9196 20476 9236 20516
rect 9196 20056 9236 20096
rect 9196 18880 9236 18920
rect 10540 32320 10580 32360
rect 10540 32068 10580 32108
rect 10636 31984 10676 32024
rect 10924 34168 10964 34208
rect 10924 33412 10964 33452
rect 10828 32656 10868 32696
rect 11308 34924 11348 34964
rect 11980 41056 12020 41096
rect 11500 40804 11540 40844
rect 12172 40636 12212 40676
rect 12076 40132 12116 40172
rect 12172 39964 12212 40004
rect 12076 39796 12116 39836
rect 11596 39124 11636 39164
rect 11500 37612 11540 37652
rect 11500 37360 11540 37400
rect 11980 39460 12020 39500
rect 11692 38200 11732 38240
rect 11596 36940 11636 36980
rect 11500 36520 11540 36560
rect 11596 36100 11636 36140
rect 12172 39292 12212 39332
rect 11980 38452 12020 38492
rect 11788 36772 11828 36812
rect 11788 36016 11828 36056
rect 11404 34756 11444 34796
rect 11500 34672 11540 34712
rect 11500 34420 11540 34460
rect 11404 34336 11444 34376
rect 11308 33832 11348 33872
rect 11692 34000 11732 34040
rect 11596 32824 11636 32864
rect 11212 32488 11252 32528
rect 10828 32236 10868 32276
rect 10732 31480 10772 31520
rect 10348 31228 10388 31268
rect 10444 31144 10484 31184
rect 10348 30556 10388 30596
rect 9964 28708 10004 28748
rect 9964 27280 10004 27320
rect 9868 26104 9908 26144
rect 10540 30388 10580 30428
rect 10348 27952 10388 27992
rect 10156 26944 10196 26984
rect 9676 24424 9716 24464
rect 10060 25684 10100 25724
rect 9964 25264 10004 25304
rect 10924 31228 10964 31268
rect 12076 36856 12116 36896
rect 12748 40804 12788 40844
rect 12364 40132 12404 40172
rect 12364 39964 12404 40004
rect 12556 39964 12596 40004
rect 12844 40132 12884 40172
rect 13324 42148 13364 42188
rect 13516 42064 13556 42104
rect 13900 42232 13940 42272
rect 13708 41980 13748 42020
rect 13132 40552 13172 40592
rect 12556 39712 12596 39752
rect 12460 39460 12500 39500
rect 12556 39292 12596 39332
rect 12364 39124 12404 39164
rect 12268 38284 12308 38324
rect 12364 38200 12404 38240
rect 12556 38200 12596 38240
rect 12364 37948 12404 37988
rect 12268 37360 12308 37400
rect 12172 36688 12212 36728
rect 12076 36520 12116 36560
rect 11980 36100 12020 36140
rect 11980 34588 12020 34628
rect 11980 34336 12020 34376
rect 12172 36352 12212 36392
rect 12172 34588 12212 34628
rect 12460 37696 12500 37736
rect 12364 36688 12404 36728
rect 12364 36184 12404 36224
rect 13036 39712 13076 39752
rect 12748 38368 12788 38408
rect 12748 38032 12788 38072
rect 12844 37612 12884 37652
rect 12940 37444 12980 37484
rect 12652 37276 12692 37316
rect 12652 37108 12692 37148
rect 12556 36688 12596 36728
rect 13132 38872 13172 38912
rect 13132 37948 13172 37988
rect 13132 37360 13172 37400
rect 12556 36352 12596 36392
rect 12844 36100 12884 36140
rect 12556 36016 12596 36056
rect 12268 34504 12308 34544
rect 12364 34000 12404 34040
rect 12076 33832 12116 33872
rect 11788 33683 11828 33704
rect 11788 33664 11828 33683
rect 11884 33664 11924 33704
rect 12364 33160 12404 33200
rect 11404 32404 11444 32444
rect 11116 32320 11156 32360
rect 11212 31564 11252 31604
rect 11308 31312 11348 31352
rect 11020 31144 11060 31184
rect 10924 31060 10964 31100
rect 11116 30724 11156 30764
rect 11212 30556 11252 30596
rect 11212 30220 11252 30260
rect 11116 29632 11156 29672
rect 11500 32152 11540 32192
rect 11692 32068 11732 32108
rect 12844 35848 12884 35888
rect 13132 36352 13172 36392
rect 13036 35596 13076 35636
rect 13324 37192 13364 37232
rect 13804 40972 13844 41012
rect 13612 40300 13652 40340
rect 13516 39544 13556 39584
rect 14092 40468 14132 40508
rect 14668 42904 14708 42944
rect 14476 41644 14516 41684
rect 14476 41140 14516 41180
rect 14284 40384 14324 40424
rect 13996 40300 14036 40340
rect 13900 40048 13940 40088
rect 13708 39040 13748 39080
rect 13897 39054 13937 39080
rect 13897 39040 13900 39054
rect 13900 39040 13937 39054
rect 13516 38956 13556 38996
rect 13612 38620 13652 38660
rect 13516 38452 13556 38492
rect 13516 37948 13556 37988
rect 13708 37612 13748 37652
rect 13516 37444 13556 37484
rect 13708 37360 13748 37400
rect 14188 39964 14228 40004
rect 14092 38452 14132 38492
rect 15052 41896 15092 41936
rect 15244 41476 15284 41516
rect 14860 40804 14900 40844
rect 14860 40384 14900 40424
rect 14668 40300 14708 40340
rect 14572 39964 14612 40004
rect 14476 39460 14516 39500
rect 14572 39376 14612 39416
rect 14284 39292 14324 39332
rect 14284 39124 14324 39164
rect 14380 38788 14420 38828
rect 14765 39376 14805 39416
rect 14764 39124 14804 39164
rect 14668 38872 14708 38912
rect 15148 40216 15188 40256
rect 14956 39964 14996 40004
rect 15628 41560 15668 41600
rect 15532 41392 15572 41432
rect 15436 41140 15476 41180
rect 15436 40972 15476 41012
rect 15628 41056 15668 41096
rect 15052 39796 15092 39836
rect 14956 39712 14996 39752
rect 14860 38872 14900 38912
rect 15052 38704 15092 38744
rect 14476 38452 14516 38492
rect 14860 38452 14900 38492
rect 14668 38368 14708 38408
rect 13900 37612 13940 37652
rect 14284 38200 14324 38240
rect 14572 38200 14612 38240
rect 14188 38032 14228 38072
rect 13804 37108 13844 37148
rect 13420 35596 13460 35636
rect 13708 36100 13748 36140
rect 13900 36184 13940 36224
rect 13612 36016 13652 36056
rect 13612 35596 13652 35636
rect 13228 35176 13268 35216
rect 13132 35092 13172 35132
rect 13036 34252 13076 34292
rect 12652 33244 12692 33284
rect 11884 32404 11924 32444
rect 12076 32824 12116 32864
rect 12268 32824 12308 32864
rect 12172 32740 12212 32780
rect 12364 32656 12404 32696
rect 11980 32236 12020 32276
rect 11500 31228 11540 31268
rect 11500 30724 11540 30764
rect 11404 30640 11444 30680
rect 11692 31480 11732 31520
rect 11884 31060 11924 31100
rect 12556 32656 12596 32696
rect 13324 35092 13364 35132
rect 13228 34084 13268 34124
rect 13516 35344 13556 35384
rect 13516 34924 13556 34964
rect 14092 37360 14132 37400
rect 14668 38032 14708 38072
rect 14572 37948 14612 37988
rect 14380 37612 14420 37652
rect 14284 37360 14324 37400
rect 15244 39712 15284 39752
rect 15244 39460 15284 39500
rect 15532 40384 15572 40424
rect 16204 42484 16244 42524
rect 16396 42316 16436 42356
rect 16492 41308 16532 41348
rect 16300 41224 16340 41264
rect 16012 41056 16052 41096
rect 16108 40972 16148 41012
rect 15820 40384 15860 40424
rect 15436 40300 15476 40340
rect 15532 40216 15572 40256
rect 15436 39964 15476 40004
rect 15340 39292 15380 39332
rect 15340 39040 15380 39080
rect 15148 38368 15188 38408
rect 15052 38200 15092 38240
rect 14956 38032 14996 38072
rect 16300 40636 16340 40676
rect 16588 40972 16628 41012
rect 16876 41392 16916 41432
rect 17548 42820 17588 42860
rect 17356 42652 17396 42692
rect 17644 42148 17684 42188
rect 17164 41476 17204 41516
rect 17260 41308 17300 41348
rect 17068 41224 17108 41264
rect 17068 40972 17108 41012
rect 16972 40720 17012 40760
rect 17836 42736 17876 42776
rect 17740 41392 17780 41432
rect 18124 42568 18164 42608
rect 18028 41644 18068 41684
rect 17932 41476 17972 41516
rect 17548 40972 17588 41012
rect 16012 40300 16052 40340
rect 15916 39964 15956 40004
rect 16300 39880 16340 39920
rect 15820 39460 15860 39500
rect 15628 39376 15668 39416
rect 15532 39040 15572 39080
rect 15244 37696 15284 37736
rect 15436 38200 15476 38240
rect 16204 39712 16244 39752
rect 16012 39628 16052 39668
rect 16684 40384 16724 40424
rect 16588 39796 16628 39836
rect 16492 39460 16532 39500
rect 15916 38872 15956 38912
rect 15724 38452 15764 38492
rect 16396 38620 16436 38660
rect 15628 38116 15668 38156
rect 15820 38032 15860 38072
rect 15532 37948 15572 37988
rect 16012 37948 16052 37988
rect 15340 37612 15380 37652
rect 15532 37612 15572 37652
rect 14764 37444 14804 37484
rect 14668 37360 14708 37400
rect 14188 37192 14228 37232
rect 14380 37192 14420 37232
rect 14092 37024 14132 37064
rect 13708 35344 13748 35384
rect 13612 34588 13652 34628
rect 13708 34504 13748 34544
rect 13708 34252 13748 34292
rect 13420 33832 13460 33872
rect 13324 33244 13364 33284
rect 12844 32992 12884 33032
rect 12748 32488 12788 32528
rect 13036 32824 13076 32864
rect 13132 32740 13172 32780
rect 13036 32488 13076 32528
rect 12940 32404 12980 32444
rect 12172 32068 12212 32108
rect 12460 31732 12500 31772
rect 12652 32152 12692 32192
rect 12748 32068 12788 32108
rect 12172 31396 12212 31436
rect 12556 31396 12596 31436
rect 12748 31312 12788 31352
rect 12268 31060 12308 31100
rect 12172 30892 12212 30932
rect 11884 30556 11924 30596
rect 11404 30388 11444 30428
rect 11980 30388 12020 30428
rect 12364 30808 12404 30848
rect 12556 30724 12596 30764
rect 11404 30220 11444 30260
rect 11788 30220 11828 30260
rect 11596 29632 11636 29672
rect 11404 29128 11444 29168
rect 11596 29128 11636 29168
rect 10636 27952 10676 27992
rect 10348 27112 10388 27152
rect 10252 26524 10292 26564
rect 10252 26272 10292 26312
rect 10156 24676 10196 24716
rect 10060 24592 10100 24632
rect 9964 24424 10004 24464
rect 9868 23920 9908 23960
rect 9772 23836 9812 23876
rect 9676 22744 9716 22784
rect 9676 21568 9716 21608
rect 9580 21316 9620 21356
rect 9676 21232 9716 21272
rect 9676 20728 9716 20768
rect 9484 20392 9524 20432
rect 9388 19552 9428 19592
rect 9580 20056 9620 20096
rect 9772 19636 9812 19676
rect 9772 19468 9812 19508
rect 9292 18544 9332 18584
rect 9196 17704 9236 17744
rect 9100 17536 9140 17576
rect 9004 17368 9044 17408
rect 9004 17032 9044 17072
rect 8908 16696 8948 16736
rect 9580 17704 9620 17744
rect 9484 17536 9524 17576
rect 9292 16864 9332 16904
rect 9388 16612 9428 16652
rect 9100 16360 9140 16400
rect 8524 13168 8564 13208
rect 8332 12328 8372 12368
rect 8332 11488 8372 11528
rect 8908 15604 8948 15644
rect 8908 15352 8948 15392
rect 8812 14848 8852 14888
rect 8716 14596 8756 14636
rect 8812 14512 8852 14552
rect 9100 16192 9140 16232
rect 9292 15604 9332 15644
rect 9100 15352 9140 15392
rect 9004 15184 9044 15224
rect 9388 15520 9428 15560
rect 9196 14680 9236 14720
rect 9196 14344 9236 14384
rect 8716 14176 8756 14216
rect 8716 12076 8756 12116
rect 8716 11908 8756 11948
rect 8620 11656 8660 11696
rect 8620 11320 8660 11360
rect 8044 11068 8084 11108
rect 8236 10984 8276 11024
rect 8044 10900 8084 10940
rect 7852 10144 7892 10184
rect 7756 9976 7796 10016
rect 7756 9472 7796 9512
rect 8044 10144 8084 10184
rect 7660 8632 7700 8672
rect 7468 8212 7508 8252
rect 7372 7708 7412 7748
rect 7564 7372 7604 7412
rect 7276 7120 7316 7160
rect 7276 6952 7316 6992
rect 7468 6952 7508 6992
rect 7180 5104 7220 5144
rect 6892 5020 6932 5060
rect 6796 4936 6836 4976
rect 6508 4852 6548 4892
rect 6220 4264 6260 4304
rect 6124 3340 6164 3380
rect 6988 4852 7028 4892
rect 6988 4348 7028 4388
rect 7084 4096 7124 4136
rect 6700 3928 6740 3968
rect 6412 3760 6452 3800
rect 6316 3676 6356 3716
rect 6316 3508 6356 3548
rect 6412 3256 6452 3296
rect 6220 3004 6260 3044
rect 6124 2752 6164 2792
rect 5932 2584 5972 2624
rect 6316 2584 6356 2624
rect 5836 2500 5876 2540
rect 6028 2500 6068 2540
rect 5452 2416 5492 2456
rect 5740 2248 5780 2288
rect 5548 2080 5588 2120
rect 5644 1240 5684 1280
rect 5452 1156 5492 1196
rect 5932 2164 5972 2204
rect 5356 1072 5396 1112
rect 7372 6196 7412 6236
rect 7372 5692 7412 5732
rect 7372 5188 7412 5228
rect 7948 8800 7988 8840
rect 7852 7120 7892 7160
rect 8140 8800 8180 8840
rect 8044 8464 8084 8504
rect 8044 7960 8084 8000
rect 8524 11068 8564 11108
rect 8428 10396 8468 10436
rect 8524 10144 8564 10184
rect 8332 8464 8372 8504
rect 8524 9388 8564 9428
rect 8620 9136 8660 9176
rect 8524 8968 8564 9008
rect 8620 8716 8660 8756
rect 8332 7708 8372 7748
rect 8236 7372 8276 7412
rect 8428 7456 8468 7496
rect 8044 7120 8084 7160
rect 8332 6868 8372 6908
rect 8044 6616 8084 6656
rect 7564 6448 7604 6488
rect 7660 6364 7700 6404
rect 7564 6280 7604 6320
rect 8044 6280 8084 6320
rect 7948 5104 7988 5144
rect 7756 4936 7796 4976
rect 7756 4768 7796 4808
rect 7948 4516 7988 4556
rect 7660 4264 7700 4304
rect 7372 3844 7412 3884
rect 6796 3592 6836 3632
rect 6988 2584 7028 2624
rect 6508 1912 6548 1952
rect 6988 1912 7028 1952
rect 6892 1828 6932 1868
rect 6796 1744 6836 1784
rect 6124 1660 6164 1700
rect 6220 1240 6260 1280
rect 6604 1240 6644 1280
rect 6796 1240 6836 1280
rect 6988 1240 7028 1280
rect 6124 1156 6164 1196
rect 4876 988 4916 1028
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 4876 568 4916 608
rect 5260 568 5300 608
rect 5068 64 5108 104
rect 5452 652 5492 692
rect 5356 232 5396 272
rect 5548 400 5588 440
rect 5836 652 5876 692
rect 6028 904 6068 944
rect 5932 484 5972 524
rect 6124 148 6164 188
rect 6412 568 6452 608
rect 7468 3004 7508 3044
rect 7372 2920 7412 2960
rect 7564 2500 7604 2540
rect 7468 2332 7508 2372
rect 7276 1324 7316 1364
rect 7180 1240 7220 1280
rect 7084 1072 7124 1112
rect 7468 1156 7508 1196
rect 8140 5860 8180 5900
rect 8908 14092 8948 14132
rect 10156 24340 10196 24380
rect 10060 22912 10100 22952
rect 10636 27280 10676 27320
rect 10444 26776 10484 26816
rect 10444 25852 10484 25892
rect 10636 26860 10676 26900
rect 10636 25936 10676 25976
rect 10540 25684 10580 25724
rect 10540 25516 10580 25556
rect 10540 23668 10580 23708
rect 10348 23584 10388 23624
rect 10348 23416 10388 23456
rect 10252 22744 10292 22784
rect 10060 22660 10100 22700
rect 10252 22576 10292 22616
rect 10060 22240 10100 22280
rect 9964 20056 10004 20096
rect 10060 19636 10100 19676
rect 9964 19468 10004 19508
rect 9868 18880 9908 18920
rect 9580 17116 9620 17156
rect 9772 17116 9812 17156
rect 9676 16276 9716 16316
rect 9772 16024 9812 16064
rect 9676 15856 9716 15896
rect 9964 17200 10004 17240
rect 9964 16192 10004 16232
rect 9964 15940 10004 15980
rect 9772 15352 9812 15392
rect 9484 15100 9524 15140
rect 9388 13840 9428 13880
rect 9772 15184 9812 15224
rect 9676 14680 9716 14720
rect 10251 19132 10291 19172
rect 10252 16192 10292 16232
rect 10156 15856 10196 15896
rect 9964 14932 10004 14972
rect 9964 14764 10004 14804
rect 9676 14428 9716 14468
rect 9676 13588 9716 13628
rect 9772 13420 9812 13460
rect 9292 12160 9332 12200
rect 9772 12664 9812 12704
rect 9676 12412 9716 12452
rect 9964 14512 10004 14552
rect 9964 14344 10004 14384
rect 9964 14176 10004 14216
rect 10444 23080 10484 23120
rect 10540 22660 10580 22700
rect 10732 25348 10772 25388
rect 11308 28708 11348 28748
rect 11212 28624 11252 28664
rect 11020 28456 11060 28496
rect 10924 28288 10964 28328
rect 11308 28288 11348 28328
rect 12460 30388 12500 30428
rect 12364 29884 12404 29924
rect 12076 29716 12116 29756
rect 11788 28960 11828 29000
rect 11692 28456 11732 28496
rect 11980 28456 12020 28496
rect 11404 27616 11444 27656
rect 11116 26692 11156 26732
rect 10924 26272 10964 26312
rect 10828 25264 10868 25304
rect 11212 26104 11252 26144
rect 11116 26020 11156 26060
rect 10924 24508 10964 24548
rect 10828 24340 10868 24380
rect 10732 23920 10772 23960
rect 11116 24508 11156 24548
rect 11596 28288 11636 28328
rect 11788 28120 11828 28160
rect 11692 27868 11732 27908
rect 11500 27112 11540 27152
rect 11500 26944 11540 26984
rect 11500 26524 11540 26564
rect 11404 25852 11444 25892
rect 11596 25348 11636 25388
rect 10924 23500 10964 23540
rect 10732 23080 10772 23120
rect 11404 23668 11444 23708
rect 11404 22828 11444 22868
rect 11404 22576 11444 22616
rect 11308 22408 11348 22448
rect 10732 21736 10772 21776
rect 10444 21568 10484 21608
rect 10444 19804 10484 19844
rect 10540 19636 10580 19676
rect 10924 21568 10964 21608
rect 10444 19132 10484 19172
rect 10444 18796 10484 18836
rect 11308 21988 11348 22028
rect 11404 20728 11444 20768
rect 11596 23668 11636 23708
rect 12556 30220 12596 30260
rect 12364 29464 12404 29504
rect 12460 29212 12500 29252
rect 12268 29044 12308 29084
rect 12172 28792 12212 28832
rect 12748 29884 12788 29924
rect 13132 32404 13172 32444
rect 12940 32068 12980 32108
rect 13036 31480 13076 31520
rect 12940 30556 12980 30596
rect 13324 32152 13364 32192
rect 13228 32068 13268 32108
rect 13612 33664 13652 33704
rect 13804 33076 13844 33116
rect 13708 32824 13748 32864
rect 13708 31984 13748 32024
rect 13612 31564 13652 31604
rect 13228 31228 13268 31268
rect 13228 30892 13268 30932
rect 13516 31312 13556 31352
rect 13420 30472 13460 30512
rect 13132 29632 13172 29672
rect 12076 28288 12116 28328
rect 12268 28288 12308 28328
rect 12556 28288 12596 28328
rect 11980 28120 12020 28160
rect 11980 27784 12020 27824
rect 11788 27700 11828 27740
rect 11788 27364 11828 27404
rect 11884 27196 11924 27236
rect 11788 26524 11828 26564
rect 11788 24676 11828 24716
rect 11788 22660 11828 22700
rect 11692 22492 11732 22532
rect 12364 28120 12404 28160
rect 12268 28036 12308 28076
rect 12076 27280 12116 27320
rect 11980 27028 12020 27068
rect 11980 26776 12020 26816
rect 11980 25852 12020 25892
rect 12076 25600 12116 25640
rect 12556 28120 12596 28160
rect 12460 27868 12500 27908
rect 12460 27700 12500 27740
rect 12940 28708 12980 28748
rect 13132 28624 13172 28664
rect 12940 28288 12980 28328
rect 13228 28456 13268 28496
rect 13420 28792 13460 28832
rect 13420 28624 13460 28664
rect 13708 31480 13748 31520
rect 13708 31228 13748 31268
rect 13804 30724 13844 30764
rect 14380 36856 14420 36896
rect 14284 35932 14324 35972
rect 14284 35680 14324 35720
rect 14188 34336 14228 34376
rect 14092 34252 14132 34292
rect 13996 34000 14036 34040
rect 14284 33916 14324 33956
rect 14284 33664 14324 33704
rect 14188 33496 14228 33536
rect 14188 33076 14228 33116
rect 13996 32824 14036 32864
rect 14284 32908 14324 32948
rect 14188 32740 14228 32780
rect 14476 35596 14516 35636
rect 14572 35260 14612 35300
rect 14476 34588 14516 34628
rect 14764 37192 14804 37232
rect 14860 35596 14900 35636
rect 15436 37360 15476 37400
rect 15724 37528 15764 37568
rect 15052 37108 15092 37148
rect 15052 36520 15092 36560
rect 15628 37192 15668 37232
rect 15436 36520 15476 36560
rect 15244 36184 15284 36224
rect 15436 36100 15476 36140
rect 15148 35596 15188 35636
rect 15340 35596 15380 35636
rect 14956 35092 14996 35132
rect 15244 35092 15284 35132
rect 14956 34924 14996 34964
rect 15148 34924 15188 34964
rect 15052 34588 15092 34628
rect 14860 34168 14900 34208
rect 14380 32404 14420 32444
rect 15148 34168 15188 34208
rect 14764 33664 14804 33704
rect 14668 33496 14708 33536
rect 15244 33916 15284 33956
rect 15148 33244 15188 33284
rect 14668 32488 14708 32528
rect 13996 32152 14036 32192
rect 14572 32152 14612 32192
rect 14956 32656 14996 32696
rect 14764 32320 14804 32360
rect 14764 32152 14804 32192
rect 14284 32068 14324 32108
rect 15052 32152 15092 32192
rect 16204 38116 16244 38156
rect 16108 37780 16148 37820
rect 16108 37612 16148 37652
rect 16396 37948 16436 37988
rect 16300 37528 16340 37568
rect 16012 36688 16052 36728
rect 15724 36520 15764 36560
rect 16300 37360 16340 37400
rect 16588 38536 16628 38576
rect 17068 40300 17108 40340
rect 16972 39880 17012 39920
rect 16876 39040 16916 39080
rect 17068 39040 17108 39080
rect 16876 37444 16916 37484
rect 17356 40552 17396 40592
rect 18316 41308 18356 41348
rect 18124 40552 18164 40592
rect 17260 40384 17300 40424
rect 17356 40216 17396 40256
rect 17356 39292 17396 39332
rect 17740 39796 17780 39836
rect 18124 39712 18164 39752
rect 17932 39628 17972 39668
rect 18316 40972 18356 41012
rect 18316 40468 18356 40508
rect 18508 42064 18548 42104
rect 18892 42652 18932 42692
rect 18700 41896 18740 41936
rect 19276 42904 19316 42944
rect 19276 42232 19316 42272
rect 19084 41812 19124 41852
rect 18892 41140 18932 41180
rect 19564 42484 19604 42524
rect 19468 41644 19508 41684
rect 19372 41560 19412 41600
rect 18508 40636 18548 40676
rect 18412 40300 18452 40340
rect 18508 40048 18548 40088
rect 18316 39292 18356 39332
rect 17644 38788 17684 38828
rect 17836 38788 17876 38828
rect 17836 38620 17876 38660
rect 17740 38536 17780 38576
rect 17452 38032 17492 38072
rect 17740 38200 17780 38240
rect 17260 37444 17300 37484
rect 17068 37276 17108 37316
rect 16876 37192 16916 37232
rect 17164 37192 17204 37232
rect 16492 36940 16532 36980
rect 16396 36772 16436 36812
rect 16300 36688 16340 36728
rect 16204 36604 16244 36644
rect 15916 36352 15956 36392
rect 15724 36100 15764 36140
rect 15628 34924 15668 34964
rect 15532 34588 15572 34628
rect 15436 34252 15476 34292
rect 15628 33748 15668 33788
rect 15436 33496 15476 33536
rect 15340 32908 15380 32948
rect 15244 32740 15284 32780
rect 15628 33328 15668 33368
rect 16012 36268 16052 36308
rect 16108 35764 16148 35804
rect 16012 35260 16052 35300
rect 16108 34588 16148 34628
rect 15916 33412 15956 33452
rect 15820 33244 15860 33284
rect 15628 32824 15668 32864
rect 15820 32740 15860 32780
rect 15820 32488 15860 32528
rect 13996 31984 14036 32024
rect 14380 31984 14420 32024
rect 14956 31984 14996 32024
rect 14668 31900 14708 31940
rect 14476 31816 14516 31856
rect 13804 29884 13844 29924
rect 13708 29128 13748 29168
rect 13036 27784 13076 27824
rect 12364 25852 12404 25892
rect 12268 25432 12308 25472
rect 12364 25348 12404 25388
rect 11980 25180 12020 25220
rect 12364 25096 12404 25136
rect 12940 27448 12980 27488
rect 12652 27112 12692 27152
rect 12556 26188 12596 26228
rect 12556 25516 12596 25556
rect 12556 25180 12596 25220
rect 12364 24508 12404 24548
rect 12556 23836 12596 23876
rect 12940 27028 12980 27068
rect 12748 26776 12788 26816
rect 12844 26188 12884 26228
rect 13132 27616 13172 27656
rect 13324 26776 13364 26816
rect 13228 26524 13268 26564
rect 12748 25768 12788 25808
rect 12940 25348 12980 25388
rect 12748 25264 12788 25304
rect 13420 25012 13460 25052
rect 12076 23164 12116 23204
rect 11884 22324 11924 22364
rect 11788 22156 11828 22196
rect 11692 22072 11732 22112
rect 11596 21988 11636 22028
rect 11884 21736 11924 21776
rect 11692 21400 11732 21440
rect 12652 23752 12692 23792
rect 12652 22744 12692 22784
rect 12268 22324 12308 22364
rect 12268 21568 12308 21608
rect 13228 24508 13268 24548
rect 13612 27448 13652 27488
rect 13612 26524 13652 26564
rect 13228 24256 13268 24296
rect 13228 24004 13268 24044
rect 13036 23920 13076 23960
rect 13612 24256 13652 24296
rect 13900 26860 13940 26900
rect 13996 26608 14036 26648
rect 13900 26440 13940 26480
rect 13996 26188 14036 26228
rect 13900 25684 13940 25724
rect 13900 25432 13940 25472
rect 13804 25012 13844 25052
rect 13996 25180 14036 25220
rect 13900 24424 13940 24464
rect 13804 23836 13844 23876
rect 13324 23248 13364 23288
rect 13132 22996 13172 23036
rect 13228 22660 13268 22700
rect 12940 22324 12980 22364
rect 13132 22324 13172 22364
rect 12940 22072 12980 22112
rect 12844 21820 12884 21860
rect 12652 21316 12692 21356
rect 12652 20812 12692 20852
rect 12748 20644 12788 20684
rect 11692 20560 11732 20600
rect 12076 20560 12116 20600
rect 12556 20560 12596 20600
rect 11500 20476 11540 20516
rect 12652 20224 12692 20264
rect 11116 20056 11156 20096
rect 11500 20091 11540 20096
rect 11500 20056 11540 20091
rect 11980 20056 12020 20096
rect 11212 19804 11252 19844
rect 11692 19804 11732 19844
rect 11500 19720 11540 19760
rect 11212 19468 11252 19508
rect 11692 19552 11732 19592
rect 11596 19300 11636 19340
rect 10924 18544 10964 18584
rect 10924 17788 10964 17828
rect 10828 17704 10868 17744
rect 10828 17536 10868 17576
rect 10732 17116 10772 17156
rect 11020 17536 11060 17576
rect 10924 17032 10964 17072
rect 10636 15940 10676 15980
rect 10444 15520 10484 15560
rect 10348 15100 10388 15140
rect 10540 15100 10580 15140
rect 10348 14848 10388 14888
rect 10444 14596 10484 14636
rect 10156 14176 10196 14216
rect 10060 13840 10100 13880
rect 9964 12496 10004 12536
rect 9676 12244 9716 12284
rect 9580 12076 9620 12116
rect 9676 11992 9716 12032
rect 9004 11572 9044 11612
rect 9196 11572 9236 11612
rect 9100 11068 9140 11108
rect 8812 10732 8852 10772
rect 9100 10732 9140 10772
rect 9004 10396 9044 10436
rect 9292 11068 9332 11108
rect 9004 10144 9044 10184
rect 8812 9388 8852 9428
rect 8716 8632 8756 8672
rect 8716 8212 8756 8252
rect 8620 8044 8660 8084
rect 8716 7708 8756 7748
rect 8716 7288 8756 7328
rect 8524 7204 8564 7244
rect 8428 6616 8468 6656
rect 8332 6532 8372 6572
rect 7948 3760 7988 3800
rect 8044 3424 8084 3464
rect 7948 3172 7988 3212
rect 7852 3088 7892 3128
rect 7756 2752 7796 2792
rect 8428 6448 8468 6488
rect 8428 6028 8468 6068
rect 8428 5692 8468 5732
rect 9484 11572 9524 11612
rect 9100 9892 9140 9932
rect 9196 9388 9236 9428
rect 9004 8800 9044 8840
rect 9196 8716 9236 8756
rect 9100 8632 9140 8672
rect 9004 8128 9044 8168
rect 8908 8044 8948 8084
rect 8908 7876 8948 7916
rect 9772 11656 9812 11696
rect 9964 11488 10004 11528
rect 9772 11404 9812 11444
rect 9964 11236 10004 11276
rect 9292 8548 9332 8588
rect 9580 9472 9620 9512
rect 10156 13504 10196 13544
rect 10348 14344 10388 14384
rect 11404 18376 11444 18416
rect 11788 18544 11828 18584
rect 11788 18124 11828 18164
rect 11692 17956 11732 17996
rect 11596 17788 11636 17828
rect 11500 17620 11540 17660
rect 11404 16864 11444 16904
rect 11308 16780 11348 16820
rect 11020 16360 11060 16400
rect 10636 14932 10676 14972
rect 11116 15184 11156 15224
rect 10540 14008 10580 14048
rect 10540 13840 10580 13880
rect 10348 13588 10388 13628
rect 11020 14848 11060 14888
rect 10924 14764 10964 14804
rect 10828 14344 10868 14384
rect 11500 16360 11540 16400
rect 11404 16276 11444 16316
rect 11500 15856 11540 15896
rect 11500 15688 11540 15728
rect 12268 20056 12308 20096
rect 12460 19804 12500 19844
rect 12364 19636 12404 19676
rect 12268 18880 12308 18920
rect 12172 18712 12212 18752
rect 11788 15856 11828 15896
rect 11692 15688 11732 15728
rect 11596 15520 11636 15560
rect 11500 15352 11540 15392
rect 11404 14932 11444 14972
rect 11308 14764 11348 14804
rect 10924 14260 10964 14300
rect 11116 14260 11156 14300
rect 10732 14092 10772 14132
rect 12460 18208 12500 18248
rect 13036 20728 13076 20768
rect 13324 22324 13364 22364
rect 13228 21652 13268 21692
rect 12844 19216 12884 19256
rect 12748 18796 12788 18836
rect 12652 18208 12692 18248
rect 12556 18124 12596 18164
rect 12460 17368 12500 17408
rect 12844 17620 12884 17660
rect 13324 21400 13364 21440
rect 13228 20308 13268 20348
rect 13228 20140 13268 20180
rect 13132 19636 13172 19676
rect 13324 19972 13364 20012
rect 13516 23080 13556 23120
rect 13996 24004 14036 24044
rect 13900 23752 13940 23792
rect 13996 23668 14036 23708
rect 13612 22660 13652 22700
rect 13516 22492 13556 22532
rect 13612 22408 13652 22448
rect 13516 21820 13556 21860
rect 13900 22156 13940 22196
rect 13996 21736 14036 21776
rect 13900 21652 13940 21692
rect 14188 30640 14228 30680
rect 14476 30640 14516 30680
rect 14572 29800 14612 29840
rect 14380 29128 14420 29168
rect 14284 28708 14324 28748
rect 14380 28288 14420 28328
rect 14284 27448 14324 27488
rect 14572 27532 14612 27572
rect 14476 27196 14516 27236
rect 14380 26524 14420 26564
rect 14380 25852 14420 25892
rect 14764 31816 14804 31856
rect 14860 31228 14900 31268
rect 14860 30892 14900 30932
rect 14956 30220 14996 30260
rect 14764 30052 14804 30092
rect 14956 29884 14996 29924
rect 14764 29212 14804 29252
rect 14860 29128 14900 29168
rect 15148 31480 15188 31520
rect 15436 31984 15476 32024
rect 15244 31312 15284 31352
rect 15340 31228 15380 31268
rect 15148 30556 15188 30596
rect 15052 29800 15092 29840
rect 14764 28288 14804 28328
rect 14764 27952 14804 27992
rect 15532 31900 15572 31940
rect 15532 31480 15572 31520
rect 15532 30976 15572 31016
rect 15436 30640 15476 30680
rect 15724 32152 15764 32192
rect 16300 36352 16340 36392
rect 16972 36688 17012 36728
rect 17068 36604 17108 36644
rect 16780 36352 16820 36392
rect 17260 37108 17300 37148
rect 17836 37612 17876 37652
rect 19084 40972 19124 41012
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 19180 40636 19220 40676
rect 19468 41392 19508 41432
rect 19756 42316 19796 42356
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 19852 41476 19892 41516
rect 21388 41392 21428 41432
rect 19660 41140 19700 41180
rect 19756 41056 19796 41096
rect 18988 40552 19028 40592
rect 18700 40216 18740 40256
rect 18892 40132 18932 40172
rect 18700 39880 18740 39920
rect 19468 39964 19508 40004
rect 19084 39796 19124 39836
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18123 38956 18163 38996
rect 18508 38956 18548 38996
rect 18412 38704 18452 38744
rect 18316 38620 18356 38660
rect 18604 38620 18644 38660
rect 18892 39040 18932 39080
rect 18796 38872 18836 38912
rect 18412 38536 18452 38576
rect 18700 38536 18740 38576
rect 18604 38368 18644 38408
rect 18508 38200 18548 38240
rect 19180 38956 19220 38996
rect 18891 38284 18931 38324
rect 19084 38284 19124 38324
rect 19276 38872 19316 38912
rect 19276 38704 19316 38744
rect 19276 38368 19316 38408
rect 20044 41140 20084 41180
rect 19948 40888 19988 40928
rect 20140 40300 20180 40340
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 19660 39628 19700 39668
rect 19564 39208 19604 39248
rect 20044 39628 20084 39668
rect 19468 38956 19508 38996
rect 19564 38872 19604 38912
rect 20044 38788 20084 38828
rect 19564 38368 19604 38408
rect 19372 38200 19412 38240
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 19084 37948 19124 37988
rect 18412 37864 18452 37904
rect 17932 37528 17972 37568
rect 18316 37612 18356 37652
rect 17452 37192 17492 37232
rect 17356 36772 17396 36812
rect 17644 36772 17684 36812
rect 17260 36520 17300 36560
rect 17164 36184 17204 36224
rect 16780 36100 16820 36140
rect 16972 36100 17012 36140
rect 16492 36016 16532 36056
rect 16396 35764 16436 35804
rect 16300 34000 16340 34040
rect 16300 33244 16340 33284
rect 16300 32824 16340 32864
rect 16492 33916 16532 33956
rect 16300 32572 16340 32612
rect 16012 32320 16052 32360
rect 16204 32320 16244 32360
rect 15724 31480 15764 31520
rect 15628 30052 15668 30092
rect 15628 29800 15668 29840
rect 15340 29296 15380 29336
rect 15340 28960 15380 29000
rect 15052 28288 15092 28328
rect 15148 28120 15188 28160
rect 15340 27952 15380 27992
rect 15532 29296 15572 29336
rect 15532 29044 15572 29084
rect 15628 28876 15668 28916
rect 15340 26860 15380 26900
rect 14956 26188 14996 26228
rect 14764 25852 14804 25892
rect 14668 25516 14708 25556
rect 14284 25432 14324 25472
rect 14476 25348 14516 25388
rect 14284 24424 14324 24464
rect 14188 23080 14228 23120
rect 14188 22492 14228 22532
rect 14572 25264 14612 25304
rect 15244 26440 15284 26480
rect 15244 25516 15284 25556
rect 15148 25180 15188 25220
rect 14956 24760 14996 24800
rect 14380 23920 14420 23960
rect 14284 22408 14324 22448
rect 14284 22240 14324 22280
rect 14188 22156 14228 22196
rect 13708 20812 13748 20852
rect 13612 20140 13652 20180
rect 13612 19972 13652 20012
rect 13612 19636 13652 19676
rect 13516 19468 13556 19508
rect 13324 19132 13364 19172
rect 13324 18796 13364 18836
rect 13228 18712 13268 18752
rect 13036 18208 13076 18248
rect 13228 18208 13268 18248
rect 13132 18124 13172 18164
rect 13036 17620 13076 17660
rect 13420 18124 13460 18164
rect 13420 17956 13460 17996
rect 13228 17872 13268 17912
rect 13324 17620 13364 17660
rect 12364 16780 12404 16820
rect 12268 16108 12308 16148
rect 12172 15688 12212 15728
rect 11884 15436 11924 15476
rect 11788 15268 11828 15308
rect 11980 15100 12020 15140
rect 11596 14848 11636 14888
rect 11308 14596 11348 14636
rect 11596 14428 11636 14468
rect 11404 14260 11444 14300
rect 10732 13840 10772 13880
rect 10540 13168 10580 13208
rect 11116 14008 11156 14048
rect 11212 13924 11252 13964
rect 11116 13756 11156 13796
rect 10156 12664 10196 12704
rect 10252 12580 10292 12620
rect 10156 12412 10196 12452
rect 10252 12328 10292 12368
rect 10252 11236 10292 11276
rect 10444 10900 10484 10940
rect 10252 10060 10292 10100
rect 10060 9976 10100 10016
rect 10156 9892 10196 9932
rect 9868 9556 9908 9596
rect 9580 9052 9620 9092
rect 9484 8212 9524 8252
rect 9868 9220 9908 9260
rect 10060 9472 10100 9512
rect 9772 8548 9812 8588
rect 9676 8296 9716 8336
rect 9772 8212 9812 8252
rect 9676 8044 9716 8084
rect 9100 7456 9140 7496
rect 9004 7372 9044 7412
rect 8908 7288 8948 7328
rect 9004 7120 9044 7160
rect 8908 6952 8948 6992
rect 8620 6616 8660 6656
rect 8812 6364 8852 6404
rect 8620 6028 8660 6068
rect 8524 5608 8564 5648
rect 8236 5104 8276 5144
rect 8332 4852 8372 4892
rect 8140 2584 8180 2624
rect 8428 3760 8468 3800
rect 8908 5944 8948 5984
rect 9580 7708 9620 7748
rect 9388 7540 9428 7580
rect 9196 6448 9236 6488
rect 9484 7372 9524 7412
rect 9580 7288 9620 7328
rect 9964 8632 10004 8672
rect 9964 8296 10004 8336
rect 10156 9052 10196 9092
rect 10348 9220 10388 9260
rect 10348 9052 10388 9092
rect 10348 8884 10388 8924
rect 11308 12832 11348 12872
rect 11884 14176 11924 14216
rect 11788 14092 11828 14132
rect 11500 14008 11540 14048
rect 11980 14008 12020 14048
rect 12268 15268 12308 15308
rect 12364 14260 12404 14300
rect 12364 14008 12404 14048
rect 11596 13840 11636 13880
rect 12652 17200 12692 17240
rect 12556 16948 12596 16988
rect 12940 16696 12980 16736
rect 12844 16612 12884 16652
rect 12748 14680 12788 14720
rect 12844 14596 12884 14636
rect 12652 14512 12692 14552
rect 12556 14428 12596 14468
rect 12556 14260 12596 14300
rect 12844 14260 12884 14300
rect 13612 18460 13652 18500
rect 13612 18292 13652 18332
rect 13708 18124 13748 18164
rect 13708 17620 13748 17660
rect 13612 17452 13652 17492
rect 13996 21232 14036 21272
rect 14092 20476 14132 20516
rect 13996 20224 14036 20264
rect 13996 19972 14036 20012
rect 13996 19300 14036 19340
rect 14284 21736 14324 21776
rect 14284 21148 14324 21188
rect 14284 20812 14324 20852
rect 14284 19468 14324 19508
rect 13996 18796 14036 18836
rect 13996 17956 14036 17996
rect 13900 17116 13940 17156
rect 13708 16612 13748 16652
rect 14572 22744 14612 22784
rect 15148 24592 15188 24632
rect 14764 24424 14804 24464
rect 14764 23920 14804 23960
rect 14860 23752 14900 23792
rect 14764 23416 14804 23456
rect 15148 23500 15188 23540
rect 15532 27028 15572 27068
rect 15052 22492 15092 22532
rect 14764 21820 14804 21860
rect 14764 21484 14804 21524
rect 14668 21232 14708 21272
rect 14764 20560 14804 20600
rect 14764 20140 14804 20180
rect 14572 19216 14612 19256
rect 15244 22996 15284 23036
rect 15916 31312 15956 31352
rect 15820 31228 15860 31268
rect 15820 30724 15860 30764
rect 16876 35680 16916 35720
rect 16684 35176 16724 35216
rect 16684 34252 16724 34292
rect 18124 37276 18164 37316
rect 17836 36940 17876 36980
rect 18220 37024 18260 37064
rect 18124 36856 18164 36896
rect 18028 36772 18068 36812
rect 17644 35680 17684 35720
rect 17164 35260 17204 35300
rect 17068 34756 17108 34796
rect 16972 34252 17012 34292
rect 17164 34252 17204 34292
rect 16876 34168 16916 34208
rect 16876 32992 16916 33032
rect 16780 32824 16820 32864
rect 16684 32740 16724 32780
rect 16588 32572 16628 32612
rect 16396 32488 16436 32528
rect 16396 32068 16436 32108
rect 16108 31228 16148 31268
rect 16684 31564 16724 31604
rect 16300 31480 16340 31520
rect 16492 31312 16532 31352
rect 15916 30052 15956 30092
rect 16108 30388 16148 30428
rect 15916 29548 15956 29588
rect 15820 29212 15860 29252
rect 15820 28204 15860 28244
rect 16012 29128 16052 29168
rect 16780 31312 16820 31352
rect 17068 33076 17108 33116
rect 16972 32404 17012 32444
rect 17068 32152 17108 32192
rect 17452 35176 17492 35216
rect 17548 34336 17588 34376
rect 17548 34168 17588 34208
rect 17644 33916 17684 33956
rect 17644 33664 17684 33704
rect 17356 33496 17396 33536
rect 17548 33496 17588 33536
rect 17932 35512 17972 35552
rect 17932 34420 17972 34460
rect 18028 34084 18068 34124
rect 18028 33496 18068 33536
rect 17740 33244 17780 33284
rect 17452 32572 17492 32612
rect 17548 32404 17588 32444
rect 16972 31900 17012 31940
rect 17068 31732 17108 31772
rect 16684 31228 16724 31268
rect 16684 30052 16724 30092
rect 16588 29800 16628 29840
rect 16876 29884 16916 29924
rect 17164 30976 17204 31016
rect 17452 31900 17492 31940
rect 19564 38116 19604 38156
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 19276 37780 19316 37820
rect 19756 37612 19796 37652
rect 19180 37528 19220 37568
rect 18412 36856 18452 36896
rect 18892 37192 18932 37232
rect 19084 37024 19124 37064
rect 18508 36688 18548 36728
rect 18412 36604 18452 36644
rect 18316 36520 18356 36560
rect 19468 37360 19508 37400
rect 19660 37360 19700 37400
rect 19276 36856 19316 36896
rect 19180 36772 19220 36812
rect 19660 37024 19700 37064
rect 19564 36688 19604 36728
rect 19468 36604 19508 36644
rect 18892 36520 18932 36560
rect 18700 36436 18740 36476
rect 18604 36268 18644 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 18700 36184 18740 36224
rect 18604 35932 18644 35972
rect 18412 35512 18452 35552
rect 18316 35176 18356 35216
rect 18412 34672 18452 34712
rect 18316 34252 18356 34292
rect 19468 36100 19508 36140
rect 18988 36016 19028 36056
rect 19180 35260 19220 35300
rect 18892 35176 18932 35216
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18700 34504 18740 34544
rect 18412 33076 18452 33116
rect 17932 32320 17972 32360
rect 17836 32152 17876 32192
rect 17356 30556 17396 30596
rect 17548 30724 17588 30764
rect 17356 30388 17396 30428
rect 17164 29884 17204 29924
rect 16396 29296 16436 29336
rect 16588 29128 16628 29168
rect 16108 28540 16148 28580
rect 16108 28204 16148 28244
rect 15724 27028 15764 27068
rect 15916 26860 15956 26900
rect 15724 26608 15764 26648
rect 15436 25180 15476 25220
rect 15628 24508 15668 24548
rect 15724 23836 15764 23876
rect 15436 22744 15476 22784
rect 15628 22996 15668 23036
rect 15532 22660 15572 22700
rect 15148 21484 15188 21524
rect 15052 20224 15092 20264
rect 15532 22156 15572 22196
rect 15532 21652 15572 21692
rect 15532 20728 15572 20768
rect 16300 28288 16340 28328
rect 16300 27028 16340 27068
rect 16204 26356 16244 26396
rect 16012 25600 16052 25640
rect 15916 23164 15956 23204
rect 16204 23668 16244 23708
rect 16108 22912 16148 22952
rect 15916 22828 15956 22868
rect 15820 22324 15860 22364
rect 15916 21904 15956 21944
rect 16204 21316 16244 21356
rect 15724 21064 15764 21104
rect 15628 20560 15668 20600
rect 15244 20140 15284 20180
rect 14956 19216 14996 19256
rect 14764 18964 14804 19004
rect 14956 19048 14996 19088
rect 15148 19804 15188 19844
rect 15148 19384 15188 19424
rect 15052 18796 15092 18836
rect 14284 18544 14324 18584
rect 14668 18544 14708 18584
rect 14476 18208 14516 18248
rect 14380 17872 14420 17912
rect 14764 17956 14804 17996
rect 14572 17788 14612 17828
rect 14956 18460 14996 18500
rect 15052 18292 15092 18332
rect 13900 16864 13940 16904
rect 13516 16192 13556 16232
rect 13420 15772 13460 15812
rect 13804 15772 13844 15812
rect 13324 15688 13364 15728
rect 13132 15604 13172 15644
rect 13036 15520 13076 15560
rect 13132 15184 13172 15224
rect 13420 15604 13460 15644
rect 13132 14680 13172 14720
rect 13036 14512 13076 14552
rect 12940 14092 12980 14132
rect 12844 14008 12884 14048
rect 12556 13840 12596 13880
rect 12460 13672 12500 13712
rect 11788 13420 11828 13460
rect 11596 13000 11636 13040
rect 11980 12832 12020 12872
rect 10732 12496 10772 12536
rect 10828 12412 10868 12452
rect 11020 12412 11060 12452
rect 11212 12451 11252 12452
rect 11212 12412 11252 12451
rect 10924 11740 10964 11780
rect 10732 11656 10772 11696
rect 10732 10816 10772 10856
rect 10540 10144 10580 10184
rect 10636 9556 10676 9596
rect 10636 9052 10676 9092
rect 10156 8548 10196 8588
rect 10444 8548 10484 8588
rect 10636 8632 10676 8672
rect 10540 8296 10580 8336
rect 10156 8212 10196 8252
rect 10444 7960 10484 8000
rect 10060 7624 10100 7664
rect 10156 7456 10196 7496
rect 10060 6868 10100 6908
rect 10540 7288 10580 7328
rect 11308 11908 11348 11948
rect 11596 12076 11636 12116
rect 11500 11992 11540 12032
rect 11212 11572 11252 11612
rect 11404 11488 11444 11528
rect 11212 11236 11252 11276
rect 11020 11068 11060 11108
rect 11308 11152 11348 11192
rect 11596 11656 11636 11696
rect 11500 10900 11540 10940
rect 11596 10816 11636 10856
rect 11308 10732 11348 10772
rect 11020 10312 11060 10352
rect 11020 10144 11060 10184
rect 10924 10060 10964 10100
rect 11884 12412 11924 12452
rect 11980 12244 12020 12284
rect 11980 11992 12020 12032
rect 11980 11572 12020 11612
rect 12268 13168 12308 13208
rect 13036 13756 13076 13796
rect 12652 13672 12692 13712
rect 12172 13000 12212 13040
rect 12172 12832 12212 12872
rect 12172 12580 12212 12620
rect 12172 11572 12212 11612
rect 12076 11488 12116 11528
rect 11788 11152 11828 11192
rect 12076 11152 12116 11192
rect 13036 13168 13076 13208
rect 12844 13000 12884 13040
rect 12940 12832 12980 12872
rect 12748 12496 12788 12536
rect 12652 11908 12692 11948
rect 12844 11908 12884 11948
rect 12556 11488 12596 11528
rect 12364 10816 12404 10856
rect 11692 10648 11732 10688
rect 11308 10480 11348 10520
rect 11980 10480 12020 10520
rect 11404 10312 11444 10352
rect 12364 10396 12404 10436
rect 10828 9724 10868 9764
rect 11020 9640 11060 9680
rect 10828 8632 10868 8672
rect 11116 8632 11156 8672
rect 11020 8128 11060 8168
rect 11212 8044 11252 8084
rect 10156 6784 10196 6824
rect 9676 6616 9716 6656
rect 10636 7036 10676 7076
rect 10444 6448 10484 6488
rect 10060 6196 10100 6236
rect 10156 5944 10196 5984
rect 10348 5944 10388 5984
rect 9868 5860 9908 5900
rect 9484 5272 9524 5312
rect 9676 5188 9716 5228
rect 9388 5104 9428 5144
rect 9004 4936 9044 4976
rect 9196 4852 9236 4892
rect 8908 4264 8948 4304
rect 9004 4096 9044 4136
rect 9292 4600 9332 4640
rect 8620 3844 8660 3884
rect 8428 2668 8468 2708
rect 9004 3340 9044 3380
rect 8620 2500 8660 2540
rect 7852 2416 7892 2456
rect 7660 2164 7700 2204
rect 7852 1912 7892 1952
rect 7756 1240 7796 1280
rect 7372 904 7412 944
rect 7564 904 7604 944
rect 8236 1324 8276 1364
rect 8140 1240 8180 1280
rect 8044 988 8084 1028
rect 7948 820 7988 860
rect 7852 568 7892 608
rect 8332 1240 8372 1280
rect 8236 988 8276 1028
rect 8721 2500 8761 2540
rect 8524 1912 8564 1952
rect 8524 1240 8564 1280
rect 8428 1156 8468 1196
rect 8812 2164 8852 2204
rect 8812 1408 8852 1448
rect 9196 3424 9236 3464
rect 9580 4936 9620 4976
rect 9484 4852 9524 4892
rect 9292 2752 9332 2792
rect 9964 4936 10004 4976
rect 9772 4600 9812 4640
rect 10060 4432 10100 4472
rect 9580 4264 9620 4304
rect 9676 3844 9716 3884
rect 9772 3340 9812 3380
rect 9772 2584 9812 2624
rect 9676 2164 9716 2204
rect 9580 2080 9620 2120
rect 9292 1156 9332 1196
rect 8908 988 8948 1028
rect 8812 652 8852 692
rect 8908 316 8948 356
rect 9772 1912 9812 1952
rect 9772 1744 9812 1784
rect 9772 1324 9812 1364
rect 9484 904 9524 944
rect 9292 652 9332 692
rect 10444 5608 10484 5648
rect 10156 4096 10196 4136
rect 9964 2500 10004 2540
rect 9964 2080 10004 2120
rect 9964 1072 10004 1112
rect 9772 148 9812 188
rect 10348 5356 10388 5396
rect 10444 5272 10484 5312
rect 10540 5020 10580 5060
rect 11596 10144 11636 10184
rect 11788 10060 11828 10100
rect 11980 9976 12020 10016
rect 11500 9640 11540 9680
rect 11404 9052 11444 9092
rect 11884 9220 11924 9260
rect 11500 8464 11540 8504
rect 11404 8212 11444 8252
rect 11404 7876 11444 7916
rect 11308 7540 11348 7580
rect 11692 8548 11732 8588
rect 11884 8548 11924 8588
rect 11785 8464 11825 8504
rect 12652 10312 12692 10352
rect 12460 10144 12500 10184
rect 12563 10144 12596 10184
rect 12596 10144 12603 10184
rect 12364 9976 12404 10016
rect 12076 9640 12116 9680
rect 12268 9640 12308 9680
rect 13132 13000 13172 13040
rect 13132 12580 13172 12620
rect 13708 15520 13748 15560
rect 13612 15352 13652 15392
rect 13612 14008 13652 14048
rect 13612 13840 13652 13880
rect 14092 16864 14132 16904
rect 14476 17620 14516 17660
rect 14860 17452 14900 17492
rect 15052 17284 15092 17324
rect 14284 16612 14324 16652
rect 13996 16024 14036 16064
rect 13996 15436 14036 15476
rect 13900 14680 13940 14720
rect 13996 14596 14036 14636
rect 13996 13924 14036 13964
rect 13900 13840 13940 13880
rect 13516 12832 13556 12872
rect 13324 12748 13364 12788
rect 13612 12580 13652 12620
rect 13324 11908 13364 11948
rect 13420 11824 13460 11864
rect 13036 10984 13076 11024
rect 12844 10312 12884 10352
rect 12844 10060 12884 10100
rect 12940 9892 12980 9932
rect 12940 9724 12980 9764
rect 12748 9640 12788 9680
rect 12172 9388 12212 9428
rect 12268 9220 12308 9260
rect 12172 9052 12212 9092
rect 11692 8296 11732 8336
rect 11980 8296 12020 8336
rect 11692 8128 11732 8168
rect 11980 8044 12020 8084
rect 11884 7960 11924 8000
rect 11692 7792 11732 7832
rect 11596 7036 11636 7076
rect 11212 6784 11252 6824
rect 11212 6448 11252 6488
rect 10924 5104 10964 5144
rect 11116 5020 11156 5060
rect 10348 3760 10388 3800
rect 10156 3424 10196 3464
rect 10348 3424 10388 3464
rect 10348 2332 10388 2372
rect 10252 2080 10292 2120
rect 10252 1660 10292 1700
rect 10156 988 10196 1028
rect 10924 4516 10964 4556
rect 10828 4264 10868 4304
rect 10924 4096 10964 4136
rect 11500 6700 11540 6740
rect 11308 5188 11348 5228
rect 11308 4852 11348 4892
rect 11692 6700 11732 6740
rect 11692 6364 11732 6404
rect 11692 5440 11732 5480
rect 12076 7960 12116 8000
rect 12364 9052 12404 9092
rect 12268 8716 12308 8756
rect 12268 8044 12308 8084
rect 12460 8884 12500 8924
rect 12652 9388 12692 9428
rect 14092 13672 14132 13712
rect 14284 15520 14324 15560
rect 14276 15016 14316 15056
rect 14476 16948 14516 16988
rect 14764 16192 14804 16232
rect 14956 16024 14996 16064
rect 15244 17704 15284 17744
rect 15436 20056 15476 20096
rect 15436 19300 15476 19340
rect 15340 16612 15380 16652
rect 15148 16276 15188 16316
rect 15532 18880 15572 18920
rect 15916 20812 15956 20852
rect 16012 20560 16052 20600
rect 15724 19300 15764 19340
rect 15916 19972 15956 20012
rect 15820 19216 15860 19256
rect 15628 17620 15668 17660
rect 15724 17116 15764 17156
rect 15820 17032 15860 17072
rect 16012 19804 16052 19844
rect 16204 20728 16244 20768
rect 16204 20308 16244 20348
rect 16204 19720 16244 19760
rect 16684 28120 16724 28160
rect 16588 26776 16628 26816
rect 16492 26440 16532 26480
rect 16396 26356 16436 26396
rect 16588 26188 16628 26228
rect 16684 26020 16724 26060
rect 16396 24256 16436 24296
rect 17068 29128 17108 29168
rect 17740 30388 17780 30428
rect 17644 30220 17684 30260
rect 17740 30052 17780 30092
rect 18028 31984 18068 32024
rect 18220 32152 18260 32192
rect 18124 31396 18164 31436
rect 18124 31144 18164 31184
rect 17932 30724 17972 30764
rect 17452 29212 17492 29252
rect 17548 29128 17588 29168
rect 17548 28876 17588 28916
rect 17164 27700 17204 27740
rect 16972 26776 17012 26816
rect 16972 26356 17012 26396
rect 17644 28288 17684 28328
rect 17356 27784 17396 27824
rect 17548 27784 17588 27824
rect 17164 26944 17204 26984
rect 17164 26356 17204 26396
rect 17068 26272 17108 26312
rect 17260 25852 17300 25892
rect 17836 28204 17876 28244
rect 17740 28120 17780 28160
rect 17836 27448 17876 27488
rect 17452 27364 17492 27404
rect 18028 29464 18068 29504
rect 17932 27196 17972 27236
rect 17452 26944 17492 26984
rect 17548 26692 17588 26732
rect 17356 25768 17396 25808
rect 17740 26356 17780 26396
rect 17644 26188 17684 26228
rect 17644 25768 17684 25808
rect 17164 25096 17204 25136
rect 17356 25096 17396 25136
rect 17260 24760 17300 24800
rect 16684 24256 16724 24296
rect 16492 23416 16532 23456
rect 17164 24508 17204 24548
rect 16780 23332 16820 23372
rect 17260 23757 17300 23792
rect 17260 23752 17300 23757
rect 17452 24676 17492 24716
rect 17836 25852 17876 25892
rect 17740 25600 17780 25640
rect 17740 25348 17780 25388
rect 18028 26776 18068 26816
rect 18220 30724 18260 30764
rect 18220 30472 18260 30512
rect 18220 28708 18260 28748
rect 18604 33664 18644 33704
rect 18604 33496 18644 33536
rect 19084 34168 19124 34208
rect 19372 35932 19412 35972
rect 19564 35680 19604 35720
rect 20236 37780 20276 37820
rect 19948 37360 19988 37400
rect 20044 37276 20084 37316
rect 19948 37192 19988 37232
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 19948 36940 19988 36980
rect 19852 36772 19892 36812
rect 19756 36100 19796 36140
rect 19468 35008 19508 35048
rect 19372 33832 19412 33872
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 19468 33580 19508 33620
rect 18892 32908 18932 32948
rect 19084 32824 19124 32864
rect 19660 34840 19700 34880
rect 20236 35764 20276 35804
rect 19852 35512 19892 35552
rect 19852 35092 19892 35132
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 19948 34504 19988 34544
rect 19852 34252 19892 34292
rect 20140 34168 20180 34208
rect 19756 33832 19796 33872
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 19756 33160 19796 33200
rect 19660 32992 19700 33032
rect 19372 32740 19412 32780
rect 18604 32488 18644 32528
rect 18412 31564 18452 31604
rect 18412 31396 18452 31436
rect 18604 32236 18644 32276
rect 18604 31816 18644 31856
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18796 31564 18836 31604
rect 18700 31480 18740 31520
rect 18604 31228 18644 31268
rect 18892 31396 18932 31436
rect 18508 30724 18548 30764
rect 18220 28204 18260 28244
rect 18412 27196 18452 27236
rect 18316 25684 18356 25724
rect 17740 25180 17780 25220
rect 17932 25180 17972 25220
rect 17836 25096 17876 25136
rect 17932 24256 17972 24296
rect 17740 23668 17780 23708
rect 17740 23500 17780 23540
rect 16876 22660 16916 22700
rect 16588 22240 16628 22280
rect 16780 22240 16820 22280
rect 16492 20728 16532 20768
rect 16396 20644 16436 20684
rect 16396 20392 16436 20432
rect 16492 20308 16532 20348
rect 16300 19384 16340 19424
rect 16396 18880 16436 18920
rect 16300 18712 16340 18752
rect 16204 18544 16244 18584
rect 16108 18376 16148 18416
rect 16300 17956 16340 17996
rect 16972 21484 17012 21524
rect 16972 20896 17012 20936
rect 17164 22492 17204 22532
rect 17164 22240 17204 22280
rect 17164 21568 17204 21608
rect 16876 20728 16916 20768
rect 16780 20476 16820 20516
rect 16684 20224 16724 20264
rect 16588 19552 16628 19592
rect 16684 19132 16724 19172
rect 16588 18796 16628 18836
rect 17356 23080 17396 23120
rect 17356 22156 17396 22196
rect 17548 22072 17588 22112
rect 17644 21736 17684 21776
rect 17356 21400 17396 21440
rect 17260 20476 17300 20516
rect 17260 20224 17300 20264
rect 16876 20056 16916 20096
rect 17260 19552 17300 19592
rect 16972 19300 17012 19340
rect 16876 19216 16916 19256
rect 16492 18376 16532 18416
rect 16300 17704 16340 17744
rect 16108 17536 16148 17576
rect 15628 16444 15668 16484
rect 15244 15940 15284 15980
rect 15052 15772 15092 15812
rect 14764 15688 14804 15728
rect 14860 15268 14900 15308
rect 14764 15100 14804 15140
rect 14572 15016 14612 15056
rect 14668 14848 14708 14888
rect 14092 12832 14132 12872
rect 13996 12580 14036 12620
rect 13804 12496 13844 12536
rect 13804 11404 13844 11444
rect 13708 11320 13748 11360
rect 13324 11236 13364 11276
rect 13612 11152 13652 11192
rect 13324 11068 13364 11108
rect 13324 10144 13364 10184
rect 13228 9892 13268 9932
rect 13228 9724 13268 9764
rect 13516 9556 13556 9596
rect 13324 9388 13364 9428
rect 12652 9052 12692 9092
rect 12556 8128 12596 8168
rect 12460 7960 12500 8000
rect 13420 8968 13460 9008
rect 12748 8716 12788 8756
rect 13324 8716 13364 8756
rect 12748 8464 12788 8504
rect 12844 8380 12884 8420
rect 13708 10732 13748 10772
rect 13708 10228 13748 10268
rect 13900 11236 13940 11276
rect 13804 10060 13844 10100
rect 13708 9892 13748 9932
rect 13420 8632 13460 8672
rect 13036 8548 13076 8588
rect 13612 8632 13652 8672
rect 13612 8464 13652 8504
rect 12268 7624 12308 7664
rect 12076 7456 12116 7496
rect 12364 7540 12404 7580
rect 12268 7120 12308 7160
rect 12172 6952 12212 6992
rect 12076 6364 12116 6404
rect 12172 6280 12212 6320
rect 11980 5608 12020 5648
rect 12172 5524 12212 5564
rect 11884 4936 11924 4976
rect 11500 4852 11540 4892
rect 11404 4516 11444 4556
rect 11308 4264 11348 4304
rect 11212 4180 11252 4220
rect 11404 4096 11444 4136
rect 10828 4012 10868 4052
rect 10732 3844 10772 3884
rect 10732 3340 10772 3380
rect 10636 2836 10676 2876
rect 10732 2752 10772 2792
rect 10540 1912 10580 1952
rect 10540 1576 10580 1616
rect 11212 3928 11252 3968
rect 11692 4516 11732 4556
rect 11596 4180 11636 4220
rect 11980 4768 12020 4808
rect 12076 4684 12116 4724
rect 11884 4096 11924 4136
rect 11692 4012 11732 4052
rect 12076 4096 12116 4136
rect 11596 3928 11636 3968
rect 10828 2500 10868 2540
rect 11020 2500 11060 2540
rect 11020 2164 11060 2204
rect 11212 2752 11252 2792
rect 11212 2500 11252 2540
rect 10924 1576 10964 1616
rect 11692 3760 11732 3800
rect 11788 3424 11828 3464
rect 11788 3172 11828 3212
rect 11596 2836 11636 2876
rect 11500 2584 11540 2624
rect 11404 2080 11444 2120
rect 11980 3928 12020 3968
rect 12076 3760 12116 3800
rect 12076 3424 12116 3464
rect 12652 7120 12692 7160
rect 13804 8296 13844 8336
rect 13324 7120 13364 7160
rect 12556 7036 12596 7076
rect 13516 7456 13556 7496
rect 13612 7372 13652 7412
rect 13516 7288 13556 7328
rect 13708 7288 13748 7328
rect 13420 7036 13460 7076
rect 12940 6616 12980 6656
rect 14572 14764 14612 14804
rect 15148 15604 15188 15644
rect 15052 15436 15092 15476
rect 15148 15100 15188 15140
rect 15436 15016 15476 15056
rect 15820 16276 15860 16316
rect 15724 16024 15764 16064
rect 15916 15940 15956 15980
rect 15820 15520 15860 15560
rect 15628 14764 15668 14804
rect 15052 14596 15092 14636
rect 14476 14260 14516 14300
rect 15052 14260 15092 14300
rect 14764 14176 14804 14216
rect 14476 14008 14516 14048
rect 14860 14008 14900 14048
rect 14668 13924 14708 13964
rect 14476 13588 14516 13628
rect 14284 12748 14324 12788
rect 15244 13924 15284 13964
rect 15244 13588 15284 13628
rect 15436 13420 15476 13460
rect 16492 17200 16532 17240
rect 16780 18544 16820 18584
rect 17164 18796 17204 18836
rect 17068 18628 17108 18668
rect 17164 18544 17204 18584
rect 17068 18460 17108 18500
rect 17164 18376 17204 18416
rect 16972 17872 17012 17912
rect 16781 17704 16821 17744
rect 16876 17620 16916 17660
rect 16780 17452 16820 17492
rect 16684 17200 16724 17240
rect 16396 16864 16436 16904
rect 16300 16192 16340 16232
rect 17548 21316 17588 21356
rect 17452 20728 17492 20768
rect 17644 21148 17684 21188
rect 17548 20140 17588 20180
rect 17548 19552 17588 19592
rect 17452 19300 17492 19340
rect 17548 19216 17588 19256
rect 17452 18796 17492 18836
rect 17356 18460 17396 18500
rect 17452 18208 17492 18248
rect 17356 17200 17396 17240
rect 17356 16948 17396 16988
rect 16876 16360 16916 16400
rect 17260 16360 17300 16400
rect 16780 16024 16820 16064
rect 16876 15856 16916 15896
rect 16204 15520 16244 15560
rect 16684 15436 16724 15476
rect 16396 15352 16436 15392
rect 16300 15268 16340 15308
rect 16396 15184 16436 15224
rect 16300 15100 16340 15140
rect 16588 14932 16628 14972
rect 16492 14680 16532 14720
rect 16300 14344 16340 14384
rect 15628 14008 15668 14048
rect 15724 13840 15764 13880
rect 15628 13420 15668 13460
rect 15436 13252 15476 13292
rect 15340 13168 15380 13208
rect 14860 13000 14900 13040
rect 15244 12832 15284 12872
rect 14572 12748 14612 12788
rect 14476 12496 14516 12536
rect 14284 11992 14324 12032
rect 14284 11824 14324 11864
rect 14188 11152 14228 11192
rect 14572 12412 14612 12452
rect 14572 12076 14612 12116
rect 15052 11908 15092 11948
rect 14476 11320 14516 11360
rect 15148 11656 15188 11696
rect 15052 11320 15092 11360
rect 14860 10984 14900 11024
rect 14284 10732 14324 10772
rect 14092 10228 14132 10268
rect 14284 10060 14324 10100
rect 14188 9724 14228 9764
rect 13996 8716 14036 8756
rect 14092 8296 14132 8336
rect 14092 8128 14132 8168
rect 14188 7960 14228 8000
rect 13996 7372 14036 7412
rect 13996 7120 14036 7160
rect 13612 7036 13652 7076
rect 13900 7036 13940 7076
rect 12844 6448 12884 6488
rect 12364 6112 12404 6152
rect 12460 5860 12500 5900
rect 12460 5356 12500 5396
rect 12364 5188 12404 5228
rect 13516 6532 13556 6572
rect 13324 6448 13364 6488
rect 13228 6364 13268 6404
rect 13036 5608 13076 5648
rect 12652 5188 12692 5228
rect 12844 5440 12884 5480
rect 13420 6196 13460 6236
rect 13324 5860 13364 5900
rect 13324 5692 13364 5732
rect 13132 5356 13172 5396
rect 12364 4936 12404 4976
rect 12652 4936 12692 4976
rect 12844 4936 12884 4976
rect 12460 4852 12500 4892
rect 12748 4852 12788 4892
rect 12556 4768 12596 4808
rect 12364 4684 12404 4724
rect 12268 3340 12308 3380
rect 12172 3172 12212 3212
rect 12172 2668 12212 2708
rect 12460 4516 12500 4556
rect 12460 2668 12500 2708
rect 11500 1744 11540 1784
rect 11596 1576 11636 1616
rect 11308 1408 11348 1448
rect 11020 1240 11060 1280
rect 10732 1156 10772 1196
rect 11212 904 11252 944
rect 11020 484 11060 524
rect 10924 316 10964 356
rect 10636 232 10676 272
rect 10828 64 10868 104
rect 11500 232 11540 272
rect 11404 148 11444 188
rect 11980 2248 12020 2288
rect 11788 1492 11828 1532
rect 12172 2332 12212 2372
rect 13132 4684 13172 4724
rect 13132 4348 13172 4388
rect 13516 5692 13556 5732
rect 13708 6616 13748 6656
rect 13804 6448 13844 6488
rect 13900 6364 13940 6404
rect 13708 6196 13748 6236
rect 13900 5860 13940 5900
rect 13420 5440 13460 5480
rect 14860 10732 14900 10772
rect 14764 10396 14804 10436
rect 14572 10060 14612 10100
rect 14476 9556 14516 9596
rect 14764 9892 14804 9932
rect 14668 9556 14708 9596
rect 14668 9136 14708 9176
rect 16012 13840 16052 13880
rect 15916 13588 15956 13628
rect 15532 12412 15572 12452
rect 16108 13168 16148 13208
rect 16108 13000 16148 13040
rect 16780 14596 16820 14636
rect 16972 15352 17012 15392
rect 16972 15100 17012 15140
rect 17260 15940 17300 15980
rect 17260 15352 17300 15392
rect 17164 14932 17204 14972
rect 17452 15772 17492 15812
rect 17836 21988 17876 22028
rect 18220 25432 18260 25472
rect 18124 25096 18164 25136
rect 18028 23500 18068 23540
rect 18508 26356 18548 26396
rect 18508 26188 18548 26228
rect 18508 25432 18548 25472
rect 18700 30640 18740 30680
rect 19372 31984 19412 32024
rect 19180 30808 19220 30848
rect 19276 30724 19316 30764
rect 18892 30388 18932 30428
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 19468 31396 19508 31436
rect 19756 32320 19796 32360
rect 20140 33496 20180 33536
rect 19948 33412 19988 33452
rect 20140 33076 20180 33116
rect 21196 40384 21236 40424
rect 20812 40048 20852 40088
rect 20812 39544 20852 39584
rect 21004 37192 21044 37232
rect 20716 37108 20756 37148
rect 20716 36856 20756 36896
rect 20812 35932 20852 35972
rect 20812 34000 20852 34040
rect 20716 33664 20756 33704
rect 20620 33328 20660 33368
rect 20524 32992 20564 33032
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 19852 31984 19892 32024
rect 19756 31648 19796 31688
rect 19660 31396 19700 31436
rect 19756 31312 19796 31352
rect 19660 31144 19700 31184
rect 19564 31060 19604 31100
rect 19660 30808 19700 30848
rect 19948 31396 19988 31436
rect 20044 31312 20084 31352
rect 19852 30724 19892 30764
rect 19756 30640 19796 30680
rect 19468 30556 19508 30596
rect 19372 30052 19412 30092
rect 19372 29884 19412 29924
rect 19756 29884 19796 29924
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 19948 29800 19988 29840
rect 21196 35596 21236 35636
rect 21196 33412 21236 33452
rect 21004 30304 21044 30344
rect 18604 25348 18644 25388
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18988 28456 19028 28496
rect 18892 28204 18932 28244
rect 19372 29044 19412 29084
rect 19468 28456 19508 28496
rect 19276 28372 19316 28412
rect 18796 27700 18836 27740
rect 19276 27700 19316 27740
rect 18892 27616 18932 27656
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 19468 27532 19508 27572
rect 19372 27028 19412 27068
rect 19660 28036 19700 28076
rect 19660 27364 19700 27404
rect 20044 29632 20084 29672
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 21388 30136 21428 30176
rect 19948 29212 19988 29252
rect 19948 28960 19988 29000
rect 19948 28120 19988 28160
rect 20908 28120 20948 28160
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 19852 27700 19892 27740
rect 19852 27364 19892 27404
rect 19564 26944 19604 26984
rect 19180 26608 19220 26648
rect 19660 26692 19700 26732
rect 19564 26608 19604 26648
rect 19372 26440 19412 26480
rect 18892 26188 18932 26228
rect 19276 26104 19316 26144
rect 19383 26104 19412 26144
rect 19412 26104 19423 26144
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18892 25432 18932 25472
rect 18412 24844 18452 24884
rect 18316 24592 18356 24632
rect 18220 23332 18260 23372
rect 18124 22576 18164 22616
rect 18124 21652 18164 21692
rect 18028 21568 18068 21608
rect 17932 21148 17972 21188
rect 17836 21064 17876 21104
rect 17836 20812 17876 20852
rect 18412 23080 18452 23120
rect 18796 24760 18836 24800
rect 19372 25936 19412 25976
rect 19276 25348 19316 25388
rect 19756 26020 19796 26060
rect 19948 27028 19988 27068
rect 19948 26776 19988 26816
rect 20044 26608 20084 26648
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20908 26272 20948 26312
rect 19756 25348 19796 25388
rect 19276 24760 19316 24800
rect 19468 24424 19508 24464
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 21004 25936 21044 25976
rect 21292 29128 21332 29168
rect 21196 25180 21236 25220
rect 19852 24760 19892 24800
rect 19756 24592 19796 24632
rect 19564 24088 19604 24128
rect 18700 23668 18740 23708
rect 18988 23080 19028 23120
rect 18412 22240 18452 22280
rect 18604 22240 18644 22280
rect 19180 23752 19220 23792
rect 19851 24508 19891 24548
rect 20044 25096 20084 25136
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20044 24592 20084 24632
rect 19948 24256 19988 24296
rect 19948 23836 19988 23876
rect 19180 23080 19220 23120
rect 19660 23248 19700 23288
rect 19276 22996 19316 23036
rect 19084 22912 19124 22952
rect 19372 22912 19412 22952
rect 18796 22828 18836 22868
rect 19276 22828 19316 22868
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 19276 22492 19316 22532
rect 19084 22240 19124 22280
rect 18700 22156 18740 22196
rect 19564 22828 19604 22868
rect 19756 22996 19796 23036
rect 19660 22660 19700 22700
rect 19660 22492 19700 22532
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 19948 22996 19988 23036
rect 19948 22828 19988 22868
rect 20140 22912 20180 22952
rect 20236 22744 20276 22784
rect 20524 22576 20564 22616
rect 19468 22156 19508 22196
rect 20140 22072 20180 22112
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 19372 21736 19412 21776
rect 20044 21736 20084 21776
rect 18796 21652 18836 21692
rect 18604 21568 18644 21608
rect 18316 21316 18356 21356
rect 18508 20728 18548 20768
rect 18220 20644 18260 20684
rect 18028 20224 18068 20264
rect 18508 20308 18548 20348
rect 17932 20056 17972 20096
rect 18124 20056 18164 20096
rect 18028 19972 18068 20012
rect 17740 19720 17780 19760
rect 17836 18628 17876 18668
rect 17932 18292 17972 18332
rect 17740 18124 17780 18164
rect 17740 17116 17780 17156
rect 17356 14848 17396 14888
rect 17644 15352 17684 15392
rect 17548 14932 17588 14972
rect 16780 14344 16820 14384
rect 17356 14512 17396 14552
rect 16876 14092 16916 14132
rect 17164 14092 17204 14132
rect 16492 13504 16532 13544
rect 15436 12244 15476 12284
rect 15628 10984 15668 11024
rect 15244 10480 15284 10520
rect 15436 10480 15476 10520
rect 15052 10228 15092 10268
rect 14572 8296 14612 8336
rect 14476 8128 14516 8168
rect 14860 8296 14900 8336
rect 14860 8128 14900 8168
rect 14764 7960 14804 8000
rect 15148 9724 15188 9764
rect 15244 9556 15284 9596
rect 15148 9472 15188 9512
rect 15244 9304 15284 9344
rect 15340 8968 15380 9008
rect 15148 8716 15188 8756
rect 14668 7540 14708 7580
rect 14380 7456 14420 7496
rect 14188 7036 14228 7076
rect 14092 5776 14132 5816
rect 14284 6532 14324 6572
rect 14476 6448 14516 6488
rect 14668 6448 14708 6488
rect 14380 6280 14420 6320
rect 14284 6196 14324 6236
rect 14188 5692 14228 5732
rect 13804 5440 13844 5480
rect 13324 4936 13364 4976
rect 13516 5356 13556 5396
rect 13708 5356 13748 5396
rect 13900 5188 13940 5228
rect 13612 4852 13652 4892
rect 13516 4768 13556 4808
rect 14188 5020 14228 5060
rect 13996 4936 14036 4976
rect 13804 4684 13844 4724
rect 12844 4264 12884 4304
rect 13132 3760 13172 3800
rect 13324 3760 13364 3800
rect 13228 3340 13268 3380
rect 12748 2920 12788 2960
rect 12652 2584 12692 2624
rect 12556 2332 12596 2372
rect 12460 2164 12500 2204
rect 13036 2164 13076 2204
rect 12172 2080 12212 2120
rect 12556 2080 12596 2120
rect 12172 1744 12212 1784
rect 12364 1492 12404 1532
rect 12748 1744 12788 1784
rect 12940 1240 12980 1280
rect 13132 2080 13172 2120
rect 13612 3676 13652 3716
rect 13516 3424 13556 3464
rect 14092 4432 14132 4472
rect 13996 4180 14036 4220
rect 13900 3676 13940 3716
rect 13996 3424 14036 3464
rect 13516 3004 13556 3044
rect 13420 2416 13460 2456
rect 13132 1576 13172 1616
rect 13324 1576 13364 1616
rect 13324 1240 13364 1280
rect 13132 1072 13172 1112
rect 13228 988 13268 1028
rect 12556 904 12596 944
rect 12940 904 12980 944
rect 12460 148 12500 188
rect 12748 484 12788 524
rect 13132 820 13172 860
rect 13420 1072 13460 1112
rect 13708 2668 13748 2708
rect 13612 2080 13652 2120
rect 14188 4180 14228 4220
rect 13900 2752 13940 2792
rect 13804 1744 13844 1784
rect 14284 2920 14324 2960
rect 14188 1660 14228 1700
rect 13708 1576 13748 1616
rect 15340 8632 15380 8672
rect 15148 8296 15188 8336
rect 14860 7624 14900 7664
rect 14764 5860 14804 5900
rect 15052 7288 15092 7328
rect 14956 6868 14996 6908
rect 15532 10060 15572 10100
rect 16300 11572 16340 11612
rect 16972 13336 17012 13376
rect 16684 13168 16724 13208
rect 17068 12664 17108 12704
rect 17260 14008 17300 14048
rect 17260 12496 17300 12536
rect 16780 11908 16820 11948
rect 16492 11488 16532 11528
rect 16108 11320 16148 11360
rect 15820 10144 15860 10184
rect 16012 10648 16052 10688
rect 16108 10312 16148 10352
rect 16780 11488 16820 11528
rect 16780 10984 16820 11024
rect 16684 10900 16724 10940
rect 16396 10732 16436 10772
rect 17452 14428 17492 14468
rect 17452 12580 17492 12620
rect 17452 11740 17492 11780
rect 17644 14596 17684 14636
rect 17644 14260 17684 14300
rect 17644 12916 17684 12956
rect 17644 12664 17684 12704
rect 17548 11656 17588 11696
rect 17356 11488 17396 11528
rect 17932 15352 17972 15392
rect 17836 13084 17876 13124
rect 19276 21484 19316 21524
rect 19468 21568 19508 21608
rect 19948 21484 19988 21524
rect 19756 21400 19796 21440
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 19372 21316 19412 21356
rect 19372 20980 19412 21020
rect 18604 20224 18644 20264
rect 19564 20980 19604 21020
rect 19084 20812 19124 20852
rect 18316 19804 18356 19844
rect 18508 19636 18548 19676
rect 18220 19216 18260 19256
rect 18988 20056 19028 20096
rect 19276 20308 19316 20348
rect 19276 20140 19316 20180
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18700 18880 18740 18920
rect 18604 18712 18644 18752
rect 18412 18628 18452 18668
rect 18220 18376 18260 18416
rect 18124 18040 18164 18080
rect 18316 16696 18356 16736
rect 19180 19216 19220 19256
rect 19564 20392 19604 20432
rect 19468 19384 19508 19424
rect 20236 20728 20276 20768
rect 20044 20644 20084 20684
rect 19756 20560 19796 20600
rect 19852 20392 19892 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 19948 19972 19988 20012
rect 19948 19804 19988 19844
rect 20812 19888 20852 19928
rect 19660 19552 19700 19592
rect 19660 19384 19700 19424
rect 19468 19216 19508 19256
rect 19372 18964 19412 19004
rect 19564 18880 19604 18920
rect 19276 18796 19316 18836
rect 19180 18712 19220 18752
rect 19372 18712 19412 18752
rect 20236 19216 20276 19256
rect 19756 19132 19796 19172
rect 19852 19048 19892 19088
rect 20140 19048 20180 19088
rect 19756 18964 19796 19004
rect 19660 18544 19700 18584
rect 19948 18880 19988 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 19852 18712 19892 18752
rect 20332 18712 20372 18752
rect 19468 18292 19508 18332
rect 19756 18292 19796 18332
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 20236 18292 20276 18332
rect 20140 18040 20180 18080
rect 19180 17956 19220 17996
rect 19948 17956 19988 17996
rect 19372 17788 19412 17828
rect 19756 17788 19796 17828
rect 19948 17620 19988 17660
rect 19180 17368 19220 17408
rect 18604 17284 18644 17324
rect 18988 17284 19028 17324
rect 18796 17116 18836 17156
rect 18508 16192 18548 16232
rect 19084 16864 19124 16904
rect 18988 16780 19028 16820
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18508 16024 18548 16064
rect 18412 15268 18452 15308
rect 18412 15100 18452 15140
rect 20620 18544 20660 18584
rect 20332 17704 20372 17744
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20127 17116 20167 17156
rect 19468 16528 19508 16568
rect 19948 17032 19988 17072
rect 19660 16948 19700 16988
rect 19756 16864 19796 16904
rect 19660 16444 19700 16484
rect 19372 15856 19412 15896
rect 19276 15520 19316 15560
rect 19564 16192 19604 16232
rect 19468 15436 19508 15476
rect 18604 15100 18644 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18604 14848 18644 14888
rect 19084 14764 19124 14804
rect 18412 13504 18452 13544
rect 18316 13168 18356 13208
rect 18028 12664 18068 12704
rect 18028 12496 18068 12536
rect 17836 11656 17876 11696
rect 18220 11572 18260 11612
rect 16972 10900 17012 10940
rect 16876 10732 16916 10772
rect 16300 10396 16340 10436
rect 16684 10564 16724 10604
rect 16588 10312 16628 10352
rect 16492 10144 16532 10184
rect 16012 9724 16052 9764
rect 15436 8296 15476 8336
rect 15436 8044 15476 8084
rect 15244 7372 15284 7412
rect 15436 7624 15476 7664
rect 15916 9556 15956 9596
rect 15820 9472 15860 9512
rect 15724 9220 15764 9260
rect 15628 9136 15668 9176
rect 16300 9976 16340 10016
rect 16300 9640 16340 9680
rect 16588 9640 16628 9680
rect 16300 9472 16340 9512
rect 16492 9472 16532 9512
rect 16204 9388 16244 9428
rect 16396 9304 16436 9344
rect 16204 8968 16244 9008
rect 15628 7624 15668 7664
rect 15340 7288 15380 7328
rect 15628 7288 15668 7328
rect 15436 7204 15476 7244
rect 15148 6616 15188 6656
rect 15052 5860 15092 5900
rect 14860 5020 14900 5060
rect 14476 4936 14516 4976
rect 14476 3760 14516 3800
rect 15148 3592 15188 3632
rect 15052 3340 15092 3380
rect 15148 3256 15188 3296
rect 14956 2752 14996 2792
rect 15148 2752 15188 2792
rect 13900 1156 13940 1196
rect 13516 904 13556 944
rect 13708 904 13748 944
rect 13900 652 13940 692
rect 14284 1240 14324 1280
rect 14476 1240 14516 1280
rect 14188 568 14228 608
rect 14668 1240 14708 1280
rect 14380 1156 14420 1196
rect 14380 148 14420 188
rect 14860 1156 14900 1196
rect 15532 6952 15572 6992
rect 16012 7120 16052 7160
rect 15916 7036 15956 7076
rect 16108 6700 16148 6740
rect 15820 6280 15860 6320
rect 15916 6196 15956 6236
rect 15532 5860 15572 5900
rect 16780 10480 16820 10520
rect 17164 10816 17204 10856
rect 17068 10480 17108 10520
rect 16972 10396 17012 10436
rect 16876 10312 16916 10352
rect 16780 9808 16820 9848
rect 16876 9472 16916 9512
rect 16780 9220 16820 9260
rect 16300 8044 16340 8084
rect 16300 7792 16340 7832
rect 17260 10144 17300 10184
rect 17164 9892 17204 9932
rect 17836 10984 17876 11024
rect 17644 10900 17684 10940
rect 17644 10732 17684 10772
rect 17740 10648 17780 10688
rect 17644 10480 17684 10520
rect 17452 10312 17492 10352
rect 17644 10312 17684 10352
rect 18124 11152 18164 11192
rect 17836 10060 17876 10100
rect 17548 9976 17588 10016
rect 16972 9220 17012 9260
rect 16588 8380 16628 8420
rect 16780 8632 16820 8672
rect 16780 8380 16820 8420
rect 16684 8044 16724 8084
rect 16876 8044 16916 8084
rect 16780 7792 16820 7832
rect 17164 8968 17204 9008
rect 17068 8632 17108 8672
rect 17260 8380 17300 8420
rect 17164 8044 17204 8084
rect 17068 7960 17108 8000
rect 17452 8632 17492 8672
rect 17644 9724 17684 9764
rect 17548 8212 17588 8252
rect 17740 9472 17780 9512
rect 17932 9976 17972 10016
rect 18220 10984 18260 11024
rect 18124 10144 18164 10184
rect 18028 9892 18068 9932
rect 18028 9724 18068 9764
rect 17932 9640 17972 9680
rect 18220 9640 18260 9680
rect 18124 9556 18164 9596
rect 17932 9388 17972 9428
rect 18225 9388 18265 9428
rect 18220 9220 18260 9260
rect 17356 7792 17396 7832
rect 16684 7120 16724 7160
rect 16588 7036 16628 7076
rect 16396 6784 16436 6824
rect 16300 6700 16340 6740
rect 16492 6700 16532 6740
rect 16301 6280 16341 6320
rect 16588 6280 16628 6320
rect 16204 5692 16244 5732
rect 15724 5608 15764 5648
rect 15436 5524 15476 5564
rect 15820 5440 15860 5480
rect 16012 5608 16052 5648
rect 15916 5272 15956 5312
rect 16204 5524 16244 5564
rect 16108 4936 16148 4976
rect 17836 8464 17876 8504
rect 17548 7792 17588 7832
rect 17260 6952 17300 6992
rect 17164 6532 17204 6572
rect 17356 6532 17396 6572
rect 17740 7456 17780 7496
rect 17644 6532 17684 6572
rect 17452 6448 17492 6488
rect 17068 5692 17108 5732
rect 16684 5608 16724 5648
rect 17260 5608 17300 5648
rect 18124 8548 18164 8588
rect 18028 8044 18068 8084
rect 18028 7540 18068 7580
rect 17452 6196 17492 6236
rect 16588 5188 16628 5228
rect 16492 5104 16532 5144
rect 16300 5020 16340 5060
rect 16492 4936 16532 4976
rect 15916 4432 15956 4472
rect 15820 4264 15860 4304
rect 15724 4096 15764 4136
rect 15628 3928 15668 3968
rect 15532 3592 15572 3632
rect 15628 3508 15668 3548
rect 15820 3508 15860 3548
rect 16012 4096 16052 4136
rect 17164 4684 17204 4724
rect 17068 4264 17108 4304
rect 16780 4096 16820 4136
rect 16492 3760 16532 3800
rect 16396 3676 16436 3716
rect 16204 3592 16244 3632
rect 15436 3256 15476 3296
rect 15724 3172 15764 3212
rect 15340 2920 15380 2960
rect 15916 2920 15956 2960
rect 15244 2248 15284 2288
rect 16012 2584 16052 2624
rect 15532 1996 15572 2036
rect 15436 1744 15476 1784
rect 15052 1660 15092 1700
rect 15436 1408 15476 1448
rect 14956 1072 14996 1112
rect 15244 820 15284 860
rect 14860 484 14900 524
rect 15052 400 15092 440
rect 15628 1072 15668 1112
rect 15916 1912 15956 1952
rect 16108 2500 16148 2540
rect 16300 2836 16340 2876
rect 16300 2500 16340 2540
rect 16588 3592 16628 3632
rect 16492 3256 16532 3296
rect 16204 1744 16244 1784
rect 15820 736 15860 776
rect 15820 400 15860 440
rect 15628 232 15668 272
rect 16108 400 16148 440
rect 16396 1408 16436 1448
rect 16300 1072 16340 1112
rect 16492 1156 16532 1196
rect 16684 3508 16724 3548
rect 17068 3760 17108 3800
rect 16972 3508 17012 3548
rect 16876 3088 16916 3128
rect 16780 2668 16820 2708
rect 17452 5020 17492 5060
rect 17356 4096 17396 4136
rect 18700 13840 18740 13880
rect 18988 13840 19028 13880
rect 19756 15688 19796 15728
rect 19660 15604 19700 15644
rect 19756 15352 19796 15392
rect 19660 15268 19700 15308
rect 19180 14680 19220 14720
rect 19468 14680 19508 14720
rect 19564 14596 19604 14636
rect 19756 14932 19796 14972
rect 19948 16780 19988 16820
rect 20236 16948 20276 16988
rect 20236 16024 20276 16064
rect 19948 15856 19988 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20044 15688 20084 15728
rect 19948 15604 19988 15644
rect 19372 14344 19412 14384
rect 19180 13756 19220 13796
rect 18700 13588 18740 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18796 13336 18836 13376
rect 19084 13336 19124 13376
rect 18508 13168 18548 13208
rect 18700 13168 18740 13208
rect 18604 12580 18644 12620
rect 18412 11992 18452 12032
rect 20236 14932 20276 14972
rect 20716 17200 20756 17240
rect 20620 14932 20660 14972
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 19660 13840 19700 13880
rect 19756 13756 19796 13796
rect 19660 13168 19700 13208
rect 20236 14092 20276 14132
rect 20044 13924 20084 13964
rect 19948 13168 19988 13208
rect 19372 13000 19412 13040
rect 18796 12496 18836 12536
rect 19180 12496 19220 12536
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 19756 12916 19796 12956
rect 19564 12832 19604 12872
rect 19468 12412 19508 12452
rect 19564 11992 19604 12032
rect 19372 11908 19412 11948
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20044 12664 20084 12704
rect 19948 12580 19988 12620
rect 21388 28960 21428 29000
rect 21292 19216 21332 19256
rect 20908 18880 20948 18920
rect 20812 14092 20852 14132
rect 20236 12412 20276 12452
rect 20716 12412 20756 12452
rect 21004 17704 21044 17744
rect 20524 12076 20564 12116
rect 20908 12076 20948 12116
rect 19276 10984 19316 11024
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18604 10480 18644 10520
rect 18700 10228 18740 10268
rect 18508 10060 18548 10100
rect 18604 9976 18644 10016
rect 18508 9136 18548 9176
rect 18508 8800 18548 8840
rect 18409 8716 18449 8756
rect 18412 8548 18452 8588
rect 18316 8128 18356 8168
rect 18796 9388 18836 9428
rect 19180 9472 19220 9512
rect 19468 10648 19508 10688
rect 19372 10396 19412 10436
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 19948 11236 19988 11276
rect 20620 11992 20660 12032
rect 19852 10648 19892 10688
rect 19852 10228 19892 10268
rect 19468 9556 19508 9596
rect 19276 9304 19316 9344
rect 19084 9220 19124 9260
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18796 8800 18836 8840
rect 18700 8548 18740 8588
rect 18604 8464 18644 8504
rect 18508 8380 18548 8420
rect 18988 8296 19028 8336
rect 18892 8128 18932 8168
rect 18220 8044 18260 8084
rect 18604 7876 18644 7916
rect 19084 7960 19124 8000
rect 19756 8632 19796 8672
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20524 9640 20564 9680
rect 20127 9556 20167 9596
rect 19948 9304 19988 9344
rect 20236 9388 20276 9428
rect 18988 7792 19028 7832
rect 18220 7624 18260 7664
rect 18508 7624 18548 7664
rect 18508 7120 18548 7160
rect 18508 5608 18548 5648
rect 17548 4516 17588 4556
rect 17644 4264 17684 4304
rect 17260 3592 17300 3632
rect 17644 4012 17684 4052
rect 17932 4096 17972 4136
rect 17836 3760 17876 3800
rect 17548 3592 17588 3632
rect 17740 3592 17780 3632
rect 17260 3256 17300 3296
rect 17164 2500 17204 2540
rect 17548 3004 17588 3044
rect 17548 2752 17588 2792
rect 17548 2500 17588 2540
rect 17740 3256 17780 3296
rect 18028 3340 18068 3380
rect 18316 4936 18356 4976
rect 18220 4516 18260 4556
rect 18220 4348 18260 4388
rect 18220 3760 18260 3800
rect 18220 3424 18260 3464
rect 18124 3172 18164 3212
rect 18028 2920 18068 2960
rect 17932 2752 17972 2792
rect 18028 2584 18068 2624
rect 18124 2500 18164 2540
rect 18508 4936 18548 4976
rect 18412 4768 18452 4808
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 20140 8464 20180 8504
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 20044 8128 20084 8168
rect 19468 7708 19508 7748
rect 19372 7540 19412 7580
rect 19660 7792 19700 7832
rect 19660 7540 19700 7580
rect 19276 7204 19316 7244
rect 18988 7120 19028 7160
rect 19468 7204 19508 7244
rect 19564 7120 19604 7160
rect 20812 11908 20852 11948
rect 20812 11152 20852 11192
rect 20716 11068 20756 11108
rect 20620 8464 20660 8504
rect 21100 14176 21140 14216
rect 21004 10144 21044 10184
rect 21004 9136 21044 9176
rect 19852 7456 19892 7496
rect 19756 7120 19796 7160
rect 19756 6700 19796 6740
rect 19852 6616 19892 6656
rect 19660 6448 19700 6488
rect 19564 6280 19604 6320
rect 18700 6028 18740 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18700 5608 18740 5648
rect 18796 5020 18836 5060
rect 18700 4936 18740 4976
rect 19468 5944 19508 5984
rect 19180 5272 19220 5312
rect 19276 5020 19316 5060
rect 19084 4936 19124 4976
rect 18412 4600 18452 4640
rect 18508 4264 18548 4304
rect 18412 3760 18452 3800
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 18796 4348 18836 4388
rect 19084 4348 19124 4388
rect 19276 4012 19316 4052
rect 19756 6364 19796 6404
rect 19660 5272 19700 5312
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20332 6616 20372 6656
rect 20236 6532 20276 6572
rect 19852 5440 19892 5480
rect 19756 5020 19796 5060
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 19948 4936 19988 4976
rect 20044 4768 20084 4808
rect 19564 4432 19604 4472
rect 19564 4264 19604 4304
rect 19372 3928 19412 3968
rect 19084 3844 19124 3884
rect 18412 3256 18452 3296
rect 18220 2164 18260 2204
rect 18028 2080 18068 2120
rect 17740 1996 17780 2036
rect 17932 1912 17972 1952
rect 17452 1828 17492 1868
rect 16876 1492 16916 1532
rect 16972 1240 17012 1280
rect 16876 400 16916 440
rect 16780 316 16820 356
rect 17164 1744 17204 1784
rect 17452 1660 17492 1700
rect 17356 1156 17396 1196
rect 17164 148 17204 188
rect 17548 1324 17588 1364
rect 17740 1828 17780 1868
rect 17932 1240 17972 1280
rect 17740 1072 17780 1112
rect 17548 988 17588 1028
rect 17740 904 17780 944
rect 17548 400 17588 440
rect 19468 3760 19508 3800
rect 18796 3256 18836 3296
rect 19276 3424 19316 3464
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 20122 4180 20162 4220
rect 19948 4096 19988 4136
rect 19564 3256 19604 3296
rect 19756 3256 19796 3296
rect 19276 2332 19316 2372
rect 18604 2080 18644 2120
rect 18508 1912 18548 1952
rect 19372 2248 19412 2288
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 19660 2920 19700 2960
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 19948 3592 19988 3632
rect 20044 3508 20084 3548
rect 20129 3172 20169 3212
rect 19852 2836 19892 2876
rect 20140 2500 20180 2540
rect 19948 2416 19988 2456
rect 19852 2248 19892 2288
rect 19660 2080 19700 2120
rect 19276 1408 19316 1448
rect 18508 1240 18548 1280
rect 18700 1240 18740 1280
rect 18316 652 18356 692
rect 18124 64 18164 104
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 20127 1912 20167 1952
rect 19852 1744 19892 1784
rect 21196 9976 21236 10016
rect 21100 7120 21140 7160
rect 21004 5188 21044 5228
rect 20716 4852 20756 4892
rect 20812 3928 20852 3968
rect 20716 3760 20756 3800
rect 20812 2416 20852 2456
rect 19084 904 19124 944
rect 18892 400 18932 440
rect 19468 736 19508 776
rect 19276 568 19316 608
rect 20044 904 20084 944
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 19660 484 19700 524
rect 21196 64 21236 104
<< metal3 >>
rect 15523 42944 15581 42945
rect 1219 42904 1228 42944
rect 1268 42904 14668 42944
rect 14708 42904 14717 42944
rect 15523 42904 15532 42944
rect 15572 42904 19276 42944
rect 19316 42904 19325 42944
rect 15523 42903 15581 42904
rect 1411 42860 1469 42861
rect 1411 42820 1420 42860
rect 1460 42820 17548 42860
rect 17588 42820 17597 42860
rect 1411 42819 1469 42820
rect 21091 42776 21149 42777
rect 21424 42776 21504 42796
rect 8131 42736 8140 42776
rect 8180 42736 17836 42776
rect 17876 42736 17885 42776
rect 21091 42736 21100 42776
rect 21140 42736 21504 42776
rect 21091 42735 21149 42736
rect 21424 42716 21504 42736
rect 7555 42692 7613 42693
rect 18307 42692 18365 42693
rect 7555 42652 7564 42692
rect 7604 42652 17356 42692
rect 17396 42652 17405 42692
rect 18307 42652 18316 42692
rect 18356 42652 18892 42692
rect 18932 42652 18941 42692
rect 7555 42651 7613 42652
rect 18307 42651 18365 42652
rect 9475 42608 9533 42609
rect 18019 42608 18077 42609
rect 9475 42568 9484 42608
rect 9524 42568 9676 42608
rect 9716 42568 9725 42608
rect 18019 42568 18028 42608
rect 18068 42568 18124 42608
rect 18164 42568 18173 42608
rect 9475 42567 9533 42568
rect 18019 42567 18077 42568
rect 451 42524 509 42525
rect 451 42484 460 42524
rect 500 42484 5260 42524
rect 5300 42484 5309 42524
rect 5731 42484 5740 42524
rect 5780 42484 11980 42524
rect 12020 42484 12029 42524
rect 16195 42484 16204 42524
rect 16244 42484 19564 42524
rect 19604 42484 19613 42524
rect 451 42483 509 42484
rect 1027 42440 1085 42441
rect 21424 42440 21504 42460
rect 1027 42400 1036 42440
rect 1076 42400 3916 42440
rect 3956 42400 3965 42440
rect 7267 42400 7276 42440
rect 7316 42400 21504 42440
rect 1027 42399 1085 42400
rect 21424 42380 21504 42400
rect 16387 42316 16396 42356
rect 16436 42316 19756 42356
rect 19796 42316 19805 42356
rect 13891 42232 13900 42272
rect 13940 42232 19276 42272
rect 19316 42232 19325 42272
rect 2275 42148 2284 42188
rect 2324 42148 3340 42188
rect 3380 42148 3389 42188
rect 11107 42148 11116 42188
rect 11156 42148 12556 42188
rect 12596 42148 12605 42188
rect 13315 42148 13324 42188
rect 13364 42148 17644 42188
rect 17684 42148 17693 42188
rect 21283 42104 21341 42105
rect 21424 42104 21504 42124
rect 1891 42064 1900 42104
rect 1940 42064 4684 42104
rect 4724 42064 4733 42104
rect 13507 42064 13516 42104
rect 13556 42064 18508 42104
rect 18548 42064 18557 42104
rect 21283 42064 21292 42104
rect 21332 42064 21504 42104
rect 21283 42063 21341 42064
rect 21424 42044 21504 42064
rect 6403 42020 6461 42021
rect 16291 42020 16349 42021
rect 6403 41980 6412 42020
rect 6452 41980 6796 42020
rect 6836 41980 6845 42020
rect 10627 41980 10636 42020
rect 10676 41980 10924 42020
rect 10964 41980 10973 42020
rect 13699 41980 13708 42020
rect 13748 41980 16300 42020
rect 16340 41980 16349 42020
rect 6403 41979 6461 41980
rect 16291 41979 16349 41980
rect 5443 41936 5501 41937
rect 17923 41936 17981 41937
rect 2563 41896 2572 41936
rect 2612 41896 5452 41936
rect 5492 41896 5501 41936
rect 9379 41896 9388 41936
rect 9428 41896 15052 41936
rect 15092 41896 15101 41936
rect 17923 41896 17932 41936
rect 17972 41896 18700 41936
rect 18740 41896 18749 41936
rect 5443 41895 5501 41896
rect 17923 41895 17981 41896
rect 5539 41852 5597 41853
rect 7843 41852 7901 41853
rect 18211 41852 18269 41853
rect 5539 41812 5548 41852
rect 5588 41812 7564 41852
rect 7604 41812 7613 41852
rect 7843 41812 7852 41852
rect 7892 41812 8524 41852
rect 8564 41812 8573 41852
rect 18211 41812 18220 41852
rect 18260 41812 19084 41852
rect 19124 41812 19133 41852
rect 5539 41811 5597 41812
rect 7843 41811 7901 41812
rect 18211 41811 18269 41812
rect 16387 41768 16445 41769
rect 21424 41768 21504 41788
rect 4780 41728 5068 41768
rect 5108 41728 5117 41768
rect 7651 41728 7660 41768
rect 7700 41728 8908 41768
rect 8948 41728 8957 41768
rect 16387 41728 16396 41768
rect 16436 41728 21504 41768
rect 3139 41600 3197 41601
rect 1123 41560 1132 41600
rect 1172 41560 2380 41600
rect 2420 41560 2429 41600
rect 3054 41560 3148 41600
rect 3188 41560 3197 41600
rect 3331 41560 3340 41600
rect 3380 41560 4492 41600
rect 4532 41560 4541 41600
rect 3139 41559 3197 41560
rect 1123 41516 1181 41517
rect 4780 41516 4820 41728
rect 16387 41727 16445 41728
rect 21424 41708 21504 41728
rect 5827 41684 5885 41685
rect 11395 41684 11453 41685
rect 19459 41684 19517 41685
rect 5742 41644 5836 41684
rect 5876 41644 5885 41684
rect 8323 41644 8332 41684
rect 8372 41644 10444 41684
rect 10484 41644 10493 41684
rect 11395 41644 11404 41684
rect 11444 41644 11538 41684
rect 14467 41644 14476 41684
rect 14516 41644 18028 41684
rect 18068 41644 18077 41684
rect 19374 41644 19468 41684
rect 19508 41644 19517 41684
rect 5827 41643 5885 41644
rect 11395 41643 11453 41644
rect 19459 41643 19517 41644
rect 6595 41600 6653 41601
rect 4919 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 5305 41600
rect 6510 41560 6604 41600
rect 6644 41560 6653 41600
rect 6595 41559 6653 41560
rect 6787 41600 6845 41601
rect 7171 41600 7229 41601
rect 6787 41560 6796 41600
rect 6836 41560 6930 41600
rect 7086 41560 7180 41600
rect 7220 41560 7229 41600
rect 6787 41559 6845 41560
rect 7171 41559 7229 41560
rect 7363 41600 7421 41601
rect 7939 41600 7997 41601
rect 9283 41600 9341 41601
rect 9859 41600 9917 41601
rect 10243 41600 10301 41601
rect 11011 41600 11069 41601
rect 7363 41560 7372 41600
rect 7412 41560 7506 41600
rect 7854 41560 7948 41600
rect 7988 41560 7997 41600
rect 9198 41560 9292 41600
rect 9332 41560 9341 41600
rect 9774 41560 9868 41600
rect 9908 41560 9917 41600
rect 10158 41560 10252 41600
rect 10292 41560 10301 41600
rect 10926 41560 11020 41600
rect 11060 41560 11069 41600
rect 7363 41559 7421 41560
rect 7939 41559 7997 41560
rect 9283 41559 9341 41560
rect 9859 41559 9917 41560
rect 10243 41559 10301 41560
rect 11011 41559 11069 41560
rect 11491 41600 11549 41601
rect 11779 41600 11837 41601
rect 12259 41600 12317 41601
rect 11491 41560 11500 41600
rect 11540 41560 11596 41600
rect 11636 41560 11645 41600
rect 11779 41560 11788 41600
rect 11828 41560 11922 41600
rect 12259 41560 12268 41600
rect 12308 41560 12364 41600
rect 12404 41560 12413 41600
rect 15619 41560 15628 41600
rect 15668 41560 19372 41600
rect 19412 41560 19421 41600
rect 20039 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20425 41600
rect 11491 41559 11549 41560
rect 11779 41559 11837 41560
rect 12259 41559 12317 41560
rect 15715 41516 15773 41517
rect 17155 41516 17213 41517
rect 1123 41476 1132 41516
rect 1172 41476 4820 41516
rect 5635 41476 5644 41516
rect 5684 41476 7468 41516
rect 7508 41476 7517 41516
rect 15235 41476 15244 41516
rect 15284 41476 15724 41516
rect 15764 41476 15773 41516
rect 17070 41476 17164 41516
rect 17204 41476 17213 41516
rect 17923 41476 17932 41516
rect 17972 41476 19852 41516
rect 19892 41476 19901 41516
rect 1123 41475 1181 41476
rect 15715 41475 15773 41476
rect 17155 41475 17213 41476
rect 17251 41432 17309 41433
rect 21424 41432 21504 41452
rect 5059 41392 5068 41432
rect 5108 41392 15532 41432
rect 15572 41392 15581 41432
rect 16867 41392 16876 41432
rect 16916 41392 17260 41432
rect 17300 41392 17309 41432
rect 17731 41392 17740 41432
rect 17780 41392 19468 41432
rect 19508 41392 19517 41432
rect 21379 41392 21388 41432
rect 21428 41392 21504 41432
rect 17251 41391 17309 41392
rect 21424 41372 21504 41392
rect 18307 41348 18365 41349
rect 2500 41308 6412 41348
rect 6452 41308 6461 41348
rect 16483 41308 16492 41348
rect 16532 41308 17260 41348
rect 17300 41308 17309 41348
rect 18222 41308 18316 41348
rect 18356 41308 18365 41348
rect 2500 41096 2540 41308
rect 18307 41307 18365 41308
rect 3043 41264 3101 41265
rect 2851 41224 2860 41264
rect 2900 41224 3052 41264
rect 3092 41224 4492 41264
rect 4532 41224 4541 41264
rect 4963 41224 4972 41264
rect 5012 41224 5021 41264
rect 5251 41224 5260 41264
rect 5300 41224 11360 41264
rect 16291 41224 16300 41264
rect 16340 41224 17068 41264
rect 17108 41224 17117 41264
rect 3043 41223 3101 41224
rect 4972 41180 5012 41224
rect 7459 41180 7517 41181
rect 4972 41140 7468 41180
rect 7508 41140 7517 41180
rect 11320 41180 11360 41224
rect 15619 41180 15677 41181
rect 11320 41140 14476 41180
rect 14516 41140 14525 41180
rect 15427 41140 15436 41180
rect 15476 41140 15628 41180
rect 15668 41140 15677 41180
rect 7459 41139 7517 41140
rect 15619 41139 15677 41140
rect 16387 41180 16445 41181
rect 19651 41180 19709 41181
rect 16387 41140 16396 41180
rect 16436 41140 18892 41180
rect 18932 41140 18941 41180
rect 19566 41140 19660 41180
rect 19700 41140 19709 41180
rect 16387 41139 16445 41140
rect 19651 41139 19709 41140
rect 19843 41180 19901 41181
rect 19843 41140 19852 41180
rect 19892 41140 20044 41180
rect 20084 41140 20093 41180
rect 19843 41139 19901 41140
rect 20131 41096 20189 41097
rect 21424 41096 21504 41116
rect 2371 41056 2380 41096
rect 2420 41056 2540 41096
rect 3043 41056 3052 41096
rect 3092 41056 6412 41096
rect 6452 41056 6461 41096
rect 11971 41056 11980 41096
rect 12020 41056 15628 41096
rect 15668 41056 15677 41096
rect 16003 41056 16012 41096
rect 16052 41056 19756 41096
rect 19796 41056 19805 41096
rect 20131 41056 20140 41096
rect 20180 41056 21504 41096
rect 20131 41055 20189 41056
rect 21424 41036 21504 41056
rect 10819 41012 10877 41013
rect 15427 41012 15485 41013
rect 16387 41012 16445 41013
rect 16579 41012 16637 41013
rect 17059 41012 17117 41013
rect 17539 41012 17597 41013
rect 18307 41012 18365 41013
rect 19075 41012 19133 41013
rect 4675 40972 4684 41012
rect 4724 40972 5356 41012
rect 5396 40972 5405 41012
rect 8131 40972 8140 41012
rect 8180 40972 8332 41012
rect 8372 40972 10004 41012
rect 9964 40928 10004 40972
rect 10819 40972 10828 41012
rect 10868 40972 13804 41012
rect 13844 40972 13853 41012
rect 15342 40972 15436 41012
rect 15476 40972 15485 41012
rect 16099 40972 16108 41012
rect 16148 40972 16396 41012
rect 16436 40972 16445 41012
rect 16494 40972 16588 41012
rect 16628 40972 16637 41012
rect 16974 40972 17068 41012
rect 17108 40972 17117 41012
rect 17454 40972 17548 41012
rect 17588 40972 17597 41012
rect 18222 40972 18316 41012
rect 18356 40972 18365 41012
rect 18990 40972 19084 41012
rect 19124 40972 19133 41012
rect 10819 40971 10877 40972
rect 15427 40971 15485 40972
rect 16387 40971 16445 40972
rect 16579 40971 16637 40972
rect 17059 40971 17117 40972
rect 17539 40971 17597 40972
rect 18307 40971 18365 40972
rect 19075 40971 19133 40972
rect 1603 40888 1612 40928
rect 1652 40888 8716 40928
rect 8756 40888 8765 40928
rect 9955 40888 9964 40928
rect 10004 40888 10156 40928
rect 10196 40888 10732 40928
rect 10772 40888 19948 40928
rect 19988 40888 19997 40928
rect 3679 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 4065 40844
rect 4483 40804 4492 40844
rect 4532 40804 5644 40844
rect 5684 40804 5693 40844
rect 11491 40804 11500 40844
rect 11540 40804 12748 40844
rect 12788 40804 12797 40844
rect 14851 40804 14860 40844
rect 14900 40804 17876 40844
rect 18799 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 19185 40844
rect 12931 40760 12989 40761
rect 17731 40760 17789 40761
rect 1411 40720 1420 40760
rect 1460 40720 12940 40760
rect 12980 40720 12989 40760
rect 16963 40720 16972 40760
rect 17012 40720 17740 40760
rect 17780 40720 17789 40760
rect 17836 40760 17876 40804
rect 21424 40760 21504 40780
rect 17836 40720 19220 40760
rect 12931 40719 12989 40720
rect 17731 40719 17789 40720
rect 16579 40676 16637 40677
rect 19180 40676 19220 40720
rect 20140 40720 21504 40760
rect 6691 40636 6700 40676
rect 6740 40636 11360 40676
rect 12163 40636 12172 40676
rect 12212 40636 16300 40676
rect 16340 40636 16349 40676
rect 16579 40636 16588 40676
rect 16628 40636 18508 40676
rect 18548 40636 18557 40676
rect 19171 40636 19180 40676
rect 19220 40636 19229 40676
rect 11320 40592 11360 40636
rect 16579 40635 16637 40636
rect 12835 40592 12893 40593
rect 18115 40592 18173 40593
rect 19267 40592 19325 40593
rect 2092 40552 2956 40592
rect 2996 40552 3005 40592
rect 5251 40552 5260 40592
rect 5300 40552 10540 40592
rect 10580 40552 10589 40592
rect 11320 40552 12844 40592
rect 12884 40552 12893 40592
rect 13123 40552 13132 40592
rect 13172 40552 17356 40592
rect 17396 40552 17405 40592
rect 18030 40552 18124 40592
rect 18164 40552 18173 40592
rect 18979 40552 18988 40592
rect 19028 40552 19276 40592
rect 19316 40552 19325 40592
rect 259 40508 317 40509
rect 259 40468 268 40508
rect 308 40468 1804 40508
rect 1844 40468 1853 40508
rect 259 40467 317 40468
rect 1315 40424 1373 40425
rect 1230 40384 1324 40424
rect 1364 40384 1373 40424
rect 1315 40383 1373 40384
rect 1027 40300 1036 40340
rect 1076 40300 1996 40340
rect 2036 40300 2045 40340
rect 2092 40172 2132 40552
rect 12835 40551 12893 40552
rect 18115 40551 18173 40552
rect 19267 40551 19325 40552
rect 2275 40508 2333 40509
rect 5731 40508 5789 40509
rect 6499 40508 6557 40509
rect 2275 40468 2284 40508
rect 2324 40468 4780 40508
rect 4820 40468 4829 40508
rect 5731 40468 5740 40508
rect 5780 40468 6028 40508
rect 6068 40468 6077 40508
rect 6414 40468 6508 40508
rect 6548 40468 6557 40508
rect 2275 40467 2333 40468
rect 5731 40467 5789 40468
rect 6499 40467 6557 40468
rect 8803 40508 8861 40509
rect 8803 40468 8812 40508
rect 8852 40468 14036 40508
rect 14083 40468 14092 40508
rect 14132 40468 18316 40508
rect 18356 40468 18365 40508
rect 8803 40467 8861 40468
rect 2947 40424 3005 40425
rect 12643 40424 12701 40425
rect 2862 40384 2956 40424
rect 2996 40384 3005 40424
rect 3139 40384 3148 40424
rect 3188 40384 4876 40424
rect 4916 40384 4925 40424
rect 8707 40384 8716 40424
rect 8756 40384 10732 40424
rect 10772 40384 12652 40424
rect 12692 40384 12701 40424
rect 13996 40424 14036 40468
rect 16099 40424 16157 40425
rect 13996 40384 14284 40424
rect 14324 40384 14333 40424
rect 14851 40384 14860 40424
rect 14900 40384 15532 40424
rect 15572 40384 15581 40424
rect 15811 40384 15820 40424
rect 15860 40384 16108 40424
rect 16148 40384 16157 40424
rect 2947 40383 3005 40384
rect 12643 40383 12701 40384
rect 16099 40383 16157 40384
rect 16387 40424 16445 40425
rect 16963 40424 17021 40425
rect 17443 40424 17501 40425
rect 20140 40424 20180 40720
rect 21424 40700 21504 40720
rect 21424 40424 21504 40444
rect 16387 40384 16396 40424
rect 16436 40384 16628 40424
rect 16675 40384 16684 40424
rect 16724 40384 16972 40424
rect 17012 40384 17260 40424
rect 17300 40384 17309 40424
rect 17443 40384 17452 40424
rect 17492 40384 20180 40424
rect 21187 40384 21196 40424
rect 21236 40384 21504 40424
rect 16387 40383 16445 40384
rect 4195 40340 4253 40341
rect 2851 40300 2860 40340
rect 2900 40300 4204 40340
rect 4244 40300 4253 40340
rect 4195 40299 4253 40300
rect 6787 40340 6845 40341
rect 10147 40340 10205 40341
rect 16291 40340 16349 40341
rect 6787 40300 6796 40340
rect 6836 40300 6892 40340
rect 6932 40300 6941 40340
rect 10051 40300 10060 40340
rect 10100 40300 10156 40340
rect 10196 40300 10205 40340
rect 13603 40300 13612 40340
rect 13652 40300 13996 40340
rect 14036 40300 14045 40340
rect 14659 40300 14668 40340
rect 14708 40300 15436 40340
rect 15476 40300 16012 40340
rect 16052 40300 16300 40340
rect 16340 40300 16349 40340
rect 16588 40340 16628 40384
rect 16963 40383 17021 40384
rect 17443 40383 17501 40384
rect 21424 40364 21504 40384
rect 18403 40340 18461 40341
rect 16588 40300 17068 40340
rect 17108 40300 17117 40340
rect 18318 40300 18412 40340
rect 18452 40300 18461 40340
rect 6787 40299 6845 40300
rect 10147 40299 10205 40300
rect 16291 40299 16349 40300
rect 18403 40299 18461 40300
rect 18595 40340 18653 40341
rect 18595 40300 18604 40340
rect 18644 40300 20140 40340
rect 20180 40300 20189 40340
rect 18595 40299 18653 40300
rect 6979 40256 7037 40257
rect 15139 40256 15197 40257
rect 18499 40256 18557 40257
rect 6979 40216 6988 40256
rect 7028 40216 7084 40256
rect 7124 40216 7133 40256
rect 8323 40216 8332 40256
rect 8372 40216 8524 40256
rect 8564 40216 8573 40256
rect 10435 40216 10444 40256
rect 10484 40216 12884 40256
rect 15054 40216 15148 40256
rect 15188 40216 15197 40256
rect 15523 40216 15532 40256
rect 15572 40216 17356 40256
rect 17396 40216 17405 40256
rect 18499 40216 18508 40256
rect 18548 40216 18700 40256
rect 18740 40216 18749 40256
rect 6979 40215 7037 40216
rect 12844 40172 12884 40216
rect 15139 40215 15197 40216
rect 18499 40215 18557 40216
rect 15043 40172 15101 40173
rect 1987 40132 1996 40172
rect 2036 40132 2132 40172
rect 5923 40132 5932 40172
rect 5972 40132 12076 40172
rect 12116 40132 12125 40172
rect 12355 40132 12364 40172
rect 12404 40132 12788 40172
rect 12835 40132 12844 40172
rect 12884 40132 15052 40172
rect 15092 40132 15101 40172
rect 0 40088 80 40108
rect 12748 40088 12788 40132
rect 15043 40131 15101 40132
rect 15619 40172 15677 40173
rect 15619 40132 15628 40172
rect 15668 40132 18892 40172
rect 18932 40132 18941 40172
rect 15619 40131 15677 40132
rect 15715 40088 15773 40089
rect 21424 40088 21504 40108
rect 0 40048 4820 40088
rect 4919 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 5305 40088
rect 5635 40048 5644 40088
rect 5684 40048 6028 40088
rect 6068 40048 8840 40088
rect 12748 40048 13900 40088
rect 13940 40048 15092 40088
rect 0 40028 80 40048
rect 4780 40004 4820 40048
rect 8035 40004 8093 40005
rect 4780 39964 8044 40004
rect 8084 39964 8093 40004
rect 8800 40004 8840 40048
rect 15052 40004 15092 40048
rect 15715 40048 15724 40088
rect 15764 40048 18508 40088
rect 18548 40048 18557 40088
rect 20039 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20425 40088
rect 20803 40048 20812 40088
rect 20852 40048 21504 40088
rect 15715 40047 15773 40048
rect 21424 40028 21504 40048
rect 15235 40004 15293 40005
rect 16099 40004 16157 40005
rect 8800 39964 12172 40004
rect 12212 39964 12364 40004
rect 12404 39964 12413 40004
rect 12547 39964 12556 40004
rect 12596 39964 14188 40004
rect 14228 39964 14572 40004
rect 14612 39964 14956 40004
rect 14996 39964 15005 40004
rect 15052 39964 15244 40004
rect 15284 39964 15293 40004
rect 15427 39964 15436 40004
rect 15476 39964 15916 40004
rect 15956 39964 15965 40004
rect 16099 39964 16108 40004
rect 16148 39964 19468 40004
rect 19508 39964 19517 40004
rect 8035 39963 8093 39964
rect 15235 39963 15293 39964
rect 16099 39963 16157 39964
rect 16963 39920 17021 39921
rect 18691 39920 18749 39921
rect 3331 39880 3340 39920
rect 3380 39880 8908 39920
rect 8948 39880 11308 39920
rect 11348 39880 16300 39920
rect 16340 39880 16349 39920
rect 16878 39880 16972 39920
rect 17012 39880 17021 39920
rect 18606 39880 18700 39920
rect 18740 39880 18749 39920
rect 16963 39879 17021 39880
rect 18691 39879 18749 39880
rect 6787 39836 6845 39837
rect 19363 39836 19421 39837
rect 4867 39796 4876 39836
rect 4916 39796 5452 39836
rect 5492 39796 5501 39836
rect 6787 39796 6796 39836
rect 6836 39796 10636 39836
rect 10676 39796 10685 39836
rect 12067 39796 12076 39836
rect 12116 39796 15052 39836
rect 15092 39796 16588 39836
rect 16628 39796 16637 39836
rect 17731 39796 17740 39836
rect 17780 39796 19084 39836
rect 19124 39796 19372 39836
rect 19412 39796 19421 39836
rect 6787 39795 6845 39796
rect 19363 39795 19421 39796
rect 2179 39752 2237 39753
rect 1315 39712 1324 39752
rect 1364 39712 2188 39752
rect 2228 39712 2237 39752
rect 2179 39711 2237 39712
rect 2851 39752 2909 39753
rect 16387 39752 16445 39753
rect 21424 39752 21504 39772
rect 2851 39712 2860 39752
rect 2900 39712 3148 39752
rect 3188 39712 3197 39752
rect 7852 39712 12556 39752
rect 12596 39712 12605 39752
rect 13027 39712 13036 39752
rect 13076 39712 14956 39752
rect 14996 39712 15005 39752
rect 15235 39712 15244 39752
rect 15284 39712 16204 39752
rect 16244 39712 16253 39752
rect 16387 39712 16396 39752
rect 16436 39712 18068 39752
rect 18115 39712 18124 39752
rect 18164 39712 21504 39752
rect 2851 39711 2909 39712
rect 5347 39668 5405 39669
rect 7075 39668 7133 39669
rect 7852 39668 7892 39712
rect 16387 39711 16445 39712
rect 8515 39668 8573 39669
rect 2284 39628 5068 39668
rect 5108 39628 5117 39668
rect 5262 39628 5356 39668
rect 5396 39628 5405 39668
rect 6883 39628 6892 39668
rect 6932 39628 7084 39668
rect 7124 39628 7133 39668
rect 7843 39628 7852 39668
rect 7892 39628 7901 39668
rect 8419 39628 8428 39668
rect 8468 39628 8524 39668
rect 8564 39628 8573 39668
rect 0 39584 80 39604
rect 2284 39584 2324 39628
rect 5347 39627 5405 39628
rect 7075 39627 7133 39628
rect 8515 39627 8573 39628
rect 8899 39668 8957 39669
rect 17827 39668 17885 39669
rect 18028 39668 18068 39712
rect 21424 39692 21504 39712
rect 19939 39668 19997 39669
rect 8899 39628 8908 39668
rect 8948 39628 10924 39668
rect 10964 39628 16012 39668
rect 16052 39628 16061 39668
rect 17827 39628 17836 39668
rect 17876 39628 17932 39668
rect 17972 39628 17981 39668
rect 18028 39628 19660 39668
rect 19700 39628 19709 39668
rect 19939 39628 19948 39668
rect 19988 39628 20044 39668
rect 20084 39628 20093 39668
rect 8899 39627 8957 39628
rect 17827 39627 17885 39628
rect 19939 39627 19997 39628
rect 0 39544 2324 39584
rect 2371 39584 2429 39585
rect 12547 39584 12605 39585
rect 2371 39544 2380 39584
rect 2420 39544 2860 39584
rect 2900 39544 2909 39584
rect 5443 39544 5452 39584
rect 5492 39544 5972 39584
rect 7267 39544 7276 39584
rect 7316 39544 12556 39584
rect 12596 39544 12605 39584
rect 13507 39544 13516 39584
rect 13556 39544 20812 39584
rect 20852 39544 20861 39584
rect 0 39524 80 39544
rect 2371 39543 2429 39544
rect 5932 39500 5972 39544
rect 12547 39543 12605 39544
rect 8899 39500 8957 39501
rect 15811 39500 15869 39501
rect 16483 39500 16541 39501
rect 3628 39460 4972 39500
rect 5012 39460 5021 39500
rect 5932 39460 8908 39500
rect 8948 39460 8957 39500
rect 11971 39460 11980 39500
rect 12020 39460 12460 39500
rect 12500 39460 12509 39500
rect 14467 39460 14476 39500
rect 14516 39460 15244 39500
rect 15284 39460 15293 39500
rect 15726 39460 15820 39500
rect 15860 39460 15869 39500
rect 16398 39460 16492 39500
rect 16532 39460 16541 39500
rect 3628 39416 3668 39460
rect 8899 39459 8957 39460
rect 15811 39459 15869 39460
rect 16483 39459 16541 39460
rect 14563 39416 14621 39417
rect 21424 39416 21504 39436
rect 67 39376 76 39416
rect 116 39376 1420 39416
rect 1460 39376 3340 39416
rect 3380 39376 3389 39416
rect 3532 39376 3668 39416
rect 4195 39376 4204 39416
rect 4244 39376 4396 39416
rect 4436 39376 6508 39416
rect 6548 39376 6557 39416
rect 6787 39376 6796 39416
rect 6836 39376 7084 39416
rect 7124 39376 7133 39416
rect 14478 39376 14572 39416
rect 14612 39376 14621 39416
rect 14756 39376 14765 39416
rect 14805 39376 15572 39416
rect 15619 39376 15628 39416
rect 15668 39376 21504 39416
rect 2083 39248 2141 39249
rect 3532 39248 3572 39376
rect 14563 39375 14621 39376
rect 15532 39332 15572 39376
rect 21424 39356 21504 39376
rect 17635 39332 17693 39333
rect 3679 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 4065 39332
rect 4108 39292 10348 39332
rect 10388 39292 10397 39332
rect 12163 39292 12172 39332
rect 12212 39292 12556 39332
rect 12596 39292 12605 39332
rect 14275 39292 14284 39332
rect 14324 39292 15340 39332
rect 15380 39292 15389 39332
rect 15532 39292 17356 39332
rect 17396 39292 17405 39332
rect 17635 39292 17644 39332
rect 17684 39292 18316 39332
rect 18356 39292 18365 39332
rect 18799 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 19185 39332
rect 2083 39208 2092 39248
rect 2132 39208 3572 39248
rect 2083 39207 2141 39208
rect 4108 39164 4148 39292
rect 17635 39291 17693 39292
rect 16387 39248 16445 39249
rect 8035 39208 8044 39248
rect 8084 39208 16340 39248
rect 16300 39164 16340 39208
rect 16387 39208 16396 39248
rect 16436 39208 19564 39248
rect 19604 39208 19613 39248
rect 16387 39207 16445 39208
rect 17155 39164 17213 39165
rect 3619 39124 3628 39164
rect 3668 39124 4148 39164
rect 4387 39124 4396 39164
rect 4436 39124 4532 39164
rect 5059 39124 5068 39164
rect 5108 39124 5836 39164
rect 5876 39124 7276 39164
rect 7316 39124 7325 39164
rect 10627 39124 10636 39164
rect 10676 39124 11596 39164
rect 11636 39124 11645 39164
rect 12355 39124 12364 39164
rect 12404 39124 14284 39164
rect 14324 39124 14764 39164
rect 14804 39124 14813 39164
rect 16300 39124 17164 39164
rect 17204 39124 17213 39164
rect 0 39080 80 39100
rect 1315 39080 1373 39081
rect 1891 39080 1949 39081
rect 0 39040 76 39080
rect 116 39040 125 39080
rect 1315 39040 1324 39080
rect 1364 39040 1708 39080
rect 1748 39040 1757 39080
rect 1891 39040 1900 39080
rect 1940 39040 2476 39080
rect 2516 39040 2525 39080
rect 3523 39040 3532 39080
rect 3572 39040 4204 39080
rect 4244 39040 4253 39080
rect 0 39020 80 39040
rect 1315 39039 1373 39040
rect 1891 39039 1949 39040
rect 1795 38996 1853 38997
rect 4492 38996 4532 39124
rect 17155 39123 17213 39124
rect 10627 39080 10685 39081
rect 4963 39040 4972 39080
rect 5012 39040 5548 39080
rect 5588 39040 5597 39080
rect 6307 39040 6316 39080
rect 6356 39040 6604 39080
rect 6644 39040 6653 39080
rect 6883 39040 6892 39080
rect 6932 39040 7468 39080
rect 7508 39040 7517 39080
rect 10531 39040 10540 39080
rect 10580 39040 10636 39080
rect 10676 39040 10685 39080
rect 10627 39039 10685 39040
rect 12163 39080 12221 39081
rect 20131 39080 20189 39081
rect 21424 39080 21504 39100
rect 12163 39040 12172 39080
rect 12212 39040 13708 39080
rect 13748 39040 13757 39080
rect 13804 39040 13897 39080
rect 13937 39040 13946 39080
rect 15331 39040 15340 39080
rect 15380 39040 15476 39080
rect 15523 39040 15532 39080
rect 15572 39040 16876 39080
rect 16916 39040 16925 39080
rect 17059 39040 17068 39080
rect 17108 39040 18892 39080
rect 18932 39040 18941 39080
rect 20131 39040 20140 39080
rect 20180 39040 21504 39080
rect 12163 39039 12221 39040
rect 8803 38996 8861 38997
rect 13804 38996 13844 39040
rect 1315 38956 1324 38996
rect 1364 38956 1804 38996
rect 1844 38956 1853 38996
rect 3235 38956 3244 38996
rect 3284 38956 3293 38996
rect 4492 38956 8812 38996
rect 8852 38956 8861 38996
rect 13507 38956 13516 38996
rect 13556 38956 13844 38996
rect 1795 38955 1853 38956
rect 3043 38912 3101 38913
rect 2563 38872 2572 38912
rect 2612 38872 2956 38912
rect 2996 38872 3052 38912
rect 3092 38872 3101 38912
rect 3043 38871 3101 38872
rect 3244 38828 3284 38956
rect 8803 38955 8861 38956
rect 14947 38912 15005 38913
rect 3907 38872 3916 38912
rect 3956 38872 5260 38912
rect 5300 38872 5644 38912
rect 5684 38872 5693 38912
rect 6499 38872 6508 38912
rect 6548 38872 8140 38912
rect 8180 38872 8908 38912
rect 8948 38872 8957 38912
rect 9763 38872 9772 38912
rect 9812 38872 13132 38912
rect 13172 38872 13181 38912
rect 14284 38872 14668 38912
rect 14708 38872 14717 38912
rect 14851 38872 14860 38912
rect 14900 38872 14956 38912
rect 14996 38872 15005 38912
rect 14284 38828 14324 38872
rect 14947 38871 15005 38872
rect 15139 38912 15197 38913
rect 15436 38912 15476 39040
rect 20131 39039 20189 39040
rect 21424 39020 21504 39040
rect 15619 38996 15677 38997
rect 19555 38996 19613 38997
rect 15619 38956 15628 38996
rect 15668 38956 18123 38996
rect 18163 38956 18172 38996
rect 18499 38956 18508 38996
rect 18548 38956 19180 38996
rect 19220 38956 19229 38996
rect 19459 38956 19468 38996
rect 19508 38956 19564 38996
rect 19604 38956 19613 38996
rect 15619 38955 15677 38956
rect 19555 38955 19613 38956
rect 15139 38872 15148 38912
rect 15188 38872 15916 38912
rect 15956 38872 18796 38912
rect 18836 38872 18845 38912
rect 19267 38872 19276 38912
rect 19316 38872 19564 38912
rect 19604 38872 19613 38912
rect 15139 38871 15197 38872
rect 3244 38788 6892 38828
rect 6932 38788 6941 38828
rect 10339 38788 10348 38828
rect 10388 38788 14324 38828
rect 14371 38788 14380 38828
rect 14420 38788 15284 38828
rect 17635 38788 17644 38828
rect 17684 38788 17836 38828
rect 17876 38788 20044 38828
rect 20084 38788 20093 38828
rect 1987 38744 2045 38745
rect 3523 38744 3581 38745
rect 4291 38744 4349 38745
rect 4579 38744 4637 38745
rect 6307 38744 6365 38745
rect 6979 38744 7037 38745
rect 15139 38744 15197 38745
rect 1507 38704 1516 38744
rect 1556 38704 1996 38744
rect 2036 38704 2045 38744
rect 3438 38704 3532 38744
rect 3572 38704 3581 38744
rect 3811 38704 3820 38744
rect 3860 38704 4300 38744
rect 4340 38704 4349 38744
rect 4494 38704 4588 38744
rect 4628 38704 4637 38744
rect 1987 38703 2045 38704
rect 3523 38703 3581 38704
rect 4291 38703 4349 38704
rect 4579 38703 4637 38704
rect 5452 38704 6316 38744
rect 6356 38704 6988 38744
rect 7028 38704 9292 38744
rect 9332 38704 14996 38744
rect 15043 38704 15052 38744
rect 15092 38704 15148 38744
rect 15188 38704 15197 38744
rect 15244 38744 15284 38788
rect 16963 38744 17021 38745
rect 18403 38744 18461 38745
rect 20515 38744 20573 38745
rect 15244 38704 16972 38744
rect 17012 38704 17021 38744
rect 18318 38704 18412 38744
rect 18452 38704 18461 38744
rect 19267 38704 19276 38744
rect 19316 38704 20524 38744
rect 20564 38704 20573 38744
rect 5452 38660 5492 38704
rect 6307 38703 6365 38704
rect 6979 38703 7037 38704
rect 14956 38660 14996 38704
rect 15139 38703 15197 38704
rect 16963 38703 17021 38704
rect 18403 38703 18461 38704
rect 20515 38703 20573 38704
rect 20803 38744 20861 38745
rect 21424 38744 21504 38764
rect 20803 38704 20812 38744
rect 20852 38704 21504 38744
rect 20803 38703 20861 38704
rect 21424 38684 21504 38704
rect 18691 38660 18749 38661
rect 2500 38620 5492 38660
rect 5539 38620 5548 38660
rect 5588 38620 13612 38660
rect 13652 38620 13661 38660
rect 14956 38620 16396 38660
rect 16436 38620 16445 38660
rect 17827 38620 17836 38660
rect 17876 38620 18316 38660
rect 18356 38620 18365 38660
rect 18595 38620 18604 38660
rect 18644 38620 18700 38660
rect 18740 38620 18749 38660
rect 0 38576 80 38596
rect 2500 38576 2540 38620
rect 18691 38619 18749 38620
rect 18595 38576 18653 38577
rect 0 38536 2540 38576
rect 4195 38536 4204 38576
rect 4244 38536 4396 38576
rect 4436 38536 4445 38576
rect 4919 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 5305 38576
rect 5644 38536 9676 38576
rect 9716 38536 9725 38576
rect 10339 38536 10348 38576
rect 10388 38536 16588 38576
rect 16628 38536 16637 38576
rect 17731 38536 17740 38576
rect 17780 38536 18412 38576
rect 18452 38536 18461 38576
rect 18595 38536 18604 38576
rect 18644 38536 18700 38576
rect 18740 38536 18749 38576
rect 20039 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20425 38576
rect 0 38516 80 38536
rect 5644 38492 5684 38536
rect 18595 38535 18653 38536
rect 18499 38492 18557 38493
rect 4396 38452 5684 38492
rect 11971 38452 11980 38492
rect 12020 38452 13516 38492
rect 13556 38452 13565 38492
rect 14083 38452 14092 38492
rect 14132 38452 14476 38492
rect 14516 38452 14525 38492
rect 14851 38452 14860 38492
rect 14900 38452 15724 38492
rect 15764 38452 15773 38492
rect 15820 38452 18508 38492
rect 18548 38452 18557 38492
rect 1507 38368 1516 38408
rect 1556 38368 2380 38408
rect 2420 38368 2429 38408
rect 2755 38324 2813 38325
rect 2755 38284 2764 38324
rect 2804 38284 3340 38324
rect 3380 38284 3389 38324
rect 2755 38283 2813 38284
rect 4396 38240 4436 38452
rect 13315 38408 13373 38409
rect 15235 38408 15293 38409
rect 5932 38368 7660 38408
rect 7700 38368 8716 38408
rect 8756 38368 8765 38408
rect 12739 38368 12748 38408
rect 12788 38368 13324 38408
rect 13364 38368 14668 38408
rect 14708 38368 14717 38408
rect 15139 38368 15148 38408
rect 15188 38368 15244 38408
rect 15284 38368 15293 38408
rect 5827 38324 5885 38325
rect 5059 38284 5068 38324
rect 5108 38284 5836 38324
rect 5876 38284 5885 38324
rect 5827 38283 5885 38284
rect 5347 38240 5405 38241
rect 1891 38200 1900 38240
rect 1940 38200 2284 38240
rect 2324 38200 2333 38240
rect 3052 38200 3820 38240
rect 3860 38200 3869 38240
rect 4387 38200 4396 38240
rect 4436 38200 4445 38240
rect 4771 38200 4780 38240
rect 4820 38200 5356 38240
rect 5396 38200 5405 38240
rect 1507 38156 1565 38157
rect 1315 38116 1324 38156
rect 1364 38116 1516 38156
rect 1556 38116 1565 38156
rect 1507 38115 1565 38116
rect 1699 38156 1757 38157
rect 2563 38156 2621 38157
rect 3052 38156 3092 38200
rect 5347 38199 5405 38200
rect 1699 38116 1708 38156
rect 1748 38116 2188 38156
rect 2228 38116 2237 38156
rect 2563 38116 2572 38156
rect 2612 38116 3092 38156
rect 3331 38156 3389 38157
rect 3331 38116 3340 38156
rect 3380 38116 4588 38156
rect 4628 38116 4637 38156
rect 1699 38115 1757 38116
rect 2563 38115 2621 38116
rect 3331 38115 3389 38116
rect 0 38072 80 38092
rect 5932 38072 5972 38368
rect 13315 38367 13373 38368
rect 15235 38367 15293 38368
rect 13699 38324 13757 38325
rect 15820 38324 15860 38452
rect 18499 38451 18557 38452
rect 20131 38408 20189 38409
rect 21424 38408 21504 38428
rect 18595 38368 18604 38408
rect 18644 38368 19276 38408
rect 19316 38368 19564 38408
rect 19604 38368 19613 38408
rect 20131 38368 20140 38408
rect 20180 38368 21504 38408
rect 20131 38367 20189 38368
rect 21424 38348 21504 38368
rect 6019 38284 6028 38324
rect 6068 38284 12268 38324
rect 12308 38284 12317 38324
rect 13699 38284 13708 38324
rect 13748 38284 15860 38324
rect 16579 38324 16637 38325
rect 16963 38324 17021 38325
rect 19267 38324 19325 38325
rect 16579 38284 16588 38324
rect 16628 38284 16972 38324
rect 17012 38284 18891 38324
rect 18931 38284 18940 38324
rect 19075 38284 19084 38324
rect 19124 38284 19276 38324
rect 19316 38284 19325 38324
rect 13699 38283 13757 38284
rect 16579 38283 16637 38284
rect 16963 38283 17021 38284
rect 19267 38283 19325 38284
rect 6691 38240 6749 38241
rect 16099 38240 16157 38241
rect 6606 38200 6700 38240
rect 6740 38200 6749 38240
rect 8707 38200 8716 38240
rect 8756 38200 9332 38240
rect 10531 38200 10540 38240
rect 10580 38200 11692 38240
rect 11732 38200 11741 38240
rect 12355 38200 12364 38240
rect 12404 38200 12413 38240
rect 12547 38200 12556 38240
rect 12596 38200 14284 38240
rect 14324 38200 14333 38240
rect 14563 38200 14572 38240
rect 14612 38200 15052 38240
rect 15092 38200 15101 38240
rect 15427 38200 15436 38240
rect 15476 38200 16108 38240
rect 16148 38200 17740 38240
rect 17780 38200 17789 38240
rect 18499 38200 18508 38240
rect 18548 38200 19372 38240
rect 19412 38200 19421 38240
rect 6691 38199 6749 38200
rect 7459 38156 7517 38157
rect 9292 38156 9332 38200
rect 12364 38156 12404 38200
rect 16099 38199 16157 38200
rect 17251 38156 17309 38157
rect 6307 38116 6316 38156
rect 6356 38116 7468 38156
rect 7508 38116 7517 38156
rect 7459 38115 7517 38116
rect 8908 38116 9196 38156
rect 9236 38116 9245 38156
rect 9292 38116 12404 38156
rect 12748 38116 15188 38156
rect 15619 38116 15628 38156
rect 15668 38116 16204 38156
rect 16244 38116 16253 38156
rect 17251 38116 17260 38156
rect 17300 38116 19564 38156
rect 19604 38116 19613 38156
rect 6211 38072 6269 38073
rect 8908 38072 8948 38116
rect 12748 38072 12788 38116
rect 14179 38072 14237 38073
rect 15148 38072 15188 38116
rect 17251 38115 17309 38116
rect 15619 38072 15677 38073
rect 18691 38072 18749 38073
rect 0 38032 5972 38072
rect 6126 38032 6220 38072
rect 6260 38032 6269 38072
rect 6499 38032 6508 38072
rect 6548 38032 6892 38072
rect 6932 38032 6941 38072
rect 8899 38032 8908 38072
rect 8948 38032 8957 38072
rect 12739 38032 12748 38072
rect 12788 38032 12797 38072
rect 14094 38032 14188 38072
rect 14228 38032 14237 38072
rect 14659 38032 14668 38072
rect 14708 38032 14956 38072
rect 14996 38032 15005 38072
rect 15148 38032 15628 38072
rect 15668 38032 15677 38072
rect 15811 38032 15820 38072
rect 15860 38032 17452 38072
rect 17492 38032 17501 38072
rect 18412 38032 18700 38072
rect 18740 38032 18749 38072
rect 0 38012 80 38032
rect 6211 38031 6269 38032
rect 14179 38031 14237 38032
rect 15619 38031 15677 38032
rect 15043 37988 15101 37989
rect 17539 37988 17597 37989
rect 1795 37948 1804 37988
rect 1844 37948 10924 37988
rect 10964 37948 10973 37988
rect 12355 37948 12364 37988
rect 12404 37948 13132 37988
rect 13172 37948 13181 37988
rect 13507 37948 13516 37988
rect 13556 37948 14572 37988
rect 14612 37948 14621 37988
rect 15043 37948 15052 37988
rect 15092 37948 15532 37988
rect 15572 37948 16012 37988
rect 16052 37948 16061 37988
rect 16387 37948 16396 37988
rect 16436 37948 17548 37988
rect 17588 37948 17597 37988
rect 15043 37947 15101 37948
rect 17539 37947 17597 37948
rect 2467 37904 2525 37905
rect 2755 37904 2813 37905
rect 6979 37904 7037 37905
rect 12451 37904 12509 37905
rect 2467 37864 2476 37904
rect 2516 37864 2764 37904
rect 2804 37864 2813 37904
rect 6894 37864 6988 37904
rect 7028 37864 7037 37904
rect 9955 37864 9964 37904
rect 10004 37864 12460 37904
rect 12500 37864 12509 37904
rect 2467 37863 2525 37864
rect 2755 37863 2813 37864
rect 6979 37863 7037 37864
rect 12451 37863 12509 37864
rect 12643 37904 12701 37905
rect 14467 37904 14525 37905
rect 17827 37904 17885 37905
rect 18412 37904 18452 38032
rect 18691 38031 18749 38032
rect 20131 38072 20189 38073
rect 21424 38072 21504 38092
rect 20131 38032 20140 38072
rect 20180 38032 21504 38072
rect 20131 38031 20189 38032
rect 21424 38012 21504 38032
rect 18700 37948 19084 37988
rect 19124 37948 19133 37988
rect 12643 37864 12652 37904
rect 12692 37864 14036 37904
rect 12643 37863 12701 37864
rect 6307 37820 6365 37821
rect 13891 37820 13949 37821
rect 3139 37780 3148 37820
rect 3188 37780 3197 37820
rect 3679 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 4065 37820
rect 6307 37780 6316 37820
rect 6356 37780 6700 37820
rect 6740 37780 6749 37820
rect 10692 37780 10732 37820
rect 10772 37780 10781 37820
rect 13860 37780 13900 37820
rect 13940 37780 13949 37820
rect 13996 37820 14036 37864
rect 14467 37864 14476 37904
rect 14516 37864 17836 37904
rect 17876 37864 17885 37904
rect 18403 37864 18412 37904
rect 18452 37864 18461 37904
rect 14467 37863 14525 37864
rect 17827 37863 17885 37864
rect 15715 37820 15773 37821
rect 13996 37780 15724 37820
rect 15764 37780 16108 37820
rect 16148 37780 16157 37820
rect 1411 37652 1469 37653
rect 1326 37612 1420 37652
rect 1460 37612 1469 37652
rect 1411 37611 1469 37612
rect 1699 37652 1757 37653
rect 3148 37652 3188 37780
rect 6307 37779 6365 37780
rect 6979 37736 7037 37737
rect 10732 37736 10772 37780
rect 13891 37779 13949 37780
rect 15715 37779 15773 37780
rect 13900 37736 13940 37779
rect 15331 37736 15389 37737
rect 5731 37696 5740 37736
rect 5780 37696 6988 37736
rect 7028 37696 7037 37736
rect 7267 37696 7276 37736
rect 7316 37696 9524 37736
rect 10051 37696 10060 37736
rect 10100 37696 10772 37736
rect 12451 37696 12460 37736
rect 12500 37696 13940 37736
rect 15235 37696 15244 37736
rect 15284 37696 15340 37736
rect 15380 37696 15389 37736
rect 6979 37695 7037 37696
rect 1699 37612 1708 37652
rect 1748 37612 2708 37652
rect 3148 37612 3724 37652
rect 3764 37612 3773 37652
rect 4867 37612 4876 37652
rect 4916 37612 7468 37652
rect 7508 37612 7517 37652
rect 8323 37612 8332 37652
rect 8372 37612 9004 37652
rect 9044 37612 9053 37652
rect 9379 37612 9388 37652
rect 9428 37612 9437 37652
rect 1699 37611 1757 37612
rect 0 37568 80 37588
rect 2563 37568 2621 37569
rect 0 37528 2572 37568
rect 2612 37528 2621 37568
rect 2668 37568 2708 37612
rect 9388 37568 9428 37612
rect 2668 37528 4780 37568
rect 4820 37528 4829 37568
rect 4972 37528 9428 37568
rect 9484 37568 9524 37696
rect 15331 37695 15389 37696
rect 9955 37652 10013 37653
rect 13891 37652 13949 37653
rect 17827 37652 17885 37653
rect 18700 37652 18740 37948
rect 18799 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 19185 37820
rect 19267 37780 19276 37820
rect 19316 37780 19356 37820
rect 20044 37780 20236 37820
rect 20276 37780 20285 37820
rect 19276 37736 19316 37780
rect 20044 37736 20084 37780
rect 19276 37696 20084 37736
rect 20131 37736 20189 37737
rect 21424 37736 21504 37756
rect 20131 37696 20140 37736
rect 20180 37696 21504 37736
rect 20131 37695 20189 37696
rect 21424 37676 21504 37696
rect 21187 37652 21245 37653
rect 9571 37612 9580 37652
rect 9620 37612 9964 37652
rect 10004 37612 10013 37652
rect 10531 37612 10540 37652
rect 10580 37612 11500 37652
rect 11540 37612 11549 37652
rect 12835 37612 12844 37652
rect 12884 37612 13708 37652
rect 13748 37612 13757 37652
rect 13891 37612 13900 37652
rect 13940 37612 14034 37652
rect 14371 37612 14380 37652
rect 14420 37612 15340 37652
rect 15380 37612 15389 37652
rect 15523 37612 15532 37652
rect 15572 37612 16108 37652
rect 16148 37612 16157 37652
rect 17742 37612 17836 37652
rect 17876 37612 17885 37652
rect 18307 37612 18316 37652
rect 18356 37612 18740 37652
rect 19747 37612 19756 37652
rect 19796 37612 21196 37652
rect 21236 37612 21245 37652
rect 9955 37611 10013 37612
rect 13891 37611 13949 37612
rect 17827 37611 17885 37612
rect 21187 37611 21245 37612
rect 16387 37568 16445 37569
rect 9484 37528 10348 37568
rect 10388 37528 10397 37568
rect 10444 37528 15724 37568
rect 15764 37528 15773 37568
rect 16291 37528 16300 37568
rect 16340 37528 16396 37568
rect 16436 37528 16445 37568
rect 0 37508 80 37528
rect 2563 37527 2621 37528
rect 3523 37484 3581 37485
rect 4972 37484 5012 37528
rect 6019 37484 6077 37485
rect 9379 37484 9437 37485
rect 10444 37484 10484 37528
rect 16387 37527 16445 37528
rect 16771 37568 16829 37569
rect 18403 37568 18461 37569
rect 19363 37568 19421 37569
rect 16771 37528 16780 37568
rect 16820 37528 17396 37568
rect 17923 37528 17932 37568
rect 17972 37528 18412 37568
rect 18452 37528 18461 37568
rect 19171 37528 19180 37568
rect 19220 37528 19372 37568
rect 19412 37528 19421 37568
rect 16771 37527 16829 37528
rect 17356 37484 17396 37528
rect 18403 37527 18461 37528
rect 19363 37527 19421 37528
rect 20035 37484 20093 37485
rect 3523 37444 3532 37484
rect 3572 37444 3628 37484
rect 3668 37444 3677 37484
rect 4963 37444 4972 37484
rect 5012 37444 5021 37484
rect 6019 37444 6028 37484
rect 6068 37444 9100 37484
rect 9140 37444 9149 37484
rect 9294 37444 9388 37484
rect 9428 37444 9437 37484
rect 3523 37443 3581 37444
rect 6019 37443 6077 37444
rect 9379 37443 9437 37444
rect 9484 37444 10484 37484
rect 10723 37444 10732 37484
rect 10772 37444 12940 37484
rect 12980 37444 13516 37484
rect 13556 37444 13565 37484
rect 14755 37444 14764 37484
rect 14804 37444 16876 37484
rect 16916 37444 17260 37484
rect 17300 37444 17309 37484
rect 17356 37444 20044 37484
rect 20084 37444 20093 37484
rect 8995 37400 9053 37401
rect 9484 37400 9524 37444
rect 20035 37443 20093 37444
rect 20323 37400 20381 37401
rect 21424 37400 21504 37420
rect 5635 37360 5644 37400
rect 5684 37360 8812 37400
rect 8852 37360 8861 37400
rect 8995 37360 9004 37400
rect 9044 37360 9524 37400
rect 10243 37360 10252 37400
rect 10292 37360 11500 37400
rect 11540 37360 11549 37400
rect 12259 37360 12268 37400
rect 12308 37360 12317 37400
rect 13123 37360 13132 37400
rect 13172 37360 13708 37400
rect 13748 37360 13757 37400
rect 14083 37360 14092 37400
rect 14132 37360 14141 37400
rect 14275 37360 14284 37400
rect 14324 37360 14668 37400
rect 14708 37360 14717 37400
rect 15427 37360 15436 37400
rect 15476 37360 16300 37400
rect 16340 37360 19468 37400
rect 19508 37360 19517 37400
rect 19651 37360 19660 37400
rect 19700 37360 19948 37400
rect 19988 37360 19997 37400
rect 20323 37360 20332 37400
rect 20372 37360 21504 37400
rect 8995 37359 9053 37360
rect 12268 37316 12308 37360
rect 3628 37276 8620 37316
rect 8660 37276 8669 37316
rect 9004 37276 11116 37316
rect 11156 37276 12308 37316
rect 12355 37316 12413 37317
rect 14092 37316 14132 37360
rect 20323 37359 20381 37360
rect 21424 37340 21504 37360
rect 12355 37276 12364 37316
rect 12404 37276 12652 37316
rect 12692 37276 12701 37316
rect 14092 37276 17068 37316
rect 17108 37276 17117 37316
rect 18115 37276 18124 37316
rect 18164 37276 20044 37316
rect 20084 37276 20093 37316
rect 3043 37232 3101 37233
rect 3628 37232 3668 37276
rect 3811 37232 3869 37233
rect 4483 37232 4541 37233
rect 8899 37232 8957 37233
rect 931 37192 940 37232
rect 980 37192 1612 37232
rect 1652 37192 1661 37232
rect 3043 37192 3052 37232
rect 3092 37192 3244 37232
rect 3284 37192 3293 37232
rect 3619 37192 3628 37232
rect 3668 37192 3677 37232
rect 3726 37192 3820 37232
rect 3860 37192 3869 37232
rect 4398 37192 4492 37232
rect 4532 37192 4541 37232
rect 5155 37192 5164 37232
rect 5204 37192 8908 37232
rect 8948 37192 8957 37232
rect 3043 37191 3101 37192
rect 3811 37191 3869 37192
rect 4483 37191 4541 37192
rect 8899 37191 8957 37192
rect 3235 37148 3293 37149
rect 5635 37148 5693 37149
rect 9004 37148 9044 37276
rect 12355 37275 12413 37276
rect 13891 37232 13949 37233
rect 19267 37232 19325 37233
rect 9667 37192 9676 37232
rect 9716 37192 13324 37232
rect 13364 37192 13373 37232
rect 13891 37192 13900 37232
rect 13940 37192 14188 37232
rect 14228 37192 14237 37232
rect 14371 37192 14380 37232
rect 14420 37192 14764 37232
rect 14804 37192 14813 37232
rect 15619 37192 15628 37232
rect 15668 37192 16876 37232
rect 16916 37192 16925 37232
rect 17155 37192 17164 37232
rect 17204 37192 17452 37232
rect 17492 37192 17501 37232
rect 18883 37192 18892 37232
rect 18932 37192 19276 37232
rect 19316 37192 19325 37232
rect 19939 37192 19948 37232
rect 19988 37192 21004 37232
rect 21044 37192 21053 37232
rect 13891 37191 13949 37192
rect 19267 37191 19325 37192
rect 13987 37148 14045 37149
rect 17443 37148 17501 37149
rect 19276 37148 19316 37191
rect 2851 37108 2860 37148
rect 2900 37108 3244 37148
rect 3284 37108 5396 37148
rect 3235 37107 3293 37108
rect 0 37064 80 37084
rect 5356 37064 5396 37108
rect 5635 37108 5644 37148
rect 5684 37108 9044 37148
rect 9379 37108 9388 37148
rect 9428 37108 12652 37148
rect 12692 37108 12701 37148
rect 13795 37108 13804 37148
rect 13844 37108 13996 37148
rect 14036 37108 14045 37148
rect 15043 37108 15052 37148
rect 15092 37108 17260 37148
rect 17300 37108 17309 37148
rect 17443 37108 17452 37148
rect 17492 37108 19220 37148
rect 19276 37108 20716 37148
rect 20756 37108 20765 37148
rect 5635 37107 5693 37108
rect 13987 37107 14045 37108
rect 17443 37107 17501 37108
rect 15235 37064 15293 37065
rect 19180 37064 19220 37108
rect 20611 37064 20669 37065
rect 21424 37064 21504 37084
rect 0 37024 4684 37064
rect 4724 37024 4733 37064
rect 4919 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 5305 37064
rect 5356 37024 13940 37064
rect 14083 37024 14092 37064
rect 14132 37024 15244 37064
rect 15284 37024 18220 37064
rect 18260 37024 19084 37064
rect 19124 37024 19133 37064
rect 19180 37024 19660 37064
rect 19700 37024 19709 37064
rect 20039 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20425 37064
rect 20611 37024 20620 37064
rect 20660 37024 21504 37064
rect 0 37004 80 37024
rect 13900 36980 13940 37024
rect 15235 37023 15293 37024
rect 20611 37023 20669 37024
rect 21424 37004 21504 37024
rect 15331 36980 15389 36981
rect 18595 36980 18653 36981
rect 1507 36940 1516 36980
rect 1556 36940 4204 36980
rect 4244 36940 4253 36980
rect 8803 36940 8812 36980
rect 8852 36940 9772 36980
rect 9812 36940 10732 36980
rect 10772 36940 10781 36980
rect 11587 36940 11596 36980
rect 11636 36940 12692 36980
rect 13900 36940 15340 36980
rect 15380 36940 15389 36980
rect 16483 36940 16492 36980
rect 16532 36940 17836 36980
rect 17876 36940 17885 36980
rect 18595 36940 18604 36980
rect 18644 36940 19948 36980
rect 19988 36940 19997 36980
rect 2563 36896 2621 36897
rect 12652 36896 12692 36940
rect 15331 36939 15389 36940
rect 18595 36939 18653 36940
rect 14467 36896 14525 36897
rect 17923 36896 17981 36897
rect 2563 36856 2572 36896
rect 2612 36856 3052 36896
rect 3092 36856 3101 36896
rect 3235 36856 3244 36896
rect 3284 36856 12076 36896
rect 12116 36856 12125 36896
rect 12652 36856 14380 36896
rect 14420 36856 14476 36896
rect 14516 36856 14544 36896
rect 14668 36856 17932 36896
rect 17972 36856 17981 36896
rect 18115 36856 18124 36896
rect 18164 36856 18412 36896
rect 18452 36856 18461 36896
rect 19267 36856 19276 36896
rect 19316 36856 20716 36896
rect 20756 36856 20765 36896
rect 2563 36855 2621 36856
rect 14467 36855 14525 36856
rect 2659 36812 2717 36813
rect 12643 36812 12701 36813
rect 2659 36772 2668 36812
rect 2708 36772 3532 36812
rect 3572 36772 3581 36812
rect 3907 36772 3916 36812
rect 3956 36772 4588 36812
rect 4628 36772 4637 36812
rect 5155 36772 5164 36812
rect 5204 36772 5644 36812
rect 5684 36772 5693 36812
rect 8995 36772 9004 36812
rect 9044 36772 11360 36812
rect 11779 36772 11788 36812
rect 11828 36772 12652 36812
rect 12692 36772 12701 36812
rect 2659 36771 2717 36772
rect 10339 36728 10397 36729
rect 11320 36728 11360 36772
rect 12643 36771 12701 36772
rect 2467 36688 2476 36728
rect 2516 36688 3052 36728
rect 3092 36688 3340 36728
rect 3380 36688 3389 36728
rect 8131 36688 8140 36728
rect 8180 36688 10156 36728
rect 10196 36688 10205 36728
rect 10339 36688 10348 36728
rect 10388 36688 10444 36728
rect 10484 36688 10493 36728
rect 11320 36688 12172 36728
rect 12212 36688 12221 36728
rect 12355 36688 12364 36728
rect 12404 36688 12556 36728
rect 12596 36688 12605 36728
rect 10339 36687 10397 36688
rect 6979 36644 7037 36645
rect 9571 36644 9629 36645
rect 14668 36644 14708 36856
rect 17923 36855 17981 36856
rect 17059 36812 17117 36813
rect 16108 36772 16396 36812
rect 16436 36772 16445 36812
rect 17059 36772 17068 36812
rect 17108 36772 17356 36812
rect 17396 36772 17405 36812
rect 17635 36772 17644 36812
rect 17684 36772 18028 36812
rect 18068 36772 19180 36812
rect 19220 36772 19229 36812
rect 19843 36772 19852 36812
rect 19892 36772 19901 36812
rect 15331 36728 15389 36729
rect 15331 36688 15340 36728
rect 15380 36688 16012 36728
rect 16052 36688 16061 36728
rect 15331 36687 15389 36688
rect 16003 36644 16061 36645
rect 4003 36604 4012 36644
rect 4052 36604 4204 36644
rect 4244 36604 4628 36644
rect 5539 36604 5548 36644
rect 5588 36604 6988 36644
rect 7028 36604 7037 36644
rect 8803 36604 8812 36644
rect 8852 36604 9332 36644
rect 9486 36604 9580 36644
rect 9620 36604 9629 36644
rect 0 36560 80 36580
rect 3043 36560 3101 36561
rect 4588 36560 4628 36604
rect 6979 36603 7037 36604
rect 9292 36560 9332 36604
rect 9571 36603 9629 36604
rect 11320 36604 14708 36644
rect 14764 36604 16012 36644
rect 16052 36604 16061 36644
rect 11320 36560 11360 36604
rect 12451 36560 12509 36561
rect 14764 36560 14804 36604
rect 16003 36603 16061 36604
rect 16108 36560 16148 36772
rect 17059 36771 17117 36772
rect 19852 36728 19892 36772
rect 21424 36728 21504 36748
rect 16291 36688 16300 36728
rect 16340 36688 16972 36728
rect 17012 36688 18508 36728
rect 18548 36688 19564 36728
rect 19604 36688 19613 36728
rect 19852 36688 21504 36728
rect 21424 36668 21504 36688
rect 19459 36644 19517 36645
rect 16195 36604 16204 36644
rect 16244 36604 17068 36644
rect 17108 36604 18412 36644
rect 18452 36604 18461 36644
rect 19374 36604 19468 36644
rect 19508 36604 19517 36644
rect 19459 36603 19517 36604
rect 20131 36560 20189 36561
rect 0 36520 3052 36560
rect 3092 36520 3101 36560
rect 3427 36520 3436 36560
rect 3476 36520 4492 36560
rect 4532 36520 4541 36560
rect 4588 36520 8908 36560
rect 8948 36520 8957 36560
rect 9283 36520 9292 36560
rect 9332 36520 9341 36560
rect 9763 36520 9772 36560
rect 9812 36520 11360 36560
rect 11491 36520 11500 36560
rect 11540 36520 12076 36560
rect 12116 36520 12125 36560
rect 12451 36520 12460 36560
rect 12500 36520 14804 36560
rect 15043 36520 15052 36560
rect 15092 36520 15436 36560
rect 15476 36520 15485 36560
rect 15715 36520 15724 36560
rect 15764 36520 17260 36560
rect 17300 36520 18316 36560
rect 18356 36520 18365 36560
rect 18883 36520 18892 36560
rect 18932 36520 20140 36560
rect 20180 36520 20189 36560
rect 0 36500 80 36520
rect 3043 36519 3101 36520
rect 12451 36519 12509 36520
rect 20131 36519 20189 36520
rect 2563 36476 2621 36477
rect 2563 36436 2572 36476
rect 2612 36436 2706 36476
rect 2947 36436 2956 36476
rect 2996 36436 6028 36476
rect 6068 36436 6077 36476
rect 7363 36436 7372 36476
rect 7412 36436 8140 36476
rect 8180 36436 8189 36476
rect 8515 36436 8524 36476
rect 8564 36436 8716 36476
rect 8756 36436 10540 36476
rect 10580 36436 10589 36476
rect 11320 36436 18700 36476
rect 18740 36436 18749 36476
rect 2563 36435 2621 36436
rect 11320 36392 11360 36436
rect 15235 36392 15293 36393
rect 5539 36352 5548 36392
rect 5588 36352 11360 36392
rect 12163 36352 12172 36392
rect 12212 36352 12556 36392
rect 12596 36352 12605 36392
rect 13123 36352 13132 36392
rect 13172 36352 15244 36392
rect 15284 36352 15293 36392
rect 13132 36308 13172 36352
rect 15235 36351 15293 36352
rect 15715 36392 15773 36393
rect 17347 36392 17405 36393
rect 21424 36392 21504 36412
rect 15715 36352 15724 36392
rect 15764 36352 15916 36392
rect 15956 36352 15965 36392
rect 16291 36352 16300 36392
rect 16340 36352 16780 36392
rect 16820 36352 16829 36392
rect 17347 36352 17356 36392
rect 17396 36352 21504 36392
rect 15715 36351 15773 36352
rect 17347 36351 17405 36352
rect 21424 36332 21504 36352
rect 2179 36268 2188 36308
rect 2228 36268 2237 36308
rect 3679 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 4065 36308
rect 4588 36268 7892 36308
rect 7939 36268 7948 36308
rect 7988 36268 8236 36308
rect 8276 36268 8285 36308
rect 10243 36268 10252 36308
rect 10292 36268 13172 36308
rect 16003 36268 16012 36308
rect 16052 36268 18604 36308
rect 18644 36268 18653 36308
rect 18799 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 19185 36308
rect 0 36056 80 36076
rect 1219 36056 1277 36057
rect 2188 36056 2228 36268
rect 4588 36225 4628 36268
rect 3043 36224 3101 36225
rect 4579 36224 4637 36225
rect 3043 36184 3052 36224
rect 3092 36184 4588 36224
rect 4628 36184 4637 36224
rect 3043 36183 3101 36184
rect 4579 36183 4637 36184
rect 5068 36184 5356 36224
rect 5396 36184 5405 36224
rect 7363 36184 7372 36224
rect 7412 36184 7564 36224
rect 7604 36184 7613 36224
rect 2851 36140 2909 36141
rect 2851 36100 2860 36140
rect 2900 36100 3916 36140
rect 3956 36100 4204 36140
rect 4244 36100 4253 36140
rect 2851 36099 2909 36100
rect 5068 36056 5108 36184
rect 7852 36140 7892 36268
rect 11299 36224 11357 36225
rect 19363 36224 19421 36225
rect 8515 36184 8524 36224
rect 8564 36184 11116 36224
rect 11156 36184 11165 36224
rect 11299 36184 11308 36224
rect 11348 36184 12364 36224
rect 12404 36184 12413 36224
rect 13891 36184 13900 36224
rect 13940 36184 13949 36224
rect 15235 36184 15244 36224
rect 15284 36184 17164 36224
rect 17204 36184 17213 36224
rect 18691 36184 18700 36224
rect 18740 36184 19372 36224
rect 19412 36184 19421 36224
rect 11299 36183 11357 36184
rect 7852 36100 9196 36140
rect 9236 36100 9676 36140
rect 9716 36100 9725 36140
rect 10915 36100 10924 36140
rect 10964 36100 11212 36140
rect 11252 36100 11261 36140
rect 11587 36100 11596 36140
rect 11636 36100 11980 36140
rect 12020 36100 12029 36140
rect 12835 36100 12844 36140
rect 12884 36100 13708 36140
rect 13748 36100 13757 36140
rect 13699 36056 13757 36057
rect 0 36016 1228 36056
rect 1268 36016 1277 36056
rect 0 35996 80 36016
rect 1219 36015 1277 36016
rect 1612 36016 2228 36056
rect 2500 36016 5108 36056
rect 6787 36016 6796 36056
rect 6836 36016 7276 36056
rect 7316 36016 7325 36056
rect 10531 36016 10540 36056
rect 10580 36016 11116 36056
rect 11156 36016 11308 36056
rect 11348 36016 11357 36056
rect 11779 36016 11788 36056
rect 11828 36016 12556 36056
rect 12596 36016 13612 36056
rect 13652 36016 13708 36056
rect 13748 36016 13757 36056
rect 355 35972 413 35973
rect 1612 35972 1652 36016
rect 1891 35972 1949 35973
rect 355 35932 364 35972
rect 404 35932 1420 35972
rect 1460 35932 1469 35972
rect 1603 35932 1612 35972
rect 1652 35932 1661 35972
rect 1795 35932 1804 35972
rect 1844 35932 1900 35972
rect 1940 35932 2092 35972
rect 2132 35932 2141 35972
rect 355 35931 413 35932
rect 1891 35931 1949 35932
rect 1603 35888 1661 35889
rect 2500 35888 2540 36016
rect 13699 36015 13757 36016
rect 13900 35972 13940 36184
rect 19363 36183 19421 36184
rect 16291 36140 16349 36141
rect 17827 36140 17885 36141
rect 15427 36100 15436 36140
rect 15476 36100 15724 36140
rect 15764 36100 15773 36140
rect 16291 36100 16300 36140
rect 16340 36100 16780 36140
rect 16820 36100 16829 36140
rect 16963 36100 16972 36140
rect 17012 36100 17836 36140
rect 17876 36100 17885 36140
rect 19459 36100 19468 36140
rect 19508 36100 19756 36140
rect 19796 36100 19805 36140
rect 16291 36099 16349 36100
rect 17827 36099 17885 36100
rect 17059 36056 17117 36057
rect 16483 36016 16492 36056
rect 16532 36016 17068 36056
rect 17108 36016 17117 36056
rect 17059 36015 17117 36016
rect 18499 36056 18557 36057
rect 19939 36056 19997 36057
rect 18499 36016 18508 36056
rect 18548 36016 18557 36056
rect 18979 36016 18988 36056
rect 19028 36016 19948 36056
rect 19988 36016 19997 36056
rect 18499 36015 18557 36016
rect 19939 36015 19997 36016
rect 20131 36056 20189 36057
rect 21424 36056 21504 36076
rect 20131 36016 20140 36056
rect 20180 36016 21504 36056
rect 20131 36015 20189 36016
rect 18508 35972 18548 36015
rect 21424 35996 21504 36016
rect 2755 35932 2764 35972
rect 2804 35932 8524 35972
rect 8564 35932 8573 35972
rect 9667 35932 9676 35972
rect 9716 35932 13940 35972
rect 14275 35932 14284 35972
rect 14324 35932 18548 35972
rect 18595 35932 18604 35972
rect 18644 35932 19372 35972
rect 19412 35932 19421 35972
rect 20140 35932 20812 35972
rect 20852 35932 20861 35972
rect 1603 35848 1612 35888
rect 1652 35848 2540 35888
rect 2659 35888 2717 35889
rect 4771 35888 4829 35889
rect 8035 35888 8093 35889
rect 20140 35888 20180 35932
rect 2659 35848 2668 35888
rect 2708 35848 4396 35888
rect 4436 35848 4445 35888
rect 4771 35848 4780 35888
rect 4820 35848 5068 35888
rect 5108 35848 5117 35888
rect 5251 35848 5260 35888
rect 5300 35848 6220 35888
rect 6260 35848 6269 35888
rect 7555 35848 7564 35888
rect 7604 35848 7852 35888
rect 7892 35848 7901 35888
rect 8035 35848 8044 35888
rect 8084 35848 8236 35888
rect 8276 35848 9716 35888
rect 9763 35848 9772 35888
rect 9812 35848 10060 35888
rect 10100 35848 10109 35888
rect 10339 35848 10348 35888
rect 10388 35848 12844 35888
rect 12884 35848 12893 35888
rect 12940 35848 20180 35888
rect 1603 35847 1661 35848
rect 2659 35847 2717 35848
rect 4771 35847 4829 35848
rect 8035 35847 8093 35848
rect 2755 35804 2813 35805
rect 6019 35804 6077 35805
rect 9676 35804 9716 35848
rect 11299 35804 11357 35805
rect 1219 35764 1228 35804
rect 1268 35764 2516 35804
rect 2563 35764 2572 35804
rect 2612 35764 2764 35804
rect 2804 35764 2813 35804
rect 4003 35764 4012 35804
rect 4052 35764 4588 35804
rect 4628 35764 6028 35804
rect 6068 35764 6077 35804
rect 6979 35764 6988 35804
rect 7028 35764 8812 35804
rect 8852 35764 8861 35804
rect 9676 35764 11308 35804
rect 11348 35764 11357 35804
rect 2179 35720 2237 35721
rect 1987 35680 1996 35720
rect 2036 35680 2188 35720
rect 2228 35680 2237 35720
rect 2476 35720 2516 35764
rect 2755 35763 2813 35764
rect 6019 35763 6077 35764
rect 11299 35763 11357 35764
rect 12739 35804 12797 35805
rect 12940 35804 12980 35848
rect 16099 35804 16157 35805
rect 16387 35804 16445 35805
rect 12739 35764 12748 35804
rect 12788 35764 12980 35804
rect 16014 35764 16108 35804
rect 16148 35764 16157 35804
rect 16301 35764 16396 35804
rect 16436 35764 20236 35804
rect 20276 35764 20285 35804
rect 12739 35763 12797 35764
rect 16099 35763 16157 35764
rect 16387 35763 16445 35764
rect 3619 35720 3677 35721
rect 10819 35720 10877 35721
rect 2476 35680 3628 35720
rect 3668 35680 3677 35720
rect 4483 35680 4492 35720
rect 4532 35680 10828 35720
rect 10868 35680 10877 35720
rect 2179 35679 2237 35680
rect 3619 35679 3677 35680
rect 10819 35679 10877 35680
rect 12931 35720 12989 35721
rect 20707 35720 20765 35721
rect 12931 35680 12940 35720
rect 12980 35680 14284 35720
rect 14324 35680 14333 35720
rect 16867 35680 16876 35720
rect 16916 35680 17644 35720
rect 17684 35680 17693 35720
rect 19555 35680 19564 35720
rect 19604 35680 20716 35720
rect 20756 35680 20765 35720
rect 12931 35679 12989 35680
rect 20707 35679 20765 35680
rect 20899 35720 20957 35721
rect 21424 35720 21504 35740
rect 20899 35680 20908 35720
rect 20948 35680 21504 35720
rect 20899 35679 20957 35680
rect 21424 35660 21504 35680
rect 1411 35636 1469 35637
rect 1411 35596 1420 35636
rect 1460 35596 5548 35636
rect 5588 35596 5597 35636
rect 6019 35596 6028 35636
rect 6068 35596 7372 35636
rect 7412 35596 7421 35636
rect 10147 35596 10156 35636
rect 10196 35596 13036 35636
rect 13076 35596 13085 35636
rect 13411 35596 13420 35636
rect 13460 35596 13612 35636
rect 13652 35596 13661 35636
rect 14467 35596 14476 35636
rect 14516 35596 14860 35636
rect 14900 35596 14909 35636
rect 15139 35596 15148 35636
rect 15188 35596 15340 35636
rect 15380 35596 15389 35636
rect 15724 35596 21196 35636
rect 21236 35596 21245 35636
rect 1411 35595 1469 35596
rect 0 35552 80 35572
rect 15724 35552 15764 35596
rect 0 35512 4588 35552
rect 4628 35512 4637 35552
rect 4919 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 5305 35552
rect 6979 35512 6988 35552
rect 7028 35512 8332 35552
rect 8372 35512 8716 35552
rect 8756 35512 8765 35552
rect 9379 35512 9388 35552
rect 9428 35512 15764 35552
rect 17923 35512 17932 35552
rect 17972 35512 18412 35552
rect 18452 35512 19852 35552
rect 19892 35512 19901 35552
rect 20039 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20425 35552
rect 0 35492 80 35512
rect 7651 35468 7709 35469
rect 3331 35428 3340 35468
rect 3380 35428 5836 35468
rect 5876 35428 5885 35468
rect 7566 35428 7660 35468
rect 7700 35428 7709 35468
rect 7651 35427 7709 35428
rect 13219 35468 13277 35469
rect 16675 35468 16733 35469
rect 13219 35428 13228 35468
rect 13268 35428 16684 35468
rect 16724 35428 16733 35468
rect 13219 35427 13277 35428
rect 16675 35427 16733 35428
rect 17155 35384 17213 35385
rect 163 35344 172 35384
rect 212 35344 2380 35384
rect 2420 35344 2429 35384
rect 4003 35344 4012 35384
rect 4052 35344 6124 35384
rect 6164 35344 6173 35384
rect 7084 35344 7756 35384
rect 7796 35344 7805 35384
rect 9571 35344 9580 35384
rect 9620 35344 10964 35384
rect 11203 35344 11212 35384
rect 11252 35344 13516 35384
rect 13556 35344 13565 35384
rect 13699 35344 13708 35384
rect 13748 35344 17164 35384
rect 17204 35344 17213 35384
rect 4099 35300 4157 35301
rect 4099 35260 4108 35300
rect 4148 35260 4780 35300
rect 4820 35260 4829 35300
rect 5356 35260 5644 35300
rect 5684 35260 5693 35300
rect 5827 35260 5836 35300
rect 5876 35260 5885 35300
rect 6019 35260 6028 35300
rect 6068 35260 6077 35300
rect 6403 35260 6412 35300
rect 6452 35260 6461 35300
rect 4099 35259 4157 35260
rect 2179 35216 2237 35217
rect 4771 35216 4829 35217
rect 1315 35176 1324 35216
rect 1364 35176 1804 35216
rect 1844 35176 1853 35216
rect 2083 35176 2092 35216
rect 2132 35176 2188 35216
rect 2228 35176 2237 35216
rect 2467 35176 2476 35216
rect 2516 35176 4204 35216
rect 4244 35176 4253 35216
rect 4483 35176 4492 35216
rect 4532 35176 4780 35216
rect 4820 35176 4829 35216
rect 2179 35175 2237 35176
rect 4771 35175 4829 35176
rect 5251 35216 5309 35217
rect 5356 35216 5396 35260
rect 5836 35216 5876 35260
rect 5251 35176 5260 35216
rect 5300 35176 5396 35216
rect 5443 35176 5452 35216
rect 5492 35176 5876 35216
rect 5923 35176 5932 35216
rect 5972 35176 5981 35216
rect 5251 35175 5309 35176
rect 835 35132 893 35133
rect 4387 35132 4445 35133
rect 5932 35132 5972 35176
rect 835 35092 844 35132
rect 884 35092 1516 35132
rect 1556 35092 1565 35132
rect 2476 35092 2572 35132
rect 2612 35092 2640 35132
rect 3811 35092 3820 35132
rect 3860 35092 4396 35132
rect 4436 35092 4445 35132
rect 835 35091 893 35092
rect 0 35048 80 35068
rect 0 35008 1420 35048
rect 1460 35008 1469 35048
rect 0 34988 80 35008
rect 1891 34964 1949 34965
rect 1315 34924 1324 34964
rect 1364 34924 1900 34964
rect 1940 34924 1949 34964
rect 1891 34923 1949 34924
rect 2476 34880 2516 35092
rect 4387 35091 4445 35092
rect 4780 35092 5164 35132
rect 5204 35092 5213 35132
rect 5731 35092 5740 35132
rect 5780 35092 5972 35132
rect 3523 35048 3581 35049
rect 4780 35048 4820 35092
rect 6028 35048 6068 35260
rect 6412 35216 6452 35260
rect 6883 35216 6941 35217
rect 6412 35176 6892 35216
rect 6932 35176 6941 35216
rect 6883 35175 6941 35176
rect 7084 35133 7124 35344
rect 9955 35300 10013 35301
rect 10435 35300 10493 35301
rect 10819 35300 10877 35301
rect 9870 35260 9964 35300
rect 10004 35260 10013 35300
rect 10243 35260 10252 35300
rect 10292 35260 10444 35300
rect 10484 35260 10493 35300
rect 10734 35260 10828 35300
rect 10868 35260 10877 35300
rect 10924 35300 10964 35344
rect 17155 35343 17213 35344
rect 17635 35384 17693 35385
rect 21424 35384 21504 35404
rect 17635 35344 17644 35384
rect 17684 35344 21504 35384
rect 17635 35343 17693 35344
rect 21424 35324 21504 35344
rect 16003 35300 16061 35301
rect 18787 35300 18845 35301
rect 10924 35260 14572 35300
rect 14612 35260 14621 35300
rect 15918 35260 16012 35300
rect 16052 35260 16061 35300
rect 17155 35260 17164 35300
rect 17204 35260 17492 35300
rect 9955 35259 10013 35260
rect 10435 35259 10493 35260
rect 10819 35259 10877 35260
rect 16003 35259 16061 35260
rect 7747 35216 7805 35217
rect 14083 35216 14141 35217
rect 17452 35216 17492 35260
rect 18787 35260 18796 35300
rect 18836 35260 19180 35300
rect 19220 35260 19229 35300
rect 18787 35259 18845 35260
rect 7651 35176 7660 35216
rect 7700 35176 7756 35216
rect 7796 35176 8812 35216
rect 8852 35176 8861 35216
rect 8995 35176 9004 35216
rect 9044 35176 13228 35216
rect 13268 35176 13277 35216
rect 14083 35176 14092 35216
rect 14132 35176 16684 35216
rect 16724 35176 16733 35216
rect 17443 35176 17452 35216
rect 17492 35176 17501 35216
rect 18307 35176 18316 35216
rect 18356 35176 18892 35216
rect 18932 35176 18941 35216
rect 7747 35175 7805 35176
rect 14083 35175 14141 35176
rect 7075 35132 7133 35133
rect 14563 35132 14621 35133
rect 17827 35132 17885 35133
rect 6403 35092 6412 35132
rect 6452 35092 7084 35132
rect 7124 35092 7133 35132
rect 7843 35092 7852 35132
rect 7892 35092 13132 35132
rect 13172 35092 13324 35132
rect 13364 35092 13373 35132
rect 14563 35092 14572 35132
rect 14612 35092 14956 35132
rect 14996 35092 15244 35132
rect 15284 35092 15293 35132
rect 17827 35092 17836 35132
rect 17876 35092 19852 35132
rect 19892 35092 19901 35132
rect 7075 35091 7133 35092
rect 14563 35091 14621 35092
rect 17827 35091 17885 35092
rect 6307 35048 6365 35049
rect 9379 35048 9437 35049
rect 3438 35008 3532 35048
rect 3572 35008 4108 35048
rect 4148 35008 4820 35048
rect 5827 35008 5836 35048
rect 5876 35008 6068 35048
rect 6115 35008 6124 35048
rect 6164 35008 6316 35048
rect 6356 35008 6365 35048
rect 6499 35008 6508 35048
rect 6548 35008 7372 35048
rect 7412 35008 7421 35048
rect 7651 35008 7660 35048
rect 7700 35008 8044 35048
rect 8084 35008 8093 35048
rect 8803 35008 8812 35048
rect 8852 35008 9388 35048
rect 9428 35008 9437 35048
rect 3523 35007 3581 35008
rect 6307 35007 6365 35008
rect 9379 35007 9437 35008
rect 10051 35048 10109 35049
rect 13507 35048 13565 35049
rect 10051 35008 10060 35048
rect 10100 35008 13516 35048
rect 13556 35008 13565 35048
rect 10051 35007 10109 35008
rect 13507 35007 13565 35008
rect 17731 35048 17789 35049
rect 21424 35048 21504 35068
rect 17731 35008 17740 35048
rect 17780 35008 19468 35048
rect 19508 35008 19517 35048
rect 20140 35008 21504 35048
rect 17731 35007 17789 35008
rect 3043 34964 3101 34965
rect 16387 34964 16445 34965
rect 20140 34964 20180 35008
rect 21424 34988 21504 35008
rect 3043 34924 3052 34964
rect 3092 34924 3340 34964
rect 3380 34924 3389 34964
rect 4972 34924 11308 34964
rect 11348 34924 11357 34964
rect 13507 34924 13516 34964
rect 13556 34924 14956 34964
rect 14996 34924 15005 34964
rect 15139 34924 15148 34964
rect 15188 34924 15628 34964
rect 15668 34924 15677 34964
rect 16387 34924 16396 34964
rect 16436 34924 20180 34964
rect 3043 34923 3101 34924
rect 4972 34880 5012 34924
rect 16387 34923 16445 34924
rect 5635 34880 5693 34881
rect 10051 34880 10109 34881
rect 1891 34840 1900 34880
rect 1940 34840 5012 34880
rect 5443 34840 5452 34880
rect 5492 34840 5644 34880
rect 5684 34840 5693 34880
rect 5923 34840 5932 34880
rect 5972 34840 7084 34880
rect 7124 34840 7133 34880
rect 10051 34840 10060 34880
rect 10100 34840 19660 34880
rect 19700 34840 19709 34880
rect 5635 34839 5693 34840
rect 10051 34839 10109 34840
rect 2179 34796 2237 34797
rect 11107 34796 11165 34797
rect 11875 34796 11933 34797
rect 2179 34756 2188 34796
rect 2228 34756 2764 34796
rect 2804 34756 2813 34796
rect 3679 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 4065 34796
rect 4195 34756 4204 34796
rect 4244 34756 10924 34796
rect 10964 34756 10973 34796
rect 11022 34756 11116 34796
rect 11156 34756 11165 34796
rect 11395 34756 11404 34796
rect 11444 34756 11884 34796
rect 11924 34756 17068 34796
rect 17108 34756 17117 34796
rect 18799 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 19185 34796
rect 2179 34755 2237 34756
rect 11107 34755 11165 34756
rect 11875 34755 11933 34756
rect 2947 34712 3005 34713
rect 20131 34712 20189 34713
rect 21424 34712 21504 34732
rect 1315 34672 1324 34712
rect 1364 34672 2956 34712
rect 2996 34672 6508 34712
rect 6548 34672 6557 34712
rect 9091 34672 9100 34712
rect 9140 34672 11500 34712
rect 11540 34672 11549 34712
rect 11884 34672 18412 34712
rect 18452 34672 18461 34712
rect 20131 34672 20140 34712
rect 20180 34672 21504 34712
rect 2947 34671 3005 34672
rect 1603 34628 1661 34629
rect 4675 34628 4733 34629
rect 6691 34628 6749 34629
rect 11884 34628 11924 34672
rect 20131 34671 20189 34672
rect 21424 34652 21504 34672
rect 13411 34628 13469 34629
rect 1507 34588 1516 34628
rect 1556 34588 1612 34628
rect 1652 34588 1661 34628
rect 4387 34588 4396 34628
rect 4436 34588 4684 34628
rect 4724 34588 4733 34628
rect 5443 34588 5452 34628
rect 5492 34588 6604 34628
rect 6644 34588 6700 34628
rect 6740 34588 6768 34628
rect 10051 34588 10060 34628
rect 10100 34588 11924 34628
rect 11971 34588 11980 34628
rect 12020 34588 12172 34628
rect 12212 34588 12221 34628
rect 13411 34588 13420 34628
rect 13460 34588 13612 34628
rect 13652 34588 13661 34628
rect 14467 34588 14476 34628
rect 14516 34588 15052 34628
rect 15092 34588 15101 34628
rect 15523 34588 15532 34628
rect 15572 34588 16108 34628
rect 16148 34588 16157 34628
rect 1603 34587 1661 34588
rect 4675 34587 4733 34588
rect 6691 34587 6749 34588
rect 13411 34587 13469 34588
rect 0 34544 80 34564
rect 4483 34544 4541 34545
rect 17635 34544 17693 34545
rect 19939 34544 19997 34545
rect 0 34504 4492 34544
rect 4532 34504 4541 34544
rect 5251 34504 5260 34544
rect 5300 34504 12268 34544
rect 12308 34504 12317 34544
rect 13699 34504 13708 34544
rect 13748 34504 17644 34544
rect 17684 34504 18700 34544
rect 18740 34504 18749 34544
rect 19854 34504 19948 34544
rect 19988 34504 19997 34544
rect 0 34484 80 34504
rect 4483 34503 4541 34504
rect 17635 34503 17693 34504
rect 19939 34503 19997 34504
rect 4867 34460 4925 34461
rect 6787 34460 6845 34461
rect 4867 34420 4876 34460
rect 4916 34420 6796 34460
rect 6836 34420 6845 34460
rect 4867 34419 4925 34420
rect 6787 34419 6845 34420
rect 7555 34460 7613 34461
rect 8419 34460 8477 34461
rect 7555 34420 7564 34460
rect 7604 34420 8180 34460
rect 8334 34420 8428 34460
rect 8468 34420 8477 34460
rect 7555 34419 7613 34420
rect 4771 34376 4829 34377
rect 5635 34376 5693 34377
rect 7267 34376 7325 34377
rect 8035 34376 8093 34377
rect 2947 34336 2956 34376
rect 2996 34336 3244 34376
rect 3284 34336 3293 34376
rect 4771 34336 4780 34376
rect 4820 34336 4914 34376
rect 5635 34336 5644 34376
rect 5684 34336 6988 34376
rect 7028 34336 7037 34376
rect 7267 34336 7276 34376
rect 7316 34336 8044 34376
rect 8084 34336 8093 34376
rect 8140 34376 8180 34420
rect 8419 34419 8477 34420
rect 9772 34420 10060 34460
rect 10100 34420 10109 34460
rect 11491 34420 11500 34460
rect 11540 34420 17932 34460
rect 17972 34420 17981 34460
rect 9772 34376 9812 34420
rect 8140 34336 9812 34376
rect 9955 34376 10013 34377
rect 11683 34376 11741 34377
rect 17443 34376 17501 34377
rect 20515 34376 20573 34377
rect 21424 34376 21504 34396
rect 9955 34336 9964 34376
rect 10004 34336 10924 34376
rect 10964 34336 10973 34376
rect 11395 34336 11404 34376
rect 11444 34336 11692 34376
rect 11732 34336 11741 34376
rect 11971 34336 11980 34376
rect 12020 34336 14188 34376
rect 14228 34336 14237 34376
rect 17443 34336 17452 34376
rect 17492 34336 17548 34376
rect 17588 34336 17597 34376
rect 20515 34336 20524 34376
rect 20564 34336 21504 34376
rect 4771 34335 4829 34336
rect 5635 34335 5693 34336
rect 7267 34335 7325 34336
rect 8035 34335 8093 34336
rect 9955 34335 10013 34336
rect 11683 34335 11741 34336
rect 17443 34335 17501 34336
rect 20515 34335 20573 34336
rect 21424 34316 21504 34336
rect 3619 34292 3677 34293
rect 13027 34292 13085 34293
rect 16483 34292 16541 34293
rect 3523 34252 3532 34292
rect 3572 34252 3628 34292
rect 3668 34252 7756 34292
rect 7796 34252 7805 34292
rect 8131 34252 8140 34292
rect 8180 34252 11020 34292
rect 11060 34252 11069 34292
rect 12942 34252 13036 34292
rect 13076 34252 13708 34292
rect 13748 34252 13757 34292
rect 14083 34252 14092 34292
rect 14132 34252 15436 34292
rect 15476 34252 16492 34292
rect 16532 34252 16541 34292
rect 16675 34252 16684 34292
rect 16724 34252 16972 34292
rect 17012 34252 17164 34292
rect 17204 34252 18316 34292
rect 18356 34252 19852 34292
rect 19892 34252 19901 34292
rect 3619 34251 3677 34252
rect 13027 34251 13085 34252
rect 16483 34251 16541 34252
rect 1891 34208 1949 34209
rect 6115 34208 6173 34209
rect 10051 34208 10109 34209
rect 10723 34208 10781 34209
rect 15139 34208 15197 34209
rect 1891 34168 1900 34208
rect 1940 34168 3148 34208
rect 3188 34168 3197 34208
rect 4195 34168 4204 34208
rect 4244 34168 6124 34208
rect 6164 34168 6173 34208
rect 7363 34168 7372 34208
rect 7412 34168 8812 34208
rect 8852 34168 8861 34208
rect 9966 34168 10060 34208
rect 10100 34168 10109 34208
rect 10339 34168 10348 34208
rect 10388 34168 10732 34208
rect 10772 34168 10781 34208
rect 10915 34168 10924 34208
rect 10964 34168 14860 34208
rect 14900 34168 14909 34208
rect 15054 34168 15148 34208
rect 15188 34168 15197 34208
rect 16867 34168 16876 34208
rect 16916 34168 17548 34208
rect 17588 34168 17597 34208
rect 19075 34168 19084 34208
rect 19124 34168 20140 34208
rect 20180 34168 20189 34208
rect 1891 34167 1949 34168
rect 6115 34167 6173 34168
rect 10051 34167 10109 34168
rect 10723 34167 10781 34168
rect 15139 34167 15197 34168
rect 10627 34124 10685 34125
rect 12067 34124 12125 34125
rect 15715 34124 15773 34125
rect 460 34084 5452 34124
rect 5492 34084 5501 34124
rect 5731 34084 5740 34124
rect 5780 34084 10636 34124
rect 10676 34084 12076 34124
rect 12116 34084 12125 34124
rect 13219 34084 13228 34124
rect 13268 34084 15724 34124
rect 15764 34084 18028 34124
rect 18068 34084 18077 34124
rect 0 34040 80 34060
rect 460 34040 500 34084
rect 10627 34083 10685 34084
rect 12067 34083 12125 34084
rect 15715 34083 15773 34084
rect 3523 34040 3581 34041
rect 5923 34040 5981 34041
rect 21424 34040 21504 34060
rect 0 34000 500 34040
rect 547 34000 556 34040
rect 596 34000 3532 34040
rect 3572 34000 3581 34040
rect 4919 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 5305 34040
rect 5635 34000 5644 34040
rect 5684 34000 5932 34040
rect 5972 34000 8468 34040
rect 10531 34000 10540 34040
rect 10580 34000 11692 34040
rect 11732 34000 11741 34040
rect 12355 34000 12364 34040
rect 12404 34000 13996 34040
rect 14036 34000 16300 34040
rect 16340 34000 16349 34040
rect 20039 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20425 34040
rect 20803 34000 20812 34040
rect 20852 34000 21504 34040
rect 0 33980 80 34000
rect 3523 33999 3581 34000
rect 5923 33999 5981 34000
rect 6883 33872 6941 33873
rect 7651 33872 7709 33873
rect 1699 33832 1708 33872
rect 1748 33832 3820 33872
rect 3860 33832 3869 33872
rect 4675 33832 4684 33872
rect 4724 33832 6892 33872
rect 6932 33832 7660 33872
rect 7700 33832 7709 33872
rect 6883 33831 6941 33832
rect 7651 33831 7709 33832
rect 7555 33788 7613 33789
rect 1612 33748 5740 33788
rect 5780 33748 5789 33788
rect 7075 33748 7084 33788
rect 7124 33748 7276 33788
rect 7316 33748 7325 33788
rect 7470 33748 7564 33788
rect 7604 33748 7613 33788
rect 8428 33788 8468 34000
rect 21424 33980 21504 34000
rect 16195 33956 16253 33957
rect 8515 33916 8524 33956
rect 8564 33916 14228 33956
rect 14275 33916 14284 33956
rect 14324 33916 15244 33956
rect 15284 33916 16204 33956
rect 16244 33916 16492 33956
rect 16532 33916 16541 33956
rect 17635 33916 17644 33956
rect 17684 33916 20276 33956
rect 14188 33872 14228 33916
rect 16195 33915 16253 33916
rect 16579 33872 16637 33873
rect 20236 33872 20276 33916
rect 21379 33872 21437 33873
rect 9283 33832 9292 33872
rect 9332 33832 9580 33872
rect 9620 33832 9629 33872
rect 10147 33832 10156 33872
rect 10196 33832 10444 33872
rect 10484 33832 10493 33872
rect 10627 33832 10636 33872
rect 10676 33832 11308 33872
rect 11348 33832 11357 33872
rect 12067 33832 12076 33872
rect 12116 33832 13420 33872
rect 13460 33832 13469 33872
rect 14188 33832 16588 33872
rect 16628 33832 16637 33872
rect 19363 33832 19372 33872
rect 19412 33832 19756 33872
rect 19796 33832 19805 33872
rect 20236 33832 21388 33872
rect 21428 33832 21437 33872
rect 16579 33831 16637 33832
rect 21379 33831 21437 33832
rect 13315 33788 13373 33789
rect 19555 33788 19613 33789
rect 8428 33748 13324 33788
rect 13364 33748 13373 33788
rect 15619 33748 15628 33788
rect 15668 33748 19564 33788
rect 19604 33748 19613 33788
rect 1612 33704 1652 33748
rect 7555 33747 7613 33748
rect 13315 33747 13373 33748
rect 19555 33747 19613 33748
rect 10531 33704 10589 33705
rect 17923 33704 17981 33705
rect 21424 33704 21504 33724
rect 739 33664 748 33704
rect 788 33664 1612 33704
rect 1652 33664 1661 33704
rect 4099 33664 4108 33704
rect 4148 33664 4780 33704
rect 4820 33664 4829 33704
rect 5827 33664 5836 33704
rect 5876 33664 6508 33704
rect 6548 33664 6557 33704
rect 7363 33664 7372 33704
rect 7412 33664 8236 33704
rect 8276 33664 8285 33704
rect 8515 33664 8524 33704
rect 8564 33664 9292 33704
rect 9332 33664 9341 33704
rect 10446 33664 10540 33704
rect 10580 33664 10589 33704
rect 11760 33664 11788 33704
rect 11828 33664 11884 33704
rect 11924 33664 11933 33704
rect 13603 33664 13612 33704
rect 13652 33664 14284 33704
rect 14324 33664 14333 33704
rect 14755 33664 14764 33704
rect 14804 33664 17644 33704
rect 17684 33664 17693 33704
rect 17923 33664 17932 33704
rect 17972 33664 18604 33704
rect 18644 33664 18653 33704
rect 20707 33664 20716 33704
rect 20756 33664 21504 33704
rect 1228 33580 1900 33620
rect 1940 33580 1949 33620
rect 2947 33580 2956 33620
rect 2996 33580 3436 33620
rect 3476 33580 3485 33620
rect 0 33536 80 33556
rect 1228 33536 1268 33580
rect 4108 33536 4148 33664
rect 10531 33663 10589 33664
rect 4579 33620 4637 33621
rect 11884 33620 11924 33664
rect 17923 33663 17981 33664
rect 21424 33644 21504 33664
rect 4579 33580 4588 33620
rect 4628 33580 4876 33620
rect 4916 33580 4925 33620
rect 6211 33580 6220 33620
rect 6260 33580 6604 33620
rect 6644 33580 6653 33620
rect 7267 33580 7276 33620
rect 7316 33580 9772 33620
rect 9812 33580 10156 33620
rect 10196 33580 11924 33620
rect 13315 33620 13373 33621
rect 19459 33620 19517 33621
rect 13315 33580 13324 33620
rect 13364 33580 17588 33620
rect 19374 33580 19468 33620
rect 19508 33580 19517 33620
rect 4579 33579 4637 33580
rect 13315 33579 13373 33580
rect 0 33496 1268 33536
rect 1315 33496 1324 33536
rect 1364 33496 1996 33536
rect 2036 33496 4148 33536
rect 6691 33536 6749 33537
rect 10531 33536 10589 33537
rect 17548 33536 17588 33580
rect 19459 33579 19517 33580
rect 19843 33536 19901 33537
rect 6691 33496 6700 33536
rect 6740 33496 10540 33536
rect 10580 33496 10589 33536
rect 14179 33496 14188 33536
rect 14228 33496 14668 33536
rect 14708 33496 14717 33536
rect 15427 33496 15436 33536
rect 15476 33496 17356 33536
rect 17396 33496 17405 33536
rect 17539 33496 17548 33536
rect 17588 33496 17597 33536
rect 18019 33496 18028 33536
rect 18068 33496 18604 33536
rect 18644 33496 18653 33536
rect 19843 33496 19852 33536
rect 19892 33496 20140 33536
rect 20180 33496 20189 33536
rect 0 33476 80 33496
rect 6691 33495 6749 33496
rect 10531 33495 10589 33496
rect 19843 33495 19901 33496
rect 2563 33452 2621 33453
rect 15427 33452 15485 33453
rect 1603 33412 1612 33452
rect 1652 33412 2092 33452
rect 2132 33412 2141 33452
rect 2563 33412 2572 33452
rect 2612 33412 3148 33452
rect 3188 33412 3197 33452
rect 6307 33412 6316 33452
rect 6356 33412 8236 33452
rect 8276 33412 8285 33452
rect 10339 33412 10348 33452
rect 10388 33412 10924 33452
rect 10964 33412 10973 33452
rect 15427 33412 15436 33452
rect 15476 33412 15916 33452
rect 15956 33412 15965 33452
rect 19939 33412 19948 33452
rect 19988 33412 21196 33452
rect 21236 33412 21245 33452
rect 2563 33411 2621 33412
rect 15427 33411 15485 33412
rect 10915 33368 10973 33369
rect 21424 33368 21504 33388
rect 2500 33328 2956 33368
rect 2996 33328 8908 33368
rect 8948 33328 8957 33368
rect 10915 33328 10924 33368
rect 10964 33328 15628 33368
rect 15668 33328 15677 33368
rect 20611 33328 20620 33368
rect 20660 33328 21504 33368
rect 2500 33284 2540 33328
rect 10915 33327 10973 33328
rect 21424 33308 21504 33328
rect 6787 33284 6845 33285
rect 16291 33284 16349 33285
rect 17731 33284 17789 33285
rect 67 33244 76 33284
rect 116 33244 2540 33284
rect 3679 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 4065 33284
rect 6787 33244 6796 33284
rect 6836 33244 12652 33284
rect 12692 33244 12701 33284
rect 13315 33244 13324 33284
rect 13364 33244 15148 33284
rect 15188 33244 15820 33284
rect 15860 33244 15869 33284
rect 16206 33244 16300 33284
rect 16340 33244 16349 33284
rect 17646 33244 17740 33284
rect 17780 33244 17789 33284
rect 18799 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 19185 33284
rect 6787 33243 6845 33244
rect 16291 33243 16349 33244
rect 17731 33243 17789 33244
rect 12451 33200 12509 33201
rect 5539 33160 5548 33200
rect 5588 33160 8428 33200
rect 8468 33160 8477 33200
rect 12355 33160 12364 33200
rect 12404 33160 12460 33200
rect 12500 33160 12509 33200
rect 12451 33159 12509 33160
rect 15907 33200 15965 33201
rect 15907 33160 15916 33200
rect 15956 33160 19756 33200
rect 19796 33160 19805 33200
rect 15907 33159 15965 33160
rect 2275 33116 2333 33117
rect 6115 33116 6173 33117
rect 7747 33116 7805 33117
rect 13795 33116 13853 33117
rect 18499 33116 18557 33117
rect 2275 33076 2284 33116
rect 2324 33076 2380 33116
rect 2420 33076 2429 33116
rect 6115 33076 6124 33116
rect 6164 33076 6700 33116
rect 6740 33076 6749 33116
rect 7555 33076 7564 33116
rect 7604 33076 7756 33116
rect 7796 33076 8044 33116
rect 8084 33076 8093 33116
rect 13710 33076 13804 33116
rect 13844 33076 13853 33116
rect 14179 33076 14188 33116
rect 14228 33076 17068 33116
rect 17108 33076 17117 33116
rect 18403 33076 18412 33116
rect 18452 33076 18508 33116
rect 18548 33076 18557 33116
rect 2275 33075 2333 33076
rect 6115 33075 6173 33076
rect 7747 33075 7805 33076
rect 13795 33075 13853 33076
rect 18499 33075 18557 33076
rect 19651 33116 19709 33117
rect 19651 33076 19660 33116
rect 19700 33076 20140 33116
rect 20180 33076 20189 33116
rect 19651 33075 19709 33076
rect 0 33032 80 33052
rect 6499 33032 6557 33033
rect 11971 33032 12029 33033
rect 21424 33032 21504 33052
rect 0 32992 76 33032
rect 116 32992 125 33032
rect 1795 32992 1804 33032
rect 1844 32992 1940 33032
rect 2755 32992 2764 33032
rect 2804 32992 2900 33032
rect 3235 32992 3244 33032
rect 3284 32992 3532 33032
rect 3572 32992 3581 33032
rect 4675 32992 4684 33032
rect 4724 32992 6508 33032
rect 6548 32992 6557 33032
rect 7651 32992 7660 33032
rect 7700 32992 7709 33032
rect 11971 32992 11980 33032
rect 12020 32992 12844 33032
rect 12884 32992 16876 33032
rect 16916 32992 16925 33032
rect 19651 32992 19660 33032
rect 19700 32992 19709 33032
rect 20515 32992 20524 33032
rect 20564 32992 21504 33032
rect 0 32972 80 32992
rect 1219 32824 1228 32864
rect 1268 32824 1804 32864
rect 1844 32824 1853 32864
rect 1900 32696 1940 32992
rect 2179 32948 2237 32949
rect 2094 32908 2188 32948
rect 2228 32908 2237 32948
rect 2179 32907 2237 32908
rect 2275 32864 2333 32865
rect 2755 32864 2813 32865
rect 2275 32824 2284 32864
rect 2324 32824 2764 32864
rect 2804 32824 2813 32864
rect 2275 32823 2333 32824
rect 2755 32823 2813 32824
rect 2860 32780 2900 32992
rect 6499 32991 6557 32992
rect 6691 32948 6749 32949
rect 3139 32908 3148 32948
rect 3188 32908 6700 32948
rect 6740 32908 6749 32948
rect 7660 32948 7700 32992
rect 11971 32991 12029 32992
rect 14275 32948 14333 32949
rect 7660 32908 7948 32948
rect 7988 32908 8852 32948
rect 9859 32908 9868 32948
rect 9908 32908 12116 32948
rect 14190 32908 14284 32948
rect 14324 32908 14333 32948
rect 15331 32908 15340 32948
rect 15380 32908 18892 32948
rect 18932 32908 18941 32948
rect 6691 32907 6749 32908
rect 3235 32864 3293 32865
rect 3150 32824 3244 32864
rect 3284 32824 3293 32864
rect 3235 32823 3293 32824
rect 3523 32864 3581 32865
rect 8227 32864 8285 32865
rect 3523 32824 3532 32864
rect 3572 32824 3724 32864
rect 3764 32824 3773 32864
rect 7747 32824 7756 32864
rect 7796 32824 8236 32864
rect 8276 32824 8285 32864
rect 3523 32823 3581 32824
rect 8227 32823 8285 32824
rect 8419 32864 8477 32865
rect 8812 32864 8852 32908
rect 11587 32864 11645 32865
rect 12076 32864 12116 32908
rect 14275 32907 14333 32908
rect 8419 32824 8428 32864
rect 8468 32824 8620 32864
rect 8660 32824 8669 32864
rect 8803 32824 8812 32864
rect 8852 32824 8861 32864
rect 9187 32824 9196 32864
rect 9236 32824 10636 32864
rect 10676 32824 10685 32864
rect 11502 32824 11596 32864
rect 11636 32824 11645 32864
rect 12067 32824 12076 32864
rect 12116 32824 12125 32864
rect 12259 32824 12268 32864
rect 12308 32824 13036 32864
rect 13076 32824 13085 32864
rect 13699 32824 13708 32864
rect 13748 32824 13996 32864
rect 14036 32824 15628 32864
rect 15668 32824 16300 32864
rect 16340 32824 16349 32864
rect 16771 32824 16780 32864
rect 16820 32824 19084 32864
rect 19124 32824 19133 32864
rect 8419 32823 8477 32824
rect 11587 32823 11645 32824
rect 4675 32780 4733 32781
rect 6211 32780 6269 32781
rect 14083 32780 14141 32781
rect 2764 32740 2900 32780
rect 3052 32740 4396 32780
rect 4436 32740 4445 32780
rect 4675 32740 4684 32780
rect 4724 32740 6220 32780
rect 6260 32740 6269 32780
rect 6787 32740 6796 32780
rect 6836 32740 8276 32780
rect 12163 32740 12172 32780
rect 12212 32740 13132 32780
rect 13172 32740 13181 32780
rect 14083 32740 14092 32780
rect 14132 32740 14188 32780
rect 14228 32740 14237 32780
rect 15235 32740 15244 32780
rect 15284 32740 15820 32780
rect 15860 32740 15869 32780
rect 16675 32740 16684 32780
rect 16724 32740 19372 32780
rect 19412 32740 19421 32780
rect 1900 32656 2188 32696
rect 2228 32656 2237 32696
rect 2764 32612 2804 32740
rect 3052 32696 3092 32740
rect 4675 32739 4733 32740
rect 6211 32739 6269 32740
rect 8236 32696 8276 32740
rect 14083 32739 14141 32740
rect 19660 32696 19700 32992
rect 21424 32972 21504 32992
rect 3043 32656 3052 32696
rect 3092 32656 3101 32696
rect 4195 32656 4204 32696
rect 4244 32656 4876 32696
rect 4916 32656 4925 32696
rect 8227 32656 8236 32696
rect 8276 32656 8285 32696
rect 10435 32656 10444 32696
rect 10484 32656 10828 32696
rect 10868 32656 10877 32696
rect 12355 32656 12364 32696
rect 12404 32656 12556 32696
rect 12596 32656 12605 32696
rect 14947 32656 14956 32696
rect 14996 32656 19700 32696
rect 21187 32696 21245 32697
rect 21424 32696 21504 32716
rect 21187 32656 21196 32696
rect 21236 32656 21504 32696
rect 21187 32655 21245 32656
rect 21424 32636 21504 32656
rect 6211 32612 6269 32613
rect 11107 32612 11165 32613
rect 16003 32612 16061 32613
rect 16291 32612 16349 32613
rect 17059 32612 17117 32613
rect 2755 32572 2764 32612
rect 2804 32572 2813 32612
rect 3331 32572 3340 32612
rect 3380 32572 4492 32612
rect 4532 32572 6220 32612
rect 6260 32572 6269 32612
rect 7459 32572 7468 32612
rect 7508 32572 9004 32612
rect 9044 32572 9053 32612
rect 11107 32572 11116 32612
rect 11156 32572 16012 32612
rect 16052 32572 16061 32612
rect 16206 32572 16300 32612
rect 16340 32572 16349 32612
rect 16579 32572 16588 32612
rect 16628 32572 17068 32612
rect 17108 32572 17452 32612
rect 17492 32572 17501 32612
rect 6211 32571 6269 32572
rect 11107 32571 11165 32572
rect 16003 32571 16061 32572
rect 16291 32571 16349 32572
rect 17059 32571 17117 32572
rect 0 32528 80 32548
rect 6307 32528 6365 32529
rect 6979 32528 7037 32529
rect 7747 32528 7805 32529
rect 11299 32528 11357 32529
rect 13891 32528 13949 32529
rect 0 32488 76 32528
rect 116 32488 125 32528
rect 4919 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 5305 32528
rect 6307 32488 6316 32528
rect 6356 32488 6508 32528
rect 6548 32488 6557 32528
rect 6979 32488 6988 32528
rect 7028 32488 7756 32528
rect 7796 32488 7805 32528
rect 8131 32488 8140 32528
rect 8180 32488 8524 32528
rect 8564 32488 8573 32528
rect 11203 32488 11212 32528
rect 11252 32488 11308 32528
rect 11348 32488 11357 32528
rect 12739 32488 12748 32528
rect 12788 32488 13036 32528
rect 13076 32488 13900 32528
rect 13940 32488 13949 32528
rect 14659 32488 14668 32528
rect 14708 32488 14717 32528
rect 15811 32488 15820 32528
rect 15860 32488 16396 32528
rect 16436 32488 16445 32528
rect 16492 32488 18604 32528
rect 18644 32488 18653 32528
rect 20039 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20425 32528
rect 0 32468 80 32488
rect 6307 32487 6365 32488
rect 6979 32487 7037 32488
rect 7747 32487 7805 32488
rect 11299 32487 11357 32488
rect 13891 32487 13949 32488
rect 14275 32444 14333 32445
rect 14668 32444 14708 32488
rect 16492 32444 16532 32488
rect 1603 32404 1612 32444
rect 1652 32404 1661 32444
rect 1891 32404 1900 32444
rect 1940 32404 6124 32444
rect 6164 32404 7180 32444
rect 7220 32404 7564 32444
rect 7604 32404 7613 32444
rect 11395 32404 11404 32444
rect 11444 32404 11884 32444
rect 11924 32404 11933 32444
rect 12931 32404 12940 32444
rect 12980 32404 13132 32444
rect 13172 32404 13181 32444
rect 14275 32404 14284 32444
rect 14324 32404 14380 32444
rect 14420 32404 14429 32444
rect 14668 32404 16532 32444
rect 16963 32404 16972 32444
rect 17012 32404 17548 32444
rect 17588 32404 17597 32444
rect 20 32320 76 32360
rect 116 32320 125 32360
rect 20 32192 60 32320
rect 1315 32276 1373 32277
rect 1230 32236 1324 32276
rect 1364 32236 1373 32276
rect 1315 32235 1373 32236
rect 1612 32192 1652 32404
rect 14275 32403 14333 32404
rect 3331 32360 3389 32361
rect 7555 32360 7613 32361
rect 16003 32360 16061 32361
rect 21424 32360 21504 32380
rect 2275 32320 2284 32360
rect 2324 32320 2476 32360
rect 2516 32320 2525 32360
rect 3235 32320 3244 32360
rect 3284 32320 3340 32360
rect 3380 32320 3389 32360
rect 3907 32320 3916 32360
rect 3956 32320 7564 32360
rect 7604 32320 7613 32360
rect 9955 32320 9964 32360
rect 10004 32320 10540 32360
rect 10580 32320 10589 32360
rect 11107 32320 11116 32360
rect 11156 32320 14764 32360
rect 14804 32320 14813 32360
rect 16003 32320 16012 32360
rect 16052 32320 16146 32360
rect 16195 32320 16204 32360
rect 16244 32320 17932 32360
rect 17972 32320 17981 32360
rect 19747 32320 19756 32360
rect 19796 32320 21504 32360
rect 3331 32319 3389 32320
rect 7555 32319 7613 32320
rect 16003 32319 16061 32320
rect 21424 32300 21504 32320
rect 11971 32276 12029 32277
rect 18211 32276 18269 32277
rect 18691 32276 18749 32277
rect 5443 32236 5452 32276
rect 5492 32236 6028 32276
rect 6068 32236 6077 32276
rect 6691 32236 6700 32276
rect 6740 32236 8620 32276
rect 8660 32236 8669 32276
rect 10819 32236 10828 32276
rect 10868 32236 11980 32276
rect 12020 32236 12029 32276
rect 11971 32235 12029 32236
rect 13708 32236 18220 32276
rect 18260 32236 18269 32276
rect 18595 32236 18604 32276
rect 18644 32236 18700 32276
rect 18740 32236 18749 32276
rect 4195 32192 4253 32193
rect 8611 32192 8669 32193
rect 11107 32192 11165 32193
rect 20 32152 2132 32192
rect 1411 32108 1469 32109
rect 1315 32068 1324 32108
rect 1364 32068 1420 32108
rect 1460 32068 1469 32108
rect 1411 32067 1469 32068
rect 1603 32108 1661 32109
rect 2092 32108 2132 32152
rect 4195 32152 4204 32192
rect 4244 32152 4972 32192
rect 5012 32152 5021 32192
rect 5251 32152 5260 32192
rect 5300 32152 6988 32192
rect 7028 32152 7468 32192
rect 7508 32152 7517 32192
rect 8515 32152 8524 32192
rect 8564 32152 8620 32192
rect 8660 32152 8669 32192
rect 9091 32152 9100 32192
rect 9140 32152 9292 32192
rect 9332 32152 11116 32192
rect 11156 32152 11165 32192
rect 11491 32152 11500 32192
rect 11540 32152 12652 32192
rect 12692 32152 12701 32192
rect 13315 32152 13324 32192
rect 13364 32152 13373 32192
rect 4195 32151 4253 32152
rect 8611 32151 8669 32152
rect 11107 32151 11165 32152
rect 1603 32068 1612 32108
rect 1652 32068 1708 32108
rect 1748 32068 1757 32108
rect 2083 32068 2092 32108
rect 2132 32068 2141 32108
rect 4099 32068 4108 32108
rect 4148 32068 4492 32108
rect 4532 32068 10060 32108
rect 10100 32068 10109 32108
rect 10531 32068 10540 32108
rect 10580 32068 11692 32108
rect 11732 32068 12172 32108
rect 12212 32068 12748 32108
rect 12788 32068 12797 32108
rect 12931 32068 12940 32108
rect 12980 32068 13228 32108
rect 13268 32068 13277 32108
rect 1603 32067 1661 32068
rect 0 32024 80 32044
rect 7171 32024 7229 32025
rect 12940 32024 12980 32068
rect 0 31984 1612 32024
rect 1652 31984 1661 32024
rect 2755 31984 2764 32024
rect 2804 31984 5932 32024
rect 5972 31984 6508 32024
rect 6548 31984 6557 32024
rect 7075 31984 7084 32024
rect 7124 31984 7180 32024
rect 7220 31984 7229 32024
rect 7555 31984 7564 32024
rect 7604 31984 8332 32024
rect 8372 31984 8381 32024
rect 10627 31984 10636 32024
rect 10676 31984 12980 32024
rect 0 31964 80 31984
rect 7171 31983 7229 31984
rect 3043 31940 3101 31941
rect 3523 31940 3581 31941
rect 7555 31940 7613 31941
rect 11587 31940 11645 31941
rect 13324 31940 13364 32152
rect 13708 32024 13748 32236
rect 18211 32235 18269 32236
rect 18691 32235 18749 32236
rect 13987 32152 13996 32192
rect 14036 32152 14572 32192
rect 14612 32152 14621 32192
rect 14755 32152 14764 32192
rect 14804 32152 14813 32192
rect 15043 32152 15052 32192
rect 15092 32152 15724 32192
rect 15764 32152 15773 32192
rect 17059 32152 17068 32192
rect 17108 32152 17836 32192
rect 17876 32152 17885 32192
rect 18211 32152 18220 32192
rect 18260 32152 18269 32192
rect 14764 32108 14804 32152
rect 18220 32108 18260 32152
rect 14275 32068 14284 32108
rect 14324 32068 14333 32108
rect 14764 32068 15140 32108
rect 16387 32068 16396 32108
rect 16436 32068 18260 32108
rect 14284 32024 14324 32068
rect 15100 32024 15140 32068
rect 21424 32024 21504 32044
rect 13699 31984 13708 32024
rect 13748 31984 13757 32024
rect 13987 31984 13996 32024
rect 14036 31984 14324 32024
rect 14371 31984 14380 32024
rect 14420 31984 14956 32024
rect 14996 31984 15005 32024
rect 15100 31984 15436 32024
rect 15476 31984 15485 32024
rect 18019 31984 18028 32024
rect 18068 31984 19372 32024
rect 19412 31984 19421 32024
rect 19843 31984 19852 32024
rect 19892 31984 21504 32024
rect 21424 31964 21504 31984
rect 3043 31900 3052 31940
rect 3092 31900 3532 31940
rect 3572 31900 5356 31940
rect 5396 31900 5405 31940
rect 6979 31900 6988 31940
rect 7028 31900 7564 31940
rect 7604 31900 7613 31940
rect 8131 31900 8140 31940
rect 8180 31900 11596 31940
rect 11636 31900 13364 31940
rect 14563 31940 14621 31941
rect 16675 31940 16733 31941
rect 14563 31900 14572 31940
rect 14612 31900 14668 31940
rect 14708 31900 14717 31940
rect 15523 31900 15532 31940
rect 15572 31900 16684 31940
rect 16724 31900 16733 31940
rect 16963 31900 16972 31940
rect 17012 31900 17452 31940
rect 17492 31900 17501 31940
rect 3043 31899 3101 31900
rect 3523 31899 3581 31900
rect 7555 31899 7613 31900
rect 11587 31899 11645 31900
rect 14563 31899 14621 31900
rect 16675 31899 16733 31900
rect 4387 31816 4396 31856
rect 4436 31816 14476 31856
rect 14516 31816 14525 31856
rect 14755 31816 14764 31856
rect 14804 31816 18604 31856
rect 18644 31816 18653 31856
rect 9955 31772 10013 31773
rect 3679 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 4065 31772
rect 4867 31732 4876 31772
rect 4916 31732 9964 31772
rect 10004 31732 10013 31772
rect 12451 31732 12460 31772
rect 12500 31732 17068 31772
rect 17108 31732 17117 31772
rect 18799 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 19185 31772
rect 9955 31731 10013 31732
rect 20131 31688 20189 31689
rect 21424 31688 21504 31708
rect 652 31648 6892 31688
rect 6932 31648 6941 31688
rect 8419 31648 8428 31688
rect 8468 31648 19756 31688
rect 19796 31648 19805 31688
rect 20131 31648 20140 31688
rect 20180 31648 21504 31688
rect 0 31520 80 31540
rect 652 31520 692 31648
rect 20131 31647 20189 31648
rect 21424 31628 21504 31648
rect 13795 31604 13853 31605
rect 16387 31604 16445 31605
rect 18691 31604 18749 31605
rect 4579 31564 4588 31604
rect 4628 31564 6220 31604
rect 6260 31564 6269 31604
rect 11203 31564 11212 31604
rect 11252 31564 13612 31604
rect 13652 31564 13661 31604
rect 13795 31564 13804 31604
rect 13844 31564 16396 31604
rect 16436 31564 16445 31604
rect 16675 31564 16684 31604
rect 16724 31564 18412 31604
rect 18452 31564 18461 31604
rect 18691 31564 18700 31604
rect 18740 31564 18796 31604
rect 18836 31564 18845 31604
rect 13795 31563 13853 31564
rect 16387 31563 16445 31564
rect 5443 31520 5501 31521
rect 7555 31520 7613 31521
rect 8803 31520 8861 31521
rect 9091 31520 9149 31521
rect 10435 31520 10493 31521
rect 15715 31520 15773 31521
rect 16684 31520 16724 31564
rect 18691 31563 18749 31564
rect 20899 31520 20957 31521
rect 0 31480 364 31520
rect 404 31480 413 31520
rect 643 31480 652 31520
rect 692 31480 701 31520
rect 2467 31480 2476 31520
rect 2516 31480 3476 31520
rect 4675 31480 4684 31520
rect 4724 31480 5452 31520
rect 5492 31480 5501 31520
rect 6883 31480 6892 31520
rect 6932 31480 7372 31520
rect 7412 31480 7421 31520
rect 7555 31480 7564 31520
rect 7604 31480 7852 31520
rect 7892 31480 7901 31520
rect 8718 31480 8812 31520
rect 8852 31480 9100 31520
rect 9140 31480 9149 31520
rect 9667 31480 9676 31520
rect 9716 31480 10444 31520
rect 10484 31480 10493 31520
rect 10723 31480 10732 31520
rect 10772 31480 11692 31520
rect 11732 31480 11741 31520
rect 13027 31480 13036 31520
rect 13076 31480 13708 31520
rect 13748 31480 13757 31520
rect 15139 31480 15148 31520
rect 15188 31480 15532 31520
rect 15572 31480 15581 31520
rect 15630 31480 15724 31520
rect 15764 31480 15773 31520
rect 16291 31480 16300 31520
rect 16340 31480 16724 31520
rect 18691 31480 18700 31520
rect 18740 31480 20908 31520
rect 20948 31480 20957 31520
rect 0 31460 80 31480
rect 3436 31352 3476 31480
rect 5443 31479 5501 31480
rect 7555 31479 7613 31480
rect 8803 31479 8861 31480
rect 9091 31479 9149 31480
rect 10435 31479 10493 31480
rect 15715 31479 15773 31480
rect 20899 31479 20957 31480
rect 8419 31436 8477 31437
rect 11971 31436 12029 31437
rect 12835 31436 12893 31437
rect 6211 31396 6220 31436
rect 6260 31396 8428 31436
rect 8468 31396 10252 31436
rect 10292 31396 10301 31436
rect 11971 31396 11980 31436
rect 12020 31396 12172 31436
rect 12212 31396 12556 31436
rect 12596 31396 12844 31436
rect 12884 31396 12893 31436
rect 8419 31395 8477 31396
rect 11971 31395 12029 31396
rect 12835 31395 12893 31396
rect 17059 31436 17117 31437
rect 18499 31436 18557 31437
rect 21187 31436 21245 31437
rect 17059 31396 17068 31436
rect 17108 31396 18124 31436
rect 18164 31396 18173 31436
rect 18403 31396 18412 31436
rect 18452 31396 18508 31436
rect 18548 31396 18557 31436
rect 18883 31396 18892 31436
rect 18932 31396 19468 31436
rect 19508 31396 19517 31436
rect 19651 31396 19660 31436
rect 19700 31396 19709 31436
rect 19939 31396 19948 31436
rect 19988 31396 21196 31436
rect 21236 31396 21245 31436
rect 17059 31395 17117 31396
rect 18499 31395 18557 31396
rect 5635 31352 5693 31353
rect 10051 31352 10109 31353
rect 10339 31352 10397 31353
rect 355 31312 364 31352
rect 404 31312 1228 31352
rect 1268 31312 1277 31352
rect 1891 31312 1900 31352
rect 1940 31312 2668 31352
rect 2708 31312 2717 31352
rect 3427 31312 3436 31352
rect 3476 31312 4972 31352
rect 5012 31312 5644 31352
rect 5684 31312 5693 31352
rect 7651 31312 7660 31352
rect 7700 31312 8620 31352
rect 8660 31312 8669 31352
rect 9091 31312 9100 31352
rect 9140 31312 10060 31352
rect 10100 31312 10348 31352
rect 10388 31312 10397 31352
rect 1228 31268 1268 31312
rect 5635 31311 5693 31312
rect 10051 31311 10109 31312
rect 10339 31311 10397 31312
rect 10723 31352 10781 31353
rect 13795 31352 13853 31353
rect 10723 31312 10732 31352
rect 10772 31312 11308 31352
rect 11348 31312 12748 31352
rect 12788 31312 12797 31352
rect 13507 31312 13516 31352
rect 13556 31312 13804 31352
rect 13844 31312 13853 31352
rect 15235 31312 15244 31352
rect 15284 31312 15916 31352
rect 15956 31312 16492 31352
rect 16532 31312 16541 31352
rect 16771 31312 16780 31352
rect 16820 31312 16829 31352
rect 10723 31311 10781 31312
rect 13795 31311 13853 31312
rect 7651 31268 7709 31269
rect 10915 31268 10973 31269
rect 13699 31268 13757 31269
rect 16195 31268 16253 31269
rect 16780 31268 16820 31312
rect 19660 31268 19700 31396
rect 21187 31395 21245 31396
rect 20707 31352 20765 31353
rect 21424 31352 21504 31372
rect 19747 31312 19756 31352
rect 19796 31312 20044 31352
rect 20084 31312 20093 31352
rect 20707 31312 20716 31352
rect 20756 31312 21504 31352
rect 20707 31311 20765 31312
rect 21424 31292 21504 31312
rect 1228 31228 6508 31268
rect 6548 31228 6557 31268
rect 7651 31228 7660 31268
rect 7700 31228 7852 31268
rect 7892 31228 10156 31268
rect 10196 31228 10348 31268
rect 10388 31228 10397 31268
rect 10830 31228 10924 31268
rect 10964 31228 10973 31268
rect 11491 31228 11500 31268
rect 11540 31228 13228 31268
rect 13268 31228 13277 31268
rect 13614 31228 13708 31268
rect 13748 31228 13757 31268
rect 14851 31228 14860 31268
rect 14900 31228 15340 31268
rect 15380 31228 15389 31268
rect 15811 31228 15820 31268
rect 15860 31228 16108 31268
rect 16148 31228 16204 31268
rect 16244 31228 16272 31268
rect 16675 31228 16684 31268
rect 16724 31228 16820 31268
rect 18595 31228 18604 31268
rect 18644 31228 18653 31268
rect 19660 31228 20180 31268
rect 7651 31227 7709 31228
rect 10915 31227 10973 31228
rect 13699 31227 13757 31228
rect 12067 31184 12125 31185
rect 14275 31184 14333 31185
rect 14860 31184 14900 31228
rect 16195 31227 16253 31228
rect 17731 31184 17789 31185
rect 2947 31144 2956 31184
rect 2996 31144 4204 31184
rect 4244 31144 9388 31184
rect 9428 31144 9437 31184
rect 10435 31144 10444 31184
rect 10484 31144 11020 31184
rect 11060 31144 11069 31184
rect 12067 31144 12076 31184
rect 12116 31144 14284 31184
rect 14324 31144 14900 31184
rect 14956 31144 17740 31184
rect 17780 31144 18124 31184
rect 18164 31144 18173 31184
rect 12067 31143 12125 31144
rect 14275 31143 14333 31144
rect 3436 31060 6604 31100
rect 6644 31060 10924 31100
rect 10964 31060 10973 31100
rect 11875 31060 11884 31100
rect 11924 31060 12268 31100
rect 12308 31060 12317 31100
rect 0 31016 80 31036
rect 3436 31017 3476 31060
rect 3427 31016 3485 31017
rect 5923 31016 5981 31017
rect 11875 31016 11933 31017
rect 14956 31016 14996 31144
rect 17731 31143 17789 31144
rect 18604 31100 18644 31228
rect 19555 31184 19613 31185
rect 19555 31144 19564 31184
rect 19604 31144 19660 31184
rect 19700 31144 19709 31184
rect 19555 31143 19613 31144
rect 19651 31100 19709 31101
rect 17836 31060 18644 31100
rect 19555 31060 19564 31100
rect 19604 31060 19660 31100
rect 19700 31060 19709 31100
rect 20140 31100 20180 31228
rect 20140 31060 20564 31100
rect 16195 31016 16253 31017
rect 17836 31016 17876 31060
rect 19651 31059 19709 31060
rect 0 30976 3436 31016
rect 3476 30976 3485 31016
rect 4919 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 5305 31016
rect 5923 30976 5932 31016
rect 5972 30976 11884 31016
rect 11924 30976 11933 31016
rect 0 30956 80 30976
rect 3427 30975 3485 30976
rect 5923 30975 5981 30976
rect 11875 30975 11933 30976
rect 12268 30976 14996 31016
rect 15523 30976 15532 31016
rect 15572 30976 16204 31016
rect 16244 30976 17164 31016
rect 17204 30976 17876 31016
rect 17923 31016 17981 31017
rect 19843 31016 19901 31017
rect 20524 31016 20564 31060
rect 21424 31016 21504 31036
rect 17923 30976 17932 31016
rect 17972 30976 19852 31016
rect 19892 30976 19901 31016
rect 20039 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20425 31016
rect 20524 30976 21504 31016
rect 2563 30932 2621 30933
rect 11107 30932 11165 30933
rect 12163 30932 12221 30933
rect 2563 30892 2572 30932
rect 2612 30892 4396 30932
rect 4436 30892 4445 30932
rect 11107 30892 11116 30932
rect 11156 30892 12172 30932
rect 12212 30892 12221 30932
rect 2563 30891 2621 30892
rect 3427 30848 3485 30849
rect 2179 30808 2188 30848
rect 2228 30808 3436 30848
rect 3476 30808 3485 30848
rect 4396 30848 4436 30892
rect 11107 30891 11165 30892
rect 12163 30891 12221 30892
rect 12268 30848 12308 30976
rect 16195 30975 16253 30976
rect 17923 30975 17981 30976
rect 19843 30975 19901 30976
rect 21424 30956 21504 30976
rect 14083 30932 14141 30933
rect 13219 30892 13228 30932
rect 13268 30892 14092 30932
rect 14132 30892 14860 30932
rect 14900 30892 14909 30932
rect 14083 30891 14141 30892
rect 16867 30848 16925 30849
rect 4396 30808 5492 30848
rect 6499 30808 6508 30848
rect 6548 30808 12308 30848
rect 12355 30808 12364 30848
rect 12404 30808 16876 30848
rect 16916 30808 16925 30848
rect 19171 30808 19180 30848
rect 19220 30808 19660 30848
rect 19700 30808 19709 30848
rect 3427 30807 3485 30808
rect 5452 30680 5492 30808
rect 16867 30807 16925 30808
rect 5539 30764 5597 30765
rect 11875 30764 11933 30765
rect 12835 30764 12893 30765
rect 17731 30764 17789 30765
rect 5539 30724 5548 30764
rect 5588 30724 7372 30764
rect 7412 30724 7421 30764
rect 11107 30724 11116 30764
rect 11156 30724 11500 30764
rect 11540 30724 11549 30764
rect 11875 30724 11884 30764
rect 11924 30724 12556 30764
rect 12596 30724 12605 30764
rect 12835 30724 12844 30764
rect 12884 30724 13804 30764
rect 13844 30724 13853 30764
rect 15811 30724 15820 30764
rect 15860 30724 17548 30764
rect 17588 30724 17660 30764
rect 5539 30723 5597 30724
rect 11875 30723 11933 30724
rect 12835 30723 12893 30724
rect 7651 30680 7709 30681
rect 16003 30680 16061 30681
rect 1795 30640 1804 30680
rect 1844 30640 4684 30680
rect 4724 30640 4733 30680
rect 5452 30640 7660 30680
rect 7700 30640 7756 30680
rect 7796 30640 7805 30680
rect 8803 30640 8812 30680
rect 8852 30640 11404 30680
rect 11444 30640 11453 30680
rect 14179 30640 14188 30680
rect 14228 30640 14476 30680
rect 14516 30640 14525 30680
rect 15427 30640 15436 30680
rect 15476 30640 16012 30680
rect 16052 30640 16061 30680
rect 17620 30680 17660 30724
rect 17731 30724 17740 30764
rect 17780 30724 17932 30764
rect 17972 30724 17981 30764
rect 18211 30724 18220 30764
rect 18260 30724 18508 30764
rect 18548 30724 18557 30764
rect 19267 30724 19276 30764
rect 19316 30724 19852 30764
rect 19892 30724 19901 30764
rect 17731 30723 17789 30724
rect 21424 30680 21504 30700
rect 17620 30640 18700 30680
rect 18740 30640 18749 30680
rect 19747 30640 19756 30680
rect 19796 30640 21504 30680
rect 7651 30639 7709 30640
rect 16003 30639 16061 30640
rect 21424 30620 21504 30640
rect 6115 30596 6173 30597
rect 931 30556 940 30596
rect 980 30556 1228 30596
rect 1268 30556 1277 30596
rect 2467 30556 2476 30596
rect 2516 30556 2860 30596
rect 2900 30556 6124 30596
rect 6164 30556 6173 30596
rect 10339 30556 10348 30596
rect 10388 30556 11212 30596
rect 11252 30556 11261 30596
rect 11875 30556 11884 30596
rect 11924 30556 12940 30596
rect 12980 30556 12989 30596
rect 15139 30556 15148 30596
rect 15188 30556 17356 30596
rect 17396 30556 19468 30596
rect 19508 30556 19517 30596
rect 6115 30555 6173 30556
rect 0 30512 80 30532
rect 5923 30512 5981 30513
rect 11107 30512 11165 30513
rect 0 30472 5932 30512
rect 5972 30472 5981 30512
rect 0 30452 80 30472
rect 5923 30471 5981 30472
rect 6508 30472 9964 30512
rect 10004 30472 11116 30512
rect 11156 30472 11165 30512
rect 6508 30428 6548 30472
rect 11107 30471 11165 30472
rect 11212 30472 13420 30512
rect 13460 30472 13469 30512
rect 16108 30472 18220 30512
rect 18260 30472 18269 30512
rect 8995 30428 9053 30429
rect 11212 30428 11252 30472
rect 16108 30428 16148 30472
rect 547 30388 556 30428
rect 596 30388 940 30428
rect 980 30388 989 30428
rect 4099 30388 4108 30428
rect 4148 30388 6508 30428
rect 6548 30388 6557 30428
rect 8035 30388 8044 30428
rect 8084 30388 8620 30428
rect 8660 30388 8669 30428
rect 8910 30388 9004 30428
rect 9044 30388 9053 30428
rect 10531 30388 10540 30428
rect 10580 30388 11252 30428
rect 11395 30388 11404 30428
rect 11444 30388 11980 30428
rect 12020 30388 12460 30428
rect 12500 30388 12509 30428
rect 16099 30388 16108 30428
rect 16148 30388 16157 30428
rect 17347 30388 17356 30428
rect 17396 30388 17740 30428
rect 17780 30388 17789 30428
rect 18883 30388 18892 30428
rect 18932 30388 18941 30428
rect 8995 30387 9053 30388
rect 643 30344 701 30345
rect 5635 30344 5693 30345
rect 18892 30344 18932 30388
rect 21424 30344 21504 30364
rect 643 30304 652 30344
rect 692 30304 5068 30344
rect 5108 30304 5117 30344
rect 5635 30304 5644 30344
rect 5684 30304 8524 30344
rect 8564 30304 8573 30344
rect 9571 30304 9580 30344
rect 9620 30304 18932 30344
rect 20995 30304 21004 30344
rect 21044 30304 21504 30344
rect 643 30303 701 30304
rect 5635 30303 5693 30304
rect 21424 30284 21504 30304
rect 4771 30260 4829 30261
rect 3679 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 4065 30260
rect 4483 30220 4492 30260
rect 4532 30220 4780 30260
rect 4820 30220 4829 30260
rect 6307 30220 6316 30260
rect 6356 30220 8812 30260
rect 8852 30220 8861 30260
rect 11203 30220 11212 30260
rect 11252 30220 11404 30260
rect 11444 30220 11453 30260
rect 11779 30220 11788 30260
rect 11828 30220 12212 30260
rect 12547 30220 12556 30260
rect 12596 30220 14956 30260
rect 14996 30220 17644 30260
rect 17684 30220 17693 30260
rect 18799 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 19185 30260
rect 4771 30219 4829 30220
rect 12067 30176 12125 30177
rect 835 30136 844 30176
rect 884 30136 1132 30176
rect 1172 30136 1181 30176
rect 8236 30136 12076 30176
rect 12116 30136 12125 30176
rect 4771 30092 4829 30093
rect 8236 30092 8276 30136
rect 12067 30135 12125 30136
rect 12172 30092 12212 30220
rect 12835 30176 12893 30177
rect 12835 30136 12844 30176
rect 12884 30136 21388 30176
rect 21428 30136 21437 30176
rect 12835 30135 12893 30136
rect 16579 30092 16637 30093
rect 3139 30052 3148 30092
rect 3188 30052 3628 30092
rect 3668 30052 3677 30092
rect 4771 30052 4780 30092
rect 4820 30052 8276 30092
rect 8323 30052 8332 30092
rect 8372 30052 9580 30092
rect 9620 30052 9629 30092
rect 12172 30052 14764 30092
rect 14804 30052 14813 30092
rect 15619 30052 15628 30092
rect 15668 30052 15916 30092
rect 15956 30052 15965 30092
rect 16579 30052 16588 30092
rect 16628 30052 16684 30092
rect 16724 30052 17740 30092
rect 17780 30052 17789 30092
rect 19363 30052 19372 30092
rect 19412 30052 20180 30092
rect 4771 30051 4829 30052
rect 16579 30051 16637 30052
rect 0 30008 80 30028
rect 8131 30008 8189 30009
rect 15043 30008 15101 30009
rect 0 29968 1420 30008
rect 1460 29968 1469 30008
rect 1603 29968 1612 30008
rect 1652 29968 6700 30008
rect 6740 29968 6749 30008
rect 8131 29968 8140 30008
rect 8180 29968 8236 30008
rect 8276 29968 8285 30008
rect 8803 29968 8812 30008
rect 8852 29968 9388 30008
rect 9428 29968 9437 30008
rect 10051 29968 10060 30008
rect 10100 29968 15052 30008
rect 15092 29968 15101 30008
rect 20140 30008 20180 30052
rect 21424 30008 21504 30028
rect 20140 29968 21504 30008
rect 0 29948 80 29968
rect 8131 29967 8189 29968
rect 15043 29967 15101 29968
rect 21424 29948 21504 29968
rect 12355 29924 12413 29925
rect 12739 29924 12797 29925
rect 16675 29924 16733 29925
rect 7747 29884 7756 29924
rect 7796 29884 7948 29924
rect 7988 29884 7997 29924
rect 8899 29884 8908 29924
rect 8948 29884 9580 29924
rect 9620 29884 9629 29924
rect 12270 29884 12364 29924
rect 12404 29884 12413 29924
rect 12654 29884 12748 29924
rect 12788 29884 12797 29924
rect 13795 29884 13804 29924
rect 13844 29884 14956 29924
rect 14996 29884 15005 29924
rect 16675 29884 16684 29924
rect 16724 29884 16876 29924
rect 16916 29884 16925 29924
rect 17155 29884 17164 29924
rect 17204 29884 19372 29924
rect 19412 29884 19421 29924
rect 19747 29884 19756 29924
rect 19796 29884 19805 29924
rect 12355 29883 12413 29884
rect 12739 29883 12797 29884
rect 16675 29883 16733 29884
rect 2851 29840 2909 29841
rect 1315 29800 1324 29840
rect 1364 29800 2860 29840
rect 2900 29800 2909 29840
rect 3235 29800 3244 29840
rect 3284 29800 3916 29840
rect 3956 29800 3965 29840
rect 4579 29800 4588 29840
rect 4628 29800 13748 29840
rect 14563 29800 14572 29840
rect 14612 29800 15052 29840
rect 15092 29800 15628 29840
rect 15668 29800 16588 29840
rect 16628 29800 16637 29840
rect 2851 29799 2909 29800
rect 1987 29756 2045 29757
rect 2467 29756 2525 29757
rect 4588 29756 4628 29800
rect 8707 29756 8765 29757
rect 9187 29756 9245 29757
rect 13708 29756 13748 29800
rect 16483 29756 16541 29757
rect 1987 29716 1996 29756
rect 2036 29716 2476 29756
rect 2516 29716 4628 29756
rect 6307 29716 6316 29756
rect 6356 29716 7468 29756
rect 7508 29716 8716 29756
rect 8756 29716 8765 29756
rect 8899 29716 8908 29756
rect 8948 29716 9196 29756
rect 9236 29716 9245 29756
rect 9859 29716 9868 29756
rect 9908 29716 12076 29756
rect 12116 29716 12125 29756
rect 13708 29716 16492 29756
rect 16532 29716 16541 29756
rect 1987 29715 2045 29716
rect 2467 29715 2525 29716
rect 8707 29715 8765 29716
rect 9187 29715 9245 29716
rect 16483 29715 16541 29716
rect 3235 29672 3293 29673
rect 7171 29672 7229 29673
rect 11875 29672 11933 29673
rect 19756 29672 19796 29884
rect 19843 29840 19901 29841
rect 19843 29800 19852 29840
rect 19892 29800 19948 29840
rect 19988 29800 19997 29840
rect 19843 29799 19901 29800
rect 21424 29672 21504 29692
rect 1507 29632 1516 29672
rect 1556 29632 3244 29672
rect 3284 29632 4300 29672
rect 4340 29632 4349 29672
rect 4483 29632 4492 29672
rect 4532 29632 5068 29672
rect 5108 29632 5117 29672
rect 6691 29632 6700 29672
rect 6740 29632 6749 29672
rect 7171 29632 7180 29672
rect 7220 29632 8812 29672
rect 8852 29632 11116 29672
rect 11156 29632 11165 29672
rect 11587 29632 11596 29672
rect 11636 29632 11884 29672
rect 11924 29632 11933 29672
rect 13123 29632 13132 29672
rect 13172 29632 19796 29672
rect 20035 29632 20044 29672
rect 20084 29632 21504 29672
rect 3235 29631 3293 29632
rect 6700 29588 6740 29632
rect 7171 29631 7229 29632
rect 11875 29631 11933 29632
rect 21424 29612 21504 29632
rect 1699 29548 1708 29588
rect 1748 29548 5780 29588
rect 6700 29548 15916 29588
rect 15956 29548 15965 29588
rect 0 29504 80 29524
rect 1708 29504 1748 29548
rect 5740 29504 5780 29548
rect 9667 29504 9725 29505
rect 0 29464 1748 29504
rect 3331 29464 3340 29504
rect 3380 29464 4492 29504
rect 4532 29464 4541 29504
rect 4919 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 5305 29504
rect 5740 29464 9676 29504
rect 9716 29464 9725 29504
rect 12355 29464 12364 29504
rect 12404 29464 18028 29504
rect 18068 29464 18077 29504
rect 20039 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20425 29504
rect 0 29444 80 29464
rect 9667 29463 9725 29464
rect 6115 29420 6173 29421
rect 8995 29420 9053 29421
rect 13891 29420 13949 29421
rect 18211 29420 18269 29421
rect 3235 29380 3244 29420
rect 3284 29380 3532 29420
rect 3572 29380 3581 29420
rect 6030 29380 6124 29420
rect 6164 29380 6173 29420
rect 7843 29380 7852 29420
rect 7892 29380 8428 29420
rect 8468 29380 8477 29420
rect 8995 29380 9004 29420
rect 9044 29380 9196 29420
rect 9236 29380 9868 29420
rect 9908 29380 9917 29420
rect 13891 29380 13900 29420
rect 13940 29380 18220 29420
rect 18260 29380 18269 29420
rect 6115 29379 6173 29380
rect 8995 29379 9053 29380
rect 13891 29379 13949 29380
rect 18211 29379 18269 29380
rect 2947 29336 3005 29337
rect 8419 29336 8477 29337
rect 2947 29296 2956 29336
rect 2996 29296 6508 29336
rect 6548 29296 8428 29336
rect 8468 29296 8477 29336
rect 2947 29295 3005 29296
rect 8419 29295 8477 29296
rect 9187 29336 9245 29337
rect 21424 29336 21504 29356
rect 9187 29296 9196 29336
rect 9236 29296 15340 29336
rect 15380 29296 15389 29336
rect 15523 29296 15532 29336
rect 15572 29296 16396 29336
rect 16436 29296 16445 29336
rect 17452 29296 21504 29336
rect 9187 29295 9245 29296
rect 3235 29252 3293 29253
rect 1699 29212 1708 29252
rect 1748 29212 2668 29252
rect 2708 29212 2717 29252
rect 3150 29212 3244 29252
rect 3284 29212 3293 29252
rect 3235 29211 3293 29212
rect 7555 29252 7613 29253
rect 12259 29252 12317 29253
rect 13315 29252 13373 29253
rect 15427 29252 15485 29253
rect 17452 29252 17492 29296
rect 21424 29276 21504 29296
rect 7555 29212 7564 29252
rect 7604 29212 8140 29252
rect 8180 29212 8189 29252
rect 8419 29212 8428 29252
rect 8468 29212 9388 29252
rect 9428 29212 9437 29252
rect 11692 29212 12268 29252
rect 12308 29212 12460 29252
rect 12500 29212 12509 29252
rect 13315 29212 13324 29252
rect 13364 29212 14764 29252
rect 14804 29212 15436 29252
rect 15476 29212 15820 29252
rect 15860 29212 15869 29252
rect 17443 29212 17452 29252
rect 17492 29212 17501 29252
rect 19939 29212 19948 29252
rect 19988 29212 20180 29252
rect 7555 29211 7613 29212
rect 3331 29168 3389 29169
rect 2851 29128 2860 29168
rect 2900 29128 3340 29168
rect 3380 29128 3389 29168
rect 3331 29127 3389 29128
rect 4195 29168 4253 29169
rect 4771 29168 4829 29169
rect 8419 29168 8477 29169
rect 10723 29168 10781 29169
rect 4195 29128 4204 29168
rect 4244 29128 4492 29168
rect 4532 29128 4541 29168
rect 4771 29128 4780 29168
rect 4820 29128 4876 29168
rect 4916 29128 4925 29168
rect 5635 29128 5644 29168
rect 5684 29128 8180 29168
rect 4195 29127 4253 29128
rect 4771 29127 4829 29128
rect 5443 29084 5501 29085
rect 8140 29084 8180 29128
rect 8419 29128 8428 29168
rect 8468 29128 10732 29168
rect 10772 29128 10781 29168
rect 11395 29128 11404 29168
rect 11444 29128 11596 29168
rect 11636 29128 11645 29168
rect 8419 29127 8477 29128
rect 10723 29127 10781 29128
rect 11692 29084 11732 29212
rect 12259 29211 12317 29212
rect 12460 29084 12500 29212
rect 13315 29211 13373 29212
rect 15427 29211 15485 29212
rect 13411 29168 13469 29169
rect 17539 29168 17597 29169
rect 13411 29128 13420 29168
rect 13460 29128 13708 29168
rect 13748 29128 13757 29168
rect 14371 29128 14380 29168
rect 14420 29128 14860 29168
rect 14900 29128 16012 29168
rect 16052 29128 16061 29168
rect 16579 29128 16588 29168
rect 16628 29128 17068 29168
rect 17108 29128 17117 29168
rect 17454 29128 17548 29168
rect 17588 29128 17597 29168
rect 20140 29168 20180 29212
rect 20140 29128 21292 29168
rect 21332 29128 21341 29168
rect 13411 29127 13469 29128
rect 17539 29127 17597 29128
rect 13891 29084 13949 29085
rect 15811 29084 15869 29085
rect 19363 29084 19421 29085
rect 1123 29044 1132 29084
rect 1172 29044 3284 29084
rect 0 29000 80 29020
rect 3244 29000 3284 29044
rect 3340 29044 5452 29084
rect 5492 29044 5501 29084
rect 7555 29044 7564 29084
rect 7604 29044 7852 29084
rect 7892 29044 7901 29084
rect 8140 29044 11732 29084
rect 11788 29044 12268 29084
rect 12308 29044 12317 29084
rect 12460 29044 13900 29084
rect 13940 29044 13949 29084
rect 15523 29044 15532 29084
rect 15572 29044 15820 29084
rect 15860 29044 15869 29084
rect 19278 29044 19372 29084
rect 19412 29044 19421 29084
rect 0 28960 1516 29000
rect 1556 28960 1565 29000
rect 3043 28960 3052 29000
rect 3092 28960 3101 29000
rect 3204 28960 3244 29000
rect 3284 28960 3293 29000
rect 0 28940 80 28960
rect 3052 28916 3092 28960
rect 3340 28916 3380 29044
rect 5443 29043 5501 29044
rect 11788 29000 11828 29044
rect 13891 29043 13949 29044
rect 15811 29043 15869 29044
rect 19363 29043 19421 29044
rect 21424 29000 21504 29020
rect 11748 28960 11788 29000
rect 11828 28960 11837 29000
rect 15331 28960 15340 29000
rect 15380 28960 15389 29000
rect 19939 28960 19948 29000
rect 19988 28960 20180 29000
rect 21379 28960 21388 29000
rect 21428 28960 21504 29000
rect 6691 28916 6749 28917
rect 9955 28916 10013 28917
rect 13699 28916 13757 28917
rect 1315 28876 1324 28916
rect 1364 28876 2284 28916
rect 2324 28876 2333 28916
rect 3052 28876 3380 28916
rect 3619 28876 3628 28916
rect 3668 28876 3677 28916
rect 4675 28876 4684 28916
rect 4724 28876 5356 28916
rect 5396 28876 5405 28916
rect 6307 28876 6316 28916
rect 6356 28876 6700 28916
rect 6740 28876 6749 28916
rect 7939 28876 7948 28916
rect 7988 28876 8236 28916
rect 8276 28876 8285 28916
rect 9955 28876 9964 28916
rect 10004 28876 13708 28916
rect 13748 28876 13757 28916
rect 15340 28916 15380 28960
rect 17731 28916 17789 28917
rect 15340 28876 15628 28916
rect 15668 28876 15677 28916
rect 17539 28876 17548 28916
rect 17588 28876 17740 28916
rect 17780 28876 17789 28916
rect 20140 28916 20180 28960
rect 21424 28940 21504 28960
rect 20515 28916 20573 28917
rect 20140 28876 20524 28916
rect 20564 28876 20573 28916
rect 3235 28832 3293 28833
rect 2755 28792 2764 28832
rect 2804 28792 3244 28832
rect 3284 28792 3293 28832
rect 3628 28832 3668 28876
rect 6691 28875 6749 28876
rect 9955 28875 10013 28876
rect 13699 28875 13757 28876
rect 17731 28875 17789 28876
rect 20515 28875 20573 28876
rect 12067 28832 12125 28833
rect 3628 28792 4532 28832
rect 5539 28792 5548 28832
rect 5588 28792 5740 28832
rect 5780 28792 5789 28832
rect 6508 28792 7756 28832
rect 7796 28792 7805 28832
rect 12067 28792 12076 28832
rect 12116 28792 12172 28832
rect 12212 28792 12221 28832
rect 13411 28792 13420 28832
rect 13460 28792 13469 28832
rect 3235 28791 3293 28792
rect 4492 28748 4532 28792
rect 6508 28748 6548 28792
rect 12067 28791 12125 28792
rect 6979 28748 7037 28749
rect 9955 28748 10013 28749
rect 13420 28748 13460 28792
rect 18211 28748 18269 28749
rect 3679 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 4065 28748
rect 4483 28708 4492 28748
rect 4532 28708 4541 28748
rect 5923 28708 5932 28748
rect 5972 28708 6124 28748
rect 6164 28708 6508 28748
rect 6548 28708 6557 28748
rect 6883 28708 6892 28748
rect 6932 28708 6988 28748
rect 7028 28708 7276 28748
rect 7316 28708 7325 28748
rect 8611 28708 8620 28748
rect 8660 28708 9964 28748
rect 10004 28708 10013 28748
rect 11299 28708 11308 28748
rect 11348 28708 12940 28748
rect 12980 28708 12989 28748
rect 13420 28708 14284 28748
rect 14324 28708 14333 28748
rect 18126 28708 18220 28748
rect 18260 28708 18269 28748
rect 18799 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 19185 28748
rect 6979 28707 7037 28708
rect 9955 28707 10013 28708
rect 18211 28707 18269 28708
rect 5539 28664 5597 28665
rect 10051 28664 10109 28665
rect 10339 28664 10397 28665
rect 11875 28664 11933 28665
rect 18595 28664 18653 28665
rect 5539 28624 5548 28664
rect 5588 28624 10060 28664
rect 10100 28624 10348 28664
rect 10388 28624 10397 28664
rect 11203 28624 11212 28664
rect 11252 28624 11884 28664
rect 11924 28624 13132 28664
rect 13172 28624 13181 28664
rect 13411 28624 13420 28664
rect 13460 28624 18604 28664
rect 18644 28624 18653 28664
rect 5539 28623 5597 28624
rect 10051 28623 10109 28624
rect 10339 28623 10397 28624
rect 11875 28623 11933 28624
rect 18595 28623 18653 28624
rect 19267 28664 19325 28665
rect 21424 28664 21504 28684
rect 19267 28624 19276 28664
rect 19316 28624 21504 28664
rect 19267 28623 19325 28624
rect 21424 28604 21504 28624
rect 5731 28580 5789 28581
rect 16003 28580 16061 28581
rect 16867 28580 16925 28581
rect 20803 28580 20861 28581
rect 2371 28540 2380 28580
rect 2420 28540 3724 28580
rect 3764 28540 3773 28580
rect 4195 28540 4204 28580
rect 4244 28540 5740 28580
rect 5780 28540 5789 28580
rect 6211 28540 6220 28580
rect 6260 28540 9196 28580
rect 9236 28540 9245 28580
rect 16003 28540 16012 28580
rect 16052 28540 16108 28580
rect 16148 28540 16157 28580
rect 16867 28540 16876 28580
rect 16916 28540 20812 28580
rect 20852 28540 20861 28580
rect 5731 28539 5789 28540
rect 16003 28539 16061 28540
rect 16867 28539 16925 28540
rect 20803 28539 20861 28540
rect 0 28496 80 28516
rect 7939 28496 7997 28497
rect 17251 28496 17309 28497
rect 0 28456 1804 28496
rect 1844 28456 1853 28496
rect 2755 28456 2764 28496
rect 2804 28456 3148 28496
rect 3188 28456 3197 28496
rect 3811 28456 3820 28496
rect 3860 28456 7948 28496
rect 7988 28456 7997 28496
rect 11011 28456 11020 28496
rect 11060 28456 11692 28496
rect 11732 28456 11741 28496
rect 11971 28456 11980 28496
rect 12020 28456 13228 28496
rect 13268 28456 13277 28496
rect 14284 28456 17260 28496
rect 17300 28456 17309 28496
rect 18979 28456 18988 28496
rect 19028 28456 19468 28496
rect 19508 28456 19517 28496
rect 0 28436 80 28456
rect 7939 28455 7997 28456
rect 3619 28412 3677 28413
rect 4099 28412 4157 28413
rect 7459 28412 7517 28413
rect 1411 28372 1420 28412
rect 1460 28372 3476 28412
rect 3534 28372 3628 28412
rect 3668 28372 3677 28412
rect 4003 28372 4012 28412
rect 4052 28372 4108 28412
rect 4148 28372 4157 28412
rect 3436 28328 3476 28372
rect 3619 28371 3677 28372
rect 4099 28371 4157 28372
rect 4492 28372 6124 28412
rect 6164 28372 6173 28412
rect 6307 28372 6316 28412
rect 6356 28372 6700 28412
rect 6740 28372 6749 28412
rect 6883 28372 6892 28412
rect 6932 28372 7468 28412
rect 7508 28372 7517 28412
rect 4492 28328 4532 28372
rect 7459 28371 7517 28372
rect 8131 28412 8189 28413
rect 14284 28412 14324 28456
rect 17251 28455 17309 28456
rect 8131 28372 8140 28412
rect 8180 28372 9196 28412
rect 9236 28372 14324 28412
rect 15244 28372 19276 28412
rect 19316 28372 19325 28412
rect 8131 28371 8189 28372
rect 2500 28288 3148 28328
rect 3188 28288 3197 28328
rect 3436 28288 4532 28328
rect 4579 28288 4588 28328
rect 4628 28288 5876 28328
rect 7747 28288 7756 28328
rect 7796 28288 7948 28328
rect 7988 28288 8524 28328
rect 8564 28288 8573 28328
rect 8908 28288 9004 28328
rect 9044 28288 9053 28328
rect 10915 28288 10924 28328
rect 10964 28288 11308 28328
rect 11348 28288 11357 28328
rect 11587 28288 11596 28328
rect 11636 28288 12076 28328
rect 12116 28288 12125 28328
rect 12259 28288 12268 28328
rect 12308 28288 12556 28328
rect 12596 28288 12940 28328
rect 12980 28288 12989 28328
rect 14371 28288 14380 28328
rect 14420 28288 14764 28328
rect 14804 28288 15052 28328
rect 15092 28288 15101 28328
rect 2500 28244 2540 28288
rect 5539 28244 5597 28245
rect 1507 28204 1516 28244
rect 1556 28204 2540 28244
rect 2947 28204 2956 28244
rect 2996 28204 4780 28244
rect 4820 28204 4829 28244
rect 5251 28204 5260 28244
rect 5300 28204 5548 28244
rect 5588 28204 5597 28244
rect 5836 28244 5876 28288
rect 8419 28244 8477 28245
rect 5836 28204 8428 28244
rect 8468 28204 8477 28244
rect 2956 28160 2996 28204
rect 5539 28203 5597 28204
rect 8419 28203 8477 28204
rect 1987 28120 1996 28160
rect 2036 28120 2996 28160
rect 3427 28160 3485 28161
rect 8908 28160 8948 28288
rect 15244 28160 15284 28372
rect 16003 28328 16061 28329
rect 16195 28328 16253 28329
rect 21424 28328 21504 28348
rect 16003 28288 16012 28328
rect 16052 28288 16204 28328
rect 16244 28288 16300 28328
rect 16340 28288 16349 28328
rect 17635 28288 17644 28328
rect 17684 28288 21504 28328
rect 16003 28287 16061 28288
rect 16195 28287 16253 28288
rect 21424 28268 21504 28288
rect 21091 28244 21149 28245
rect 15811 28204 15820 28244
rect 15860 28204 16108 28244
rect 16148 28204 16157 28244
rect 17827 28204 17836 28244
rect 17876 28204 18220 28244
rect 18260 28204 18269 28244
rect 18883 28204 18892 28244
rect 18932 28204 21100 28244
rect 21140 28204 21149 28244
rect 21091 28203 21149 28204
rect 3427 28120 3436 28160
rect 3476 28120 4876 28160
rect 4916 28120 4925 28160
rect 6691 28120 6700 28160
rect 6740 28120 7084 28160
rect 7124 28120 7133 28160
rect 8908 28120 11540 28160
rect 11779 28120 11788 28160
rect 11828 28120 11980 28160
rect 12020 28120 12029 28160
rect 12355 28120 12364 28160
rect 12404 28120 12556 28160
rect 12596 28120 12605 28160
rect 15139 28120 15148 28160
rect 15188 28120 15284 28160
rect 16675 28120 16684 28160
rect 16724 28120 17740 28160
rect 17780 28120 17789 28160
rect 19939 28120 19948 28160
rect 19988 28120 20908 28160
rect 20948 28120 20957 28160
rect 3427 28119 3485 28120
rect 3235 28036 3244 28076
rect 3284 28036 3724 28076
rect 3764 28036 6220 28076
rect 6260 28036 6269 28076
rect 0 27992 80 28012
rect 1987 27992 2045 27993
rect 0 27952 1996 27992
rect 2036 27952 2045 27992
rect 0 27932 80 27952
rect 1987 27951 2045 27952
rect 4579 27992 4637 27993
rect 8908 27992 8948 28120
rect 11500 27992 11540 28120
rect 11587 28076 11645 28077
rect 12739 28076 12797 28077
rect 18211 28076 18269 28077
rect 11587 28036 11596 28076
rect 11636 28036 12268 28076
rect 12308 28036 12317 28076
rect 12739 28036 12748 28076
rect 12788 28036 18220 28076
rect 18260 28036 18269 28076
rect 19651 28036 19660 28076
rect 19700 28036 20852 28076
rect 11587 28035 11645 28036
rect 12739 28035 12797 28036
rect 18211 28035 18269 28036
rect 20812 27992 20852 28036
rect 21424 27992 21504 28012
rect 4579 27952 4588 27992
rect 4628 27952 4780 27992
rect 4820 27952 4829 27992
rect 4919 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 5305 27992
rect 6115 27952 6124 27992
rect 6164 27952 6892 27992
rect 6932 27952 6941 27992
rect 7459 27952 7468 27992
rect 7508 27952 8948 27992
rect 10339 27952 10348 27992
rect 10388 27952 10636 27992
rect 10676 27952 10685 27992
rect 11500 27952 14764 27992
rect 14804 27952 15340 27992
rect 15380 27952 15389 27992
rect 20039 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20425 27992
rect 20812 27952 21504 27992
rect 4579 27951 4637 27952
rect 21424 27932 21504 27952
rect 3235 27908 3293 27909
rect 3043 27868 3052 27908
rect 3092 27868 3244 27908
rect 3284 27868 3293 27908
rect 3235 27867 3293 27868
rect 4099 27908 4157 27909
rect 5443 27908 5501 27909
rect 11011 27908 11069 27909
rect 4099 27868 4108 27908
rect 4148 27868 5452 27908
rect 5492 27868 5501 27908
rect 4099 27867 4157 27868
rect 5443 27867 5501 27868
rect 8908 27868 11020 27908
rect 11060 27868 11069 27908
rect 11683 27868 11692 27908
rect 11732 27868 12460 27908
rect 12500 27868 12509 27908
rect 4483 27740 4541 27741
rect 8908 27740 8948 27868
rect 11011 27867 11069 27868
rect 12355 27824 12413 27825
rect 8995 27784 9004 27824
rect 9044 27784 9053 27824
rect 11971 27784 11980 27824
rect 12020 27784 12364 27824
rect 12404 27784 12413 27824
rect 13027 27784 13036 27824
rect 13076 27784 17356 27824
rect 17396 27784 17548 27824
rect 17588 27784 17597 27824
rect 1795 27700 1804 27740
rect 1844 27700 2092 27740
rect 2132 27700 2141 27740
rect 4398 27700 4492 27740
rect 4532 27700 4541 27740
rect 4483 27699 4541 27700
rect 4876 27700 8948 27740
rect 9004 27740 9044 27784
rect 12355 27783 12413 27784
rect 11875 27740 11933 27741
rect 9004 27700 9140 27740
rect 11779 27700 11788 27740
rect 11828 27700 11884 27740
rect 11924 27700 12460 27740
rect 12500 27700 12509 27740
rect 13036 27700 17164 27740
rect 17204 27700 17213 27740
rect 18787 27700 18796 27740
rect 18836 27700 19276 27740
rect 19316 27700 19325 27740
rect 19843 27700 19852 27740
rect 19892 27700 19901 27740
rect 4876 27656 4916 27700
rect 6211 27656 6269 27657
rect 8515 27656 8573 27657
rect 1603 27616 1612 27656
rect 1652 27616 4684 27656
rect 4724 27616 4733 27656
rect 4867 27616 4876 27656
rect 4916 27616 4925 27656
rect 6211 27616 6220 27656
rect 6260 27616 6700 27656
rect 6740 27616 6749 27656
rect 8515 27616 8524 27656
rect 8564 27616 9004 27656
rect 9044 27616 9053 27656
rect 6211 27615 6269 27616
rect 8515 27615 8573 27616
rect 4291 27572 4349 27573
rect 9100 27572 9140 27700
rect 11875 27699 11933 27700
rect 9379 27656 9437 27657
rect 11971 27656 12029 27657
rect 9379 27616 9388 27656
rect 9428 27616 9484 27656
rect 9524 27616 9533 27656
rect 11395 27616 11404 27656
rect 11444 27616 11980 27656
rect 12020 27616 12029 27656
rect 9379 27615 9437 27616
rect 9484 27572 9524 27616
rect 11971 27615 12029 27616
rect 13036 27572 13076 27700
rect 19852 27656 19892 27700
rect 21424 27656 21504 27676
rect 13123 27616 13132 27656
rect 13172 27616 18892 27656
rect 18932 27616 18941 27656
rect 19852 27616 21504 27656
rect 21424 27596 21504 27616
rect 4206 27532 4300 27572
rect 4340 27532 4349 27572
rect 7267 27532 7276 27572
rect 7316 27532 7660 27572
rect 7700 27532 7709 27572
rect 9091 27532 9100 27572
rect 9140 27532 9149 27572
rect 9484 27532 13076 27572
rect 14563 27532 14572 27572
rect 14612 27532 19468 27572
rect 19508 27532 19517 27572
rect 4291 27531 4349 27532
rect 0 27488 80 27508
rect 3427 27488 3485 27489
rect 7363 27488 7421 27489
rect 0 27448 1268 27488
rect 1315 27448 1324 27488
rect 1364 27448 1460 27488
rect 3342 27448 3436 27488
rect 3476 27448 3916 27488
rect 3956 27448 3965 27488
rect 6595 27448 6604 27488
rect 6644 27448 7372 27488
rect 7412 27448 7421 27488
rect 7660 27488 7700 27532
rect 9283 27488 9341 27489
rect 7660 27448 9292 27488
rect 9332 27448 9341 27488
rect 0 27428 80 27448
rect 1228 27404 1268 27448
rect 1315 27404 1373 27405
rect 1228 27364 1324 27404
rect 1364 27364 1373 27404
rect 1420 27404 1460 27448
rect 3427 27447 3485 27448
rect 7363 27447 7421 27448
rect 9283 27447 9341 27448
rect 11320 27448 12940 27488
rect 12980 27448 13612 27488
rect 13652 27448 13661 27488
rect 14275 27448 14284 27488
rect 14324 27448 17836 27488
rect 17876 27448 17885 27488
rect 3523 27404 3581 27405
rect 6691 27404 6749 27405
rect 1420 27364 3532 27404
rect 3572 27364 4108 27404
rect 4148 27364 6412 27404
rect 6452 27364 6461 27404
rect 6606 27364 6700 27404
rect 6740 27364 6749 27404
rect 1315 27363 1373 27364
rect 3523 27363 3581 27364
rect 6691 27363 6749 27364
rect 6979 27404 7037 27405
rect 11320 27404 11360 27448
rect 20515 27404 20573 27405
rect 6979 27364 6988 27404
rect 7028 27364 11360 27404
rect 11779 27364 11788 27404
rect 11828 27364 17452 27404
rect 17492 27364 17501 27404
rect 19651 27364 19660 27404
rect 19700 27364 19852 27404
rect 19892 27364 19901 27404
rect 20515 27364 20524 27404
rect 20564 27364 21428 27404
rect 6979 27363 7037 27364
rect 20515 27363 20573 27364
rect 21388 27340 21428 27364
rect 5635 27320 5693 27321
rect 12067 27320 12125 27321
rect 4291 27280 4300 27320
rect 4340 27280 5644 27320
rect 5684 27280 5693 27320
rect 8803 27280 8812 27320
rect 8852 27280 9964 27320
rect 10004 27280 10636 27320
rect 10676 27280 10685 27320
rect 11982 27280 12076 27320
rect 12116 27280 12125 27320
rect 5635 27279 5693 27280
rect 12067 27279 12125 27280
rect 17251 27320 17309 27321
rect 21283 27320 21341 27321
rect 17251 27280 17260 27320
rect 17300 27280 21292 27320
rect 21332 27280 21341 27320
rect 21388 27280 21504 27340
rect 17251 27279 17309 27280
rect 21283 27279 21341 27280
rect 21424 27260 21504 27280
rect 19363 27236 19421 27237
rect 3679 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 4065 27236
rect 5539 27196 5548 27236
rect 5588 27196 11884 27236
rect 11924 27196 14476 27236
rect 14516 27196 14525 27236
rect 17923 27196 17932 27236
rect 17972 27196 18412 27236
rect 18452 27196 18461 27236
rect 18799 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 19185 27236
rect 19363 27196 19372 27236
rect 19412 27196 19421 27236
rect 19363 27195 19421 27196
rect 11299 27152 11357 27153
rect 19372 27152 19412 27195
rect 3532 27112 6796 27152
rect 6836 27112 7180 27152
rect 7220 27112 7229 27152
rect 10339 27112 10348 27152
rect 10388 27112 11308 27152
rect 11348 27112 11357 27152
rect 11491 27112 11500 27152
rect 11540 27112 12596 27152
rect 12643 27112 12652 27152
rect 12692 27112 19412 27152
rect 1219 27028 1228 27068
rect 1268 27028 3340 27068
rect 3380 27028 3389 27068
rect 0 26984 80 27004
rect 1411 26984 1469 26985
rect 1795 26984 1853 26985
rect 3532 26984 3572 27112
rect 11299 27111 11357 27112
rect 4099 27068 4157 27069
rect 12556 27068 12596 27112
rect 15523 27068 15581 27069
rect 19363 27068 19421 27069
rect 4003 27028 4012 27068
rect 4052 27028 4108 27068
rect 4148 27028 4157 27068
rect 4675 27028 4684 27068
rect 4724 27028 5548 27068
rect 5588 27028 5597 27068
rect 6115 27028 6124 27068
rect 6164 27028 8332 27068
rect 8372 27028 8381 27068
rect 9187 27028 9196 27068
rect 9236 27028 9676 27068
rect 9716 27028 9725 27068
rect 9772 27028 11980 27068
rect 12020 27028 12029 27068
rect 12556 27028 12940 27068
rect 12980 27028 12989 27068
rect 15438 27028 15532 27068
rect 15572 27028 15581 27068
rect 15715 27028 15724 27068
rect 15764 27028 16300 27068
rect 16340 27028 16349 27068
rect 19278 27028 19372 27068
rect 19412 27028 19421 27068
rect 4099 27027 4157 27028
rect 9772 26984 9812 27028
rect 15523 27027 15581 27028
rect 19363 27027 19421 27028
rect 19468 27028 19948 27068
rect 19988 27028 19997 27068
rect 0 26944 1420 26984
rect 1460 26944 1804 26984
rect 1844 26944 1853 26984
rect 1896 26944 1905 26984
rect 1945 26944 3572 26984
rect 3619 26944 3628 26984
rect 3668 26944 7756 26984
rect 7796 26944 7805 26984
rect 9763 26944 9772 26984
rect 9812 26944 9821 26984
rect 10147 26944 10156 26984
rect 10196 26944 11500 26984
rect 11540 26944 11549 26984
rect 17155 26944 17164 26984
rect 17204 26944 17452 26984
rect 17492 26944 17501 26984
rect 0 26924 80 26944
rect 1411 26943 1469 26944
rect 1795 26943 1853 26944
rect 15523 26900 15581 26901
rect 19468 26900 19508 27028
rect 21424 26984 21504 27004
rect 19555 26944 19564 26984
rect 19604 26944 21504 26984
rect 21424 26924 21504 26944
rect 1411 26860 1420 26900
rect 1460 26860 9100 26900
rect 9140 26860 9388 26900
rect 9428 26860 9437 26900
rect 9667 26860 9676 26900
rect 9716 26860 10580 26900
rect 10627 26860 10636 26900
rect 10676 26860 13900 26900
rect 13940 26860 13949 26900
rect 15331 26860 15340 26900
rect 15380 26860 15532 26900
rect 15572 26860 15581 26900
rect 15907 26860 15916 26900
rect 15956 26860 19508 26900
rect 10540 26816 10580 26860
rect 15523 26859 15581 26860
rect 11971 26816 12029 26817
rect 17443 26816 17501 26817
rect 20803 26816 20861 26817
rect 1603 26776 1612 26816
rect 1652 26776 4204 26816
rect 4244 26776 4253 26816
rect 5347 26776 5356 26816
rect 5396 26776 6220 26816
rect 6260 26776 6269 26816
rect 6499 26776 6508 26816
rect 6548 26776 7276 26816
rect 7316 26776 7325 26816
rect 7747 26776 7756 26816
rect 7796 26776 8140 26816
rect 8180 26776 9772 26816
rect 9812 26776 10444 26816
rect 10484 26776 10493 26816
rect 10540 26776 11828 26816
rect 11886 26776 11980 26816
rect 12020 26776 12029 26816
rect 12739 26776 12748 26816
rect 12788 26776 13324 26816
rect 13364 26776 13373 26816
rect 16579 26776 16588 26816
rect 16628 26776 16972 26816
rect 17012 26776 17021 26816
rect 17443 26776 17452 26816
rect 17492 26776 18028 26816
rect 18068 26776 18077 26816
rect 19939 26776 19948 26816
rect 19988 26776 20812 26816
rect 20852 26776 20861 26816
rect 2275 26732 2333 26733
rect 11788 26732 11828 26776
rect 11971 26775 12029 26776
rect 17443 26775 17501 26776
rect 20803 26775 20861 26776
rect 2190 26692 2284 26732
rect 2324 26692 2333 26732
rect 2851 26692 2860 26732
rect 2900 26692 3476 26732
rect 3523 26692 3532 26732
rect 3572 26692 11116 26732
rect 11156 26692 11165 26732
rect 11788 26692 17548 26732
rect 17588 26692 17597 26732
rect 19180 26692 19660 26732
rect 19700 26692 19709 26732
rect 2275 26691 2333 26692
rect 3436 26648 3476 26692
rect 6691 26648 6749 26649
rect 10915 26648 10973 26649
rect 19180 26648 19220 26692
rect 21424 26648 21504 26668
rect 2371 26608 2380 26648
rect 2420 26608 2540 26648
rect 2755 26608 2764 26648
rect 2804 26608 3340 26648
rect 3380 26608 3389 26648
rect 3436 26608 3628 26648
rect 3668 26608 3677 26648
rect 4012 26608 6356 26648
rect 1315 26564 1373 26565
rect 2275 26564 2333 26565
rect 1315 26524 1324 26564
rect 1364 26524 2284 26564
rect 2324 26524 2333 26564
rect 2500 26564 2540 26608
rect 4012 26564 4052 26608
rect 6316 26564 6356 26608
rect 6691 26608 6700 26648
rect 6740 26608 7180 26648
rect 7220 26608 7564 26648
rect 7604 26608 7988 26648
rect 8419 26608 8428 26648
rect 8468 26608 10924 26648
rect 10964 26608 13996 26648
rect 14036 26608 15724 26648
rect 15764 26608 15773 26648
rect 19171 26608 19180 26648
rect 19220 26608 19229 26648
rect 19555 26608 19564 26648
rect 19604 26608 19613 26648
rect 20035 26608 20044 26648
rect 20084 26608 21504 26648
rect 6691 26607 6749 26608
rect 7948 26564 7988 26608
rect 10915 26607 10973 26608
rect 11299 26564 11357 26565
rect 12835 26564 12893 26565
rect 17731 26564 17789 26565
rect 19459 26564 19517 26565
rect 2500 26524 4052 26564
rect 4099 26524 4108 26564
rect 4148 26524 4780 26564
rect 4820 26524 4829 26564
rect 6316 26524 6508 26564
rect 6548 26524 6557 26564
rect 6691 26524 6700 26564
rect 6740 26524 7852 26564
rect 7892 26524 7901 26564
rect 7948 26524 9292 26564
rect 9332 26524 9341 26564
rect 10243 26524 10252 26564
rect 10292 26524 11308 26564
rect 11348 26524 11357 26564
rect 11491 26524 11500 26564
rect 11540 26524 11788 26564
rect 11828 26524 11837 26564
rect 12835 26524 12844 26564
rect 12884 26524 13228 26564
rect 13268 26524 13612 26564
rect 13652 26524 14380 26564
rect 14420 26524 14429 26564
rect 17731 26524 17740 26564
rect 17780 26524 19468 26564
rect 19508 26524 19517 26564
rect 19564 26564 19604 26608
rect 21424 26588 21504 26608
rect 20899 26564 20957 26565
rect 19564 26524 20908 26564
rect 20948 26524 20957 26564
rect 1315 26523 1373 26524
rect 2275 26523 2333 26524
rect 11299 26523 11357 26524
rect 12835 26523 12893 26524
rect 17731 26523 17789 26524
rect 19459 26523 19517 26524
rect 20899 26523 20957 26524
rect 0 26480 80 26500
rect 3523 26480 3581 26481
rect 6499 26480 6557 26481
rect 8611 26480 8669 26481
rect 8803 26480 8861 26481
rect 0 26440 1268 26480
rect 1315 26440 1324 26480
rect 1364 26440 3532 26480
rect 3572 26440 3581 26480
rect 3811 26440 3820 26480
rect 3860 26440 4396 26480
rect 4436 26440 4445 26480
rect 4919 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 5305 26480
rect 6499 26440 6508 26480
rect 6548 26440 6604 26480
rect 6644 26440 6653 26480
rect 7171 26440 7180 26480
rect 7220 26440 7468 26480
rect 7508 26440 7517 26480
rect 8526 26440 8620 26480
rect 8660 26440 8669 26480
rect 8718 26440 8812 26480
rect 8852 26440 8861 26480
rect 0 26420 80 26440
rect 1228 26396 1268 26440
rect 3523 26439 3581 26440
rect 6499 26439 6557 26440
rect 8611 26439 8669 26440
rect 8803 26439 8861 26440
rect 8995 26480 9053 26481
rect 9571 26480 9629 26481
rect 13891 26480 13949 26481
rect 15235 26480 15293 26481
rect 16483 26480 16541 26481
rect 8995 26440 9004 26480
rect 9044 26440 9100 26480
rect 9140 26440 9149 26480
rect 9486 26440 9580 26480
rect 9620 26440 9629 26480
rect 13806 26440 13900 26480
rect 13940 26440 13949 26480
rect 15150 26440 15244 26480
rect 15284 26440 15293 26480
rect 16398 26440 16492 26480
rect 16532 26440 16541 26480
rect 8995 26439 9053 26440
rect 9571 26439 9629 26440
rect 13891 26439 13949 26440
rect 15235 26439 15293 26440
rect 16483 26439 16541 26440
rect 17620 26440 19372 26480
rect 19412 26440 19421 26480
rect 20039 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20425 26480
rect 1891 26396 1949 26397
rect 17620 26396 17660 26440
rect 1228 26356 1900 26396
rect 1940 26356 16204 26396
rect 16244 26356 16253 26396
rect 16387 26356 16396 26396
rect 16436 26356 16972 26396
rect 17012 26356 17021 26396
rect 17155 26356 17164 26396
rect 17204 26356 17660 26396
rect 17731 26356 17740 26396
rect 17780 26356 18508 26396
rect 18548 26356 18557 26396
rect 1891 26355 1949 26356
rect 21424 26312 21504 26332
rect 1411 26272 1420 26312
rect 1460 26272 2956 26312
rect 2996 26272 3005 26312
rect 3139 26272 3148 26312
rect 3188 26272 5164 26312
rect 5204 26272 5213 26312
rect 7075 26272 7084 26312
rect 7124 26272 10252 26312
rect 10292 26272 10301 26312
rect 10915 26272 10924 26312
rect 10964 26272 17068 26312
rect 17108 26272 17117 26312
rect 20899 26272 20908 26312
rect 20948 26272 21504 26312
rect 21424 26252 21504 26272
rect 1219 26228 1277 26229
rect 4291 26228 4349 26229
rect 1123 26188 1132 26228
rect 1172 26188 1228 26228
rect 1268 26188 1277 26228
rect 1219 26187 1277 26188
rect 1324 26188 1996 26228
rect 2036 26188 2045 26228
rect 4291 26188 4300 26228
rect 4340 26188 4684 26228
rect 4724 26188 4733 26228
rect 7267 26188 7276 26228
rect 7316 26188 9196 26228
rect 9236 26188 9245 26228
rect 12547 26188 12556 26228
rect 12596 26188 12844 26228
rect 12884 26188 12893 26228
rect 13987 26188 13996 26228
rect 14036 26188 14956 26228
rect 14996 26188 16588 26228
rect 16628 26188 17644 26228
rect 17684 26188 18508 26228
rect 18548 26188 18892 26228
rect 18932 26188 19412 26228
rect 1324 26144 1364 26188
rect 4291 26187 4349 26188
rect 2851 26144 2909 26145
rect 19372 26144 19412 26188
rect 1315 26104 1324 26144
rect 1364 26104 1373 26144
rect 1507 26104 1516 26144
rect 1556 26104 2860 26144
rect 2900 26104 2909 26144
rect 6883 26104 6892 26144
rect 6932 26104 7468 26144
rect 7508 26104 7517 26144
rect 8707 26104 8716 26144
rect 8756 26104 9388 26144
rect 9428 26104 9868 26144
rect 9908 26104 9917 26144
rect 11203 26104 11212 26144
rect 11252 26104 19276 26144
rect 19316 26104 19325 26144
rect 19372 26104 19383 26144
rect 19423 26104 19432 26144
rect 2851 26103 2909 26104
rect 12259 26060 12317 26061
rect 739 26020 748 26060
rect 788 26020 1268 26060
rect 4195 26020 4204 26060
rect 4244 26020 8044 26060
rect 8084 26020 8093 26060
rect 8332 26020 11116 26060
rect 11156 26020 12268 26060
rect 12308 26020 12317 26060
rect 16675 26020 16684 26060
rect 16724 26020 19756 26060
rect 19796 26020 19805 26060
rect 0 25977 80 25996
rect 0 25976 125 25977
rect 1228 25976 1268 26020
rect 1411 25976 1469 25977
rect 8332 25976 8372 26020
rect 12259 26019 12317 26020
rect 21424 25976 21504 25996
rect 0 25936 76 25976
rect 116 25936 125 25976
rect 1219 25936 1228 25976
rect 1268 25936 1277 25976
rect 1411 25936 1420 25976
rect 1460 25936 8372 25976
rect 8800 25936 10580 25976
rect 10627 25936 10636 25976
rect 10676 25936 19372 25976
rect 19412 25936 19421 25976
rect 20995 25936 21004 25976
rect 21044 25936 21504 25976
rect 0 25935 125 25936
rect 1411 25935 1469 25936
rect 0 25916 80 25935
rect 7939 25892 7997 25893
rect 8800 25892 8840 25936
rect 10540 25892 10580 25936
rect 21424 25916 21504 25936
rect 11011 25892 11069 25893
rect 739 25852 748 25892
rect 788 25852 3820 25892
rect 3860 25852 3869 25892
rect 5827 25852 5836 25892
rect 5876 25852 7660 25892
rect 7700 25852 7709 25892
rect 7920 25852 7948 25892
rect 7988 25852 8044 25892
rect 8084 25852 8840 25892
rect 8899 25852 8908 25892
rect 8948 25852 10444 25892
rect 10484 25852 10493 25892
rect 10540 25852 11020 25892
rect 11060 25852 11069 25892
rect 11395 25852 11404 25892
rect 11444 25852 11980 25892
rect 12020 25852 12364 25892
rect 12404 25852 12413 25892
rect 14371 25852 14380 25892
rect 14420 25852 14764 25892
rect 14804 25852 14813 25892
rect 17251 25852 17260 25892
rect 17300 25852 17836 25892
rect 17876 25852 17885 25892
rect 7939 25851 7997 25852
rect 11011 25851 11069 25852
rect 5731 25808 5789 25809
rect 17443 25808 17501 25809
rect 17635 25808 17693 25809
rect 3043 25768 3052 25808
rect 3092 25768 5740 25808
rect 5780 25768 5789 25808
rect 8707 25768 8716 25808
rect 8756 25768 12748 25808
rect 12788 25768 12797 25808
rect 17347 25768 17356 25808
rect 17396 25768 17452 25808
rect 17492 25768 17501 25808
rect 17550 25768 17644 25808
rect 17684 25768 17693 25808
rect 5731 25767 5789 25768
rect 17443 25767 17501 25768
rect 17635 25767 17693 25768
rect 13987 25724 14045 25725
rect 3679 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 4065 25724
rect 4675 25684 4684 25724
rect 4724 25684 7564 25724
rect 7604 25684 7613 25724
rect 10051 25684 10060 25724
rect 10100 25684 10540 25724
rect 10580 25684 10589 25724
rect 13891 25684 13900 25724
rect 13940 25684 13996 25724
rect 14036 25684 14045 25724
rect 13987 25683 14045 25684
rect 16003 25724 16061 25725
rect 16003 25684 16012 25724
rect 16052 25684 18316 25724
rect 18356 25684 18365 25724
rect 18799 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 19185 25724
rect 16003 25683 16061 25684
rect 5827 25640 5885 25641
rect 17539 25640 17597 25641
rect 20899 25640 20957 25641
rect 21424 25640 21504 25660
rect 1315 25600 1324 25640
rect 1364 25600 2476 25640
rect 2516 25600 4052 25640
rect 835 25516 844 25556
rect 884 25516 2860 25556
rect 2900 25516 2909 25556
rect 0 25472 80 25492
rect 4012 25472 4052 25600
rect 4108 25600 5260 25640
rect 5300 25600 5836 25640
rect 5876 25600 12076 25640
rect 12116 25600 16012 25640
rect 16052 25600 17548 25640
rect 17588 25600 17740 25640
rect 17780 25600 17789 25640
rect 20899 25600 20908 25640
rect 20948 25600 21504 25640
rect 4108 25556 4148 25600
rect 5827 25599 5885 25600
rect 17539 25599 17597 25600
rect 20899 25599 20957 25600
rect 21424 25580 21504 25600
rect 6403 25556 6461 25557
rect 10531 25556 10589 25557
rect 12547 25556 12605 25557
rect 14755 25556 14813 25557
rect 4099 25516 4108 25556
rect 4148 25516 4157 25556
rect 6211 25516 6220 25556
rect 6260 25516 6412 25556
rect 6452 25516 6461 25556
rect 10446 25516 10540 25556
rect 10580 25516 10589 25556
rect 12462 25516 12556 25556
rect 12596 25516 12605 25556
rect 14659 25516 14668 25556
rect 14708 25516 14764 25556
rect 14804 25516 14813 25556
rect 15235 25516 15244 25556
rect 15284 25516 20180 25556
rect 6403 25515 6461 25516
rect 10531 25515 10589 25516
rect 12547 25515 12605 25516
rect 14755 25515 14813 25516
rect 12259 25472 12317 25473
rect 18019 25472 18077 25473
rect 0 25432 1324 25472
rect 1364 25432 1373 25472
rect 2083 25432 2092 25472
rect 2132 25432 2668 25472
rect 2708 25432 2717 25472
rect 4012 25432 8716 25472
rect 8756 25432 8765 25472
rect 12174 25432 12268 25472
rect 12308 25432 12317 25472
rect 13891 25432 13900 25472
rect 13940 25432 14284 25472
rect 14324 25432 14333 25472
rect 18019 25432 18028 25472
rect 18068 25432 18220 25472
rect 18260 25432 18269 25472
rect 18499 25432 18508 25472
rect 18548 25432 18892 25472
rect 18932 25432 18941 25472
rect 0 25412 80 25432
rect 12259 25431 12317 25432
rect 18019 25431 18077 25432
rect 3523 25388 3581 25389
rect 4579 25388 4637 25389
rect 7459 25388 7517 25389
rect 9667 25388 9725 25389
rect 10723 25388 10781 25389
rect 3523 25348 3532 25388
rect 3572 25348 4588 25388
rect 4628 25348 4684 25388
rect 4724 25348 4733 25388
rect 6019 25348 6028 25388
rect 6068 25348 7468 25388
rect 7508 25348 7517 25388
rect 9187 25348 9196 25388
rect 9236 25348 9484 25388
rect 9524 25348 9533 25388
rect 9667 25348 9676 25388
rect 9716 25348 10732 25388
rect 10772 25348 10781 25388
rect 3523 25347 3581 25348
rect 4579 25347 4637 25348
rect 7459 25347 7517 25348
rect 9667 25347 9725 25348
rect 10723 25347 10781 25348
rect 11107 25388 11165 25389
rect 12835 25388 12893 25389
rect 14563 25388 14621 25389
rect 11107 25348 11116 25388
rect 11156 25348 11596 25388
rect 11636 25348 12364 25388
rect 12404 25348 12413 25388
rect 12835 25348 12844 25388
rect 12884 25348 12940 25388
rect 12980 25348 12989 25388
rect 14467 25348 14476 25388
rect 14516 25348 14572 25388
rect 14612 25348 14621 25388
rect 17731 25348 17740 25388
rect 17780 25348 18604 25388
rect 18644 25348 18653 25388
rect 19267 25348 19276 25388
rect 19316 25348 19756 25388
rect 19796 25348 19805 25388
rect 11107 25347 11165 25348
rect 12835 25347 12893 25348
rect 14563 25347 14621 25348
rect 2659 25304 2717 25305
rect 5059 25304 5117 25305
rect 19363 25304 19421 25305
rect 2467 25264 2476 25304
rect 2516 25264 2668 25304
rect 2708 25264 2717 25304
rect 3235 25264 3244 25304
rect 3284 25264 3628 25304
rect 3668 25264 3677 25304
rect 4974 25264 5068 25304
rect 5108 25264 5117 25304
rect 9379 25264 9388 25304
rect 9428 25264 9964 25304
rect 10004 25264 10013 25304
rect 10819 25264 10828 25304
rect 10868 25264 12748 25304
rect 12788 25264 12797 25304
rect 14563 25264 14572 25304
rect 14612 25264 19372 25304
rect 19412 25264 19421 25304
rect 20140 25304 20180 25516
rect 21424 25304 21504 25324
rect 20140 25264 21504 25304
rect 2659 25263 2717 25264
rect 5059 25263 5117 25264
rect 19363 25263 19421 25264
rect 21424 25244 21504 25264
rect 163 25180 172 25220
rect 212 25180 1844 25220
rect 1804 25136 1844 25180
rect 2380 25180 3436 25220
rect 3476 25180 3485 25220
rect 4483 25180 4492 25220
rect 4532 25180 7180 25220
rect 7220 25180 7229 25220
rect 11971 25180 11980 25220
rect 12020 25180 12556 25220
rect 12596 25180 13996 25220
rect 14036 25180 14045 25220
rect 15139 25180 15148 25220
rect 15188 25180 15436 25220
rect 15476 25180 15485 25220
rect 17356 25180 17740 25220
rect 17780 25180 17789 25220
rect 17923 25180 17932 25220
rect 17972 25180 21196 25220
rect 21236 25180 21245 25220
rect 2380 25136 2420 25180
rect 17356 25136 17396 25180
rect 1804 25096 2420 25136
rect 12355 25096 12364 25136
rect 12404 25096 17164 25136
rect 17204 25096 17213 25136
rect 17347 25096 17356 25136
rect 17396 25096 17405 25136
rect 17827 25096 17836 25136
rect 17876 25096 18124 25136
rect 18164 25096 18173 25136
rect 20035 25096 20044 25136
rect 20084 25096 20180 25136
rect 2371 25052 2429 25053
rect 20140 25052 20180 25096
rect 1891 25012 1900 25052
rect 1940 25012 2380 25052
rect 2420 25012 2429 25052
rect 3139 25012 3148 25052
rect 3188 25012 13420 25052
rect 13460 25012 13804 25052
rect 13844 25012 13853 25052
rect 20140 25012 20756 25052
rect 2371 25011 2429 25012
rect 0 24968 80 24988
rect 6883 24968 6941 24969
rect 18691 24968 18749 24969
rect 0 24928 1324 24968
rect 1364 24928 1373 24968
rect 4919 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 5305 24968
rect 6883 24928 6892 24968
rect 6932 24928 6988 24968
rect 7028 24928 7037 24968
rect 7171 24928 7180 24968
rect 7220 24928 18700 24968
rect 18740 24928 18749 24968
rect 20039 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20425 24968
rect 0 24908 80 24928
rect 6883 24927 6941 24928
rect 18691 24927 18749 24928
rect 5635 24844 5644 24884
rect 5684 24844 6124 24884
rect 6164 24844 10196 24884
rect 739 24800 797 24801
rect 6403 24800 6461 24801
rect 6691 24800 6749 24801
rect 8515 24800 8573 24801
rect 739 24760 748 24800
rect 788 24760 3052 24800
rect 3092 24760 3101 24800
rect 6318 24760 6412 24800
rect 6452 24760 6461 24800
rect 6606 24760 6700 24800
rect 6740 24760 6988 24800
rect 7028 24760 7037 24800
rect 7459 24760 7468 24800
rect 7508 24760 8524 24800
rect 8564 24760 8573 24800
rect 10156 24800 10196 24844
rect 14764 24844 18412 24884
rect 18452 24844 18461 24884
rect 14764 24800 14804 24844
rect 14947 24800 15005 24801
rect 17251 24800 17309 24801
rect 19843 24800 19901 24801
rect 10156 24760 14804 24800
rect 14862 24760 14956 24800
rect 14996 24760 15005 24800
rect 17166 24760 17260 24800
rect 17300 24760 17309 24800
rect 18787 24760 18796 24800
rect 18836 24760 19276 24800
rect 19316 24760 19325 24800
rect 19758 24760 19852 24800
rect 19892 24760 19901 24800
rect 739 24759 797 24760
rect 6403 24759 6461 24760
rect 6691 24759 6749 24760
rect 8515 24759 8573 24760
rect 14947 24759 15005 24760
rect 17251 24759 17309 24760
rect 19843 24759 19901 24760
rect 6796 24676 10156 24716
rect 10196 24676 10205 24716
rect 11779 24676 11788 24716
rect 11828 24676 17452 24716
rect 17492 24676 17501 24716
rect 2467 24632 2525 24633
rect 4195 24632 4253 24633
rect 6796 24632 6836 24676
rect 10339 24632 10397 24633
rect 15235 24632 15293 24633
rect 2467 24592 2476 24632
rect 2516 24592 2540 24632
rect 3523 24592 3532 24632
rect 3572 24592 4204 24632
rect 4244 24592 4300 24632
rect 4340 24592 5548 24632
rect 5588 24592 5932 24632
rect 5972 24592 5981 24632
rect 6595 24592 6604 24632
rect 6644 24592 6796 24632
rect 6836 24592 6845 24632
rect 7171 24592 7180 24632
rect 7220 24592 7468 24632
rect 7508 24592 10060 24632
rect 10100 24592 10109 24632
rect 10339 24592 10348 24632
rect 10388 24592 15148 24632
rect 15188 24592 15244 24632
rect 15284 24592 15293 24632
rect 2467 24591 2540 24592
rect 4195 24591 4253 24592
rect 10339 24591 10397 24592
rect 15235 24591 15293 24592
rect 18019 24632 18077 24633
rect 20716 24632 20756 25012
rect 20803 24968 20861 24969
rect 21424 24968 21504 24988
rect 20803 24928 20812 24968
rect 20852 24928 21504 24968
rect 20803 24927 20861 24928
rect 21424 24908 21504 24928
rect 21424 24632 21504 24652
rect 18019 24592 18028 24632
rect 18068 24592 18316 24632
rect 18356 24592 18365 24632
rect 19747 24592 19756 24632
rect 19796 24592 20044 24632
rect 20084 24592 20093 24632
rect 20716 24592 21504 24632
rect 18019 24591 18077 24592
rect 2500 24548 2540 24591
rect 21424 24572 21504 24592
rect 8131 24548 8189 24549
rect 10915 24548 10973 24549
rect 2500 24508 3052 24548
rect 3092 24508 5836 24548
rect 5876 24508 5885 24548
rect 5932 24508 8140 24548
rect 8180 24508 8189 24548
rect 10830 24508 10924 24548
rect 10964 24508 10973 24548
rect 11107 24508 11116 24548
rect 11156 24508 12364 24548
rect 12404 24508 12413 24548
rect 13219 24508 13228 24548
rect 13268 24508 15628 24548
rect 15668 24508 15677 24548
rect 17155 24508 17164 24548
rect 17204 24508 19851 24548
rect 19891 24508 19900 24548
rect 0 24464 80 24484
rect 5932 24464 5972 24508
rect 8131 24507 8189 24508
rect 10915 24507 10973 24508
rect 15427 24464 15485 24465
rect 0 24404 116 24464
rect 1315 24424 1324 24464
rect 1364 24424 4684 24464
rect 4724 24424 5972 24464
rect 8131 24424 8140 24464
rect 8180 24424 9676 24464
rect 9716 24424 9964 24464
rect 10004 24424 10013 24464
rect 13891 24424 13900 24464
rect 13940 24424 14284 24464
rect 14324 24424 14764 24464
rect 14804 24424 14813 24464
rect 15427 24424 15436 24464
rect 15476 24424 19468 24464
rect 19508 24424 19517 24464
rect 15427 24423 15485 24424
rect 76 24380 116 24404
rect 2467 24380 2525 24381
rect 4195 24380 4253 24381
rect 13027 24380 13085 24381
rect 76 24340 2476 24380
rect 2516 24340 2525 24380
rect 3715 24340 3724 24380
rect 3764 24340 4204 24380
rect 4244 24340 4253 24380
rect 4483 24340 4492 24380
rect 4532 24340 6028 24380
rect 6068 24340 6077 24380
rect 6979 24340 6988 24380
rect 7028 24340 7276 24380
rect 7316 24340 7325 24380
rect 10147 24340 10156 24380
rect 10196 24340 10828 24380
rect 10868 24340 10877 24380
rect 13027 24340 13036 24380
rect 13076 24340 17972 24380
rect 2467 24339 2525 24340
rect 4195 24339 4253 24340
rect 13027 24339 13085 24340
rect 4204 24296 4244 24339
rect 14755 24296 14813 24297
rect 17932 24296 17972 24340
rect 21424 24296 21504 24316
rect 4204 24256 13228 24296
rect 13268 24256 13277 24296
rect 13603 24256 13612 24296
rect 13652 24256 14764 24296
rect 14804 24256 14813 24296
rect 16387 24256 16396 24296
rect 16436 24256 16684 24296
rect 16724 24256 16733 24296
rect 17923 24256 17932 24296
rect 17972 24256 17981 24296
rect 19939 24256 19948 24296
rect 19988 24256 21504 24296
rect 14755 24255 14813 24256
rect 21424 24236 21504 24256
rect 1795 24212 1853 24213
rect 11779 24212 11837 24213
rect 16483 24212 16541 24213
rect 1795 24172 1804 24212
rect 1844 24172 1996 24212
rect 2036 24172 2045 24212
rect 3679 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 4065 24212
rect 7459 24172 7468 24212
rect 7508 24172 11788 24212
rect 11828 24172 11837 24212
rect 1795 24171 1853 24172
rect 11779 24171 11837 24172
rect 13132 24172 16492 24212
rect 16532 24172 16541 24212
rect 18799 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 19185 24212
rect 1507 24128 1565 24129
rect 7267 24128 7325 24129
rect 1507 24088 1516 24128
rect 1556 24088 7276 24128
rect 7316 24088 7325 24128
rect 1507 24087 1565 24088
rect 7267 24087 7325 24088
rect 7363 24044 7421 24045
rect 7278 24004 7372 24044
rect 7412 24004 7421 24044
rect 7363 24003 7421 24004
rect 10051 24044 10109 24045
rect 13132 24044 13172 24172
rect 16483 24171 16541 24172
rect 15331 24128 15389 24129
rect 15331 24088 15340 24128
rect 15380 24088 19412 24128
rect 19555 24088 19564 24128
rect 19604 24088 21044 24128
rect 15331 24087 15389 24088
rect 10051 24004 10060 24044
rect 10100 24004 13172 24044
rect 13219 24044 13277 24045
rect 19267 24044 19325 24045
rect 13219 24004 13228 24044
rect 13268 24004 13362 24044
rect 13987 24004 13996 24044
rect 14036 24004 19276 24044
rect 19316 24004 19325 24044
rect 19372 24044 19412 24088
rect 20899 24044 20957 24045
rect 19372 24004 20908 24044
rect 20948 24004 20957 24044
rect 10051 24003 10109 24004
rect 13219 24003 13277 24004
rect 19267 24003 19325 24004
rect 20899 24003 20957 24004
rect 0 23961 80 23980
rect 0 23960 125 23961
rect 547 23960 605 23961
rect 8131 23960 8189 23961
rect 12643 23960 12701 23961
rect 13027 23960 13085 23961
rect 0 23920 76 23960
rect 116 23920 125 23960
rect 462 23920 556 23960
rect 596 23920 605 23960
rect 1507 23920 1516 23960
rect 1556 23920 2092 23960
rect 2132 23920 2141 23960
rect 6115 23920 6124 23960
rect 6164 23920 7660 23960
rect 7700 23920 7709 23960
rect 7939 23920 7948 23960
rect 7988 23920 8140 23960
rect 8180 23920 8189 23960
rect 9859 23920 9868 23960
rect 9908 23920 10732 23960
rect 10772 23920 11360 23960
rect 0 23919 125 23920
rect 547 23919 605 23920
rect 8131 23919 8189 23920
rect 0 23900 80 23919
rect 6691 23876 6749 23877
rect 11320 23876 11360 23920
rect 12643 23920 12652 23960
rect 12692 23920 12701 23960
rect 12942 23920 13036 23960
rect 13076 23920 13085 23960
rect 12643 23919 12701 23920
rect 13027 23919 13085 23920
rect 13603 23960 13661 23961
rect 16771 23960 16829 23961
rect 13603 23920 13612 23960
rect 13652 23920 14380 23960
rect 14420 23920 14429 23960
rect 14755 23920 14764 23960
rect 14804 23920 16780 23960
rect 16820 23920 16829 23960
rect 21004 23960 21044 24088
rect 21424 23960 21504 23980
rect 21004 23920 21504 23960
rect 13603 23919 13661 23920
rect 16771 23919 16829 23920
rect 12652 23876 12692 23919
rect 21424 23900 21504 23920
rect 6606 23836 6700 23876
rect 6740 23836 6749 23876
rect 9763 23836 9772 23876
rect 9812 23836 10388 23876
rect 11320 23836 12556 23876
rect 12596 23836 12605 23876
rect 12652 23836 13804 23876
rect 13844 23836 13853 23876
rect 15715 23836 15724 23876
rect 15764 23836 19948 23876
rect 19988 23836 19997 23876
rect 6691 23835 6749 23836
rect 10348 23792 10388 23836
rect 11779 23792 11837 23793
rect 12643 23792 12701 23793
rect 1411 23752 1420 23792
rect 1460 23752 2860 23792
rect 2900 23752 3340 23792
rect 3380 23752 3389 23792
rect 7075 23752 7084 23792
rect 7124 23752 8620 23792
rect 8660 23752 8669 23792
rect 8995 23752 9004 23792
rect 9044 23752 9388 23792
rect 9428 23752 10292 23792
rect 10348 23752 11788 23792
rect 11828 23752 11837 23792
rect 12558 23752 12652 23792
rect 12692 23752 12701 23792
rect 13891 23752 13900 23792
rect 13940 23752 14860 23792
rect 14900 23752 14909 23792
rect 17251 23752 17260 23792
rect 17300 23752 19180 23792
rect 19220 23752 19229 23792
rect 6403 23708 6461 23709
rect 7363 23708 7421 23709
rect 10252 23708 10292 23752
rect 11779 23751 11837 23752
rect 12643 23751 12701 23752
rect 6403 23668 6412 23708
rect 6452 23668 7372 23708
rect 7412 23668 9484 23708
rect 9524 23668 9533 23708
rect 10252 23668 10540 23708
rect 10580 23668 10589 23708
rect 11395 23668 11404 23708
rect 11444 23668 11596 23708
rect 11636 23668 11645 23708
rect 6403 23667 6461 23668
rect 7363 23667 7421 23668
rect 1891 23624 1949 23625
rect 8803 23624 8861 23625
rect 11299 23624 11357 23625
rect 13900 23624 13940 23752
rect 13987 23708 14045 23709
rect 18691 23708 18749 23709
rect 13987 23668 13996 23708
rect 14036 23668 14130 23708
rect 16195 23668 16204 23708
rect 16244 23668 17740 23708
rect 17780 23668 17789 23708
rect 18606 23668 18700 23708
rect 18740 23668 18749 23708
rect 13987 23667 14045 23668
rect 18691 23667 18749 23668
rect 1315 23584 1324 23624
rect 1364 23584 1708 23624
rect 1748 23584 1757 23624
rect 1806 23584 1900 23624
rect 1940 23584 1949 23624
rect 2083 23584 2092 23624
rect 2132 23584 2380 23624
rect 2420 23584 2429 23624
rect 6595 23584 6604 23624
rect 6644 23584 7180 23624
rect 7220 23584 7229 23624
rect 7555 23584 7564 23624
rect 7604 23584 8812 23624
rect 8852 23584 8861 23624
rect 10339 23584 10348 23624
rect 10388 23584 11308 23624
rect 11348 23584 13940 23624
rect 19843 23624 19901 23625
rect 21424 23624 21504 23644
rect 19843 23584 19852 23624
rect 19892 23584 21504 23624
rect 1891 23583 1949 23584
rect 8803 23583 8861 23584
rect 11299 23583 11357 23584
rect 19843 23583 19901 23584
rect 21424 23564 21504 23584
rect 9187 23540 9245 23541
rect 3043 23500 3052 23540
rect 3092 23500 9196 23540
rect 9236 23500 9245 23540
rect 9187 23499 9245 23500
rect 10243 23540 10301 23541
rect 10243 23500 10252 23540
rect 10292 23500 10301 23540
rect 10243 23499 10301 23500
rect 10348 23500 10924 23540
rect 10964 23500 15148 23540
rect 15188 23500 15197 23540
rect 17731 23500 17740 23540
rect 17780 23500 18028 23540
rect 18068 23500 18077 23540
rect 0 23456 80 23476
rect 7459 23456 7517 23457
rect 10252 23456 10292 23499
rect 10348 23456 10388 23500
rect 14755 23456 14813 23457
rect 0 23416 4204 23456
rect 4244 23416 4253 23456
rect 4919 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 5305 23456
rect 7459 23416 7468 23456
rect 7508 23416 10292 23456
rect 10339 23416 10348 23456
rect 10388 23416 10397 23456
rect 14670 23416 14764 23456
rect 14804 23416 16492 23456
rect 16532 23416 16541 23456
rect 20039 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20425 23456
rect 0 23396 80 23416
rect 7459 23415 7517 23416
rect 14755 23415 14813 23416
rect 7468 23372 7508 23415
rect 9283 23372 9341 23373
rect 1315 23332 1324 23372
rect 1364 23332 3956 23372
rect 4003 23332 4012 23372
rect 4052 23332 4684 23372
rect 4724 23332 7508 23372
rect 8323 23332 8332 23372
rect 8372 23332 9292 23372
rect 9332 23332 16780 23372
rect 16820 23332 18220 23372
rect 18260 23332 18269 23372
rect 3916 23288 3956 23332
rect 9283 23331 9341 23332
rect 6307 23288 6365 23289
rect 7843 23288 7901 23289
rect 1027 23248 1036 23288
rect 1076 23248 1516 23288
rect 1556 23248 1565 23288
rect 1987 23248 1996 23288
rect 2036 23248 3628 23288
rect 3668 23248 3677 23288
rect 3916 23248 6316 23288
rect 6356 23248 6365 23288
rect 6595 23248 6604 23288
rect 6644 23248 7852 23288
rect 7892 23248 7901 23288
rect 6307 23247 6365 23248
rect 7843 23247 7901 23248
rect 8515 23288 8573 23289
rect 16867 23288 16925 23289
rect 19939 23288 19997 23289
rect 21424 23288 21504 23308
rect 8515 23248 8524 23288
rect 8564 23248 11360 23288
rect 13315 23248 13324 23288
rect 13364 23248 16876 23288
rect 16916 23248 16925 23288
rect 19651 23248 19660 23288
rect 19700 23248 19709 23288
rect 19939 23248 19948 23288
rect 19988 23248 21504 23288
rect 8515 23247 8573 23248
rect 2467 23204 2525 23205
rect 5923 23204 5981 23205
rect 2382 23164 2476 23204
rect 2516 23164 2956 23204
rect 2996 23164 3005 23204
rect 5923 23164 5932 23204
rect 5972 23164 8908 23204
rect 8948 23164 8957 23204
rect 2467 23163 2525 23164
rect 5923 23163 5981 23164
rect 1219 23120 1277 23121
rect 11320 23120 11360 23248
rect 16867 23247 16925 23248
rect 19660 23204 19700 23248
rect 19939 23247 19997 23248
rect 21424 23228 21504 23248
rect 12067 23164 12076 23204
rect 12116 23164 15916 23204
rect 15956 23164 15965 23204
rect 19660 23164 20852 23204
rect 1219 23080 1228 23120
rect 1268 23080 1708 23120
rect 1748 23080 1757 23120
rect 2851 23080 2860 23120
rect 2900 23080 3148 23120
rect 3188 23080 3197 23120
rect 3715 23080 3724 23120
rect 3764 23080 4108 23120
rect 4148 23080 4157 23120
rect 5155 23080 5164 23120
rect 5204 23080 7468 23120
rect 7508 23080 7517 23120
rect 10435 23080 10444 23120
rect 10484 23080 10732 23120
rect 10772 23080 10781 23120
rect 11320 23080 13516 23120
rect 13556 23080 13565 23120
rect 14179 23080 14188 23120
rect 14228 23080 17356 23120
rect 17396 23080 17405 23120
rect 18403 23080 18412 23120
rect 18452 23080 18988 23120
rect 19028 23080 19037 23120
rect 19171 23080 19180 23120
rect 19220 23080 19988 23120
rect 1219 23079 1277 23080
rect 2179 23036 2237 23037
rect 3331 23036 3389 23037
rect 4579 23036 4637 23037
rect 2179 22996 2188 23036
rect 2228 22996 3340 23036
rect 3380 22996 4300 23036
rect 4340 22996 4349 23036
rect 4494 22996 4588 23036
rect 4628 22996 4637 23036
rect 2179 22995 2237 22996
rect 3331 22995 3389 22996
rect 4579 22995 4637 22996
rect 5923 23036 5981 23037
rect 6403 23036 6461 23037
rect 5923 22996 5932 23036
rect 5972 22996 6028 23036
rect 6068 22996 6077 23036
rect 6318 22996 6412 23036
rect 6452 22996 6461 23036
rect 5923 22995 5981 22996
rect 6403 22995 6461 22996
rect 10723 23036 10781 23037
rect 19948 23036 19988 23080
rect 10723 22996 10732 23036
rect 10772 22996 13132 23036
rect 13172 22996 15244 23036
rect 15284 22996 15628 23036
rect 15668 22996 15677 23036
rect 19267 22996 19276 23036
rect 19316 22996 19756 23036
rect 19796 22996 19805 23036
rect 19939 22996 19948 23036
rect 19988 22996 19997 23036
rect 10723 22995 10781 22996
rect 0 22952 80 22972
rect 19756 22952 19796 22996
rect 20812 22952 20852 23164
rect 21424 22952 21504 22972
rect 0 22912 1804 22952
rect 1844 22912 1853 22952
rect 5827 22912 5836 22952
rect 5876 22912 10060 22952
rect 10100 22912 16108 22952
rect 16148 22912 16157 22952
rect 19075 22912 19084 22952
rect 19124 22912 19372 22952
rect 19412 22912 19421 22952
rect 19756 22912 20140 22952
rect 20180 22912 20189 22952
rect 20812 22912 21504 22952
rect 0 22892 80 22912
rect 21424 22892 21504 22912
rect 6211 22868 6269 22869
rect 3139 22828 3148 22868
rect 3188 22828 4204 22868
rect 4244 22828 4253 22868
rect 4387 22828 4396 22868
rect 4436 22828 4972 22868
rect 5012 22828 5021 22868
rect 6126 22828 6220 22868
rect 6260 22828 6269 22868
rect 6211 22827 6269 22828
rect 6691 22868 6749 22869
rect 12067 22868 12125 22869
rect 6691 22828 6700 22868
rect 6740 22828 11404 22868
rect 11444 22828 12076 22868
rect 12116 22828 12125 22868
rect 6691 22827 6749 22828
rect 12067 22827 12125 22828
rect 13027 22868 13085 22869
rect 13027 22828 13036 22868
rect 13076 22828 15916 22868
rect 15956 22828 15965 22868
rect 18787 22828 18796 22868
rect 18836 22828 19276 22868
rect 19316 22828 19325 22868
rect 19555 22828 19564 22868
rect 19604 22828 19948 22868
rect 19988 22828 19997 22868
rect 13027 22827 13085 22828
rect 2755 22784 2813 22785
rect 7171 22784 7229 22785
rect 19459 22784 19517 22785
rect 1603 22744 1612 22784
rect 1652 22744 2764 22784
rect 2804 22744 7180 22784
rect 7220 22744 7229 22784
rect 7843 22744 7852 22784
rect 7892 22744 9676 22784
rect 9716 22744 10252 22784
rect 10292 22744 10301 22784
rect 12643 22744 12652 22784
rect 12692 22744 14572 22784
rect 14612 22744 14621 22784
rect 15427 22744 15436 22784
rect 15476 22744 19468 22784
rect 19508 22744 20236 22784
rect 20276 22744 20285 22784
rect 2755 22743 2813 22744
rect 7171 22743 7229 22744
rect 19459 22743 19517 22744
rect 16291 22700 16349 22701
rect 3679 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 4065 22700
rect 7267 22660 7276 22700
rect 7316 22660 7756 22700
rect 7796 22660 7805 22700
rect 10051 22660 10060 22700
rect 10100 22660 10540 22700
rect 10580 22660 10589 22700
rect 11404 22660 11788 22700
rect 11828 22660 11837 22700
rect 13219 22660 13228 22700
rect 13268 22660 13612 22700
rect 13652 22660 13661 22700
rect 15523 22660 15532 22700
rect 15572 22660 16300 22700
rect 16340 22660 16349 22700
rect 259 22616 317 22617
rect 10252 22616 10292 22660
rect 11404 22616 11444 22660
rect 16291 22659 16349 22660
rect 16771 22700 16829 22701
rect 19363 22700 19421 22701
rect 16771 22660 16780 22700
rect 16820 22660 16876 22700
rect 16916 22660 16925 22700
rect 18799 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 19185 22700
rect 19363 22660 19372 22700
rect 19412 22660 19660 22700
rect 19700 22660 19709 22700
rect 16771 22659 16829 22660
rect 19363 22659 19421 22660
rect 21424 22616 21504 22636
rect 259 22576 268 22616
rect 308 22576 1708 22616
rect 1748 22576 1757 22616
rect 3724 22576 9196 22616
rect 9236 22576 9245 22616
rect 10243 22576 10252 22616
rect 10292 22576 10301 22616
rect 11395 22576 11404 22616
rect 11444 22576 11453 22616
rect 11692 22576 18124 22616
rect 18164 22576 18173 22616
rect 20515 22576 20524 22616
rect 20564 22576 21504 22616
rect 259 22575 317 22576
rect 931 22532 989 22533
rect 3724 22532 3764 22576
rect 6595 22532 6653 22533
rect 11692 22532 11732 22576
rect 21424 22556 21504 22576
rect 13603 22532 13661 22533
rect 931 22492 940 22532
rect 980 22492 1516 22532
rect 1556 22492 1565 22532
rect 3715 22492 3724 22532
rect 3764 22492 3773 22532
rect 4483 22492 4492 22532
rect 4532 22492 6604 22532
rect 6644 22492 6653 22532
rect 7363 22492 7372 22532
rect 7412 22492 11692 22532
rect 11732 22492 11741 22532
rect 13507 22492 13516 22532
rect 13556 22492 13612 22532
rect 13652 22492 13661 22532
rect 14179 22492 14188 22532
rect 14228 22492 15052 22532
rect 15092 22492 15101 22532
rect 17155 22492 17164 22532
rect 17204 22492 19276 22532
rect 19316 22492 19660 22532
rect 19700 22492 19709 22532
rect 931 22491 989 22492
rect 6595 22491 6653 22492
rect 13603 22491 13661 22492
rect 0 22448 80 22468
rect 1219 22448 1277 22449
rect 4675 22448 4733 22449
rect 13987 22448 14045 22449
rect 0 22408 1228 22448
rect 1268 22408 1277 22448
rect 4590 22408 4684 22448
rect 4724 22408 4733 22448
rect 6691 22408 6700 22448
rect 6740 22408 6988 22448
rect 7028 22408 7276 22448
rect 7316 22408 7325 22448
rect 11299 22408 11308 22448
rect 11348 22408 13612 22448
rect 13652 22408 13661 22448
rect 13987 22408 13996 22448
rect 14036 22408 14284 22448
rect 14324 22408 14333 22448
rect 0 22388 80 22408
rect 1219 22407 1277 22408
rect 4675 22407 4733 22408
rect 13987 22407 14045 22408
rect 2659 22364 2717 22365
rect 7843 22364 7901 22365
rect 13411 22364 13469 22365
rect 2371 22324 2380 22364
rect 2420 22324 2668 22364
rect 2708 22324 2717 22364
rect 4291 22324 4300 22364
rect 4340 22324 7852 22364
rect 7892 22324 7901 22364
rect 11875 22324 11884 22364
rect 11924 22324 12268 22364
rect 12308 22324 12317 22364
rect 12931 22324 12940 22364
rect 12980 22324 13132 22364
rect 13172 22324 13181 22364
rect 13315 22324 13324 22364
rect 13364 22324 13420 22364
rect 13460 22324 15820 22364
rect 15860 22324 15869 22364
rect 2659 22323 2717 22324
rect 7843 22323 7901 22324
rect 13411 22323 13469 22324
rect 19651 22280 19709 22281
rect 21424 22280 21504 22300
rect 3619 22240 3628 22280
rect 3668 22240 6220 22280
rect 6260 22240 6892 22280
rect 6932 22240 6941 22280
rect 10051 22240 10060 22280
rect 10100 22240 14284 22280
rect 14324 22240 14333 22280
rect 16579 22240 16588 22280
rect 16628 22240 16780 22280
rect 16820 22240 17164 22280
rect 17204 22240 18412 22280
rect 18452 22240 18604 22280
rect 18644 22240 19084 22280
rect 19124 22240 19133 22280
rect 19651 22240 19660 22280
rect 19700 22240 21504 22280
rect 4483 22196 4541 22197
rect 6892 22196 6932 22240
rect 19651 22239 19709 22240
rect 21424 22220 21504 22240
rect 15907 22196 15965 22197
rect 2179 22156 2188 22196
rect 2228 22156 4492 22196
rect 4532 22156 5932 22196
rect 5972 22156 5981 22196
rect 6892 22156 8140 22196
rect 8180 22156 8189 22196
rect 11779 22156 11788 22196
rect 11828 22156 13900 22196
rect 13940 22156 14188 22196
rect 14228 22156 14237 22196
rect 15523 22156 15532 22196
rect 15572 22156 15916 22196
rect 15956 22156 15965 22196
rect 17347 22156 17356 22196
rect 17396 22156 18700 22196
rect 18740 22156 19468 22196
rect 19508 22156 19517 22196
rect 4483 22155 4541 22156
rect 15907 22155 15965 22156
rect 12643 22112 12701 22113
rect 16579 22112 16637 22113
rect 17539 22112 17597 22113
rect 6403 22072 6412 22112
rect 6452 22072 7660 22112
rect 7700 22072 7709 22112
rect 8419 22072 8428 22112
rect 8468 22072 11692 22112
rect 11732 22072 11741 22112
rect 12643 22072 12652 22112
rect 12692 22072 12940 22112
rect 12980 22072 12989 22112
rect 16579 22072 16588 22112
rect 16628 22072 17548 22112
rect 17588 22072 17597 22112
rect 20131 22072 20140 22112
rect 20180 22072 21332 22112
rect 12643 22071 12701 22072
rect 16579 22071 16637 22072
rect 17539 22071 17597 22072
rect 451 22028 509 22029
rect 9187 22028 9245 22029
rect 12739 22028 12797 22029
rect 451 21988 460 22028
rect 500 21988 2284 22028
rect 2324 21988 2333 22028
rect 3139 21988 3148 22028
rect 3188 21988 9196 22028
rect 9236 21988 9292 22028
rect 9332 21988 11308 22028
rect 11348 21988 11357 22028
rect 11587 21988 11596 22028
rect 11636 21988 12748 22028
rect 12788 21988 17836 22028
rect 17876 21988 17885 22028
rect 451 21987 509 21988
rect 9187 21987 9245 21988
rect 12739 21987 12797 21988
rect 0 21944 80 21964
rect 1027 21944 1085 21945
rect 6883 21944 6941 21945
rect 15907 21944 15965 21945
rect 21292 21944 21332 22072
rect 21424 21944 21504 21964
rect 0 21904 1036 21944
rect 1076 21904 1085 21944
rect 4919 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 5305 21944
rect 6499 21904 6508 21944
rect 6548 21904 6892 21944
rect 6932 21904 6941 21944
rect 15822 21904 15916 21944
rect 15956 21904 15965 21944
rect 20039 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20425 21944
rect 21292 21904 21504 21944
rect 0 21884 80 21904
rect 1027 21903 1085 21904
rect 6883 21903 6941 21904
rect 15907 21903 15965 21904
rect 21424 21884 21504 21904
rect 259 21820 268 21860
rect 308 21820 3148 21860
rect 3188 21820 3197 21860
rect 6403 21820 6412 21860
rect 6452 21820 6796 21860
rect 6836 21820 6845 21860
rect 12835 21820 12844 21860
rect 12884 21820 13516 21860
rect 13556 21820 14764 21860
rect 14804 21820 14813 21860
rect 1123 21776 1181 21777
rect 1891 21776 1949 21777
rect 3523 21776 3581 21777
rect 3715 21776 3773 21777
rect 4483 21776 4541 21777
rect 6979 21776 7037 21777
rect 1123 21736 1132 21776
rect 1172 21736 1516 21776
rect 1556 21736 1565 21776
rect 1806 21736 1900 21776
rect 1940 21736 1949 21776
rect 1123 21735 1181 21736
rect 1891 21735 1949 21736
rect 2500 21736 3532 21776
rect 3572 21736 3724 21776
rect 3764 21736 3773 21776
rect 4291 21736 4300 21776
rect 4340 21736 4349 21776
rect 4483 21736 4492 21776
rect 4532 21736 6988 21776
rect 7028 21736 7037 21776
rect 10723 21736 10732 21776
rect 10772 21736 11884 21776
rect 11924 21736 11933 21776
rect 13987 21736 13996 21776
rect 14036 21736 14284 21776
rect 14324 21736 14333 21776
rect 17635 21736 17644 21776
rect 17684 21736 19372 21776
rect 19412 21736 20044 21776
rect 20084 21736 20093 21776
rect 2500 21692 2540 21736
rect 3523 21735 3581 21736
rect 3715 21735 3773 21736
rect 4300 21692 4340 21736
rect 4483 21735 4541 21736
rect 6979 21735 7037 21736
rect 1315 21652 1324 21692
rect 1364 21652 2540 21692
rect 2755 21652 2764 21692
rect 2804 21652 4108 21692
rect 4148 21652 4157 21692
rect 4300 21652 4876 21692
rect 4916 21652 4925 21692
rect 6019 21652 6028 21692
rect 6068 21652 9620 21692
rect 13219 21652 13228 21692
rect 13268 21652 13900 21692
rect 13940 21652 15532 21692
rect 15572 21652 15581 21692
rect 18115 21652 18124 21692
rect 18164 21652 18796 21692
rect 18836 21652 18845 21692
rect 9580 21609 9620 21652
rect 3043 21608 3101 21609
rect 9571 21608 9629 21609
rect 20611 21608 20669 21609
rect 21424 21608 21504 21628
rect 1027 21568 1036 21608
rect 1076 21568 2668 21608
rect 2708 21568 2717 21608
rect 2958 21568 3052 21608
rect 3092 21568 3101 21608
rect 3811 21568 3820 21608
rect 3860 21568 6124 21608
rect 6164 21568 6173 21608
rect 6595 21568 6604 21608
rect 6644 21568 7124 21608
rect 7171 21568 7180 21608
rect 7220 21568 7756 21608
rect 7796 21568 7805 21608
rect 9091 21568 9100 21608
rect 9140 21568 9388 21608
rect 9428 21568 9437 21608
rect 9571 21568 9580 21608
rect 9620 21568 9676 21608
rect 9716 21568 9725 21608
rect 10435 21568 10444 21608
rect 10484 21568 10924 21608
rect 10964 21568 10973 21608
rect 11320 21568 12268 21608
rect 12308 21568 17164 21608
rect 17204 21568 17213 21608
rect 18019 21568 18028 21608
rect 18068 21568 18604 21608
rect 18644 21568 19468 21608
rect 19508 21568 19517 21608
rect 20611 21568 20620 21608
rect 20660 21568 21504 21608
rect 3043 21567 3101 21568
rect 451 21524 509 21525
rect 1411 21524 1469 21525
rect 2083 21524 2141 21525
rect 3235 21524 3293 21525
rect 7084 21524 7124 21568
rect 9571 21567 9629 21568
rect 11320 21524 11360 21568
rect 20611 21567 20669 21568
rect 21424 21548 21504 21568
rect 16195 21524 16253 21525
rect 451 21484 460 21524
rect 500 21484 1268 21524
rect 451 21483 509 21484
rect 0 21440 80 21460
rect 1228 21440 1268 21484
rect 1411 21484 1420 21524
rect 1460 21484 1554 21524
rect 1997 21484 2092 21524
rect 2132 21484 3244 21524
rect 3284 21484 3436 21524
rect 3476 21484 3485 21524
rect 6691 21484 6700 21524
rect 6740 21484 6988 21524
rect 7028 21484 7037 21524
rect 7084 21484 7276 21524
rect 7316 21484 7468 21524
rect 7508 21484 7517 21524
rect 8515 21484 8524 21524
rect 8564 21484 11360 21524
rect 11596 21484 13460 21524
rect 14755 21484 14764 21524
rect 14804 21484 15148 21524
rect 15188 21484 16204 21524
rect 16244 21484 16253 21524
rect 16963 21484 16972 21524
rect 17012 21484 19276 21524
rect 19316 21484 19948 21524
rect 19988 21484 19997 21524
rect 1411 21483 1469 21484
rect 2083 21483 2141 21484
rect 3235 21483 3293 21484
rect 11596 21440 11636 21484
rect 13420 21440 13460 21484
rect 16195 21483 16253 21484
rect 0 21400 1132 21440
rect 1172 21400 1181 21440
rect 1228 21400 3628 21440
rect 3668 21400 3677 21440
rect 5251 21400 5260 21440
rect 5300 21400 11636 21440
rect 11683 21400 11692 21440
rect 11732 21400 13324 21440
rect 13364 21400 13373 21440
rect 13420 21400 17300 21440
rect 17347 21400 17356 21440
rect 17396 21400 19756 21440
rect 19796 21400 19805 21440
rect 0 21380 80 21400
rect 5347 21356 5405 21357
rect 9667 21356 9725 21357
rect 13219 21356 13277 21357
rect 5155 21316 5164 21356
rect 5204 21316 5356 21356
rect 5396 21316 5405 21356
rect 6307 21316 6316 21356
rect 6356 21316 7084 21356
rect 7124 21316 7133 21356
rect 9571 21316 9580 21356
rect 9620 21316 9676 21356
rect 9716 21316 9725 21356
rect 5347 21315 5405 21316
rect 9667 21315 9725 21316
rect 11320 21316 12652 21356
rect 12692 21316 12701 21356
rect 13219 21316 13228 21356
rect 13268 21316 16204 21356
rect 16244 21316 16253 21356
rect 1891 21272 1949 21273
rect 7267 21272 7325 21273
rect 11320 21272 11360 21316
rect 13219 21315 13277 21316
rect 17260 21272 17300 21400
rect 19363 21356 19421 21357
rect 17539 21316 17548 21356
rect 17588 21316 18316 21356
rect 18356 21316 18365 21356
rect 19278 21316 19372 21356
rect 19412 21316 19421 21356
rect 19363 21315 19421 21316
rect 17635 21272 17693 21273
rect 1891 21232 1900 21272
rect 1940 21232 5356 21272
rect 5396 21232 5405 21272
rect 7267 21232 7276 21272
rect 7316 21232 9004 21272
rect 9044 21232 9053 21272
rect 9667 21232 9676 21272
rect 9716 21232 11360 21272
rect 13987 21232 13996 21272
rect 14036 21232 14668 21272
rect 14708 21232 14717 21272
rect 17260 21232 17644 21272
rect 17684 21232 17693 21272
rect 1891 21231 1949 21232
rect 7267 21231 7325 21232
rect 17635 21231 17693 21232
rect 21283 21272 21341 21273
rect 21424 21272 21504 21292
rect 21283 21232 21292 21272
rect 21332 21232 21504 21272
rect 21283 21231 21341 21232
rect 21424 21212 21504 21232
rect 3679 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 4065 21188
rect 4108 21148 5548 21188
rect 5588 21148 5597 21188
rect 6595 21148 6604 21188
rect 6644 21148 6892 21188
rect 6932 21148 6941 21188
rect 7747 21148 7756 21188
rect 7796 21148 14284 21188
rect 14324 21148 14333 21188
rect 17635 21148 17644 21188
rect 17684 21148 17932 21188
rect 17972 21148 17981 21188
rect 18799 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 19185 21188
rect 4108 21104 4148 21148
rect 12835 21104 12893 21105
rect 2947 21064 2956 21104
rect 2996 21064 4148 21104
rect 4195 21064 4204 21104
rect 4244 21064 12844 21104
rect 12884 21064 12893 21104
rect 12835 21063 12893 21064
rect 15619 21104 15677 21105
rect 17443 21104 17501 21105
rect 15619 21064 15628 21104
rect 15668 21064 15724 21104
rect 15764 21064 15773 21104
rect 17443 21064 17452 21104
rect 17492 21064 17836 21104
rect 17876 21064 17885 21104
rect 15619 21063 15677 21064
rect 17443 21063 17501 21064
rect 1507 21020 1565 21021
rect 11587 21020 11645 21021
rect 1422 20980 1516 21020
rect 1556 20980 1565 21020
rect 2275 20980 2284 21020
rect 2324 20980 4148 21020
rect 1507 20979 1565 20980
rect 0 20936 80 20956
rect 4108 20936 4148 20980
rect 4300 20980 11596 21020
rect 11636 20980 11645 21020
rect 4300 20936 4340 20980
rect 11587 20979 11645 20980
rect 17740 20980 19372 21020
rect 19412 20980 19564 21020
rect 19604 20980 19613 21020
rect 0 20896 76 20936
rect 116 20896 125 20936
rect 4108 20896 4340 20936
rect 4483 20896 4492 20936
rect 4532 20896 8812 20936
rect 8852 20896 8861 20936
rect 8995 20896 9004 20936
rect 9044 20896 16972 20936
rect 17012 20896 17021 20936
rect 0 20876 80 20896
rect 1411 20852 1469 20853
rect 4291 20852 4349 20853
rect 12163 20852 12221 20853
rect 17740 20852 17780 20980
rect 19939 20936 19997 20937
rect 21424 20936 21504 20956
rect 19939 20896 19948 20936
rect 19988 20896 21504 20936
rect 19939 20895 19997 20896
rect 21424 20876 21504 20896
rect 1315 20812 1324 20852
rect 1364 20812 1420 20852
rect 1460 20812 1469 20852
rect 2947 20812 2956 20852
rect 2996 20812 3340 20852
rect 3380 20812 3389 20852
rect 4206 20812 4300 20852
rect 4340 20812 4349 20852
rect 5347 20812 5356 20852
rect 5396 20812 6028 20852
rect 6068 20812 6077 20852
rect 6211 20812 6220 20852
rect 6260 20812 12172 20852
rect 12212 20812 12221 20852
rect 12643 20812 12652 20852
rect 12692 20812 13708 20852
rect 13748 20812 13757 20852
rect 14275 20812 14284 20852
rect 14324 20812 15916 20852
rect 15956 20812 17780 20852
rect 17827 20812 17836 20852
rect 17876 20812 19084 20852
rect 19124 20812 19133 20852
rect 1411 20811 1469 20812
rect 4291 20811 4349 20812
rect 12163 20811 12221 20812
rect 5539 20768 5597 20769
rect 2467 20728 2476 20768
rect 2516 20728 5548 20768
rect 5588 20728 5597 20768
rect 5539 20727 5597 20728
rect 5923 20768 5981 20769
rect 11587 20768 11645 20769
rect 5923 20728 5932 20768
rect 5972 20728 9676 20768
rect 9716 20728 9725 20768
rect 11395 20728 11404 20768
rect 11444 20728 11596 20768
rect 11636 20728 11645 20768
rect 13027 20728 13036 20768
rect 13076 20728 13085 20768
rect 15523 20728 15532 20768
rect 15572 20728 16204 20768
rect 16244 20728 16253 20768
rect 16483 20728 16492 20768
rect 16532 20728 16876 20768
rect 16916 20728 16925 20768
rect 17443 20728 17452 20768
rect 17492 20728 18508 20768
rect 18548 20728 20236 20768
rect 20276 20728 20285 20768
rect 5923 20727 5981 20728
rect 11587 20727 11645 20728
rect 9859 20684 9917 20685
rect 13036 20684 13076 20728
rect 4099 20644 4108 20684
rect 4148 20644 4972 20684
rect 5012 20644 5021 20684
rect 6115 20644 6124 20684
rect 6164 20644 9868 20684
rect 9908 20644 9917 20684
rect 12739 20644 12748 20684
rect 12788 20644 13076 20684
rect 9859 20643 9917 20644
rect 14179 20600 14237 20601
rect 15427 20600 15485 20601
rect 1699 20560 1708 20600
rect 1748 20560 3820 20600
rect 3860 20560 3869 20600
rect 11683 20560 11692 20600
rect 11732 20560 12076 20600
rect 12116 20560 12125 20600
rect 12547 20560 12556 20600
rect 12596 20560 14188 20600
rect 14228 20560 14237 20600
rect 14755 20560 14764 20600
rect 14804 20560 15436 20600
rect 15476 20560 15485 20600
rect 15619 20560 15628 20600
rect 15668 20560 16012 20600
rect 16052 20560 16061 20600
rect 14179 20559 14237 20560
rect 15427 20559 15485 20560
rect 2371 20516 2429 20517
rect 2286 20476 2380 20516
rect 2420 20476 2429 20516
rect 9187 20476 9196 20516
rect 9236 20476 11500 20516
rect 11540 20476 14092 20516
rect 14132 20476 14141 20516
rect 2371 20475 2429 20476
rect 0 20432 80 20452
rect 259 20432 317 20433
rect 0 20392 268 20432
rect 308 20392 317 20432
rect 0 20372 80 20392
rect 259 20391 317 20392
rect 2563 20432 2621 20433
rect 16204 20432 16244 20728
rect 16387 20684 16445 20685
rect 16387 20644 16396 20684
rect 16436 20644 16530 20684
rect 18211 20644 18220 20684
rect 18260 20644 20044 20684
rect 20084 20644 20093 20684
rect 16387 20643 16445 20644
rect 19747 20600 19805 20601
rect 21424 20600 21504 20620
rect 19662 20560 19756 20600
rect 19796 20560 19805 20600
rect 19747 20559 19805 20560
rect 19852 20560 21504 20600
rect 19852 20517 19892 20560
rect 21424 20540 21504 20560
rect 19843 20516 19901 20517
rect 16771 20476 16780 20516
rect 16820 20476 17260 20516
rect 17300 20476 17309 20516
rect 19843 20476 19852 20516
rect 19892 20476 19901 20516
rect 19843 20475 19901 20476
rect 2563 20392 2572 20432
rect 2612 20392 3244 20432
rect 3284 20392 3293 20432
rect 4919 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 5305 20432
rect 6019 20392 6028 20432
rect 6068 20392 9484 20432
rect 9524 20392 9533 20432
rect 16204 20392 16396 20432
rect 16436 20392 16445 20432
rect 19555 20392 19564 20432
rect 19604 20392 19852 20432
rect 19892 20392 19901 20432
rect 20039 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20425 20432
rect 2563 20391 2621 20392
rect 3139 20348 3197 20349
rect 9484 20348 9524 20392
rect 14179 20348 14237 20349
rect 3054 20308 3148 20348
rect 3188 20308 3436 20348
rect 3476 20308 3485 20348
rect 9484 20308 13228 20348
rect 13268 20308 13277 20348
rect 14179 20308 14188 20348
rect 14228 20308 16148 20348
rect 16195 20308 16204 20348
rect 16244 20308 16492 20348
rect 16532 20308 16541 20348
rect 18499 20308 18508 20348
rect 18548 20308 19276 20348
rect 19316 20308 19325 20348
rect 3139 20307 3197 20308
rect 14179 20307 14237 20308
rect 12355 20264 12413 20265
rect 12643 20264 12701 20265
rect 16108 20264 16148 20308
rect 21424 20264 21504 20284
rect 67 20224 76 20264
rect 116 20224 12364 20264
rect 12404 20224 12413 20264
rect 12558 20224 12652 20264
rect 12692 20224 12701 20264
rect 12355 20223 12413 20224
rect 12643 20223 12701 20224
rect 13228 20224 13996 20264
rect 14036 20224 14045 20264
rect 14956 20224 15052 20264
rect 15092 20224 15101 20264
rect 16108 20224 16684 20264
rect 16724 20224 17260 20264
rect 17300 20224 17309 20264
rect 18019 20224 18028 20264
rect 18068 20224 18604 20264
rect 18644 20224 18653 20264
rect 19948 20224 21504 20264
rect 13228 20180 13268 20224
rect 13603 20180 13661 20181
rect 14755 20180 14813 20181
rect 2916 20140 2956 20180
rect 2996 20140 3005 20180
rect 13219 20140 13228 20180
rect 13268 20140 13277 20180
rect 13518 20140 13612 20180
rect 13652 20140 13661 20180
rect 14670 20140 14764 20180
rect 14804 20140 14813 20180
rect 2956 20096 2996 20140
rect 13603 20139 13661 20140
rect 14755 20139 14813 20140
rect 12259 20096 12317 20097
rect 2956 20056 5164 20096
rect 5204 20056 5213 20096
rect 6883 20056 6892 20096
rect 6932 20056 9196 20096
rect 9236 20056 9245 20096
rect 9571 20056 9580 20096
rect 9620 20056 9964 20096
rect 10004 20056 10013 20096
rect 11107 20056 11116 20096
rect 11156 20056 11500 20096
rect 11540 20056 11549 20096
rect 11971 20056 11980 20096
rect 12020 20056 12268 20096
rect 12308 20056 12317 20096
rect 12259 20055 12317 20056
rect 8227 20012 8285 20013
rect 14956 20012 14996 20224
rect 17539 20180 17597 20181
rect 15235 20140 15244 20180
rect 15284 20140 15293 20180
rect 17454 20140 17548 20180
rect 17588 20140 17597 20180
rect 15244 20012 15284 20140
rect 17539 20139 17597 20140
rect 18691 20180 18749 20181
rect 18691 20140 18700 20180
rect 18740 20140 19276 20180
rect 19316 20140 19325 20180
rect 18691 20139 18749 20140
rect 16387 20096 16445 20097
rect 19948 20096 19988 20224
rect 21424 20204 21504 20224
rect 15427 20056 15436 20096
rect 15476 20056 16396 20096
rect 16436 20056 16445 20096
rect 16867 20056 16876 20096
rect 16916 20056 17932 20096
rect 17972 20056 17981 20096
rect 18115 20056 18124 20096
rect 18164 20056 18988 20096
rect 19028 20056 19037 20096
rect 19084 20056 19988 20096
rect 16387 20055 16445 20056
rect 15331 20012 15389 20013
rect 4867 19972 4876 20012
rect 4916 19972 5740 20012
rect 5780 19972 8180 20012
rect 0 19928 80 19948
rect 1219 19928 1277 19929
rect 2947 19928 3005 19929
rect 3139 19928 3197 19929
rect 7363 19928 7421 19929
rect 0 19888 1228 19928
rect 1268 19888 1277 19928
rect 2862 19888 2956 19928
rect 2996 19888 3005 19928
rect 3054 19888 3148 19928
rect 3188 19888 3197 19928
rect 4579 19888 4588 19928
rect 4628 19888 6700 19928
rect 6740 19888 6749 19928
rect 6883 19888 6892 19928
rect 6932 19888 7372 19928
rect 7412 19888 7421 19928
rect 8140 19928 8180 19972
rect 8227 19972 8236 20012
rect 8276 19972 8332 20012
rect 8372 19972 8381 20012
rect 13315 19972 13324 20012
rect 13364 19972 13612 20012
rect 13652 19972 13661 20012
rect 13987 19972 13996 20012
rect 14036 19972 15092 20012
rect 15244 19972 15340 20012
rect 15380 19972 15389 20012
rect 8227 19971 8285 19972
rect 10819 19928 10877 19929
rect 8140 19888 10828 19928
rect 10868 19888 10877 19928
rect 15052 19928 15092 19972
rect 15331 19971 15389 19972
rect 15619 20012 15677 20013
rect 19084 20012 19124 20056
rect 15619 19972 15628 20012
rect 15668 19972 15916 20012
rect 15956 19972 15965 20012
rect 18019 19972 18028 20012
rect 18068 19972 19124 20012
rect 19651 20012 19709 20013
rect 19651 19972 19660 20012
rect 19700 19972 19948 20012
rect 19988 19972 19997 20012
rect 15619 19971 15677 19972
rect 19651 19971 19709 19972
rect 21424 19928 21504 19948
rect 15052 19888 16148 19928
rect 20803 19888 20812 19928
rect 20852 19888 21504 19928
rect 0 19868 80 19888
rect 1219 19887 1277 19888
rect 2947 19887 3005 19888
rect 3139 19887 3197 19888
rect 7363 19887 7421 19888
rect 10819 19887 10877 19888
rect 2563 19844 2621 19845
rect 3427 19844 3485 19845
rect 6595 19844 6653 19845
rect 16108 19844 16148 19888
rect 21424 19868 21504 19888
rect 1411 19804 1420 19844
rect 1460 19804 2572 19844
rect 2612 19804 3436 19844
rect 3476 19804 3485 19844
rect 3811 19804 3820 19844
rect 3860 19804 6604 19844
rect 6644 19804 6653 19844
rect 7843 19804 7852 19844
rect 7892 19804 10444 19844
rect 10484 19804 11212 19844
rect 11252 19804 11261 19844
rect 11404 19804 11692 19844
rect 11732 19804 11741 19844
rect 12451 19804 12460 19844
rect 12500 19804 15148 19844
rect 15188 19804 16012 19844
rect 16052 19804 16061 19844
rect 16108 19804 17780 19844
rect 18307 19804 18316 19844
rect 18356 19804 19948 19844
rect 19988 19804 19997 19844
rect 2563 19803 2621 19804
rect 3427 19803 3485 19804
rect 6595 19803 6653 19804
rect 11404 19760 11444 19804
rect 15331 19760 15389 19761
rect 16195 19760 16253 19761
rect 17740 19760 17780 19804
rect 1507 19720 1516 19760
rect 1556 19720 2572 19760
rect 2612 19720 2621 19760
rect 2755 19720 2764 19760
rect 2804 19720 3532 19760
rect 3572 19720 4396 19760
rect 4436 19720 4445 19760
rect 8227 19720 8236 19760
rect 8276 19720 11444 19760
rect 11491 19720 11500 19760
rect 11540 19720 15340 19760
rect 15380 19720 15389 19760
rect 16110 19720 16204 19760
rect 16244 19720 16253 19760
rect 17731 19720 17740 19760
rect 17780 19720 17789 19760
rect 15331 19719 15389 19720
rect 16195 19719 16253 19720
rect 13603 19676 13661 19677
rect 3679 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 4065 19676
rect 9763 19636 9772 19676
rect 9812 19636 10060 19676
rect 10100 19636 10109 19676
rect 10531 19636 10540 19676
rect 10580 19636 12364 19676
rect 12404 19636 13132 19676
rect 13172 19636 13181 19676
rect 13518 19636 13612 19676
rect 13652 19636 13661 19676
rect 13603 19635 13661 19636
rect 14947 19676 15005 19677
rect 14947 19636 14956 19676
rect 14996 19636 18508 19676
rect 18548 19636 18557 19676
rect 18799 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 19185 19676
rect 14947 19635 15005 19636
rect 835 19592 893 19593
rect 10051 19592 10109 19593
rect 20995 19592 21053 19593
rect 21424 19592 21504 19612
rect 835 19552 844 19592
rect 884 19552 7084 19592
rect 7124 19552 7133 19592
rect 9379 19552 9388 19592
rect 9428 19552 10060 19592
rect 10100 19552 10109 19592
rect 11683 19552 11692 19592
rect 11732 19552 16588 19592
rect 16628 19552 17260 19592
rect 17300 19552 17309 19592
rect 17539 19552 17548 19592
rect 17588 19552 19660 19592
rect 19700 19552 19709 19592
rect 20995 19552 21004 19592
rect 21044 19552 21504 19592
rect 835 19551 893 19552
rect 10051 19551 10109 19552
rect 20995 19551 21053 19552
rect 21424 19532 21504 19552
rect 10819 19508 10877 19509
rect 11011 19508 11069 19509
rect 547 19468 556 19508
rect 596 19468 1708 19508
rect 1748 19468 1757 19508
rect 9763 19468 9772 19508
rect 9812 19468 9964 19508
rect 10004 19468 10013 19508
rect 10819 19468 10828 19508
rect 10868 19468 11020 19508
rect 11060 19468 11069 19508
rect 11203 19468 11212 19508
rect 11252 19468 13516 19508
rect 13556 19468 14284 19508
rect 14324 19468 14333 19508
rect 10819 19467 10877 19468
rect 11011 19467 11069 19468
rect 0 19424 80 19444
rect 1315 19424 1373 19425
rect 8227 19424 8285 19425
rect 0 19384 1324 19424
rect 1364 19384 1373 19424
rect 0 19364 80 19384
rect 1315 19383 1373 19384
rect 2500 19384 6124 19424
rect 6164 19384 6173 19424
rect 8227 19384 8236 19424
rect 8276 19384 15092 19424
rect 15139 19384 15148 19424
rect 15188 19384 16300 19424
rect 16340 19384 16349 19424
rect 19459 19384 19468 19424
rect 19508 19384 19660 19424
rect 19700 19384 19709 19424
rect 2500 19340 2540 19384
rect 8227 19383 8285 19384
rect 15052 19340 15092 19384
rect 1315 19300 1324 19340
rect 1364 19300 2540 19340
rect 4771 19300 4780 19340
rect 4820 19300 5740 19340
rect 5780 19300 8044 19340
rect 8084 19300 11596 19340
rect 11636 19300 13996 19340
rect 14036 19300 14045 19340
rect 15052 19300 15436 19340
rect 15476 19300 15485 19340
rect 15715 19300 15724 19340
rect 15764 19300 16972 19340
rect 17012 19300 17452 19340
rect 17492 19300 17501 19340
rect 2851 19256 2909 19257
rect 10723 19256 10781 19257
rect 12835 19256 12893 19257
rect 451 19216 460 19256
rect 500 19216 1516 19256
rect 1556 19216 1565 19256
rect 2766 19216 2860 19256
rect 2900 19216 2909 19256
rect 3523 19216 3532 19256
rect 3572 19216 7124 19256
rect 7363 19216 7372 19256
rect 7412 19216 7564 19256
rect 7604 19216 7613 19256
rect 8611 19216 8620 19256
rect 8660 19216 8812 19256
rect 8852 19216 10732 19256
rect 10772 19216 10781 19256
rect 12750 19216 12844 19256
rect 12884 19216 12893 19256
rect 2851 19215 2909 19216
rect 4387 19172 4445 19173
rect 5347 19172 5405 19173
rect 7084 19172 7124 19216
rect 10723 19215 10781 19216
rect 12835 19215 12893 19216
rect 14179 19256 14237 19257
rect 14947 19256 15005 19257
rect 20515 19256 20573 19257
rect 21424 19256 21504 19276
rect 14179 19216 14188 19256
rect 14228 19216 14572 19256
rect 14612 19216 14621 19256
rect 14862 19216 14956 19256
rect 14996 19216 15005 19256
rect 15811 19216 15820 19256
rect 15860 19216 16876 19256
rect 16916 19216 16925 19256
rect 17539 19216 17548 19256
rect 17588 19216 18220 19256
rect 18260 19216 18269 19256
rect 19171 19216 19180 19256
rect 19220 19216 19468 19256
rect 19508 19216 20236 19256
rect 20276 19216 20524 19256
rect 20564 19216 20573 19256
rect 21283 19216 21292 19256
rect 21332 19216 21504 19256
rect 14179 19215 14237 19216
rect 14947 19215 15005 19216
rect 20515 19215 20573 19216
rect 21424 19196 21504 19216
rect 16675 19172 16733 19173
rect 2563 19132 2572 19172
rect 2612 19132 3628 19172
rect 3668 19132 4396 19172
rect 4436 19132 4445 19172
rect 5251 19132 5260 19172
rect 5300 19132 5356 19172
rect 5396 19132 5405 19172
rect 4387 19131 4445 19132
rect 5347 19131 5405 19132
rect 5740 19132 6988 19172
rect 7028 19132 7037 19172
rect 7084 19132 10251 19172
rect 10291 19132 10300 19172
rect 10435 19132 10444 19172
rect 10484 19132 13324 19172
rect 13364 19132 13373 19172
rect 16590 19132 16684 19172
rect 16724 19132 16733 19172
rect 163 19088 221 19089
rect 5740 19088 5780 19132
rect 6403 19088 6461 19089
rect 12067 19088 12125 19089
rect 163 19048 172 19088
rect 212 19048 3820 19088
rect 3860 19048 4204 19088
rect 4244 19048 4253 19088
rect 5731 19048 5740 19088
rect 5780 19048 5789 19088
rect 6403 19048 6412 19088
rect 6452 19048 12076 19088
rect 12116 19048 12125 19088
rect 13324 19088 13364 19132
rect 16675 19131 16733 19132
rect 19459 19172 19517 19173
rect 19459 19132 19468 19172
rect 19508 19132 19756 19172
rect 19796 19132 19805 19172
rect 19459 19131 19517 19132
rect 18691 19088 18749 19089
rect 13324 19048 14956 19088
rect 14996 19048 15005 19088
rect 17620 19048 18700 19088
rect 18740 19048 18749 19088
rect 163 19047 221 19048
rect 6403 19047 6461 19048
rect 12067 19047 12125 19048
rect 2083 19004 2141 19005
rect 11875 19004 11933 19005
rect 1795 18964 1804 19004
rect 1844 18964 2092 19004
rect 2132 18964 2141 19004
rect 2083 18963 2141 18964
rect 2500 18964 11884 19004
rect 11924 18964 11933 19004
rect 0 18920 80 18940
rect 2500 18920 2540 18964
rect 11875 18963 11933 18964
rect 12163 19004 12221 19005
rect 16867 19004 16925 19005
rect 17620 19004 17660 19048
rect 18691 19047 18749 19048
rect 19276 19048 19852 19088
rect 19892 19048 19901 19088
rect 20131 19048 20140 19088
rect 20180 19048 20189 19088
rect 19276 19004 19316 19048
rect 20140 19004 20180 19048
rect 12163 18964 12172 19004
rect 12212 18964 14764 19004
rect 14804 18964 14813 19004
rect 16867 18964 16876 19004
rect 16916 18964 17660 19004
rect 18604 18964 19316 19004
rect 19363 18964 19372 19004
rect 19412 18964 19756 19004
rect 19796 18964 19805 19004
rect 19948 18964 20180 19004
rect 12163 18963 12221 18964
rect 16867 18963 16925 18964
rect 0 18880 2540 18920
rect 3139 18920 3197 18921
rect 4387 18920 4445 18921
rect 6115 18920 6173 18921
rect 11491 18920 11549 18921
rect 13891 18920 13949 18921
rect 14083 18920 14141 18921
rect 17155 18920 17213 18921
rect 18604 18920 18644 18964
rect 19948 18920 19988 18964
rect 21424 18920 21504 18940
rect 3139 18880 3148 18920
rect 3188 18880 3340 18920
rect 3380 18880 3389 18920
rect 4302 18880 4396 18920
rect 4436 18880 4445 18920
rect 4919 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 5305 18920
rect 6030 18880 6124 18920
rect 6164 18880 6173 18920
rect 9187 18880 9196 18920
rect 9236 18880 9868 18920
rect 9908 18880 9917 18920
rect 11491 18880 11500 18920
rect 11540 18880 12268 18920
rect 12308 18880 12317 18920
rect 13891 18880 13900 18920
rect 13940 18880 14092 18920
rect 14132 18880 14141 18920
rect 15523 18880 15532 18920
rect 15572 18880 16396 18920
rect 16436 18880 16445 18920
rect 17155 18880 17164 18920
rect 17204 18880 18644 18920
rect 18691 18880 18700 18920
rect 18740 18880 19564 18920
rect 19604 18880 19613 18920
rect 19939 18880 19948 18920
rect 19988 18880 19997 18920
rect 20039 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20425 18920
rect 20899 18880 20908 18920
rect 20948 18880 21504 18920
rect 0 18860 80 18880
rect 3139 18879 3197 18880
rect 4387 18879 4445 18880
rect 6115 18879 6173 18880
rect 11491 18879 11549 18880
rect 13891 18879 13949 18880
rect 14083 18879 14141 18880
rect 17155 18879 17213 18880
rect 21424 18860 21504 18880
rect 6403 18836 6461 18837
rect 1603 18796 1612 18836
rect 1652 18796 6412 18836
rect 6452 18796 6461 18836
rect 6403 18795 6461 18796
rect 9955 18836 10013 18837
rect 16387 18836 16445 18837
rect 9955 18796 9964 18836
rect 10004 18796 10444 18836
rect 10484 18796 10493 18836
rect 12739 18796 12748 18836
rect 12788 18796 13324 18836
rect 13364 18796 13373 18836
rect 13987 18796 13996 18836
rect 14036 18796 15052 18836
rect 15092 18796 15101 18836
rect 16387 18796 16396 18836
rect 16436 18796 16588 18836
rect 16628 18796 16637 18836
rect 17155 18796 17164 18836
rect 17204 18796 17452 18836
rect 17492 18796 17501 18836
rect 19267 18796 19276 18836
rect 19316 18796 20372 18836
rect 9955 18795 10013 18796
rect 16387 18795 16445 18796
rect 5635 18752 5693 18753
rect 14371 18752 14429 18753
rect 20332 18752 20372 18796
rect 2947 18712 2956 18752
rect 2996 18712 5204 18752
rect 5539 18712 5548 18752
rect 5588 18712 5644 18752
rect 5684 18712 5693 18752
rect 6979 18712 6988 18752
rect 7028 18712 8908 18752
rect 8948 18712 8957 18752
rect 12163 18712 12172 18752
rect 12212 18712 13228 18752
rect 13268 18712 14380 18752
rect 14420 18712 14429 18752
rect 16291 18712 16300 18752
rect 16340 18712 16349 18752
rect 18595 18712 18604 18752
rect 18644 18712 19180 18752
rect 19220 18712 19372 18752
rect 19412 18712 19421 18752
rect 19843 18712 19852 18752
rect 19892 18712 20180 18752
rect 20323 18712 20332 18752
rect 20372 18712 20381 18752
rect 5164 18668 5204 18712
rect 5635 18711 5693 18712
rect 14371 18711 14429 18712
rect 10147 18668 10205 18669
rect 4387 18628 4396 18668
rect 4436 18628 5068 18668
rect 5108 18628 5117 18668
rect 5164 18628 10156 18668
rect 10196 18628 10205 18668
rect 10147 18627 10205 18628
rect 12451 18584 12509 18585
rect 451 18544 460 18584
rect 500 18544 2764 18584
rect 2804 18544 7084 18584
rect 7124 18544 7133 18584
rect 7555 18544 7564 18584
rect 7604 18544 8044 18584
rect 8084 18544 8524 18584
rect 8564 18544 8573 18584
rect 9283 18544 9292 18584
rect 9332 18544 10924 18584
rect 10964 18544 10973 18584
rect 11779 18544 11788 18584
rect 11828 18544 12460 18584
rect 12500 18544 12509 18584
rect 12451 18543 12509 18544
rect 12643 18584 12701 18585
rect 16300 18584 16340 18712
rect 16483 18668 16541 18669
rect 20140 18668 20180 18712
rect 20995 18668 21053 18669
rect 16483 18628 16492 18668
rect 16532 18628 17068 18668
rect 17108 18628 17117 18668
rect 17827 18628 17836 18668
rect 17876 18628 18412 18668
rect 18452 18628 18461 18668
rect 20140 18628 21004 18668
rect 21044 18628 21053 18668
rect 16483 18627 16541 18628
rect 20995 18627 21053 18628
rect 17155 18584 17213 18585
rect 18499 18584 18557 18585
rect 19459 18584 19517 18585
rect 21424 18584 21504 18604
rect 12643 18544 12652 18584
rect 12692 18544 14284 18584
rect 14324 18544 14333 18584
rect 14659 18544 14668 18584
rect 14708 18544 16204 18584
rect 16244 18544 16253 18584
rect 16300 18544 16780 18584
rect 16820 18544 16829 18584
rect 17070 18544 17164 18584
rect 17204 18544 17213 18584
rect 12643 18543 12701 18544
rect 12259 18500 12317 18501
rect 1795 18460 1804 18500
rect 1844 18460 2284 18500
rect 2324 18460 2333 18500
rect 2851 18460 2860 18500
rect 2900 18460 3148 18500
rect 3188 18460 3532 18500
rect 3572 18460 3581 18500
rect 3628 18460 12268 18500
rect 12308 18460 13612 18500
rect 13652 18460 13661 18500
rect 14947 18460 14956 18500
rect 14996 18460 16628 18500
rect 0 18416 80 18436
rect 1219 18416 1277 18417
rect 3628 18416 3668 18460
rect 12259 18459 12317 18460
rect 0 18376 1228 18416
rect 1268 18376 1277 18416
rect 1507 18376 1516 18416
rect 1556 18376 2956 18416
rect 2996 18376 3005 18416
rect 3235 18376 3244 18416
rect 3284 18376 3668 18416
rect 5731 18416 5789 18417
rect 13411 18416 13469 18417
rect 5731 18376 5740 18416
rect 5780 18376 6796 18416
rect 6836 18376 7372 18416
rect 7412 18376 7421 18416
rect 11395 18376 11404 18416
rect 11444 18376 13420 18416
rect 13460 18376 13469 18416
rect 16099 18376 16108 18416
rect 16148 18376 16492 18416
rect 16532 18376 16541 18416
rect 0 18356 80 18376
rect 1219 18375 1277 18376
rect 5731 18375 5789 18376
rect 13411 18375 13469 18376
rect 1699 18332 1757 18333
rect 4771 18332 4829 18333
rect 1699 18292 1708 18332
rect 1748 18292 3436 18332
rect 3476 18292 3724 18332
rect 3764 18292 3773 18332
rect 4686 18292 4780 18332
rect 4820 18292 4829 18332
rect 1699 18291 1757 18292
rect 4771 18291 4829 18292
rect 11683 18332 11741 18333
rect 14947 18332 15005 18333
rect 11683 18292 11692 18332
rect 11732 18292 13612 18332
rect 13652 18292 13661 18332
rect 14947 18292 14956 18332
rect 14996 18292 15052 18332
rect 15092 18292 15101 18332
rect 11683 18291 11741 18292
rect 14947 18291 15005 18292
rect 16492 18248 16532 18376
rect 16588 18332 16628 18460
rect 16780 18416 16820 18544
rect 17155 18543 17213 18544
rect 17260 18544 18508 18584
rect 18548 18544 19468 18584
rect 19508 18544 19517 18584
rect 19651 18544 19660 18584
rect 19700 18544 20620 18584
rect 20660 18544 20669 18584
rect 20812 18544 21504 18584
rect 17260 18500 17300 18544
rect 18499 18543 18557 18544
rect 19459 18543 19517 18544
rect 20812 18500 20852 18544
rect 21424 18524 21504 18544
rect 17059 18460 17068 18500
rect 17108 18460 17300 18500
rect 17347 18460 17356 18500
rect 17396 18460 20852 18500
rect 20611 18416 20669 18417
rect 16780 18376 17164 18416
rect 17204 18376 17213 18416
rect 18211 18376 18220 18416
rect 18260 18376 20620 18416
rect 20660 18376 20669 18416
rect 20611 18375 20669 18376
rect 19363 18332 19421 18333
rect 16588 18292 17932 18332
rect 17972 18292 17981 18332
rect 19363 18292 19372 18332
rect 19412 18292 19468 18332
rect 19508 18292 19517 18332
rect 19747 18292 19756 18332
rect 19796 18292 20236 18332
rect 20276 18292 20285 18332
rect 19363 18291 19421 18292
rect 21187 18248 21245 18249
rect 21424 18248 21504 18268
rect 1123 18208 1132 18248
rect 1172 18208 12460 18248
rect 12500 18208 12509 18248
rect 12643 18208 12652 18248
rect 12692 18208 13036 18248
rect 13076 18208 13085 18248
rect 13219 18208 13228 18248
rect 13268 18208 14476 18248
rect 14516 18208 14525 18248
rect 16492 18208 17452 18248
rect 17492 18208 17501 18248
rect 21187 18208 21196 18248
rect 21236 18208 21504 18248
rect 21187 18207 21245 18208
rect 21424 18188 21504 18208
rect 11587 18164 11645 18165
rect 3679 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 4065 18164
rect 4108 18124 4340 18164
rect 7747 18124 7756 18164
rect 7796 18124 7948 18164
rect 7988 18124 7997 18164
rect 11587 18124 11596 18164
rect 11636 18124 11788 18164
rect 11828 18124 11837 18164
rect 12547 18124 12556 18164
rect 12596 18124 13132 18164
rect 13172 18124 13181 18164
rect 13411 18124 13420 18164
rect 13460 18124 13708 18164
rect 13748 18124 17740 18164
rect 17780 18124 17789 18164
rect 18799 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 19185 18164
rect 835 18080 893 18081
rect 4108 18080 4148 18124
rect 835 18040 844 18080
rect 884 18040 4148 18080
rect 4195 18040 4204 18080
rect 4244 18040 4253 18080
rect 835 18039 893 18040
rect 4204 17996 4244 18040
rect 2659 17956 2668 17996
rect 2708 17956 4244 17996
rect 4300 17996 4340 18124
rect 11587 18123 11645 18124
rect 4387 18080 4445 18081
rect 19651 18080 19709 18081
rect 4387 18040 4396 18080
rect 4436 18040 4684 18080
rect 4724 18040 4733 18080
rect 5347 18040 5356 18080
rect 5396 18040 18124 18080
rect 18164 18040 18173 18080
rect 19180 18040 19660 18080
rect 19700 18040 20140 18080
rect 20180 18040 20189 18080
rect 4387 18039 4445 18040
rect 16387 17996 16445 17997
rect 19180 17996 19220 18040
rect 19651 18039 19709 18040
rect 19939 17996 19997 17997
rect 4300 17956 6316 17996
rect 6356 17956 6796 17996
rect 6836 17956 6845 17996
rect 11683 17956 11692 17996
rect 11732 17956 13420 17996
rect 13460 17956 13996 17996
rect 14036 17956 14045 17996
rect 14188 17956 14764 17996
rect 14804 17956 14813 17996
rect 16291 17956 16300 17996
rect 16340 17956 16396 17996
rect 16436 17956 17012 17996
rect 19171 17956 19180 17996
rect 19220 17956 19229 17996
rect 19854 17956 19948 17996
rect 19988 17956 19997 17996
rect 0 17912 80 17932
rect 547 17912 605 17913
rect 0 17872 556 17912
rect 596 17872 605 17912
rect 0 17852 80 17872
rect 547 17871 605 17872
rect 1315 17912 1373 17913
rect 1315 17872 1324 17912
rect 1364 17872 13228 17912
rect 13268 17872 13277 17912
rect 1315 17871 1373 17872
rect 2467 17828 2525 17829
rect 4099 17828 4157 17829
rect 5443 17828 5501 17829
rect 14188 17828 14228 17956
rect 16387 17955 16445 17956
rect 14371 17912 14429 17913
rect 16972 17912 17012 17956
rect 19939 17955 19997 17956
rect 19555 17912 19613 17913
rect 21424 17912 21504 17932
rect 14286 17872 14380 17912
rect 14420 17872 14429 17912
rect 16963 17872 16972 17912
rect 17012 17872 17021 17912
rect 19555 17872 19564 17912
rect 19604 17872 21504 17912
rect 14371 17871 14429 17872
rect 19555 17871 19613 17872
rect 21424 17852 21504 17872
rect 17635 17828 17693 17829
rect 19747 17828 19805 17829
rect 2382 17788 2476 17828
rect 2516 17788 4052 17828
rect 2467 17787 2525 17788
rect 1795 17744 1853 17745
rect 1710 17704 1804 17744
rect 1844 17704 1853 17744
rect 1795 17703 1853 17704
rect 2371 17744 2429 17745
rect 2659 17744 2717 17745
rect 4012 17744 4052 17788
rect 4099 17788 4108 17828
rect 4148 17788 4396 17828
rect 4436 17788 4445 17828
rect 4579 17788 4588 17828
rect 4628 17788 5452 17828
rect 5492 17788 5501 17828
rect 8131 17788 8140 17828
rect 8180 17788 10924 17828
rect 10964 17788 10973 17828
rect 11587 17788 11596 17828
rect 11636 17788 14228 17828
rect 14563 17788 14572 17828
rect 14612 17788 16340 17828
rect 4099 17787 4157 17788
rect 5443 17787 5501 17788
rect 4483 17744 4541 17745
rect 4771 17744 4829 17745
rect 8995 17744 9053 17745
rect 9187 17744 9245 17745
rect 9571 17744 9629 17745
rect 14179 17744 14237 17745
rect 14947 17744 15005 17745
rect 16300 17744 16340 17788
rect 17635 17788 17644 17828
rect 17684 17788 19372 17828
rect 19412 17788 19421 17828
rect 19662 17788 19756 17828
rect 19796 17788 19805 17828
rect 17635 17787 17693 17788
rect 19747 17787 19805 17788
rect 2371 17704 2380 17744
rect 2420 17704 2668 17744
rect 2708 17704 2860 17744
rect 2900 17704 2909 17744
rect 4012 17704 4108 17744
rect 4148 17704 4300 17744
rect 4340 17704 4349 17744
rect 4398 17704 4492 17744
rect 4532 17704 4780 17744
rect 4820 17704 4829 17744
rect 7171 17704 7180 17744
rect 7220 17704 9004 17744
rect 9044 17704 9053 17744
rect 9102 17704 9196 17744
rect 9236 17704 9245 17744
rect 9486 17704 9580 17744
rect 9620 17704 9629 17744
rect 10819 17704 10828 17744
rect 10868 17704 14188 17744
rect 14228 17704 14420 17744
rect 2371 17703 2429 17704
rect 2659 17703 2717 17704
rect 4483 17703 4541 17704
rect 4771 17703 4829 17704
rect 8995 17703 9053 17704
rect 9187 17703 9245 17704
rect 9571 17703 9629 17704
rect 14179 17703 14237 17704
rect 547 17660 605 17661
rect 835 17660 893 17661
rect 9955 17660 10013 17661
rect 547 17620 556 17660
rect 596 17620 844 17660
rect 884 17620 893 17660
rect 1603 17620 1612 17660
rect 1652 17620 2284 17660
rect 2324 17620 2333 17660
rect 5923 17620 5932 17660
rect 5972 17620 7756 17660
rect 7796 17620 7805 17660
rect 7939 17620 7948 17660
rect 7988 17620 8564 17660
rect 8707 17620 8716 17660
rect 8756 17620 9964 17660
rect 10004 17620 10013 17660
rect 547 17619 605 17620
rect 835 17619 893 17620
rect 2755 17576 2813 17577
rect 8524 17576 8564 17620
rect 9955 17619 10013 17620
rect 10147 17660 10205 17661
rect 10339 17660 10397 17661
rect 13699 17660 13757 17661
rect 13891 17660 13949 17661
rect 10147 17620 10156 17660
rect 10196 17620 10348 17660
rect 10388 17620 10397 17660
rect 11491 17620 11500 17660
rect 11540 17620 12844 17660
rect 12884 17620 13036 17660
rect 13076 17620 13085 17660
rect 13315 17620 13324 17660
rect 13364 17620 13556 17660
rect 13614 17620 13708 17660
rect 13748 17620 13757 17660
rect 10147 17619 10205 17620
rect 10339 17619 10397 17620
rect 13516 17576 13556 17620
rect 13699 17619 13757 17620
rect 13804 17620 13900 17660
rect 13940 17620 13949 17660
rect 14380 17660 14420 17704
rect 14947 17704 14956 17744
rect 14996 17704 15244 17744
rect 15284 17704 15572 17744
rect 16291 17704 16300 17744
rect 16340 17704 16349 17744
rect 16772 17704 16781 17744
rect 16821 17704 20332 17744
rect 20372 17704 21004 17744
rect 21044 17704 21053 17744
rect 14947 17703 15005 17704
rect 14380 17620 14476 17660
rect 14516 17620 14525 17660
rect 13804 17576 13844 17620
rect 13891 17619 13949 17620
rect 931 17536 940 17576
rect 980 17536 2764 17576
rect 2804 17536 2813 17576
rect 8515 17536 8524 17576
rect 8564 17536 8573 17576
rect 9091 17536 9100 17576
rect 9140 17536 9484 17576
rect 9524 17536 9533 17576
rect 10819 17536 10828 17576
rect 10868 17536 11020 17576
rect 11060 17536 11069 17576
rect 13516 17536 13844 17576
rect 15532 17576 15572 17704
rect 16867 17660 16925 17661
rect 19843 17660 19901 17661
rect 15619 17620 15628 17660
rect 15668 17620 16820 17660
rect 15532 17536 16108 17576
rect 16148 17536 16157 17576
rect 2755 17535 2813 17536
rect 4579 17492 4637 17493
rect 6979 17492 7037 17493
rect 13603 17492 13661 17493
rect 2092 17452 2956 17492
rect 2996 17452 4588 17492
rect 4628 17452 4637 17492
rect 5731 17452 5740 17492
rect 5780 17452 6988 17492
rect 7028 17452 7037 17492
rect 7939 17452 7948 17492
rect 7988 17452 8620 17492
rect 8660 17452 8669 17492
rect 13518 17452 13612 17492
rect 13652 17452 13661 17492
rect 0 17408 80 17428
rect 2092 17408 2132 17452
rect 4579 17451 4637 17452
rect 6979 17451 7037 17452
rect 13603 17451 13661 17452
rect 14083 17492 14141 17493
rect 16780 17492 16820 17620
rect 16867 17620 16876 17660
rect 16916 17620 17010 17660
rect 19843 17620 19852 17660
rect 19892 17620 19948 17660
rect 19988 17620 19997 17660
rect 16867 17619 16925 17620
rect 19843 17619 19901 17620
rect 20611 17576 20669 17577
rect 21424 17576 21504 17596
rect 20611 17536 20620 17576
rect 20660 17536 21504 17576
rect 20611 17535 20669 17536
rect 21424 17516 21504 17536
rect 14083 17452 14092 17492
rect 14132 17452 14860 17492
rect 14900 17452 14909 17492
rect 16771 17452 16780 17492
rect 16820 17452 16829 17492
rect 14083 17451 14141 17452
rect 6883 17408 6941 17409
rect 9187 17408 9245 17409
rect 0 17368 76 17408
rect 116 17368 125 17408
rect 460 17368 2132 17408
rect 2179 17368 2188 17408
rect 2228 17368 2860 17408
rect 2900 17368 2909 17408
rect 4919 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 5305 17408
rect 6019 17368 6028 17408
rect 6068 17368 6892 17408
rect 6932 17368 6941 17408
rect 8995 17368 9004 17408
rect 9044 17368 9196 17408
rect 9236 17368 9245 17408
rect 12451 17368 12460 17408
rect 12500 17368 19180 17408
rect 19220 17368 19229 17408
rect 20039 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20425 17408
rect 0 17348 80 17368
rect 460 17324 500 17368
rect 6883 17367 6941 17368
rect 9187 17367 9245 17368
rect 163 17284 172 17324
rect 212 17284 500 17324
rect 1027 17324 1085 17325
rect 5635 17324 5693 17325
rect 6403 17324 6461 17325
rect 1027 17284 1036 17324
rect 1076 17284 2092 17324
rect 2132 17284 2141 17324
rect 2275 17284 2284 17324
rect 2324 17284 5644 17324
rect 5684 17284 6412 17324
rect 6452 17284 6461 17324
rect 6883 17284 6892 17324
rect 6932 17284 15052 17324
rect 15092 17284 15101 17324
rect 16396 17284 18604 17324
rect 18644 17284 18988 17324
rect 19028 17284 19037 17324
rect 1027 17283 1085 17284
rect 5635 17283 5693 17284
rect 6403 17283 6461 17284
rect 2275 17240 2333 17241
rect 5731 17240 5789 17241
rect 16396 17240 16436 17284
rect 17443 17240 17501 17241
rect 21424 17240 21504 17260
rect 1987 17200 1996 17240
rect 2036 17200 2284 17240
rect 2324 17200 2333 17240
rect 5539 17200 5548 17240
rect 5588 17200 5740 17240
rect 5780 17200 5789 17240
rect 2275 17199 2333 17200
rect 5731 17199 5789 17200
rect 6316 17200 9964 17240
rect 10004 17200 10013 17240
rect 12643 17200 12652 17240
rect 12692 17200 16436 17240
rect 16483 17200 16492 17240
rect 16532 17200 16684 17240
rect 16724 17200 16733 17240
rect 17347 17200 17356 17240
rect 17396 17200 17452 17240
rect 17492 17200 17501 17240
rect 20707 17200 20716 17240
rect 20756 17200 21504 17240
rect 4099 17156 4157 17157
rect 1411 17116 1420 17156
rect 1460 17116 3860 17156
rect 3907 17116 3916 17156
rect 3956 17116 4108 17156
rect 4148 17116 4157 17156
rect 1315 17072 1373 17073
rect 3820 17072 3860 17116
rect 4099 17115 4157 17116
rect 5539 17156 5597 17157
rect 6316 17156 6356 17200
rect 17443 17199 17501 17200
rect 21424 17180 21504 17200
rect 15907 17156 15965 17157
rect 5539 17116 5548 17156
rect 5588 17116 6316 17156
rect 6356 17116 6365 17156
rect 6691 17116 6700 17156
rect 6740 17116 8276 17156
rect 8707 17116 8716 17156
rect 8756 17116 9580 17156
rect 9620 17116 9629 17156
rect 9763 17116 9772 17156
rect 9812 17116 10732 17156
rect 10772 17116 10781 17156
rect 13891 17116 13900 17156
rect 13940 17116 15724 17156
rect 15764 17116 15773 17156
rect 15907 17116 15916 17156
rect 15956 17116 17740 17156
rect 17780 17116 17789 17156
rect 18787 17116 18796 17156
rect 18836 17116 20127 17156
rect 20167 17116 20176 17156
rect 5539 17115 5597 17116
rect 6403 17072 6461 17073
rect 8236 17072 8276 17116
rect 15907 17115 15965 17116
rect 1230 17032 1324 17072
rect 1364 17032 1373 17072
rect 1603 17032 1612 17072
rect 1652 17032 2188 17072
rect 2228 17032 2237 17072
rect 3820 17032 6124 17072
rect 6164 17032 6173 17072
rect 6403 17032 6412 17072
rect 6452 17032 7220 17072
rect 8227 17032 8236 17072
rect 8276 17032 8285 17072
rect 8995 17032 9004 17072
rect 9044 17032 10924 17072
rect 10964 17032 10973 17072
rect 15811 17032 15820 17072
rect 15860 17032 19948 17072
rect 19988 17032 19997 17072
rect 1315 17031 1373 17032
rect 6403 17031 6461 17032
rect 7180 16988 7220 17032
rect 16963 16988 17021 16989
rect 739 16948 748 16988
rect 788 16948 2092 16988
rect 2132 16948 3436 16988
rect 3476 16948 5876 16988
rect 6691 16948 6700 16988
rect 6740 16948 7084 16988
rect 7124 16948 7133 16988
rect 7180 16948 11360 16988
rect 12547 16948 12556 16988
rect 12596 16948 14476 16988
rect 14516 16948 14525 16988
rect 16963 16948 16972 16988
rect 17012 16948 17356 16988
rect 17396 16948 17405 16988
rect 19651 16948 19660 16988
rect 19700 16948 20236 16988
rect 20276 16948 20285 16988
rect 0 16904 80 16924
rect 1219 16904 1277 16905
rect 5836 16904 5876 16948
rect 11320 16904 11360 16948
rect 16963 16947 17021 16948
rect 13891 16904 13949 16905
rect 21424 16904 21504 16924
rect 0 16864 1228 16904
rect 1268 16864 1277 16904
rect 2851 16864 2860 16904
rect 2900 16864 5740 16904
rect 5780 16864 5789 16904
rect 5836 16864 9292 16904
rect 9332 16864 9341 16904
rect 11320 16864 11404 16904
rect 11444 16864 11453 16904
rect 13806 16864 13900 16904
rect 13940 16864 13949 16904
rect 14083 16864 14092 16904
rect 14132 16864 16396 16904
rect 16436 16864 16445 16904
rect 19075 16864 19084 16904
rect 19124 16864 19756 16904
rect 19796 16864 19805 16904
rect 20140 16864 21504 16904
rect 0 16844 80 16864
rect 1219 16863 1277 16864
rect 13891 16863 13949 16864
rect 1123 16820 1181 16821
rect 16003 16820 16061 16821
rect 1123 16780 1132 16820
rect 1172 16780 3340 16820
rect 3380 16780 6796 16820
rect 6836 16780 6845 16820
rect 8227 16780 8236 16820
rect 8276 16780 11308 16820
rect 11348 16780 12364 16820
rect 12404 16780 16012 16820
rect 16052 16780 16061 16820
rect 18979 16780 18988 16820
rect 19028 16780 19948 16820
rect 19988 16780 19997 16820
rect 1123 16779 1181 16780
rect 16003 16779 16061 16780
rect 4387 16736 4445 16737
rect 20140 16736 20180 16864
rect 21424 16844 21504 16864
rect 1891 16696 1900 16736
rect 1940 16696 4396 16736
rect 4436 16696 4445 16736
rect 8899 16696 8908 16736
rect 8948 16696 12940 16736
rect 12980 16696 12989 16736
rect 18307 16696 18316 16736
rect 18356 16696 20180 16736
rect 4387 16695 4445 16696
rect 12835 16652 12893 16653
rect 14179 16652 14237 16653
rect 15331 16652 15389 16653
rect 67 16612 76 16652
rect 116 16612 3572 16652
rect 3679 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 4065 16652
rect 6499 16612 6508 16652
rect 6548 16612 7372 16652
rect 7412 16612 7421 16652
rect 9379 16612 9388 16652
rect 9428 16612 9437 16652
rect 12750 16612 12844 16652
rect 12884 16612 12893 16652
rect 13699 16612 13708 16652
rect 13748 16612 14188 16652
rect 14228 16612 14284 16652
rect 14324 16612 14352 16652
rect 15246 16612 15340 16652
rect 15380 16612 15389 16652
rect 18799 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 19185 16652
rect 1795 16568 1853 16569
rect 1699 16528 1708 16568
rect 1748 16528 1804 16568
rect 1844 16528 1853 16568
rect 1987 16528 1996 16568
rect 2036 16528 3148 16568
rect 3188 16528 3197 16568
rect 1795 16527 1853 16528
rect 1315 16484 1373 16485
rect 3532 16484 3572 16612
rect 4291 16568 4349 16569
rect 9388 16568 9428 16612
rect 12835 16611 12893 16612
rect 14179 16611 14237 16612
rect 15331 16611 15389 16612
rect 17635 16568 17693 16569
rect 21424 16568 21504 16588
rect 4206 16528 4300 16568
rect 4340 16528 4349 16568
rect 6595 16528 6604 16568
rect 6644 16528 8428 16568
rect 8468 16528 8477 16568
rect 9388 16528 17644 16568
rect 17684 16528 17693 16568
rect 19459 16528 19468 16568
rect 19508 16528 21504 16568
rect 4291 16527 4349 16528
rect 17635 16527 17693 16528
rect 21424 16508 21504 16528
rect 1230 16444 1324 16484
rect 1364 16444 1373 16484
rect 2851 16444 2860 16484
rect 2900 16444 3244 16484
rect 3284 16444 3293 16484
rect 3532 16444 15628 16484
rect 15668 16444 15677 16484
rect 19651 16444 19660 16484
rect 19700 16444 19709 16484
rect 1315 16443 1373 16444
rect 0 16400 80 16420
rect 931 16400 989 16401
rect 4099 16400 4157 16401
rect 0 16360 940 16400
rect 980 16360 989 16400
rect 1507 16360 1516 16400
rect 1556 16360 2092 16400
rect 2132 16360 2141 16400
rect 3811 16360 3820 16400
rect 3860 16360 4108 16400
rect 4148 16360 4157 16400
rect 0 16340 80 16360
rect 931 16359 989 16360
rect 4099 16359 4157 16360
rect 4483 16400 4541 16401
rect 6403 16400 6461 16401
rect 8707 16400 8765 16401
rect 11491 16400 11549 16401
rect 4483 16360 4492 16400
rect 4532 16360 5836 16400
rect 5876 16360 5885 16400
rect 6318 16360 6412 16400
rect 6452 16360 6461 16400
rect 7651 16360 7660 16400
rect 7700 16360 8716 16400
rect 8756 16360 8765 16400
rect 9091 16360 9100 16400
rect 9140 16360 11020 16400
rect 11060 16360 11069 16400
rect 11406 16360 11500 16400
rect 11540 16360 11549 16400
rect 4483 16359 4541 16360
rect 6403 16359 6461 16360
rect 8707 16359 8765 16360
rect 11491 16359 11549 16360
rect 12547 16400 12605 16401
rect 19555 16400 19613 16401
rect 12547 16360 12556 16400
rect 12596 16360 16876 16400
rect 16916 16360 16925 16400
rect 17251 16360 17260 16400
rect 17300 16360 19564 16400
rect 19604 16360 19613 16400
rect 12547 16359 12605 16360
rect 19555 16359 19613 16360
rect 1507 16316 1565 16317
rect 3427 16316 3485 16317
rect 19660 16316 19700 16444
rect 1507 16276 1516 16316
rect 1556 16276 2380 16316
rect 2420 16276 3052 16316
rect 3092 16276 3101 16316
rect 3427 16276 3436 16316
rect 3476 16276 3532 16316
rect 3572 16276 3581 16316
rect 7171 16276 7180 16316
rect 7220 16276 9676 16316
rect 9716 16276 9725 16316
rect 11395 16276 11404 16316
rect 11444 16276 15148 16316
rect 15188 16276 15820 16316
rect 15860 16276 15869 16316
rect 19564 16276 19700 16316
rect 1507 16275 1565 16276
rect 3427 16275 3485 16276
rect 13315 16232 13373 16233
rect 13891 16232 13949 16233
rect 14947 16232 15005 16233
rect 16579 16232 16637 16233
rect 19564 16232 19604 16276
rect 21424 16232 21504 16252
rect 1315 16192 1324 16232
rect 1364 16192 1373 16232
rect 1699 16192 1708 16232
rect 1748 16192 4300 16232
rect 4340 16192 4349 16232
rect 4579 16192 4588 16232
rect 4628 16192 4637 16232
rect 5539 16192 5548 16232
rect 5588 16192 5836 16232
rect 5876 16192 5885 16232
rect 6019 16192 6028 16232
rect 6068 16192 6311 16232
rect 6351 16192 6360 16232
rect 6403 16192 6412 16232
rect 6452 16192 8140 16232
rect 8180 16192 8189 16232
rect 9091 16192 9100 16232
rect 9140 16192 9964 16232
rect 10004 16192 10252 16232
rect 10292 16192 10301 16232
rect 13315 16192 13324 16232
rect 13364 16192 13516 16232
rect 13556 16192 13565 16232
rect 13891 16192 13900 16232
rect 13940 16192 14764 16232
rect 14804 16192 14813 16232
rect 14947 16192 14956 16232
rect 14996 16192 16300 16232
rect 16340 16192 16588 16232
rect 16628 16192 18508 16232
rect 18548 16192 18557 16232
rect 19555 16192 19564 16232
rect 19604 16192 19613 16232
rect 20812 16192 21504 16232
rect 1324 16148 1364 16192
rect 4588 16148 4628 16192
rect 13315 16191 13373 16192
rect 13891 16191 13949 16192
rect 14947 16191 15005 16192
rect 16579 16191 16637 16192
rect 15619 16148 15677 16149
rect 1324 16108 1900 16148
rect 1940 16108 3532 16148
rect 3572 16108 3581 16148
rect 4195 16108 4204 16148
rect 4244 16108 4253 16148
rect 4588 16108 6892 16148
rect 6932 16108 6941 16148
rect 12259 16108 12268 16148
rect 12308 16108 15628 16148
rect 15668 16108 15677 16148
rect 4204 16064 4244 16108
rect 15619 16107 15677 16108
rect 9571 16064 9629 16065
rect 1507 16024 1516 16064
rect 1556 16024 3052 16064
rect 3092 16024 4244 16064
rect 7075 16024 7084 16064
rect 7124 16024 9580 16064
rect 9620 16024 9629 16064
rect 9763 16024 9772 16064
rect 9812 16024 13996 16064
rect 14036 16024 14045 16064
rect 14947 16024 14956 16064
rect 14996 16024 15724 16064
rect 15764 16024 16780 16064
rect 16820 16024 16829 16064
rect 18499 16024 18508 16064
rect 18548 16024 20236 16064
rect 20276 16024 20285 16064
rect 9571 16023 9629 16024
rect 20812 15980 20852 16192
rect 21424 16172 21504 16192
rect 1123 15940 1132 15980
rect 1172 15940 3340 15980
rect 3380 15940 7276 15980
rect 7316 15940 9964 15980
rect 10004 15940 10013 15980
rect 10060 15940 10636 15980
rect 10676 15940 10685 15980
rect 15235 15940 15244 15980
rect 15284 15940 15916 15980
rect 15956 15940 17260 15980
rect 17300 15940 17309 15980
rect 17620 15940 20852 15980
rect 0 15896 80 15916
rect 10060 15896 10100 15940
rect 10531 15896 10589 15897
rect 13411 15896 13469 15897
rect 0 15856 2540 15896
rect 4919 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 5305 15896
rect 9667 15856 9676 15896
rect 9716 15856 10100 15896
rect 10147 15856 10156 15896
rect 10196 15856 10540 15896
rect 10580 15856 10589 15896
rect 11491 15856 11500 15896
rect 11540 15856 11788 15896
rect 11828 15856 13420 15896
rect 13460 15856 13469 15896
rect 0 15836 80 15856
rect 835 15812 893 15813
rect 643 15772 652 15812
rect 692 15772 844 15812
rect 884 15772 893 15812
rect 2500 15812 2540 15856
rect 10531 15855 10589 15856
rect 13411 15855 13469 15856
rect 14563 15896 14621 15897
rect 16003 15896 16061 15897
rect 17620 15896 17660 15940
rect 20707 15896 20765 15897
rect 21424 15896 21504 15916
rect 14563 15856 14572 15896
rect 14612 15856 16012 15896
rect 16052 15856 16061 15896
rect 16867 15856 16876 15896
rect 16916 15856 17660 15896
rect 19363 15856 19372 15896
rect 19412 15856 19948 15896
rect 19988 15856 19997 15896
rect 20039 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20425 15896
rect 20707 15856 20716 15896
rect 20756 15856 21504 15896
rect 14563 15855 14621 15856
rect 16003 15855 16061 15856
rect 20707 15855 20765 15856
rect 21424 15836 21504 15856
rect 12547 15812 12605 15813
rect 17347 15812 17405 15813
rect 2500 15772 12556 15812
rect 12596 15772 12605 15812
rect 13411 15772 13420 15812
rect 13460 15772 13804 15812
rect 13844 15772 13853 15812
rect 15043 15772 15052 15812
rect 15092 15772 17356 15812
rect 17396 15772 17452 15812
rect 17492 15772 17501 15812
rect 835 15771 893 15772
rect 12547 15771 12605 15772
rect 17347 15771 17405 15772
rect 4099 15728 4157 15729
rect 931 15688 940 15728
rect 980 15688 1228 15728
rect 1268 15688 1277 15728
rect 3811 15688 3820 15728
rect 3860 15688 4108 15728
rect 4148 15688 4396 15728
rect 4436 15688 4445 15728
rect 5443 15688 5452 15728
rect 5492 15688 5932 15728
rect 5972 15688 5981 15728
rect 7660 15688 11500 15728
rect 11540 15688 11549 15728
rect 11683 15688 11692 15728
rect 11732 15688 12172 15728
rect 12212 15688 13324 15728
rect 13364 15688 14764 15728
rect 14804 15688 14813 15728
rect 19747 15688 19756 15728
rect 19796 15688 20044 15728
rect 20084 15688 20093 15728
rect 4099 15687 4157 15688
rect 3331 15604 3340 15644
rect 3380 15604 4012 15644
rect 4052 15604 4061 15644
rect 6883 15604 6892 15644
rect 6932 15604 7180 15644
rect 7220 15604 7229 15644
rect 6979 15560 7037 15561
rect 3235 15520 3244 15560
rect 3284 15520 4108 15560
rect 4148 15520 4157 15560
rect 4579 15520 4588 15560
rect 4628 15520 5068 15560
rect 5108 15520 5548 15560
rect 5588 15520 5597 15560
rect 6691 15520 6700 15560
rect 6740 15520 6988 15560
rect 7028 15520 7037 15560
rect 6979 15519 7037 15520
rect 7171 15560 7229 15561
rect 7171 15520 7180 15560
rect 7220 15520 7276 15560
rect 7316 15520 7325 15560
rect 7171 15519 7229 15520
rect 1795 15476 1853 15477
rect 1219 15436 1228 15476
rect 1268 15436 1804 15476
rect 1844 15436 4204 15476
rect 4244 15436 4253 15476
rect 5251 15436 5260 15476
rect 5300 15436 6604 15476
rect 6644 15436 6988 15476
rect 7028 15436 7037 15476
rect 1795 15435 1853 15436
rect 0 15392 80 15412
rect 7555 15392 7613 15393
rect 0 15352 7564 15392
rect 7604 15352 7613 15392
rect 0 15332 80 15352
rect 7555 15351 7613 15352
rect 3619 15308 3677 15309
rect 5539 15308 5597 15309
rect 7660 15308 7700 15688
rect 8899 15644 8957 15645
rect 10915 15644 10973 15645
rect 19651 15644 19709 15645
rect 20515 15644 20573 15645
rect 8814 15604 8908 15644
rect 8948 15604 8957 15644
rect 9283 15604 9292 15644
rect 9332 15604 10924 15644
rect 10964 15604 13132 15644
rect 13172 15604 13181 15644
rect 13411 15604 13420 15644
rect 13460 15604 15148 15644
rect 15188 15604 15197 15644
rect 15820 15604 19660 15644
rect 19700 15604 19709 15644
rect 19939 15604 19948 15644
rect 19988 15604 20524 15644
rect 20564 15604 20573 15644
rect 8899 15603 8957 15604
rect 10915 15603 10973 15604
rect 15820 15561 15860 15604
rect 19651 15603 19709 15604
rect 20515 15603 20573 15604
rect 11587 15560 11645 15561
rect 15811 15560 15869 15561
rect 19363 15560 19421 15561
rect 9379 15520 9388 15560
rect 9428 15520 10444 15560
rect 10484 15520 10493 15560
rect 11502 15520 11596 15560
rect 11636 15520 11645 15560
rect 13027 15520 13036 15560
rect 13076 15520 13708 15560
rect 13748 15520 14284 15560
rect 14324 15520 14333 15560
rect 15726 15520 15820 15560
rect 15860 15520 15869 15560
rect 16195 15520 16204 15560
rect 16244 15520 19276 15560
rect 19316 15520 19372 15560
rect 19412 15520 19421 15560
rect 11587 15519 11645 15520
rect 15811 15519 15869 15520
rect 19363 15519 19421 15520
rect 19747 15560 19805 15561
rect 21424 15560 21504 15580
rect 19747 15520 19756 15560
rect 19796 15520 21504 15560
rect 19747 15519 19805 15520
rect 21424 15500 21504 15520
rect 14179 15476 14237 15477
rect 15043 15476 15101 15477
rect 15907 15476 15965 15477
rect 7747 15436 7756 15476
rect 7796 15436 11884 15476
rect 11924 15436 13940 15476
rect 13987 15436 13996 15476
rect 14036 15436 14188 15476
rect 14228 15436 14237 15476
rect 14958 15436 15052 15476
rect 15092 15436 15916 15476
rect 15956 15436 15965 15476
rect 16675 15436 16684 15476
rect 16724 15436 19468 15476
rect 19508 15436 19517 15476
rect 9475 15392 9533 15393
rect 13900 15392 13940 15436
rect 14179 15435 14237 15436
rect 15043 15435 15101 15436
rect 15907 15435 15965 15436
rect 19267 15392 19325 15393
rect 19555 15392 19613 15393
rect 8899 15352 8908 15392
rect 8948 15352 9100 15392
rect 9140 15352 9149 15392
rect 9475 15352 9484 15392
rect 9524 15352 9772 15392
rect 9812 15352 9821 15392
rect 11491 15352 11500 15392
rect 11540 15352 13612 15392
rect 13652 15352 13661 15392
rect 13900 15352 16396 15392
rect 16436 15352 16445 15392
rect 16963 15352 16972 15392
rect 17012 15352 17260 15392
rect 17300 15352 17309 15392
rect 17635 15352 17644 15392
rect 17684 15352 17932 15392
rect 17972 15352 17981 15392
rect 19267 15352 19276 15392
rect 19316 15352 19564 15392
rect 19604 15352 19756 15392
rect 19796 15352 19805 15392
rect 9475 15351 9533 15352
rect 19267 15351 19325 15352
rect 19555 15351 19613 15352
rect 1987 15268 1996 15308
rect 2036 15268 3244 15308
rect 3284 15268 3293 15308
rect 3534 15268 3628 15308
rect 3668 15268 3677 15308
rect 4195 15268 4204 15308
rect 4244 15268 5452 15308
rect 5492 15268 5548 15308
rect 5588 15268 5597 15308
rect 6691 15268 6700 15308
rect 6740 15268 7700 15308
rect 11779 15268 11788 15308
rect 11828 15268 12268 15308
rect 12308 15268 14860 15308
rect 14900 15268 14909 15308
rect 16291 15268 16300 15308
rect 16340 15268 18412 15308
rect 18452 15268 19660 15308
rect 19700 15268 19709 15308
rect 3619 15267 3677 15268
rect 5539 15267 5597 15268
rect 7651 15224 7709 15225
rect 8035 15224 8093 15225
rect 15811 15224 15869 15225
rect 21424 15224 21504 15244
rect 3139 15184 3148 15224
rect 3188 15184 4300 15224
rect 4340 15184 4349 15224
rect 7566 15184 7660 15224
rect 7700 15184 8044 15224
rect 8084 15184 8093 15224
rect 8995 15184 9004 15224
rect 9044 15184 9772 15224
rect 9812 15184 11116 15224
rect 11156 15184 11165 15224
rect 13123 15184 13132 15224
rect 13172 15184 15820 15224
rect 15860 15184 15869 15224
rect 16387 15184 16396 15224
rect 16436 15184 21504 15224
rect 7651 15183 7709 15184
rect 8035 15183 8093 15184
rect 15811 15183 15869 15184
rect 21424 15164 21504 15184
rect 13411 15140 13469 15141
rect 3679 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 4065 15140
rect 6499 15100 6508 15140
rect 6548 15100 9484 15140
rect 9524 15100 9533 15140
rect 10339 15100 10348 15140
rect 10388 15100 10540 15140
rect 10580 15100 10589 15140
rect 11971 15100 11980 15140
rect 12020 15100 13420 15140
rect 13460 15100 13469 15140
rect 14755 15100 14764 15140
rect 14804 15100 15148 15140
rect 15188 15100 15197 15140
rect 16291 15100 16300 15140
rect 16340 15100 16972 15140
rect 17012 15100 17021 15140
rect 18403 15100 18412 15140
rect 18452 15100 18604 15140
rect 18644 15100 18653 15140
rect 18799 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 19185 15140
rect 13411 15099 13469 15100
rect 11299 15056 11357 15057
rect 19843 15056 19901 15057
rect 1987 15016 1996 15056
rect 2036 15016 7564 15056
rect 7604 15016 7613 15056
rect 7660 15016 11308 15056
rect 11348 15016 11357 15056
rect 14267 15016 14276 15056
rect 14316 15016 14572 15056
rect 14612 15016 14621 15056
rect 15427 15016 15436 15056
rect 15476 15016 19852 15056
rect 19892 15016 19901 15056
rect 7660 14972 7700 15016
rect 11299 15015 11357 15016
rect 19843 15015 19901 15016
rect 10147 14972 10205 14973
rect 13891 14972 13949 14973
rect 3331 14932 3340 14972
rect 3380 14932 4108 14972
rect 4148 14932 4157 14972
rect 4675 14932 4684 14972
rect 4724 14932 5452 14972
rect 5492 14932 7700 14972
rect 9955 14932 9964 14972
rect 10004 14932 10156 14972
rect 10196 14932 10205 14972
rect 10627 14932 10636 14972
rect 10676 14932 11404 14972
rect 11444 14932 11453 14972
rect 13891 14932 13900 14972
rect 13940 14932 16588 14972
rect 16628 14932 16637 14972
rect 17155 14932 17164 14972
rect 17204 14932 17548 14972
rect 17588 14932 19756 14972
rect 19796 14932 19805 14972
rect 20227 14932 20236 14972
rect 20276 14932 20620 14972
rect 20660 14932 20669 14972
rect 10147 14931 10205 14932
rect 13891 14931 13949 14932
rect 0 14888 80 14908
rect 1507 14888 1565 14889
rect 4291 14888 4349 14889
rect 11011 14888 11069 14889
rect 14659 14888 14717 14889
rect 0 14848 1268 14888
rect 1422 14848 1516 14888
rect 1556 14848 1565 14888
rect 2467 14848 2476 14888
rect 2516 14848 3148 14888
rect 3188 14848 3724 14888
rect 3764 14848 4300 14888
rect 4340 14848 8332 14888
rect 8372 14848 8381 14888
rect 8803 14848 8812 14888
rect 8852 14848 10348 14888
rect 10388 14848 10397 14888
rect 10926 14848 11020 14888
rect 11060 14848 11069 14888
rect 11587 14848 11596 14888
rect 11636 14848 11645 14888
rect 14574 14848 14668 14888
rect 14708 14848 14717 14888
rect 0 14828 80 14848
rect 1228 14804 1268 14848
rect 1507 14847 1565 14848
rect 3715 14804 3773 14805
rect 4108 14804 4148 14848
rect 4291 14847 4349 14848
rect 11011 14847 11069 14848
rect 11107 14804 11165 14805
rect 11596 14804 11636 14848
rect 14659 14847 14717 14848
rect 15427 14888 15485 14889
rect 16579 14888 16637 14889
rect 20803 14888 20861 14889
rect 21424 14888 21504 14908
rect 15427 14848 15436 14888
rect 15476 14848 16588 14888
rect 16628 14848 16637 14888
rect 17347 14848 17356 14888
rect 17396 14848 18604 14888
rect 18644 14848 18653 14888
rect 20803 14848 20812 14888
rect 20852 14848 21504 14888
rect 15427 14847 15485 14848
rect 16579 14847 16637 14848
rect 20803 14847 20861 14848
rect 21424 14828 21504 14848
rect 1228 14764 3724 14804
rect 3764 14764 3773 14804
rect 4099 14764 4108 14804
rect 4148 14764 4188 14804
rect 9955 14764 9964 14804
rect 10004 14764 10924 14804
rect 10964 14764 10973 14804
rect 11107 14764 11116 14804
rect 11156 14764 11308 14804
rect 11348 14764 11357 14804
rect 11596 14764 14572 14804
rect 14612 14764 14621 14804
rect 15619 14764 15628 14804
rect 15668 14764 19084 14804
rect 19124 14764 19133 14804
rect 3715 14763 3773 14764
rect 11107 14763 11165 14764
rect 1891 14720 1949 14721
rect 13699 14720 13757 14721
rect 14371 14720 14429 14721
rect 19747 14720 19805 14721
rect 1806 14680 1900 14720
rect 1940 14680 1949 14720
rect 4291 14680 4300 14720
rect 4340 14680 5836 14720
rect 5876 14680 5885 14720
rect 6019 14680 6028 14720
rect 6068 14680 7084 14720
rect 7124 14680 9196 14720
rect 9236 14680 9245 14720
rect 9667 14680 9676 14720
rect 9716 14680 12748 14720
rect 12788 14680 12797 14720
rect 13123 14680 13132 14720
rect 13172 14680 13212 14720
rect 13699 14680 13708 14720
rect 13748 14680 13900 14720
rect 13940 14680 14380 14720
rect 14420 14680 14429 14720
rect 16483 14680 16492 14720
rect 16532 14680 19180 14720
rect 19220 14680 19229 14720
rect 19459 14680 19468 14720
rect 19508 14680 19756 14720
rect 19796 14680 19805 14720
rect 1891 14679 1949 14680
rect 4771 14636 4829 14637
rect 8899 14636 8957 14637
rect 13132 14636 13172 14680
rect 13699 14679 13757 14680
rect 14371 14679 14429 14680
rect 19747 14679 19805 14680
rect 13315 14636 13373 14637
rect 1507 14596 1516 14636
rect 1556 14596 1804 14636
rect 1844 14596 1853 14636
rect 4771 14596 4780 14636
rect 4820 14596 7564 14636
rect 7604 14596 7613 14636
rect 8707 14596 8716 14636
rect 8756 14596 8908 14636
rect 8948 14596 8957 14636
rect 10435 14596 10444 14636
rect 10484 14596 11308 14636
rect 11348 14596 11357 14636
rect 12835 14596 12844 14636
rect 12884 14596 13324 14636
rect 13364 14596 13373 14636
rect 4771 14595 4829 14596
rect 8899 14595 8957 14596
rect 13315 14595 13373 14596
rect 13603 14636 13661 14637
rect 19459 14636 19517 14637
rect 13603 14596 13612 14636
rect 13652 14596 13996 14636
rect 14036 14596 15052 14636
rect 15092 14596 15101 14636
rect 16771 14596 16780 14636
rect 16820 14596 17644 14636
rect 17684 14596 17693 14636
rect 19459 14596 19468 14636
rect 19508 14596 19564 14636
rect 19604 14596 19613 14636
rect 13603 14595 13661 14596
rect 19459 14595 19517 14596
rect 5731 14552 5789 14553
rect 6403 14552 6461 14553
rect 16099 14552 16157 14553
rect 21091 14552 21149 14553
rect 21424 14552 21504 14572
rect 5731 14512 5740 14552
rect 5780 14512 6220 14552
rect 6260 14512 6269 14552
rect 6403 14512 6412 14552
rect 6452 14512 6892 14552
rect 6932 14512 6941 14552
rect 8323 14512 8332 14552
rect 8372 14512 8812 14552
rect 8852 14512 9964 14552
rect 10004 14512 10013 14552
rect 12643 14512 12652 14552
rect 12692 14512 13036 14552
rect 13076 14512 13085 14552
rect 16099 14512 16108 14552
rect 16148 14512 17356 14552
rect 17396 14512 17405 14552
rect 21091 14512 21100 14552
rect 21140 14512 21504 14552
rect 5731 14511 5789 14512
rect 6403 14511 6461 14512
rect 16099 14511 16157 14512
rect 21091 14511 21149 14512
rect 21424 14492 21504 14512
rect 3139 14468 3197 14469
rect 12163 14468 12221 14469
rect 17155 14468 17213 14469
rect 1804 14428 3148 14468
rect 3188 14428 9676 14468
rect 9716 14428 9725 14468
rect 9772 14428 11596 14468
rect 11636 14428 12172 14468
rect 12212 14428 12556 14468
rect 12596 14428 12605 14468
rect 17155 14428 17164 14468
rect 17204 14428 17452 14468
rect 17492 14428 17501 14468
rect 0 14384 80 14404
rect 1804 14384 1844 14428
rect 3139 14427 3197 14428
rect 9187 14384 9245 14385
rect 0 14344 1132 14384
rect 1172 14344 1181 14384
rect 1795 14344 1804 14384
rect 1844 14344 1853 14384
rect 1987 14344 1996 14384
rect 2036 14344 2045 14384
rect 2755 14344 2764 14384
rect 2804 14344 2813 14384
rect 4919 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 5305 14384
rect 5539 14344 5548 14384
rect 5588 14344 7948 14384
rect 7988 14344 7997 14384
rect 9102 14344 9196 14384
rect 9236 14344 9245 14384
rect 0 14324 80 14344
rect 1996 14300 2036 14344
rect 1315 14260 1324 14300
rect 1364 14260 1900 14300
rect 1940 14260 2036 14300
rect 2764 14300 2804 14344
rect 9187 14343 9245 14344
rect 3139 14300 3197 14301
rect 9772 14300 9812 14428
rect 12163 14427 12221 14428
rect 17155 14427 17213 14428
rect 16291 14384 16349 14385
rect 9955 14344 9964 14384
rect 10004 14344 10348 14384
rect 10388 14344 10397 14384
rect 10819 14344 10828 14384
rect 10868 14344 15668 14384
rect 16206 14344 16300 14384
rect 16340 14344 16349 14384
rect 16771 14344 16780 14384
rect 16820 14344 19372 14384
rect 19412 14344 19421 14384
rect 20039 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20425 14384
rect 15628 14300 15668 14344
rect 16291 14343 16349 14344
rect 20899 14300 20957 14301
rect 2764 14260 3148 14300
rect 3188 14260 3197 14300
rect 4771 14260 4780 14300
rect 4820 14260 7180 14300
rect 7220 14260 9812 14300
rect 10915 14260 10924 14300
rect 10964 14260 11116 14300
rect 11156 14260 11165 14300
rect 11395 14260 11404 14300
rect 11444 14260 12308 14300
rect 12355 14260 12364 14300
rect 12404 14260 12556 14300
rect 12596 14260 12605 14300
rect 12835 14260 12844 14300
rect 12884 14260 14476 14300
rect 14516 14260 14525 14300
rect 15043 14260 15052 14300
rect 15092 14260 15101 14300
rect 15628 14260 17644 14300
rect 17684 14260 17693 14300
rect 20899 14260 20908 14300
rect 20948 14260 21236 14300
rect 3139 14259 3197 14260
rect 4195 14216 4253 14217
rect 5443 14216 5501 14217
rect 6979 14216 7037 14217
rect 12268 14216 12308 14260
rect 15052 14216 15092 14260
rect 20899 14259 20957 14260
rect 21196 14216 21236 14260
rect 21424 14216 21504 14236
rect 1987 14176 1996 14216
rect 2036 14176 2188 14216
rect 2228 14176 2237 14216
rect 4195 14176 4204 14216
rect 4244 14176 4876 14216
rect 4916 14176 4925 14216
rect 5443 14176 5452 14216
rect 5492 14176 5644 14216
rect 5684 14176 5693 14216
rect 6979 14176 6988 14216
rect 7028 14176 8716 14216
rect 8756 14176 8765 14216
rect 9955 14176 9964 14216
rect 10004 14176 10156 14216
rect 10196 14176 11884 14216
rect 11924 14176 11933 14216
rect 12268 14176 14764 14216
rect 14804 14176 14813 14216
rect 15052 14176 21100 14216
rect 21140 14176 21149 14216
rect 21196 14176 21504 14216
rect 4195 14175 4253 14176
rect 5443 14175 5501 14176
rect 6979 14175 7037 14176
rect 21424 14156 21504 14176
rect 8899 14132 8957 14133
rect 17155 14132 17213 14133
rect 8814 14092 8908 14132
rect 8948 14092 8957 14132
rect 10723 14092 10732 14132
rect 10772 14092 11788 14132
rect 11828 14092 11837 14132
rect 12931 14092 12940 14132
rect 12980 14092 16876 14132
rect 16916 14092 16925 14132
rect 17070 14092 17164 14132
rect 17204 14092 17213 14132
rect 20227 14092 20236 14132
rect 20276 14092 20812 14132
rect 20852 14092 20861 14132
rect 8899 14091 8957 14092
rect 17155 14091 17213 14092
rect 16099 14048 16157 14049
rect 2500 14008 7468 14048
rect 7508 14008 7517 14048
rect 10531 14008 10540 14048
rect 10580 14008 11116 14048
rect 11156 14008 11165 14048
rect 11491 14008 11500 14048
rect 11540 14008 11980 14048
rect 12020 14008 12029 14048
rect 12355 14008 12364 14048
rect 12404 14008 12844 14048
rect 12884 14008 13612 14048
rect 13652 14008 13661 14048
rect 14467 14008 14476 14048
rect 14516 14008 14860 14048
rect 14900 14008 15628 14048
rect 15668 14008 15677 14048
rect 16099 14008 16108 14048
rect 16148 14008 17260 14048
rect 17300 14008 17309 14048
rect 1315 13964 1373 13965
rect 2371 13964 2429 13965
rect 2500 13964 2540 14008
rect 16099 14007 16157 14008
rect 3427 13964 3485 13965
rect 10147 13964 10205 13965
rect 17635 13964 17693 13965
rect 1315 13924 1324 13964
rect 1364 13924 2380 13964
rect 2420 13924 2540 13964
rect 2851 13924 2860 13964
rect 2900 13924 3436 13964
rect 3476 13924 3532 13964
rect 3572 13924 3581 13964
rect 10147 13924 10156 13964
rect 10196 13924 11212 13964
rect 11252 13924 12596 13964
rect 13987 13924 13996 13964
rect 14036 13924 14668 13964
rect 14708 13924 15244 13964
rect 15284 13924 15293 13964
rect 17635 13924 17644 13964
rect 17684 13924 20044 13964
rect 20084 13924 20093 13964
rect 1315 13923 1373 13924
rect 2371 13923 2429 13924
rect 3427 13923 3485 13924
rect 10147 13923 10205 13924
rect 0 13880 80 13900
rect 1123 13880 1181 13881
rect 10051 13880 10109 13881
rect 12556 13880 12596 13924
rect 17635 13923 17693 13924
rect 18307 13880 18365 13881
rect 18691 13880 18749 13881
rect 19843 13880 19901 13881
rect 21424 13880 21504 13900
rect 0 13840 1132 13880
rect 1172 13840 1181 13880
rect 2275 13840 2284 13880
rect 2324 13840 2572 13880
rect 2612 13840 2621 13880
rect 2668 13840 4492 13880
rect 4532 13840 4541 13880
rect 4867 13840 4876 13880
rect 4916 13840 9388 13880
rect 9428 13840 9437 13880
rect 9966 13840 10060 13880
rect 10100 13840 10109 13880
rect 10531 13840 10540 13880
rect 10580 13840 10732 13880
rect 10772 13840 11596 13880
rect 11636 13840 11645 13880
rect 11692 13840 12500 13880
rect 12547 13840 12556 13880
rect 12596 13840 12605 13880
rect 12652 13840 13612 13880
rect 13652 13840 13661 13880
rect 13891 13840 13900 13880
rect 13940 13840 15724 13880
rect 15764 13840 15773 13880
rect 16003 13840 16012 13880
rect 16052 13840 18316 13880
rect 18356 13840 18365 13880
rect 18606 13840 18700 13880
rect 18740 13840 18749 13880
rect 18979 13840 18988 13880
rect 19028 13840 19660 13880
rect 19700 13840 19709 13880
rect 19756 13840 19852 13880
rect 19892 13840 21504 13880
rect 0 13820 80 13840
rect 1123 13839 1181 13840
rect 1987 13796 2045 13797
rect 2467 13796 2525 13797
rect 1315 13756 1324 13796
rect 1364 13756 1996 13796
rect 2036 13756 2476 13796
rect 2516 13756 2525 13796
rect 1987 13755 2045 13756
rect 2467 13755 2525 13756
rect 2668 13712 2708 13840
rect 10051 13839 10109 13840
rect 5827 13796 5885 13797
rect 11299 13796 11357 13797
rect 11692 13796 11732 13840
rect 5827 13756 5836 13796
rect 5876 13756 7468 13796
rect 7508 13756 7517 13796
rect 11107 13756 11116 13796
rect 11156 13756 11308 13796
rect 11348 13756 11732 13796
rect 12460 13796 12500 13840
rect 12652 13796 12692 13840
rect 18307 13839 18365 13840
rect 18691 13839 18749 13840
rect 14083 13796 14141 13797
rect 15427 13796 15485 13797
rect 12460 13756 12692 13796
rect 13027 13756 13036 13796
rect 13076 13756 14092 13796
rect 14132 13756 15436 13796
rect 15476 13756 15485 13796
rect 5827 13755 5885 13756
rect 11299 13755 11357 13756
rect 14083 13755 14141 13756
rect 15427 13755 15485 13756
rect 17059 13796 17117 13797
rect 18595 13796 18653 13797
rect 19756 13796 19796 13840
rect 19843 13839 19901 13840
rect 21424 13820 21504 13840
rect 17059 13756 17068 13796
rect 17108 13756 18604 13796
rect 18644 13756 18653 13796
rect 17059 13755 17117 13756
rect 18595 13755 18653 13756
rect 18700 13756 19180 13796
rect 19220 13756 19229 13796
rect 19747 13756 19756 13796
rect 19796 13756 19805 13796
rect 2275 13672 2284 13712
rect 2324 13672 2708 13712
rect 3532 13672 6508 13712
rect 6548 13672 6557 13712
rect 12451 13672 12460 13712
rect 12500 13672 12652 13712
rect 12692 13672 12701 13712
rect 14083 13672 14092 13712
rect 14132 13672 16628 13712
rect 1987 13628 2045 13629
rect 3532 13628 3572 13672
rect 10339 13628 10397 13629
rect 1987 13588 1996 13628
rect 2036 13588 3572 13628
rect 3679 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 4065 13628
rect 6508 13588 6892 13628
rect 6932 13588 6941 13628
rect 9667 13588 9676 13628
rect 9716 13588 10348 13628
rect 10388 13588 10397 13628
rect 1987 13587 2045 13588
rect 1795 13544 1853 13545
rect 6508 13544 6548 13588
rect 10339 13587 10397 13588
rect 11011 13628 11069 13629
rect 11011 13588 11020 13628
rect 11060 13588 14476 13628
rect 14516 13588 14525 13628
rect 15235 13588 15244 13628
rect 15284 13588 15916 13628
rect 15956 13588 15965 13628
rect 11011 13587 11069 13588
rect 12355 13544 12413 13545
rect 1795 13504 1804 13544
rect 1844 13504 6548 13544
rect 6595 13504 6604 13544
rect 6644 13504 7660 13544
rect 7700 13504 10156 13544
rect 10196 13504 10205 13544
rect 12355 13504 12364 13544
rect 12404 13504 16492 13544
rect 16532 13504 16541 13544
rect 1795 13503 1853 13504
rect 12355 13503 12413 13504
rect 9667 13460 9725 13461
rect 10531 13460 10589 13461
rect 16588 13460 16628 13672
rect 18700 13628 18740 13756
rect 18691 13588 18700 13628
rect 18740 13588 18749 13628
rect 18799 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 19185 13628
rect 21424 13544 21504 13564
rect 18403 13504 18412 13544
rect 18452 13504 21504 13544
rect 21424 13484 21504 13504
rect 19555 13460 19613 13461
rect 2179 13420 2188 13460
rect 2228 13420 6124 13460
rect 6164 13420 6173 13460
rect 9667 13420 9676 13460
rect 9716 13420 9772 13460
rect 9812 13420 9821 13460
rect 10531 13420 10540 13460
rect 10580 13420 11788 13460
rect 11828 13420 11837 13460
rect 15427 13420 15436 13460
rect 15476 13420 15628 13460
rect 15668 13420 15677 13460
rect 16588 13420 19564 13460
rect 19604 13420 19613 13460
rect 9667 13419 9725 13420
rect 10531 13419 10589 13420
rect 19555 13419 19613 13420
rect 0 13376 80 13396
rect 1699 13376 1757 13377
rect 18691 13376 18749 13377
rect 19267 13376 19325 13377
rect 0 13336 1708 13376
rect 1748 13336 1757 13376
rect 3907 13336 3916 13376
rect 3956 13336 4300 13376
rect 4340 13336 4349 13376
rect 6307 13336 6316 13376
rect 6356 13336 16972 13376
rect 17012 13336 17021 13376
rect 18691 13336 18700 13376
rect 18740 13336 18796 13376
rect 18836 13336 18845 13376
rect 19075 13336 19084 13376
rect 19124 13336 19276 13376
rect 19316 13336 19325 13376
rect 0 13316 80 13336
rect 1699 13335 1757 13336
rect 18691 13335 18749 13336
rect 19267 13335 19325 13336
rect 11587 13292 11645 13293
rect 16675 13292 16733 13293
rect 3043 13252 3052 13292
rect 3092 13252 5780 13292
rect 6979 13252 6988 13292
rect 7028 13252 7180 13292
rect 7220 13252 7852 13292
rect 7892 13252 7901 13292
rect 8800 13252 11596 13292
rect 11636 13252 15436 13292
rect 15476 13252 15485 13292
rect 16675 13252 16684 13292
rect 16724 13252 20180 13292
rect 5740 13209 5780 13252
rect 1507 13208 1565 13209
rect 4483 13208 4541 13209
rect 5731 13208 5789 13209
rect 8227 13208 8285 13209
rect 8515 13208 8573 13209
rect 1315 13168 1324 13208
rect 1364 13168 1516 13208
rect 1556 13168 1565 13208
rect 3619 13168 3628 13208
rect 3668 13168 4492 13208
rect 4532 13168 4541 13208
rect 5251 13168 5260 13208
rect 5300 13168 5548 13208
rect 5588 13168 5597 13208
rect 5731 13168 5740 13208
rect 5780 13168 6124 13208
rect 6164 13168 6173 13208
rect 6691 13168 6700 13208
rect 6740 13168 7468 13208
rect 7508 13168 7517 13208
rect 8227 13168 8236 13208
rect 8276 13168 8524 13208
rect 8564 13168 8573 13208
rect 1507 13167 1565 13168
rect 4483 13167 4541 13168
rect 5731 13167 5789 13168
rect 8227 13167 8285 13168
rect 8515 13167 8573 13168
rect 4579 13124 4637 13125
rect 4579 13084 4588 13124
rect 4628 13084 8332 13124
rect 8372 13084 8381 13124
rect 4579 13083 4637 13084
rect 2467 13040 2525 13041
rect 4483 13040 4541 13041
rect 8800 13040 8840 13252
rect 11587 13251 11645 13252
rect 16675 13251 16733 13252
rect 10435 13208 10493 13209
rect 10435 13168 10444 13208
rect 10484 13168 10540 13208
rect 10580 13168 10589 13208
rect 12259 13168 12268 13208
rect 12308 13168 13036 13208
rect 13076 13168 13085 13208
rect 15331 13168 15340 13208
rect 15380 13168 16108 13208
rect 16148 13168 16157 13208
rect 16675 13168 16684 13208
rect 16724 13168 18316 13208
rect 18356 13168 18508 13208
rect 18548 13168 18557 13208
rect 18691 13168 18700 13208
rect 18740 13168 19660 13208
rect 19700 13168 19709 13208
rect 19939 13168 19948 13208
rect 19988 13168 19997 13208
rect 10435 13167 10493 13168
rect 11107 13124 11165 13125
rect 16291 13124 16349 13125
rect 19948 13124 19988 13168
rect 11107 13084 11116 13124
rect 11156 13084 16300 13124
rect 16340 13084 16349 13124
rect 17827 13084 17836 13124
rect 17876 13084 19988 13124
rect 11107 13083 11165 13084
rect 16291 13083 16349 13084
rect 19363 13040 19421 13041
rect 2467 13000 2476 13040
rect 2516 13000 4300 13040
rect 4340 13000 4349 13040
rect 4483 13000 4492 13040
rect 4532 13000 4626 13040
rect 5155 13000 5164 13040
rect 5204 13000 5740 13040
rect 5780 13000 5789 13040
rect 6307 13000 6316 13040
rect 6356 13000 6604 13040
rect 6644 13000 6653 13040
rect 6700 13000 8840 13040
rect 11587 13000 11596 13040
rect 11636 13000 12172 13040
rect 12212 13000 12221 13040
rect 12835 13000 12844 13040
rect 12884 13000 13132 13040
rect 13172 13000 13181 13040
rect 14851 13000 14860 13040
rect 14900 13000 16108 13040
rect 16148 13000 16157 13040
rect 19278 13000 19372 13040
rect 19412 13000 19421 13040
rect 2467 12999 2525 13000
rect 4483 12999 4541 13000
rect 2179 12956 2237 12957
rect 4492 12956 4532 12999
rect 6700 12956 6740 13000
rect 19363 12999 19421 13000
rect 2179 12916 2188 12956
rect 2228 12916 4532 12956
rect 4588 12916 6740 12956
rect 7939 12956 7997 12957
rect 17155 12956 17213 12957
rect 20140 12956 20180 13252
rect 20515 13208 20573 13209
rect 21424 13208 21504 13228
rect 20515 13168 20524 13208
rect 20564 13168 21504 13208
rect 20515 13167 20573 13168
rect 21424 13148 21504 13168
rect 7939 12916 7948 12956
rect 7988 12916 17164 12956
rect 17204 12916 17213 12956
rect 17635 12916 17644 12956
rect 17684 12916 19756 12956
rect 19796 12916 19805 12956
rect 20140 12916 20852 12956
rect 2179 12915 2237 12916
rect 0 12872 80 12892
rect 4588 12872 4628 12916
rect 7939 12915 7997 12916
rect 17155 12915 17213 12916
rect 17539 12872 17597 12873
rect 0 12832 2572 12872
rect 2612 12832 3340 12872
rect 3380 12832 3389 12872
rect 3523 12832 3532 12872
rect 3572 12832 4204 12872
rect 4244 12832 4628 12872
rect 4919 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 5305 12872
rect 11299 12832 11308 12872
rect 11348 12832 11980 12872
rect 12020 12832 12029 12872
rect 12163 12832 12172 12872
rect 12212 12832 12940 12872
rect 12980 12832 12989 12872
rect 13507 12832 13516 12872
rect 13556 12832 14092 12872
rect 14132 12832 14141 12872
rect 15235 12832 15244 12872
rect 15284 12832 17548 12872
rect 17588 12832 17597 12872
rect 0 12812 80 12832
rect 17539 12831 17597 12832
rect 19459 12872 19517 12873
rect 20812 12872 20852 12916
rect 21424 12872 21504 12892
rect 19459 12832 19468 12872
rect 19508 12832 19564 12872
rect 19604 12832 19613 12872
rect 20039 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20425 12872
rect 20812 12832 21504 12872
rect 19459 12831 19517 12832
rect 21424 12812 21504 12832
rect 9571 12788 9629 12789
rect 16387 12788 16445 12789
rect 1507 12748 1516 12788
rect 1556 12748 2092 12788
rect 2132 12748 2141 12788
rect 5443 12748 5452 12788
rect 5492 12748 6028 12788
rect 6068 12748 6077 12788
rect 9571 12748 9580 12788
rect 9620 12748 11360 12788
rect 13315 12748 13324 12788
rect 13364 12748 14284 12788
rect 14324 12748 14572 12788
rect 14612 12748 14621 12788
rect 16387 12748 16396 12788
rect 16436 12748 20084 12788
rect 9571 12747 9629 12748
rect 2083 12704 2141 12705
rect 9667 12704 9725 12705
rect 11320 12704 11360 12748
rect 16387 12747 16445 12748
rect 20044 12704 20084 12748
rect 2083 12664 2092 12704
rect 2132 12664 5836 12704
rect 5876 12664 5885 12704
rect 9667 12664 9676 12704
rect 9716 12664 9772 12704
rect 9812 12664 9821 12704
rect 10147 12664 10156 12704
rect 10196 12664 10772 12704
rect 11320 12664 17068 12704
rect 17108 12664 17117 12704
rect 17635 12664 17644 12704
rect 17684 12664 18028 12704
rect 18068 12664 18077 12704
rect 20035 12664 20044 12704
rect 20084 12664 20093 12704
rect 2083 12663 2141 12664
rect 9667 12663 9725 12664
rect 8419 12620 8477 12621
rect 8899 12620 8957 12621
rect 5635 12580 5644 12620
rect 5684 12580 7564 12620
rect 7604 12580 7613 12620
rect 8419 12580 8428 12620
rect 8468 12580 8908 12620
rect 8948 12580 8957 12620
rect 9772 12620 9812 12664
rect 10732 12620 10772 12664
rect 12163 12620 12221 12621
rect 17827 12620 17885 12621
rect 9772 12580 10252 12620
rect 10292 12580 10301 12620
rect 10732 12580 10868 12620
rect 12078 12580 12172 12620
rect 12212 12580 12221 12620
rect 13123 12580 13132 12620
rect 13172 12580 13612 12620
rect 13652 12580 13996 12620
rect 14036 12580 14045 12620
rect 17443 12580 17452 12620
rect 17492 12580 17836 12620
rect 17876 12580 17885 12620
rect 8419 12579 8477 12580
rect 8899 12579 8957 12580
rect 2947 12536 3005 12537
rect 1315 12496 1324 12536
rect 1364 12496 2540 12536
rect 2500 12452 2540 12496
rect 2947 12496 2956 12536
rect 2996 12496 6412 12536
rect 6452 12496 6461 12536
rect 9955 12496 9964 12536
rect 10004 12496 10732 12536
rect 10772 12496 10781 12536
rect 2947 12495 3005 12496
rect 4099 12452 4157 12453
rect 6499 12452 6557 12453
rect 9667 12452 9725 12453
rect 10828 12452 10868 12580
rect 12163 12579 12221 12580
rect 17827 12579 17885 12580
rect 18403 12620 18461 12621
rect 20611 12620 20669 12621
rect 18403 12580 18412 12620
rect 18452 12580 18604 12620
rect 18644 12580 18653 12620
rect 19939 12580 19948 12620
rect 19988 12580 20620 12620
rect 20660 12580 20669 12620
rect 18403 12579 18461 12580
rect 20611 12579 20669 12580
rect 21424 12536 21504 12556
rect 12739 12496 12748 12536
rect 12788 12496 13804 12536
rect 13844 12496 13853 12536
rect 14467 12496 14476 12536
rect 14516 12496 17260 12536
rect 17300 12496 17309 12536
rect 18019 12496 18028 12536
rect 18068 12496 18796 12536
rect 18836 12496 19180 12536
rect 19220 12496 19229 12536
rect 19276 12496 19892 12536
rect 15907 12452 15965 12453
rect 19276 12452 19316 12496
rect 19747 12452 19805 12453
rect 2500 12412 4108 12452
rect 4148 12412 4157 12452
rect 5827 12412 5836 12452
rect 5876 12412 6508 12452
rect 6548 12412 6557 12452
rect 4099 12411 4157 12412
rect 6499 12411 6557 12412
rect 6988 12412 9524 12452
rect 0 12368 80 12388
rect 0 12328 2900 12368
rect 2947 12328 2956 12368
rect 2996 12328 6892 12368
rect 6932 12328 6941 12368
rect 0 12308 80 12328
rect 2860 12284 2900 12328
rect 3139 12284 3197 12285
rect 2860 12244 3148 12284
rect 3188 12244 3197 12284
rect 3139 12243 3197 12244
rect 3427 12284 3485 12285
rect 4099 12284 4157 12285
rect 3427 12244 3436 12284
rect 3476 12244 3628 12284
rect 3668 12244 3677 12284
rect 3907 12244 3916 12284
rect 3956 12244 4108 12284
rect 4148 12244 4157 12284
rect 3427 12243 3485 12244
rect 4099 12243 4157 12244
rect 5539 12284 5597 12285
rect 6988 12284 7028 12412
rect 9484 12368 9524 12412
rect 9667 12412 9676 12452
rect 9716 12412 10156 12452
rect 10196 12412 10205 12452
rect 10819 12412 10828 12452
rect 10868 12412 10877 12452
rect 11011 12412 11020 12452
rect 11060 12412 11212 12452
rect 11252 12412 11884 12452
rect 11924 12412 11933 12452
rect 14563 12412 14572 12452
rect 14612 12412 15532 12452
rect 15572 12412 15581 12452
rect 15907 12412 15916 12452
rect 15956 12412 19316 12452
rect 19459 12412 19468 12452
rect 19508 12412 19756 12452
rect 19796 12412 19805 12452
rect 19852 12452 19892 12496
rect 20140 12496 21504 12536
rect 20140 12452 20180 12496
rect 21424 12476 21504 12496
rect 19852 12412 20180 12452
rect 20227 12412 20236 12452
rect 20276 12412 20716 12452
rect 20756 12412 20765 12452
rect 9667 12411 9725 12412
rect 15907 12411 15965 12412
rect 19747 12411 19805 12412
rect 9571 12368 9629 12369
rect 8131 12328 8140 12368
rect 8180 12328 8332 12368
rect 8372 12328 8381 12368
rect 9484 12328 9580 12368
rect 9620 12328 9629 12368
rect 10243 12328 10252 12368
rect 10292 12328 20852 12368
rect 9571 12327 9629 12328
rect 7843 12284 7901 12285
rect 10252 12284 10292 12328
rect 5539 12244 5548 12284
rect 5588 12244 6028 12284
rect 6068 12244 6077 12284
rect 6211 12244 6220 12284
rect 6260 12244 7028 12284
rect 7075 12244 7084 12284
rect 7124 12244 7372 12284
rect 7412 12244 7421 12284
rect 7843 12244 7852 12284
rect 7892 12244 9676 12284
rect 9716 12244 9725 12284
rect 9772 12244 10292 12284
rect 10435 12284 10493 12285
rect 11491 12284 11549 12285
rect 10435 12244 10444 12284
rect 10484 12244 11500 12284
rect 11540 12244 11549 12284
rect 11971 12244 11980 12284
rect 12020 12244 15436 12284
rect 15476 12244 15485 12284
rect 5539 12243 5597 12244
rect 7843 12243 7901 12244
rect 9772 12200 9812 12244
rect 10435 12243 10493 12244
rect 11491 12243 11549 12244
rect 10339 12200 10397 12201
rect 16963 12200 17021 12201
rect 1987 12160 1996 12200
rect 2036 12160 2188 12200
rect 2228 12160 2237 12200
rect 9283 12160 9292 12200
rect 9332 12160 9812 12200
rect 9964 12160 10348 12200
rect 10388 12160 16972 12200
rect 17012 12160 17021 12200
rect 20812 12200 20852 12328
rect 21424 12200 21504 12220
rect 20812 12160 21504 12200
rect 9187 12116 9245 12117
rect 9964 12116 10004 12160
rect 10339 12159 10397 12160
rect 16963 12159 17021 12160
rect 21424 12140 21504 12160
rect 13987 12116 14045 12117
rect 355 12076 364 12116
rect 404 12076 2956 12116
rect 2996 12076 3005 12116
rect 3679 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 4065 12116
rect 8707 12076 8716 12116
rect 8756 12076 9196 12116
rect 9236 12076 9245 12116
rect 9571 12076 9580 12116
rect 9620 12076 10004 12116
rect 10060 12076 11596 12116
rect 11636 12076 11645 12116
rect 13987 12076 13996 12116
rect 14036 12076 14572 12116
rect 14612 12076 14621 12116
rect 18799 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 19185 12116
rect 20515 12076 20524 12116
rect 20564 12076 20908 12116
rect 20948 12076 20957 12116
rect 9187 12075 9245 12076
rect 7363 12032 7421 12033
rect 10060 12032 10100 12076
rect 13987 12075 14045 12076
rect 3139 11992 3148 12032
rect 3188 11992 7372 12032
rect 7412 11992 7421 12032
rect 9667 11992 9676 12032
rect 9716 11992 10100 12032
rect 11299 12032 11357 12033
rect 17347 12032 17405 12033
rect 11299 11992 11308 12032
rect 11348 11992 11500 12032
rect 11540 11992 11549 12032
rect 11971 11992 11980 12032
rect 12020 11992 12884 12032
rect 14275 11992 14284 12032
rect 14324 11992 17356 12032
rect 17396 11992 18412 12032
rect 18452 11992 18461 12032
rect 19555 11992 19564 12032
rect 19604 11992 20620 12032
rect 20660 11992 20669 12032
rect 7363 11991 7421 11992
rect 11299 11991 11357 11992
rect 8035 11948 8093 11949
rect 12844 11948 12884 11992
rect 17347 11991 17405 11992
rect 2947 11908 2956 11948
rect 2996 11908 8044 11948
rect 8084 11908 8093 11948
rect 8707 11908 8716 11948
rect 8756 11908 11308 11948
rect 11348 11908 12652 11948
rect 12692 11908 12701 11948
rect 12835 11908 12844 11948
rect 12884 11908 13324 11948
rect 13364 11908 13373 11948
rect 15043 11908 15052 11948
rect 15092 11908 16780 11948
rect 16820 11908 16829 11948
rect 19363 11908 19372 11948
rect 19412 11908 20812 11948
rect 20852 11908 20861 11948
rect 8035 11907 8093 11908
rect 0 11864 80 11884
rect 7555 11864 7613 11865
rect 8419 11864 8477 11865
rect 0 11824 460 11864
rect 500 11824 509 11864
rect 1699 11824 1708 11864
rect 1748 11824 1757 11864
rect 6979 11824 6988 11864
rect 7028 11824 7564 11864
rect 7604 11824 7613 11864
rect 7939 11824 7948 11864
rect 7988 11824 8428 11864
rect 8468 11824 8477 11864
rect 0 11804 80 11824
rect 1708 11780 1748 11824
rect 7555 11823 7613 11824
rect 8419 11823 8477 11824
rect 9187 11864 9245 11865
rect 13891 11864 13949 11865
rect 16675 11864 16733 11865
rect 21424 11864 21504 11884
rect 9187 11824 9196 11864
rect 9236 11824 13420 11864
rect 13460 11824 13900 11864
rect 13940 11824 14284 11864
rect 14324 11824 14333 11864
rect 16675 11824 16684 11864
rect 16724 11824 21504 11864
rect 9187 11823 9245 11824
rect 13891 11823 13949 11824
rect 16675 11823 16733 11824
rect 21424 11804 21504 11824
rect 5731 11780 5789 11781
rect 10435 11780 10493 11781
rect 1708 11740 2996 11780
rect 1219 11696 1277 11697
rect 1219 11656 1228 11696
rect 1268 11656 1324 11696
rect 1364 11656 1373 11696
rect 1699 11656 1708 11696
rect 1748 11656 2476 11696
rect 2516 11656 2525 11696
rect 1219 11655 1277 11656
rect 2956 11612 2996 11740
rect 4684 11740 4780 11780
rect 4820 11740 4829 11780
rect 5251 11740 5260 11780
rect 5300 11740 5740 11780
rect 5780 11740 5789 11780
rect 6595 11740 6604 11780
rect 6644 11740 10444 11780
rect 10484 11740 10493 11780
rect 10915 11740 10924 11780
rect 10964 11740 17452 11780
rect 17492 11740 17501 11780
rect 4195 11696 4253 11697
rect 4195 11656 4204 11696
rect 4244 11656 4396 11696
rect 4436 11656 4588 11696
rect 4628 11656 4637 11696
rect 4195 11655 4253 11656
rect 2947 11572 2956 11612
rect 2996 11572 3005 11612
rect 2083 11528 2141 11529
rect 2083 11488 2092 11528
rect 2132 11488 4588 11528
rect 4628 11488 4637 11528
rect 2083 11487 2141 11488
rect 1411 11444 1469 11445
rect 4684 11444 4724 11740
rect 5731 11739 5789 11740
rect 10435 11739 10493 11740
rect 7939 11696 7997 11697
rect 10723 11696 10781 11697
rect 4867 11656 4876 11696
rect 4916 11656 6988 11696
rect 7028 11656 7372 11696
rect 7412 11656 7421 11696
rect 7854 11656 7948 11696
rect 7988 11656 7997 11696
rect 8611 11656 8620 11696
rect 8660 11656 9772 11696
rect 9812 11656 9821 11696
rect 10638 11656 10732 11696
rect 10772 11656 10781 11696
rect 11587 11656 11596 11696
rect 11636 11656 15148 11696
rect 15188 11656 15197 11696
rect 17539 11656 17548 11696
rect 17588 11656 17836 11696
rect 17876 11656 17885 11696
rect 7939 11655 7997 11656
rect 10723 11655 10781 11656
rect 9283 11612 9341 11613
rect 15427 11612 15485 11613
rect 4771 11572 4780 11612
rect 4820 11572 7564 11612
rect 7604 11572 9004 11612
rect 9044 11572 9053 11612
rect 9187 11572 9196 11612
rect 9236 11572 9292 11612
rect 9332 11572 9341 11612
rect 9475 11572 9484 11612
rect 9524 11572 11212 11612
rect 11252 11572 11980 11612
rect 12020 11572 12029 11612
rect 12163 11572 12172 11612
rect 12212 11572 15140 11612
rect 9283 11571 9341 11572
rect 7267 11528 7325 11529
rect 9571 11528 9629 11529
rect 460 11404 1420 11444
rect 1460 11404 1469 11444
rect 3139 11404 3148 11444
rect 3188 11404 3436 11444
rect 3476 11404 3485 11444
rect 4483 11404 4492 11444
rect 4532 11404 4724 11444
rect 4780 11488 5068 11528
rect 5108 11488 5117 11528
rect 7182 11488 7276 11528
rect 7316 11488 7325 11528
rect 8323 11488 8332 11528
rect 8372 11488 8381 11528
rect 9571 11488 9580 11528
rect 9620 11488 9964 11528
rect 10004 11488 10013 11528
rect 11395 11488 11404 11528
rect 11444 11488 12076 11528
rect 12116 11488 12556 11528
rect 12596 11488 12605 11528
rect 0 11360 80 11380
rect 460 11360 500 11404
rect 1411 11403 1469 11404
rect 4780 11360 4820 11488
rect 7267 11487 7325 11488
rect 8332 11444 8372 11488
rect 9571 11487 9629 11488
rect 7276 11404 8372 11444
rect 8419 11444 8477 11445
rect 8419 11404 8428 11444
rect 8468 11404 8660 11444
rect 9763 11404 9772 11444
rect 9812 11404 13804 11444
rect 13844 11404 13853 11444
rect 5923 11360 5981 11361
rect 0 11320 500 11360
rect 4771 11320 4780 11360
rect 4820 11320 4829 11360
rect 4919 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 5305 11360
rect 5838 11320 5932 11360
rect 5972 11320 5981 11360
rect 0 11300 80 11320
rect 5923 11319 5981 11320
rect 6691 11360 6749 11361
rect 7276 11360 7316 11404
rect 8419 11403 8477 11404
rect 7651 11360 7709 11361
rect 8620 11360 8660 11404
rect 11299 11360 11357 11361
rect 15100 11360 15140 11572
rect 15427 11572 15436 11612
rect 15476 11572 16300 11612
rect 16340 11572 18220 11612
rect 18260 11572 18269 11612
rect 15427 11571 15485 11572
rect 16099 11528 16157 11529
rect 21424 11528 21504 11548
rect 16099 11488 16108 11528
rect 16148 11488 16492 11528
rect 16532 11488 16780 11528
rect 16820 11488 16829 11528
rect 17347 11488 17356 11528
rect 17396 11488 21504 11528
rect 16099 11487 16157 11488
rect 21424 11468 21504 11488
rect 17443 11444 17501 11445
rect 17443 11404 17452 11444
rect 17492 11404 18932 11444
rect 17443 11403 17501 11404
rect 16099 11360 16157 11361
rect 6691 11320 6700 11360
rect 6740 11320 6892 11360
rect 6932 11320 6941 11360
rect 7084 11320 7316 11360
rect 7459 11320 7468 11360
rect 7508 11320 7660 11360
rect 7700 11320 7709 11360
rect 8580 11320 8620 11360
rect 8660 11320 8669 11360
rect 11299 11320 11308 11360
rect 11348 11320 13708 11360
rect 13748 11320 13757 11360
rect 14467 11320 14476 11360
rect 14516 11320 14525 11360
rect 15043 11320 15052 11360
rect 15092 11320 15140 11360
rect 16014 11320 16108 11360
rect 16148 11320 16157 11360
rect 6691 11319 6749 11320
rect 5731 11276 5789 11277
rect 7084 11276 7124 11320
rect 7651 11319 7709 11320
rect 3715 11236 3724 11276
rect 3764 11236 5740 11276
rect 5780 11236 5789 11276
rect 6595 11236 6604 11276
rect 6644 11236 7124 11276
rect 7267 11276 7325 11277
rect 7555 11276 7613 11277
rect 8620 11276 8660 11320
rect 11299 11319 11357 11320
rect 14476 11276 14516 11320
rect 16099 11319 16157 11320
rect 7267 11236 7276 11276
rect 7316 11236 7410 11276
rect 7555 11236 7564 11276
rect 7604 11236 7660 11276
rect 7700 11236 7709 11276
rect 7939 11236 7948 11276
rect 7988 11236 8660 11276
rect 9955 11236 9964 11276
rect 10004 11236 10252 11276
rect 10292 11236 10301 11276
rect 11203 11236 11212 11276
rect 11252 11236 13324 11276
rect 13364 11236 13373 11276
rect 13891 11236 13900 11276
rect 13940 11236 14516 11276
rect 18892 11276 18932 11404
rect 20039 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20425 11360
rect 18892 11236 19948 11276
rect 19988 11236 19997 11276
rect 5731 11235 5789 11236
rect 7267 11235 7325 11236
rect 7555 11235 7613 11236
rect 11971 11192 12029 11193
rect 18115 11192 18173 11193
rect 21424 11192 21504 11212
rect 3043 11152 3052 11192
rect 3092 11152 3436 11192
rect 3476 11152 3485 11192
rect 5059 11152 5068 11192
rect 5108 11152 7180 11192
rect 7220 11152 11156 11192
rect 11299 11152 11308 11192
rect 11348 11152 11788 11192
rect 11828 11152 11837 11192
rect 11952 11152 11980 11192
rect 12020 11152 12076 11192
rect 12116 11152 13612 11192
rect 13652 11152 14188 11192
rect 14228 11152 14237 11192
rect 18030 11152 18124 11192
rect 18164 11152 18173 11192
rect 20803 11152 20812 11192
rect 20852 11152 21504 11192
rect 3043 11108 3101 11109
rect 5731 11108 5789 11109
rect 11116 11108 11156 11152
rect 11971 11151 12029 11152
rect 18115 11151 18173 11152
rect 21424 11132 21504 11152
rect 15331 11108 15389 11109
rect 3043 11068 3052 11108
rect 3092 11068 3532 11108
rect 3572 11068 3581 11108
rect 4963 11068 4972 11108
rect 5012 11068 5684 11108
rect 3043 11067 3101 11068
rect 5644 11024 5684 11068
rect 5731 11068 5740 11108
rect 5780 11068 6220 11108
rect 6260 11068 6412 11108
rect 6452 11068 6461 11108
rect 6595 11068 6604 11108
rect 6644 11068 8044 11108
rect 8084 11068 8524 11108
rect 8564 11068 8573 11108
rect 9091 11068 9100 11108
rect 9140 11068 9292 11108
rect 9332 11068 11020 11108
rect 11060 11068 11069 11108
rect 11116 11068 13324 11108
rect 13364 11068 13373 11108
rect 15331 11068 15340 11108
rect 15380 11068 20716 11108
rect 20756 11068 20765 11108
rect 5731 11067 5789 11068
rect 15331 11067 15389 11068
rect 7843 11024 7901 11025
rect 13027 11024 13085 11025
rect 931 10984 940 11024
rect 980 10984 2900 11024
rect 3139 10984 3148 11024
rect 3188 10984 5548 11024
rect 5588 10984 5597 11024
rect 5644 10984 6028 11024
rect 6068 10984 7852 11024
rect 7892 10984 7901 11024
rect 8227 10984 8236 11024
rect 8276 10984 13036 11024
rect 13076 10984 13085 11024
rect 14851 10984 14860 11024
rect 14900 10984 15628 11024
rect 15668 10984 15677 11024
rect 16771 10984 16780 11024
rect 16820 10984 17836 11024
rect 17876 10984 17885 11024
rect 18211 10984 18220 11024
rect 18260 10984 19276 11024
rect 19316 10984 19325 11024
rect 0 10856 80 10876
rect 2860 10856 2900 10984
rect 7843 10983 7901 10984
rect 13027 10983 13085 10984
rect 5539 10940 5597 10941
rect 11491 10940 11549 10941
rect 3235 10900 3244 10940
rect 3284 10900 4396 10940
rect 4436 10900 4445 10940
rect 5155 10900 5164 10940
rect 5204 10900 5548 10940
rect 5588 10900 5597 10940
rect 8035 10900 8044 10940
rect 8084 10900 10444 10940
rect 10484 10900 10493 10940
rect 11491 10900 11500 10940
rect 11540 10900 11634 10940
rect 16675 10900 16684 10940
rect 16724 10900 16733 10940
rect 16963 10900 16972 10940
rect 17012 10900 17644 10940
rect 17684 10900 17693 10940
rect 5539 10899 5597 10900
rect 11491 10899 11549 10900
rect 8803 10856 8861 10857
rect 0 10816 2540 10856
rect 2851 10816 2860 10856
rect 2900 10816 2909 10856
rect 3427 10816 3436 10856
rect 3476 10816 3724 10856
rect 3764 10816 3773 10856
rect 4099 10816 4108 10856
rect 4148 10816 8812 10856
rect 8852 10816 8861 10856
rect 0 10796 80 10816
rect 2500 10772 2540 10816
rect 8803 10815 8861 10816
rect 9571 10856 9629 10857
rect 11587 10856 11645 10857
rect 16684 10856 16724 10900
rect 21424 10856 21504 10876
rect 9571 10816 9580 10856
rect 9620 10816 10732 10856
rect 10772 10816 10781 10856
rect 11502 10816 11596 10856
rect 11636 10816 12364 10856
rect 12404 10816 12413 10856
rect 16684 10816 17164 10856
rect 17204 10816 21504 10856
rect 9571 10815 9629 10816
rect 11587 10815 11645 10816
rect 21424 10796 21504 10816
rect 2500 10732 8812 10772
rect 8852 10732 8861 10772
rect 9091 10732 9100 10772
rect 9140 10732 11308 10772
rect 11348 10732 11357 10772
rect 11596 10732 13708 10772
rect 13748 10732 13757 10772
rect 14275 10732 14284 10772
rect 14324 10732 14860 10772
rect 14900 10732 14909 10772
rect 16387 10732 16396 10772
rect 16436 10732 16876 10772
rect 16916 10732 17644 10772
rect 17684 10732 17693 10772
rect 11596 10688 11636 10732
rect 11779 10688 11837 10689
rect 1603 10648 1612 10688
rect 1652 10648 2668 10688
rect 2708 10648 4204 10688
rect 4244 10648 4253 10688
rect 7651 10648 7660 10688
rect 7700 10648 11636 10688
rect 11683 10648 11692 10688
rect 11732 10648 11788 10688
rect 11828 10648 11837 10688
rect 13708 10688 13748 10732
rect 13708 10648 16012 10688
rect 16052 10648 16061 10688
rect 17731 10648 17740 10688
rect 17780 10648 19468 10688
rect 19508 10648 19852 10688
rect 19892 10648 19901 10688
rect 11779 10647 11837 10648
rect 10531 10604 10589 10605
rect 3679 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 4065 10604
rect 7459 10564 7468 10604
rect 7508 10564 10540 10604
rect 10580 10564 10589 10604
rect 10531 10563 10589 10564
rect 16291 10604 16349 10605
rect 16291 10564 16300 10604
rect 16340 10564 16684 10604
rect 16724 10564 16733 10604
rect 18799 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 19185 10604
rect 16291 10563 16349 10564
rect 11107 10520 11165 10521
rect 15235 10520 15293 10521
rect 3331 10480 3340 10520
rect 3380 10480 11116 10520
rect 11156 10480 11165 10520
rect 11299 10480 11308 10520
rect 11348 10480 11980 10520
rect 12020 10480 12029 10520
rect 15150 10480 15244 10520
rect 15284 10480 15293 10520
rect 11107 10479 11165 10480
rect 15235 10479 15293 10480
rect 15427 10520 15485 10521
rect 20611 10520 20669 10521
rect 21424 10520 21504 10540
rect 15427 10480 15436 10520
rect 15476 10480 15570 10520
rect 16771 10480 16780 10520
rect 16820 10480 17068 10520
rect 17108 10480 17117 10520
rect 17635 10480 17644 10520
rect 17684 10480 18604 10520
rect 18644 10480 18653 10520
rect 20611 10480 20620 10520
rect 20660 10480 21504 10520
rect 15427 10479 15485 10480
rect 20611 10479 20669 10480
rect 21424 10460 21504 10480
rect 5731 10436 5789 10437
rect 2500 10396 5740 10436
rect 5780 10396 5789 10436
rect 0 10352 80 10372
rect 2500 10352 2540 10396
rect 5731 10395 5789 10396
rect 7651 10436 7709 10437
rect 17155 10436 17213 10437
rect 7651 10396 7660 10436
rect 7700 10396 8428 10436
rect 8468 10396 9004 10436
rect 9044 10396 9053 10436
rect 10540 10396 12364 10436
rect 12404 10396 12413 10436
rect 14755 10396 14764 10436
rect 14804 10396 16300 10436
rect 16340 10396 16972 10436
rect 17012 10396 17021 10436
rect 17155 10396 17164 10436
rect 17204 10396 19372 10436
rect 19412 10396 19421 10436
rect 7651 10395 7709 10396
rect 0 10312 2540 10352
rect 3523 10312 3532 10352
rect 3572 10312 4012 10352
rect 4052 10312 4061 10352
rect 4195 10312 4204 10352
rect 4244 10312 5740 10352
rect 5780 10312 5789 10352
rect 0 10292 80 10312
rect 8803 10268 8861 10269
rect 4771 10228 4780 10268
rect 4820 10228 5876 10268
rect 6019 10228 6028 10268
rect 6068 10228 8812 10268
rect 8852 10228 8861 10268
rect 3427 10184 3485 10185
rect 5836 10184 5876 10228
rect 8803 10227 8861 10228
rect 10339 10184 10397 10185
rect 10540 10184 10580 10396
rect 17155 10395 17213 10396
rect 11011 10352 11069 10353
rect 11875 10352 11933 10353
rect 10926 10312 11020 10352
rect 11060 10312 11069 10352
rect 11395 10312 11404 10352
rect 11444 10312 11884 10352
rect 11924 10312 11933 10352
rect 11011 10311 11069 10312
rect 11875 10311 11933 10312
rect 12355 10352 12413 10353
rect 13027 10352 13085 10353
rect 19459 10352 19517 10353
rect 12355 10312 12364 10352
rect 12404 10312 12652 10352
rect 12692 10312 12701 10352
rect 12835 10312 12844 10352
rect 12884 10312 13036 10352
rect 13076 10312 13085 10352
rect 16099 10312 16108 10352
rect 16148 10312 16588 10352
rect 16628 10312 16637 10352
rect 16867 10312 16876 10352
rect 16916 10312 17452 10352
rect 17492 10312 17501 10352
rect 17635 10312 17644 10352
rect 17684 10312 19468 10352
rect 19508 10312 19517 10352
rect 12355 10311 12413 10312
rect 13027 10311 13085 10312
rect 19459 10311 19517 10312
rect 12739 10268 12797 10269
rect 11320 10228 12748 10268
rect 12788 10228 12797 10268
rect 13699 10228 13708 10268
rect 13748 10228 14092 10268
rect 14132 10228 14141 10268
rect 15043 10228 15052 10268
rect 15092 10228 18164 10268
rect 18691 10228 18700 10268
rect 18740 10228 19852 10268
rect 19892 10228 19901 10268
rect 11320 10184 11360 10228
rect 12739 10227 12797 10228
rect 18124 10184 18164 10228
rect 19459 10184 19517 10185
rect 20707 10184 20765 10185
rect 21424 10184 21504 10204
rect 67 10144 76 10184
rect 116 10144 3244 10184
rect 3284 10144 3293 10184
rect 3427 10144 3436 10184
rect 3476 10144 5548 10184
rect 5588 10144 5597 10184
rect 5836 10144 7852 10184
rect 7892 10144 7901 10184
rect 8035 10144 8044 10184
rect 8084 10144 8524 10184
rect 8564 10144 8573 10184
rect 8995 10144 9004 10184
rect 9044 10144 10348 10184
rect 10388 10144 10397 10184
rect 10531 10144 10540 10184
rect 10580 10144 10589 10184
rect 11011 10144 11020 10184
rect 11060 10144 11360 10184
rect 11587 10144 11596 10184
rect 11636 10144 12460 10184
rect 12500 10144 12509 10184
rect 12554 10144 12563 10184
rect 12603 10144 12636 10184
rect 13315 10144 13324 10184
rect 13364 10144 15764 10184
rect 15811 10144 15820 10184
rect 15860 10144 16492 10184
rect 16532 10144 17260 10184
rect 17300 10144 17309 10184
rect 18115 10144 18124 10184
rect 18164 10144 18173 10184
rect 19459 10144 19468 10184
rect 19508 10144 20716 10184
rect 20756 10144 20765 10184
rect 20995 10144 21004 10184
rect 21044 10144 21504 10184
rect 3427 10143 3485 10144
rect 10339 10143 10397 10144
rect 4099 10100 4157 10101
rect 7939 10100 7997 10101
rect 11107 10100 11165 10101
rect 12067 10100 12125 10101
rect 12556 10100 12596 10144
rect 13315 10100 13373 10101
rect 15724 10100 15764 10144
rect 19459 10143 19517 10144
rect 20707 10143 20765 10144
rect 21424 10124 21504 10144
rect 3523 10060 3532 10100
rect 3572 10060 4108 10100
rect 4148 10060 4684 10100
rect 4724 10060 4733 10100
rect 5059 10060 5068 10100
rect 5108 10060 5740 10100
rect 5780 10060 5789 10100
rect 6211 10060 6220 10100
rect 6260 10060 7180 10100
rect 7220 10060 7948 10100
rect 7988 10060 7997 10100
rect 10243 10060 10252 10100
rect 10292 10060 10924 10100
rect 10964 10060 10973 10100
rect 11107 10060 11116 10100
rect 11156 10060 11788 10100
rect 11828 10060 11837 10100
rect 12067 10060 12076 10100
rect 12116 10060 12844 10100
rect 12884 10060 12893 10100
rect 13315 10060 13324 10100
rect 13364 10060 13804 10100
rect 13844 10060 13853 10100
rect 14275 10060 14284 10100
rect 14324 10060 14572 10100
rect 14612 10060 15532 10100
rect 15572 10060 15581 10100
rect 15724 10060 17836 10100
rect 17876 10060 18508 10100
rect 18548 10060 18557 10100
rect 4099 10059 4157 10060
rect 7939 10059 7997 10060
rect 11107 10059 11165 10060
rect 12067 10059 12125 10060
rect 13315 10059 13373 10060
rect 9187 10016 9245 10017
rect 11299 10016 11357 10017
rect 1219 9976 1228 10016
rect 1268 9976 1420 10016
rect 1460 9976 1469 10016
rect 3043 9976 3052 10016
rect 3092 9976 4588 10016
rect 4628 9976 4637 10016
rect 7747 9976 7756 10016
rect 7796 9976 9196 10016
rect 9236 9976 9245 10016
rect 10051 9976 10060 10016
rect 10100 9976 11308 10016
rect 11348 9976 11357 10016
rect 11971 9976 11980 10016
rect 12020 9976 12364 10016
rect 12404 9976 12413 10016
rect 16291 9976 16300 10016
rect 16340 9976 17548 10016
rect 17588 9976 17597 10016
rect 17923 9976 17932 10016
rect 17972 9976 18604 10016
rect 18644 9976 18653 10016
rect 18700 9976 21196 10016
rect 21236 9976 21245 10016
rect 9187 9975 9245 9976
rect 11299 9975 11357 9976
rect 4579 9932 4637 9933
rect 18499 9932 18557 9933
rect 2851 9892 2860 9932
rect 2900 9892 4588 9932
rect 4628 9892 4637 9932
rect 9091 9892 9100 9932
rect 9140 9892 10156 9932
rect 10196 9892 12940 9932
rect 12980 9892 12989 9932
rect 13219 9892 13228 9932
rect 13268 9892 13708 9932
rect 13748 9892 13757 9932
rect 14755 9892 14764 9932
rect 14804 9892 17164 9932
rect 17204 9892 17213 9932
rect 18019 9892 18028 9932
rect 18068 9892 18508 9932
rect 18548 9892 18557 9932
rect 4579 9891 4637 9892
rect 18499 9891 18557 9892
rect 0 9848 80 9868
rect 1219 9848 1277 9849
rect 3427 9848 3485 9849
rect 0 9808 1228 9848
rect 1268 9808 1277 9848
rect 3235 9808 3244 9848
rect 3284 9808 3436 9848
rect 3476 9808 3485 9848
rect 0 9788 80 9808
rect 1219 9807 1277 9808
rect 3427 9807 3485 9808
rect 4291 9848 4349 9849
rect 11107 9848 11165 9849
rect 4291 9808 4300 9848
rect 4340 9808 4492 9848
rect 4532 9808 4541 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 7084 9808 11116 9848
rect 11156 9808 11165 9848
rect 4291 9807 4349 9808
rect 1507 9764 1565 9765
rect 7084 9764 7124 9808
rect 11107 9807 11165 9808
rect 11779 9848 11837 9849
rect 18700 9848 18740 9976
rect 19555 9932 19613 9933
rect 19555 9892 19564 9932
rect 19604 9892 20852 9932
rect 19555 9891 19613 9892
rect 20812 9848 20852 9892
rect 21424 9848 21504 9868
rect 11779 9808 11788 9848
rect 11828 9808 13268 9848
rect 11779 9807 11837 9808
rect 10339 9764 10397 9765
rect 13228 9764 13268 9808
rect 15148 9808 16780 9848
rect 16820 9808 18740 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 20812 9808 21504 9848
rect 13891 9764 13949 9765
rect 15148 9764 15188 9808
rect 21424 9788 21504 9808
rect 1507 9724 1516 9764
rect 1556 9724 1804 9764
rect 1844 9724 1853 9764
rect 2947 9724 2956 9764
rect 2996 9724 7124 9764
rect 7267 9724 7276 9764
rect 7316 9724 10292 9764
rect 1507 9723 1565 9724
rect 3139 9680 3197 9681
rect 3054 9640 3148 9680
rect 3188 9640 3197 9680
rect 3139 9639 3197 9640
rect 4387 9680 4445 9681
rect 9571 9680 9629 9681
rect 4387 9640 4396 9680
rect 4436 9640 4492 9680
rect 4532 9640 4541 9680
rect 4867 9640 4876 9680
rect 4916 9640 9580 9680
rect 9620 9640 9629 9680
rect 10252 9680 10292 9724
rect 10339 9724 10348 9764
rect 10388 9724 10772 9764
rect 10819 9724 10828 9764
rect 10868 9724 12940 9764
rect 12980 9724 12989 9764
rect 13219 9724 13228 9764
rect 13268 9724 13277 9764
rect 13891 9724 13900 9764
rect 13940 9724 14188 9764
rect 14228 9724 14237 9764
rect 15139 9724 15148 9764
rect 15188 9724 15197 9764
rect 16003 9724 16012 9764
rect 16052 9724 17644 9764
rect 17684 9724 18028 9764
rect 18068 9724 18077 9764
rect 10339 9723 10397 9724
rect 10531 9680 10589 9681
rect 10252 9640 10540 9680
rect 10580 9640 10589 9680
rect 4387 9639 4445 9640
rect 9571 9639 9629 9640
rect 10531 9639 10589 9640
rect 1891 9596 1949 9597
rect 2179 9596 2237 9597
rect 1795 9556 1804 9596
rect 1844 9556 1900 9596
rect 1940 9556 2188 9596
rect 2228 9556 2237 9596
rect 1891 9555 1949 9556
rect 2179 9555 2237 9556
rect 3043 9596 3101 9597
rect 10627 9596 10685 9597
rect 3043 9556 3052 9596
rect 3092 9556 3532 9596
rect 3572 9556 3724 9596
rect 3764 9556 3773 9596
rect 6979 9556 6988 9596
rect 7028 9556 9868 9596
rect 9908 9556 9917 9596
rect 10542 9556 10636 9596
rect 10676 9556 10685 9596
rect 10732 9596 10772 9724
rect 13891 9723 13949 9724
rect 11011 9680 11069 9681
rect 12547 9680 12605 9681
rect 13699 9680 13757 9681
rect 10926 9640 11020 9680
rect 11060 9640 11069 9680
rect 11491 9640 11500 9680
rect 11540 9640 12076 9680
rect 12116 9640 12268 9680
rect 12308 9640 12317 9680
rect 12547 9640 12556 9680
rect 12596 9640 12748 9680
rect 12788 9640 12797 9680
rect 13699 9640 13708 9680
rect 13748 9640 16300 9680
rect 16340 9640 16349 9680
rect 16579 9640 16588 9680
rect 16628 9640 17932 9680
rect 17972 9640 17981 9680
rect 18211 9640 18220 9680
rect 18260 9640 20524 9680
rect 20564 9640 20573 9680
rect 11011 9639 11069 9640
rect 12547 9639 12605 9640
rect 13699 9639 13757 9640
rect 10732 9556 13460 9596
rect 13507 9556 13516 9596
rect 13556 9556 14476 9596
rect 14516 9556 14525 9596
rect 14659 9556 14668 9596
rect 14708 9556 15244 9596
rect 15284 9556 15293 9596
rect 15907 9556 15916 9596
rect 15956 9556 18124 9596
rect 18164 9556 18173 9596
rect 19459 9556 19468 9596
rect 19508 9556 20127 9596
rect 20167 9556 20176 9596
rect 3043 9555 3101 9556
rect 10627 9555 10685 9556
rect 3811 9512 3869 9513
rect 9571 9512 9629 9513
rect 13420 9512 13460 9556
rect 21424 9512 21504 9532
rect 1507 9472 1516 9512
rect 1556 9472 1996 9512
rect 2036 9472 2045 9512
rect 3043 9472 3052 9512
rect 3092 9472 3436 9512
rect 3476 9472 3485 9512
rect 3726 9472 3820 9512
rect 3860 9472 4300 9512
rect 4340 9472 4349 9512
rect 5635 9472 5644 9512
rect 5684 9472 6124 9512
rect 6164 9472 7756 9512
rect 7796 9472 7805 9512
rect 9486 9472 9580 9512
rect 9620 9472 9629 9512
rect 10051 9472 10060 9512
rect 10100 9472 10109 9512
rect 13420 9472 15148 9512
rect 15188 9472 15197 9512
rect 15811 9472 15820 9512
rect 15860 9472 16300 9512
rect 16340 9472 16349 9512
rect 16483 9472 16492 9512
rect 16532 9472 16876 9512
rect 16916 9472 17740 9512
rect 17780 9472 17789 9512
rect 17836 9472 19180 9512
rect 19220 9472 19229 9512
rect 20812 9472 21504 9512
rect 3811 9471 3869 9472
rect 9571 9471 9629 9472
rect 10060 9428 10100 9472
rect 1411 9388 1420 9428
rect 1460 9388 8524 9428
rect 8564 9388 8573 9428
rect 8803 9388 8812 9428
rect 8852 9388 9196 9428
rect 9236 9388 10100 9428
rect 11596 9388 12020 9428
rect 12163 9388 12172 9428
rect 12212 9388 12652 9428
rect 12692 9388 13324 9428
rect 13364 9388 13373 9428
rect 16195 9388 16204 9428
rect 16244 9388 17012 9428
rect 0 9344 80 9364
rect 11596 9344 11636 9388
rect 0 9304 11636 9344
rect 11980 9344 12020 9388
rect 15427 9344 15485 9345
rect 16387 9344 16445 9345
rect 11980 9304 12596 9344
rect 15235 9304 15244 9344
rect 15284 9304 15436 9344
rect 15476 9304 15485 9344
rect 16302 9304 16396 9344
rect 16436 9304 16445 9344
rect 0 9284 80 9304
rect 1027 9260 1085 9261
rect 9667 9260 9725 9261
rect 9859 9260 9917 9261
rect 12556 9260 12596 9304
rect 15427 9303 15485 9304
rect 16387 9303 16445 9304
rect 15235 9260 15293 9261
rect 16972 9260 17012 9388
rect 1027 9220 1036 9260
rect 1076 9220 3340 9260
rect 3380 9220 3389 9260
rect 6124 9220 9676 9260
rect 9716 9220 9725 9260
rect 9774 9220 9868 9260
rect 9908 9220 9917 9260
rect 10339 9220 10348 9260
rect 10388 9220 11884 9260
rect 11924 9220 12268 9260
rect 12308 9220 12317 9260
rect 12556 9220 15244 9260
rect 15284 9220 15293 9260
rect 15715 9220 15724 9260
rect 15764 9220 16780 9260
rect 16820 9220 16829 9260
rect 16963 9220 16972 9260
rect 17012 9220 17021 9260
rect 1027 9219 1085 9220
rect 6124 9176 6164 9220
rect 9667 9219 9725 9220
rect 9859 9219 9917 9220
rect 15235 9219 15293 9220
rect 16195 9176 16253 9177
rect 17836 9176 17876 9472
rect 18691 9428 18749 9429
rect 17923 9388 17932 9428
rect 17972 9388 18225 9428
rect 18265 9388 18274 9428
rect 18672 9388 18700 9428
rect 18740 9388 18796 9428
rect 18836 9388 20236 9428
rect 20276 9388 20285 9428
rect 18691 9387 18749 9388
rect 20812 9344 20852 9472
rect 21424 9452 21504 9472
rect 19267 9304 19276 9344
rect 19316 9304 19948 9344
rect 19988 9304 19997 9344
rect 20140 9304 20852 9344
rect 18211 9220 18220 9260
rect 18260 9220 19084 9260
rect 19124 9220 19133 9260
rect 18115 9176 18173 9177
rect 20140 9176 20180 9304
rect 21424 9176 21504 9196
rect 1987 9136 1996 9176
rect 2036 9136 6164 9176
rect 8611 9136 8620 9176
rect 8660 9136 14668 9176
rect 14708 9136 15628 9176
rect 15668 9136 15677 9176
rect 16195 9136 16204 9176
rect 16244 9136 18124 9176
rect 18164 9136 18173 9176
rect 18499 9136 18508 9176
rect 18548 9136 20180 9176
rect 20995 9136 21004 9176
rect 21044 9136 21504 9176
rect 16195 9135 16253 9136
rect 18115 9135 18173 9136
rect 21424 9116 21504 9136
rect 4195 9092 4253 9093
rect 12355 9092 12413 9093
rect 12547 9092 12605 9093
rect 13315 9092 13373 9093
rect 18019 9092 18077 9093
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 4195 9052 4204 9092
rect 4244 9052 4972 9092
rect 5012 9052 5021 9092
rect 6307 9052 6316 9092
rect 6356 9052 6700 9092
rect 6740 9052 6749 9092
rect 9571 9052 9580 9092
rect 9620 9052 10156 9092
rect 10196 9052 10205 9092
rect 10339 9052 10348 9092
rect 10388 9052 10636 9092
rect 10676 9052 10685 9092
rect 11395 9052 11404 9092
rect 11444 9052 12172 9092
rect 12212 9052 12221 9092
rect 12355 9052 12364 9092
rect 12404 9052 12498 9092
rect 12547 9052 12556 9092
rect 12596 9052 12652 9092
rect 12692 9052 12701 9092
rect 13315 9052 13324 9092
rect 13364 9052 18028 9092
rect 18068 9052 18077 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 4195 9051 4253 9052
rect 6307 9008 6365 9009
rect 547 8968 556 9008
rect 596 8968 6316 9008
rect 6356 8968 6365 9008
rect 6307 8967 6365 8968
rect 5731 8924 5789 8925
rect 2179 8884 2188 8924
rect 2228 8884 3244 8924
rect 3284 8884 3293 8924
rect 4291 8884 4300 8924
rect 4340 8884 4684 8924
rect 4724 8884 4733 8924
rect 5646 8884 5740 8924
rect 5780 8884 5789 8924
rect 5731 8883 5789 8884
rect 6115 8924 6173 8925
rect 6115 8884 6124 8924
rect 6164 8884 6173 8924
rect 6700 8924 6740 9052
rect 12355 9051 12413 9052
rect 12547 9051 12605 9052
rect 13315 9051 13373 9052
rect 18019 9051 18077 9052
rect 12643 9008 12701 9009
rect 17059 9008 17117 9009
rect 8515 8968 8524 9008
rect 8564 8968 12652 9008
rect 12692 8968 13420 9008
rect 13460 8968 13469 9008
rect 15331 8968 15340 9008
rect 15380 8968 16204 9008
rect 16244 8968 16253 9008
rect 17059 8968 17068 9008
rect 17108 8968 17164 9008
rect 17204 8968 17213 9008
rect 12643 8967 12701 8968
rect 17059 8967 17117 8968
rect 10531 8924 10589 8925
rect 20803 8924 20861 8925
rect 6700 8884 10348 8924
rect 10388 8884 10397 8924
rect 10531 8884 10540 8924
rect 10580 8884 12460 8924
rect 12500 8884 20812 8924
rect 20852 8884 20861 8924
rect 6115 8883 6173 8884
rect 10531 8883 10589 8884
rect 20803 8883 20861 8884
rect 0 8840 80 8860
rect 6124 8840 6164 8883
rect 21424 8841 21504 8860
rect 6691 8840 6749 8841
rect 9187 8840 9245 8841
rect 0 8800 76 8840
rect 116 8800 125 8840
rect 1036 8800 6028 8840
rect 6068 8800 6077 8840
rect 6124 8800 6220 8840
rect 6260 8800 6269 8840
rect 6691 8800 6700 8840
rect 6740 8800 7084 8840
rect 7124 8800 7133 8840
rect 7939 8800 7948 8840
rect 7988 8800 8140 8840
rect 8180 8800 8189 8840
rect 8995 8800 9004 8840
rect 9044 8800 9196 8840
rect 9236 8800 9245 8840
rect 0 8780 80 8800
rect 643 8756 701 8757
rect 1036 8756 1076 8800
rect 6691 8799 6749 8800
rect 9187 8799 9245 8800
rect 17539 8840 17597 8841
rect 18787 8840 18845 8841
rect 17539 8800 17548 8840
rect 17588 8800 18508 8840
rect 18548 8800 18557 8840
rect 18702 8800 18796 8840
rect 18836 8800 18845 8840
rect 17539 8799 17597 8800
rect 18787 8799 18845 8800
rect 21379 8840 21504 8841
rect 21379 8800 21388 8840
rect 21428 8800 21504 8840
rect 21379 8799 21504 8800
rect 21424 8780 21504 8799
rect 12067 8756 12125 8757
rect 12355 8756 12413 8757
rect 643 8716 652 8756
rect 692 8716 1076 8756
rect 2467 8716 2476 8756
rect 2516 8716 4972 8756
rect 5012 8716 8620 8756
rect 8660 8716 8669 8756
rect 9187 8716 9196 8756
rect 9236 8716 12076 8756
rect 12116 8716 12125 8756
rect 12259 8716 12268 8756
rect 12308 8716 12364 8756
rect 12404 8716 12413 8756
rect 643 8715 701 8716
rect 12067 8715 12125 8716
rect 12355 8715 12413 8716
rect 12643 8756 12701 8757
rect 12643 8716 12652 8756
rect 12692 8716 12748 8756
rect 12788 8716 12797 8756
rect 13315 8716 13324 8756
rect 13364 8716 13996 8756
rect 14036 8716 14045 8756
rect 15139 8716 15148 8756
rect 15188 8716 15476 8756
rect 18400 8716 18409 8756
rect 18449 8716 18458 8756
rect 12643 8715 12701 8716
rect 1219 8672 1277 8673
rect 2179 8672 2237 8673
rect 13324 8672 13364 8716
rect 15331 8672 15389 8673
rect 1134 8632 1228 8672
rect 1268 8632 1277 8672
rect 2094 8632 2188 8672
rect 2228 8632 2237 8672
rect 2563 8632 2572 8672
rect 2612 8632 3532 8672
rect 3572 8632 3581 8672
rect 4195 8632 4204 8672
rect 4244 8632 4876 8672
rect 4916 8632 4925 8672
rect 5347 8632 5356 8672
rect 5396 8632 7660 8672
rect 7700 8632 8716 8672
rect 8756 8632 8765 8672
rect 9091 8632 9100 8672
rect 9140 8632 9964 8672
rect 10004 8632 10636 8672
rect 10676 8632 10828 8672
rect 10868 8632 10877 8672
rect 11107 8632 11116 8672
rect 11156 8632 13364 8672
rect 13411 8632 13420 8672
rect 13460 8632 13612 8672
rect 13652 8632 13661 8672
rect 15246 8632 15340 8672
rect 15380 8632 15389 8672
rect 15436 8672 15476 8716
rect 17443 8672 17501 8673
rect 15436 8632 16780 8672
rect 16820 8632 16829 8672
rect 17059 8632 17068 8672
rect 17108 8632 17452 8672
rect 17492 8632 17501 8672
rect 18412 8672 18452 8716
rect 18412 8632 19756 8672
rect 19796 8632 19805 8672
rect 1219 8631 1277 8632
rect 2179 8631 2237 8632
rect 15331 8631 15389 8632
rect 17443 8631 17501 8632
rect 739 8588 797 8589
rect 12259 8588 12317 8589
rect 18115 8588 18173 8589
rect 739 8548 748 8588
rect 788 8548 2956 8588
rect 2996 8548 3005 8588
rect 4771 8548 4780 8588
rect 4820 8548 7084 8588
rect 7124 8548 7133 8588
rect 9283 8548 9292 8588
rect 9332 8548 9772 8588
rect 9812 8548 10156 8588
rect 10196 8548 10205 8588
rect 10435 8548 10444 8588
rect 10484 8548 11636 8588
rect 11683 8548 11692 8588
rect 11732 8548 11884 8588
rect 11924 8548 11933 8588
rect 12259 8548 12268 8588
rect 12308 8548 13036 8588
rect 13076 8548 13085 8588
rect 18030 8548 18124 8588
rect 18164 8548 18173 8588
rect 18403 8548 18412 8588
rect 18452 8548 18700 8588
rect 18740 8548 18749 8588
rect 739 8547 797 8548
rect 6883 8504 6941 8505
rect 11596 8504 11636 8548
rect 12259 8547 12317 8548
rect 18115 8547 18173 8548
rect 11971 8504 12029 8505
rect 12739 8504 12797 8505
rect 18691 8504 18749 8505
rect 5443 8464 5452 8504
rect 5492 8464 6892 8504
rect 6932 8464 6941 8504
rect 7171 8464 7180 8504
rect 7220 8464 8044 8504
rect 8084 8464 8093 8504
rect 8323 8464 8332 8504
rect 8372 8464 11500 8504
rect 11540 8464 11549 8504
rect 11596 8464 11732 8504
rect 11776 8464 11785 8504
rect 11825 8464 11980 8504
rect 12020 8464 12029 8504
rect 12654 8464 12748 8504
rect 12788 8464 12797 8504
rect 13603 8464 13612 8504
rect 13652 8464 17836 8504
rect 17876 8464 17885 8504
rect 18595 8464 18604 8504
rect 18644 8464 18700 8504
rect 18740 8464 18749 8504
rect 6883 8463 6941 8464
rect 2371 8420 2429 8421
rect 11692 8420 11732 8464
rect 11971 8463 12029 8464
rect 12739 8463 12797 8464
rect 18691 8463 18749 8464
rect 19939 8504 19997 8505
rect 21424 8504 21504 8524
rect 19939 8464 19948 8504
rect 19988 8464 20140 8504
rect 20180 8464 20189 8504
rect 20611 8464 20620 8504
rect 20660 8464 21504 8504
rect 19939 8463 19997 8464
rect 21424 8444 21504 8464
rect 2286 8380 2380 8420
rect 2420 8380 2429 8420
rect 4387 8380 4396 8420
rect 4436 8380 6700 8420
rect 6740 8380 11636 8420
rect 11692 8380 12844 8420
rect 12884 8380 16588 8420
rect 16628 8380 16637 8420
rect 16771 8380 16780 8420
rect 16820 8380 17260 8420
rect 17300 8380 18508 8420
rect 18548 8380 18557 8420
rect 2371 8379 2429 8380
rect 0 8336 80 8356
rect 5731 8336 5789 8337
rect 10531 8336 10589 8337
rect 0 8296 3724 8336
rect 3764 8296 3773 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 5731 8296 5740 8336
rect 5780 8296 6220 8336
rect 6260 8296 6269 8336
rect 7075 8296 7084 8336
rect 7124 8296 9140 8336
rect 9667 8296 9676 8336
rect 9716 8296 9964 8336
rect 10004 8296 10013 8336
rect 10446 8296 10540 8336
rect 10580 8296 10589 8336
rect 0 8276 80 8296
rect 5731 8295 5789 8296
rect 5635 8252 5693 8253
rect 2659 8212 2668 8252
rect 2708 8212 5457 8252
rect 5497 8212 5506 8252
rect 5635 8212 5644 8252
rect 5684 8212 5740 8252
rect 5780 8212 5789 8252
rect 6691 8212 6700 8252
rect 6740 8212 7468 8252
rect 7508 8212 8716 8252
rect 8756 8212 8765 8252
rect 5635 8211 5693 8212
rect 9100 8168 9140 8296
rect 10531 8295 10589 8296
rect 11596 8252 11636 8380
rect 13891 8336 13949 8337
rect 14083 8336 14141 8337
rect 15811 8336 15869 8337
rect 16195 8336 16253 8337
rect 11683 8296 11692 8336
rect 11732 8296 11980 8336
rect 12020 8296 12029 8336
rect 13795 8296 13804 8336
rect 13844 8296 13900 8336
rect 13940 8296 13949 8336
rect 13998 8296 14092 8336
rect 14132 8296 14141 8336
rect 14563 8296 14572 8336
rect 14612 8296 14860 8336
rect 14900 8296 14909 8336
rect 15139 8296 15148 8336
rect 15188 8296 15436 8336
rect 15476 8296 15485 8336
rect 15811 8296 15820 8336
rect 15860 8296 16204 8336
rect 16244 8296 18988 8336
rect 19028 8296 19037 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 13891 8295 13949 8296
rect 14083 8295 14141 8296
rect 15811 8295 15869 8296
rect 16195 8295 16253 8296
rect 15235 8252 15293 8253
rect 9475 8212 9484 8252
rect 9524 8212 9772 8252
rect 9812 8212 9821 8252
rect 10147 8212 10156 8252
rect 10196 8212 11404 8252
rect 11444 8212 11453 8252
rect 11596 8212 15244 8252
rect 15284 8212 15293 8252
rect 17539 8212 17548 8252
rect 17588 8212 20180 8252
rect 15235 8211 15293 8212
rect 18115 8168 18173 8169
rect 19939 8168 19997 8169
rect 20140 8168 20180 8212
rect 21424 8168 21504 8188
rect 2371 8128 2380 8168
rect 2420 8128 4972 8168
rect 5012 8128 5021 8168
rect 7075 8128 7084 8168
rect 7124 8128 9004 8168
rect 9044 8128 9053 8168
rect 9100 8128 11020 8168
rect 11060 8128 11069 8168
rect 11116 8128 11692 8168
rect 11732 8128 11741 8168
rect 12547 8128 12556 8168
rect 12596 8128 14092 8168
rect 14132 8128 14141 8168
rect 14467 8128 14476 8168
rect 14516 8128 14860 8168
rect 14900 8128 14909 8168
rect 18115 8128 18124 8168
rect 18164 8128 18316 8168
rect 18356 8128 18365 8168
rect 18883 8128 18892 8168
rect 18932 8128 18941 8168
rect 19939 8128 19948 8168
rect 19988 8128 20044 8168
rect 20084 8128 20093 8168
rect 20140 8128 21504 8168
rect 11116 8084 11156 8128
rect 18115 8127 18173 8128
rect 12835 8084 12893 8085
rect 18403 8084 18461 8085
rect 3715 8044 3724 8084
rect 3764 8044 7508 8084
rect 8611 8044 8620 8084
rect 8660 8044 8908 8084
rect 8948 8044 8957 8084
rect 9667 8044 9676 8084
rect 9716 8044 11156 8084
rect 11203 8044 11212 8084
rect 11252 8044 11980 8084
rect 12020 8044 12268 8084
rect 12308 8044 12317 8084
rect 12835 8044 12844 8084
rect 12884 8044 15436 8084
rect 15476 8044 15485 8084
rect 16291 8044 16300 8084
rect 16340 8044 16684 8084
rect 16724 8044 16733 8084
rect 16867 8044 16876 8084
rect 16916 8044 17164 8084
rect 17204 8044 18028 8084
rect 18068 8044 18077 8084
rect 18211 8044 18220 8084
rect 18260 8044 18412 8084
rect 18452 8044 18461 8084
rect 18892 8084 18932 8128
rect 19939 8127 19997 8128
rect 21424 8108 21504 8128
rect 19555 8084 19613 8085
rect 18892 8044 19564 8084
rect 19604 8044 20180 8084
rect 1315 7960 1324 8000
rect 1364 7960 2188 8000
rect 2228 7960 2237 8000
rect 2659 7960 2668 8000
rect 2708 7960 5068 8000
rect 5108 7960 5117 8000
rect 0 7832 80 7852
rect 1123 7832 1181 7833
rect 2956 7832 2996 7960
rect 4099 7916 4157 7917
rect 4387 7916 4445 7917
rect 4014 7876 4108 7916
rect 4148 7876 4157 7916
rect 4302 7876 4396 7916
rect 4436 7876 4445 7916
rect 4099 7875 4157 7876
rect 4387 7875 4445 7876
rect 4195 7832 4253 7833
rect 7468 7832 7508 8044
rect 12835 8043 12893 8044
rect 18403 8043 18461 8044
rect 19555 8043 19613 8044
rect 8035 8000 8093 8001
rect 7950 7960 8044 8000
rect 8084 7960 8093 8000
rect 8035 7959 8093 7960
rect 8227 8000 8285 8001
rect 17251 8000 17309 8001
rect 8227 7960 8236 8000
rect 8276 7960 10444 8000
rect 10484 7960 10493 8000
rect 11875 7960 11884 8000
rect 11924 7960 12076 8000
rect 12116 7960 12460 8000
rect 12500 7960 14188 8000
rect 14228 7960 14237 8000
rect 14755 7960 14764 8000
rect 14804 7960 17068 8000
rect 17108 7960 17117 8000
rect 17251 7960 17260 8000
rect 17300 7960 19084 8000
rect 19124 7960 19133 8000
rect 8227 7959 8285 7960
rect 17251 7959 17309 7960
rect 9859 7916 9917 7917
rect 13891 7916 13949 7917
rect 8899 7876 8908 7916
rect 8948 7876 9868 7916
rect 9908 7876 9917 7916
rect 11395 7876 11404 7916
rect 11444 7876 13900 7916
rect 13940 7876 16820 7916
rect 18595 7876 18604 7916
rect 18644 7876 18653 7916
rect 9859 7875 9917 7876
rect 13891 7875 13949 7876
rect 11779 7832 11837 7833
rect 16780 7832 16820 7876
rect 18604 7832 18644 7876
rect 20140 7832 20180 8044
rect 21424 7832 21504 7852
rect 0 7792 1132 7832
rect 1172 7792 1181 7832
rect 2947 7792 2956 7832
rect 2996 7792 3005 7832
rect 4110 7792 4204 7832
rect 4244 7792 4253 7832
rect 5155 7792 5164 7832
rect 5204 7792 7084 7832
rect 7124 7792 7133 7832
rect 7468 7792 11360 7832
rect 11683 7792 11692 7832
rect 11732 7792 11788 7832
rect 11828 7792 16300 7832
rect 16340 7792 16349 7832
rect 16771 7792 16780 7832
rect 16820 7792 17356 7832
rect 17396 7792 17405 7832
rect 17539 7792 17548 7832
rect 17588 7792 18644 7832
rect 18979 7792 18988 7832
rect 19028 7792 19660 7832
rect 19700 7792 19709 7832
rect 20140 7792 21504 7832
rect 0 7772 80 7792
rect 1123 7791 1181 7792
rect 4195 7791 4253 7792
rect 2179 7748 2237 7749
rect 5164 7748 5204 7792
rect 1891 7708 1900 7748
rect 1940 7708 2188 7748
rect 2228 7708 2237 7748
rect 3619 7708 3628 7748
rect 3668 7708 3820 7748
rect 3860 7708 5204 7748
rect 7363 7708 7372 7748
rect 7412 7708 8332 7748
rect 8372 7708 8381 7748
rect 8707 7708 8716 7748
rect 8756 7708 9580 7748
rect 9620 7708 9629 7748
rect 2179 7707 2237 7708
rect 9475 7664 9533 7665
rect 11320 7664 11360 7792
rect 11779 7791 11837 7792
rect 21424 7772 21504 7792
rect 12163 7748 12221 7749
rect 12163 7708 12172 7748
rect 12212 7708 19468 7748
rect 19508 7708 19517 7748
rect 12163 7707 12221 7708
rect 11587 7664 11645 7665
rect 16291 7664 16349 7665
rect 1603 7624 1612 7664
rect 1652 7624 1804 7664
rect 1844 7624 1853 7664
rect 3523 7624 3532 7664
rect 3572 7624 4300 7664
rect 4340 7624 4349 7664
rect 6499 7624 6508 7664
rect 6548 7624 9484 7664
rect 9524 7624 10060 7664
rect 10100 7624 10109 7664
rect 11320 7624 11596 7664
rect 11636 7624 12268 7664
rect 12308 7624 12317 7664
rect 14851 7624 14860 7664
rect 14900 7624 15436 7664
rect 15476 7624 15485 7664
rect 15619 7624 15628 7664
rect 15668 7624 16300 7664
rect 16340 7624 16349 7664
rect 9475 7623 9533 7624
rect 11587 7623 11645 7624
rect 16291 7623 16349 7624
rect 18115 7664 18173 7665
rect 18691 7664 18749 7665
rect 18115 7624 18124 7664
rect 18164 7624 18220 7664
rect 18260 7624 18269 7664
rect 18499 7624 18508 7664
rect 18548 7624 18700 7664
rect 18740 7624 18749 7664
rect 18115 7623 18173 7624
rect 18691 7623 18749 7624
rect 9187 7580 9245 7581
rect 11971 7580 12029 7581
rect 12835 7580 12893 7581
rect 1507 7540 1516 7580
rect 1556 7540 1900 7580
rect 1940 7540 1949 7580
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 4579 7540 4588 7580
rect 4628 7540 7316 7580
rect 7276 7496 7316 7540
rect 9187 7540 9196 7580
rect 9236 7540 9388 7580
rect 9428 7540 9437 7580
rect 11299 7540 11308 7580
rect 11348 7540 11980 7580
rect 12020 7540 12029 7580
rect 12355 7540 12364 7580
rect 12404 7540 12844 7580
rect 12884 7540 12893 7580
rect 14659 7540 14668 7580
rect 14708 7540 18028 7580
rect 18068 7540 18077 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 19363 7540 19372 7580
rect 19412 7540 19660 7580
rect 19700 7540 19709 7580
rect 9187 7539 9245 7540
rect 9283 7496 9341 7497
rect 1603 7456 1612 7496
rect 1652 7456 5260 7496
rect 5300 7456 5309 7496
rect 7276 7456 8428 7496
rect 8468 7456 9100 7496
rect 9140 7456 9149 7496
rect 9283 7456 9292 7496
rect 9332 7456 10156 7496
rect 10196 7456 10205 7496
rect 9283 7455 9341 7456
rect 2947 7412 3005 7413
rect 5635 7412 5693 7413
rect 8035 7412 8093 7413
rect 11308 7412 11348 7540
rect 11971 7539 12029 7540
rect 12835 7539 12893 7540
rect 20995 7496 21053 7497
rect 21424 7496 21504 7516
rect 12067 7456 12076 7496
rect 12116 7456 13516 7496
rect 13556 7456 13565 7496
rect 14371 7456 14380 7496
rect 14420 7456 17740 7496
rect 17780 7456 17789 7496
rect 19756 7456 19852 7496
rect 19892 7456 19901 7496
rect 20995 7456 21004 7496
rect 21044 7456 21504 7496
rect 18691 7412 18749 7413
rect 1987 7372 1996 7412
rect 2036 7372 2956 7412
rect 2996 7372 3005 7412
rect 3811 7372 3820 7412
rect 3860 7372 4492 7412
rect 4532 7372 4541 7412
rect 5550 7372 5644 7412
rect 5684 7372 5693 7412
rect 6499 7372 6508 7412
rect 6548 7372 7564 7412
rect 7604 7372 7613 7412
rect 8035 7372 8044 7412
rect 8084 7372 8236 7412
rect 8276 7372 8285 7412
rect 8995 7372 9004 7412
rect 9044 7372 9484 7412
rect 9524 7372 11348 7412
rect 13603 7372 13612 7412
rect 13652 7372 13996 7412
rect 14036 7372 14045 7412
rect 15235 7372 15244 7412
rect 15284 7372 18700 7412
rect 18740 7372 18749 7412
rect 2947 7371 3005 7372
rect 5635 7371 5693 7372
rect 8035 7371 8093 7372
rect 18691 7371 18749 7372
rect 0 7328 80 7348
rect 15331 7328 15389 7329
rect 15619 7328 15677 7329
rect 0 7288 556 7328
rect 596 7288 605 7328
rect 1507 7288 1516 7328
rect 1556 7288 3436 7328
rect 3476 7288 3485 7328
rect 4099 7288 4108 7328
rect 4148 7288 8716 7328
rect 8756 7288 8908 7328
rect 8948 7288 8957 7328
rect 9571 7288 9580 7328
rect 9620 7288 10540 7328
rect 10580 7288 10589 7328
rect 13507 7288 13516 7328
rect 13556 7288 13708 7328
rect 13748 7288 13757 7328
rect 15043 7288 15052 7328
rect 15092 7288 15101 7328
rect 15246 7288 15340 7328
rect 15380 7288 15389 7328
rect 15534 7288 15628 7328
rect 15668 7288 15677 7328
rect 0 7268 80 7288
rect 7363 7244 7421 7245
rect 8515 7244 8573 7245
rect 12643 7244 12701 7245
rect 4003 7204 4012 7244
rect 4052 7204 6796 7244
rect 6836 7204 6845 7244
rect 7276 7204 7372 7244
rect 7412 7204 8468 7244
rect 4291 7160 4349 7161
rect 172 7120 3188 7160
rect 4195 7120 4204 7160
rect 4244 7120 4300 7160
rect 4340 7120 4349 7160
rect 0 6824 80 6844
rect 0 6764 116 6824
rect 76 6740 116 6764
rect 172 6740 212 7120
rect 1315 7036 1324 7076
rect 1364 7036 2092 7076
rect 2132 7036 2141 7076
rect 1507 6992 1565 6993
rect 1507 6952 1516 6992
rect 1556 6952 1708 6992
rect 1748 6952 1757 6992
rect 1507 6951 1565 6952
rect 355 6908 413 6909
rect 355 6868 364 6908
rect 404 6868 2668 6908
rect 2708 6868 2717 6908
rect 355 6867 413 6868
rect 1699 6784 1708 6824
rect 1748 6784 2380 6824
rect 2420 6784 2429 6824
rect 76 6700 212 6740
rect 1411 6700 1420 6740
rect 1460 6700 2092 6740
rect 2132 6700 2141 6740
rect 1987 6656 2045 6657
rect 3148 6656 3188 7120
rect 4291 7119 4349 7120
rect 6499 7160 6557 7161
rect 7276 7160 7316 7204
rect 7363 7203 7421 7204
rect 8428 7160 8468 7204
rect 8515 7204 8524 7244
rect 8564 7204 8658 7244
rect 8800 7204 12652 7244
rect 12692 7204 12701 7244
rect 15052 7244 15092 7288
rect 15331 7287 15389 7288
rect 15619 7287 15677 7288
rect 15052 7204 15436 7244
rect 15476 7204 15485 7244
rect 19267 7204 19276 7244
rect 19316 7204 19468 7244
rect 19508 7204 19517 7244
rect 8515 7203 8573 7204
rect 8800 7160 8840 7204
rect 12643 7203 12701 7204
rect 8995 7160 9053 7161
rect 14563 7160 14621 7161
rect 19459 7160 19517 7161
rect 19756 7160 19796 7456
rect 20995 7455 21053 7456
rect 21424 7436 21504 7456
rect 21424 7160 21504 7180
rect 6499 7120 6508 7160
rect 6548 7120 7276 7160
rect 7316 7120 7325 7160
rect 7843 7120 7852 7160
rect 7892 7120 8044 7160
rect 8084 7120 8093 7160
rect 8428 7120 8840 7160
rect 8910 7120 9004 7160
rect 9044 7120 9053 7160
rect 12259 7120 12268 7160
rect 12308 7120 12652 7160
rect 12692 7120 12701 7160
rect 13315 7120 13324 7160
rect 13364 7120 13996 7160
rect 14036 7120 14045 7160
rect 14563 7120 14572 7160
rect 14612 7120 16012 7160
rect 16052 7120 16061 7160
rect 16108 7120 16684 7160
rect 16724 7120 18508 7160
rect 18548 7120 18988 7160
rect 19028 7120 19037 7160
rect 19459 7120 19468 7160
rect 19508 7120 19564 7160
rect 19604 7120 19613 7160
rect 19747 7120 19756 7160
rect 19796 7120 19805 7160
rect 21091 7120 21100 7160
rect 21140 7120 21504 7160
rect 6499 7119 6557 7120
rect 8995 7119 9053 7120
rect 14563 7119 14621 7120
rect 7555 7076 7613 7077
rect 11395 7076 11453 7077
rect 16108 7076 16148 7120
rect 19459 7119 19517 7120
rect 21424 7100 21504 7120
rect 5635 7036 5644 7076
rect 5684 7036 6700 7076
rect 6740 7036 6749 7076
rect 7555 7036 7564 7076
rect 7604 7036 10636 7076
rect 10676 7036 10685 7076
rect 11395 7036 11404 7076
rect 11444 7036 11596 7076
rect 11636 7036 12556 7076
rect 12596 7036 12605 7076
rect 13411 7036 13420 7076
rect 13460 7036 13612 7076
rect 13652 7036 13900 7076
rect 13940 7036 14188 7076
rect 14228 7036 14237 7076
rect 15907 7036 15916 7076
rect 15956 7036 16148 7076
rect 16579 7036 16588 7076
rect 16628 7036 20180 7076
rect 7555 7035 7613 7036
rect 11395 7035 11453 7036
rect 8035 6992 8093 6993
rect 3907 6952 3916 6992
rect 3956 6952 7276 6992
rect 7316 6952 7325 6992
rect 7459 6952 7468 6992
rect 7508 6952 8044 6992
rect 8084 6952 8093 6992
rect 8899 6952 8908 6992
rect 8948 6952 12172 6992
rect 12212 6952 12221 6992
rect 15523 6952 15532 6992
rect 15572 6952 17260 6992
rect 17300 6952 17309 6992
rect 8035 6951 8093 6952
rect 20140 6908 20180 7036
rect 3235 6868 3244 6908
rect 3284 6868 8332 6908
rect 8372 6868 8381 6908
rect 10051 6868 10060 6908
rect 10100 6868 14956 6908
rect 14996 6868 15005 6908
rect 20140 6868 20852 6908
rect 16387 6824 16445 6825
rect 20812 6824 20852 6868
rect 21424 6824 21504 6844
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 5356 6784 10156 6824
rect 10196 6784 10205 6824
rect 11203 6784 11212 6824
rect 11252 6784 15860 6824
rect 16302 6784 16396 6824
rect 16436 6784 16445 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 20812 6784 21504 6824
rect 5356 6740 5396 6784
rect 4579 6700 4588 6740
rect 4628 6700 5396 6740
rect 5452 6700 11360 6740
rect 11491 6700 11500 6740
rect 11540 6700 11692 6740
rect 11732 6700 11741 6740
rect 12460 6700 15764 6740
rect 5452 6656 5492 6700
rect 11320 6656 11360 6700
rect 11587 6656 11645 6657
rect 12355 6656 12413 6657
rect 1987 6616 1996 6656
rect 2036 6616 2380 6656
rect 2420 6616 2429 6656
rect 3148 6616 5492 6656
rect 6019 6616 6028 6656
rect 6068 6616 6508 6656
rect 6548 6616 6557 6656
rect 8035 6616 8044 6656
rect 8084 6616 8428 6656
rect 8468 6616 8477 6656
rect 8611 6616 8620 6656
rect 8660 6616 9676 6656
rect 9716 6616 9725 6656
rect 11320 6616 11596 6656
rect 11636 6616 12364 6656
rect 12404 6616 12413 6656
rect 1987 6615 2045 6616
rect 8428 6572 8468 6616
rect 11587 6615 11645 6616
rect 12355 6615 12413 6616
rect 12460 6572 12500 6700
rect 15331 6656 15389 6657
rect 12931 6616 12940 6656
rect 12980 6616 13708 6656
rect 13748 6616 13757 6656
rect 15139 6616 15148 6656
rect 15188 6616 15340 6656
rect 15380 6616 15389 6656
rect 15331 6615 15389 6616
rect 14563 6572 14621 6573
rect 15724 6572 15764 6700
rect 15820 6656 15860 6784
rect 16387 6783 16445 6784
rect 21424 6764 21504 6784
rect 16675 6740 16733 6741
rect 16099 6700 16108 6740
rect 16148 6700 16300 6740
rect 16340 6700 16349 6740
rect 16483 6700 16492 6740
rect 16532 6700 16684 6740
rect 16724 6700 16733 6740
rect 19747 6700 19756 6740
rect 19796 6700 19805 6740
rect 16675 6699 16733 6700
rect 16579 6656 16637 6657
rect 15820 6616 16588 6656
rect 16628 6616 16637 6656
rect 16579 6615 16637 6616
rect 16483 6572 16541 6573
rect 19756 6572 19796 6700
rect 19843 6616 19852 6656
rect 19892 6616 20332 6656
rect 20372 6616 20381 6656
rect 1891 6532 1900 6572
rect 1940 6532 2476 6572
rect 2516 6532 2525 6572
rect 4675 6532 4684 6572
rect 4724 6532 8332 6572
rect 8372 6532 8381 6572
rect 8428 6532 12500 6572
rect 13507 6532 13516 6572
rect 13556 6532 14284 6572
rect 14324 6532 14333 6572
rect 14563 6532 14572 6572
rect 14612 6532 14708 6572
rect 15724 6532 16492 6572
rect 16532 6532 17164 6572
rect 17204 6532 17213 6572
rect 17347 6532 17356 6572
rect 17396 6532 17644 6572
rect 17684 6532 17693 6572
rect 19756 6532 20236 6572
rect 20276 6532 20285 6572
rect 14563 6531 14621 6532
rect 3811 6488 3869 6489
rect 7555 6488 7613 6489
rect 13027 6488 13085 6489
rect 14668 6488 14708 6532
rect 16483 6531 16541 6532
rect 15043 6488 15101 6489
rect 20611 6488 20669 6489
rect 21424 6488 21504 6508
rect 1795 6448 1804 6488
rect 1844 6448 3724 6488
rect 3764 6448 3820 6488
rect 3860 6448 3869 6488
rect 7470 6448 7564 6488
rect 7604 6448 7613 6488
rect 8419 6448 8428 6488
rect 8468 6448 9196 6488
rect 9236 6448 9245 6488
rect 10435 6448 10444 6488
rect 10484 6448 11212 6488
rect 11252 6448 11261 6488
rect 11320 6448 12116 6488
rect 12835 6448 12844 6488
rect 12884 6448 13036 6488
rect 13076 6448 13324 6488
rect 13364 6448 13373 6488
rect 13795 6448 13804 6488
rect 13844 6448 14476 6488
rect 14516 6448 14525 6488
rect 14659 6448 14668 6488
rect 14708 6448 14717 6488
rect 15043 6448 15052 6488
rect 15092 6448 17452 6488
rect 17492 6448 17501 6488
rect 19651 6448 19660 6488
rect 19700 6448 20620 6488
rect 20660 6448 20669 6488
rect 3811 6447 3869 6448
rect 7555 6447 7613 6448
rect 7651 6404 7709 6405
rect 8803 6404 8861 6405
rect 11320 6404 11360 6448
rect 11779 6404 11837 6405
rect 12076 6404 12116 6448
rect 13027 6447 13085 6448
rect 15043 6447 15101 6448
rect 20611 6447 20669 6448
rect 21292 6448 21504 6488
rect 7566 6364 7660 6404
rect 7700 6364 7709 6404
rect 8718 6364 8812 6404
rect 8852 6364 11360 6404
rect 11683 6364 11692 6404
rect 11732 6364 11788 6404
rect 11828 6364 11837 6404
rect 12067 6364 12076 6404
rect 12116 6364 12125 6404
rect 13219 6364 13228 6404
rect 13268 6364 13900 6404
rect 13940 6364 13949 6404
rect 14284 6364 19756 6404
rect 19796 6364 19805 6404
rect 7651 6363 7709 6364
rect 8803 6363 8861 6364
rect 11779 6363 11837 6364
rect 0 6320 80 6340
rect 8515 6320 8573 6321
rect 14284 6320 14324 6364
rect 14851 6320 14909 6321
rect 16579 6320 16637 6321
rect 19555 6320 19613 6321
rect 21292 6320 21332 6448
rect 21424 6428 21504 6448
rect 0 6280 364 6320
rect 404 6280 413 6320
rect 931 6280 940 6320
rect 980 6280 6412 6320
rect 6452 6280 6461 6320
rect 6595 6280 6604 6320
rect 6644 6280 7564 6320
rect 7604 6280 7613 6320
rect 8035 6280 8044 6320
rect 8084 6280 8524 6320
rect 8564 6280 8573 6320
rect 12163 6280 12172 6320
rect 12212 6280 14324 6320
rect 14371 6280 14380 6320
rect 14420 6280 14860 6320
rect 14900 6280 14909 6320
rect 15811 6280 15820 6320
rect 15860 6280 16301 6320
rect 16341 6280 16350 6320
rect 16494 6280 16588 6320
rect 16628 6280 19412 6320
rect 19470 6280 19564 6320
rect 19604 6280 19613 6320
rect 0 6260 80 6280
rect 8515 6279 8573 6280
rect 14851 6279 14909 6280
rect 16579 6279 16637 6280
rect 2563 6236 2621 6237
rect 10339 6236 10397 6237
rect 14179 6236 14237 6237
rect 15715 6236 15773 6237
rect 16099 6236 16157 6237
rect 19372 6236 19412 6280
rect 19555 6279 19613 6280
rect 19660 6280 21332 6320
rect 19660 6236 19700 6280
rect 1411 6196 1420 6236
rect 1460 6196 2188 6236
rect 2228 6196 2237 6236
rect 2563 6196 2572 6236
rect 2612 6196 2668 6236
rect 2708 6196 2717 6236
rect 3043 6196 3052 6236
rect 3092 6196 3436 6236
rect 3476 6196 5548 6236
rect 5588 6196 5597 6236
rect 7363 6196 7372 6236
rect 7412 6196 10060 6236
rect 10100 6196 10348 6236
rect 10388 6196 10397 6236
rect 13411 6196 13420 6236
rect 13460 6196 13708 6236
rect 13748 6196 13757 6236
rect 14179 6196 14188 6236
rect 14228 6196 14284 6236
rect 14324 6196 14333 6236
rect 15715 6196 15724 6236
rect 15764 6196 15916 6236
rect 15956 6196 15965 6236
rect 16099 6196 16108 6236
rect 16148 6196 17452 6236
rect 17492 6196 17501 6236
rect 19372 6196 19700 6236
rect 2563 6195 2621 6196
rect 10339 6195 10397 6196
rect 14179 6195 14237 6196
rect 15715 6195 15773 6196
rect 16099 6195 16157 6196
rect 15907 6152 15965 6153
rect 21424 6152 21504 6172
rect 1891 6112 1900 6152
rect 1940 6112 2956 6152
rect 2996 6112 3005 6152
rect 3235 6112 3244 6152
rect 3284 6112 4148 6152
rect 4483 6112 4492 6152
rect 4532 6112 12364 6152
rect 12404 6112 12413 6152
rect 15907 6112 15916 6152
rect 15956 6112 21504 6152
rect 2371 6068 2429 6069
rect 4108 6068 4148 6112
rect 15907 6111 15965 6112
rect 21424 6092 21504 6112
rect 11971 6068 12029 6069
rect 1603 6028 1612 6068
rect 1652 6028 2092 6068
rect 2132 6028 2380 6068
rect 2420 6028 2429 6068
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 4108 6028 4780 6068
rect 4820 6028 8428 6068
rect 8468 6028 8477 6068
rect 8611 6028 8620 6068
rect 8660 6028 10292 6068
rect 2371 6027 2429 6028
rect 4195 5944 4204 5984
rect 4244 5944 5356 5984
rect 5396 5944 8908 5984
rect 8948 5944 10156 5984
rect 10196 5944 10205 5984
rect 10147 5900 10205 5901
rect 5923 5860 5932 5900
rect 5972 5860 8140 5900
rect 8180 5860 8189 5900
rect 9859 5860 9868 5900
rect 9908 5860 10156 5900
rect 10196 5860 10205 5900
rect 10252 5900 10292 6028
rect 11971 6028 11980 6068
rect 12020 6028 18700 6068
rect 18740 6028 18749 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 11971 6027 12029 6028
rect 10339 5944 10348 5984
rect 10388 5944 19468 5984
rect 19508 5944 19517 5984
rect 10252 5860 12460 5900
rect 12500 5860 12509 5900
rect 13315 5860 13324 5900
rect 13364 5860 13900 5900
rect 13940 5860 14764 5900
rect 14804 5860 14813 5900
rect 15043 5860 15052 5900
rect 15092 5860 15532 5900
rect 15572 5860 15581 5900
rect 10147 5859 10205 5860
rect 0 5816 80 5836
rect 451 5816 509 5817
rect 18883 5816 18941 5817
rect 19267 5816 19325 5817
rect 21424 5816 21504 5836
rect 0 5776 460 5816
rect 500 5776 509 5816
rect 1507 5776 1516 5816
rect 1556 5776 2284 5816
rect 2324 5776 3532 5816
rect 3572 5776 3581 5816
rect 6115 5776 6124 5816
rect 6164 5776 14092 5816
rect 14132 5776 14141 5816
rect 18883 5776 18892 5816
rect 18932 5776 19276 5816
rect 19316 5776 21504 5816
rect 0 5756 80 5776
rect 451 5775 509 5776
rect 18883 5775 18941 5776
rect 19267 5775 19325 5776
rect 21424 5756 21504 5776
rect 5731 5692 5740 5732
rect 5780 5692 7372 5732
rect 7412 5692 7421 5732
rect 8419 5692 8428 5732
rect 8468 5692 13324 5732
rect 13364 5692 13373 5732
rect 13507 5692 13516 5732
rect 13556 5692 14188 5732
rect 14228 5692 14237 5732
rect 16195 5692 16204 5732
rect 16244 5692 17068 5732
rect 17108 5692 17117 5732
rect 10435 5648 10493 5649
rect 11779 5648 11837 5649
rect 1315 5608 1324 5648
rect 1364 5608 2380 5648
rect 2420 5608 2429 5648
rect 2563 5608 2572 5648
rect 2612 5608 8524 5648
rect 8564 5608 8573 5648
rect 10350 5608 10444 5648
rect 10484 5608 11788 5648
rect 11828 5608 11837 5648
rect 11971 5608 11980 5648
rect 12020 5608 13036 5648
rect 13076 5608 13085 5648
rect 13132 5608 15724 5648
rect 15764 5608 15773 5648
rect 16003 5608 16012 5648
rect 16052 5608 16684 5648
rect 16724 5608 17260 5648
rect 17300 5608 17309 5648
rect 18499 5608 18508 5648
rect 18548 5608 18700 5648
rect 18740 5608 18749 5648
rect 10435 5607 10493 5608
rect 11779 5607 11837 5608
rect 7459 5564 7517 5565
rect 12451 5564 12509 5565
rect 13132 5564 13172 5608
rect 2179 5524 2188 5564
rect 2228 5524 6028 5564
rect 6068 5524 6077 5564
rect 7459 5524 7468 5564
rect 7508 5524 12172 5564
rect 12212 5524 12221 5564
rect 12451 5524 12460 5564
rect 12500 5524 13172 5564
rect 15427 5524 15436 5564
rect 15476 5524 16204 5564
rect 16244 5524 16253 5564
rect 7459 5523 7517 5524
rect 12451 5523 12509 5524
rect 1795 5480 1853 5481
rect 10243 5480 10301 5481
rect 12067 5480 12125 5481
rect 21424 5480 21504 5500
rect 1795 5440 1804 5480
rect 1844 5440 1900 5480
rect 1940 5440 1949 5480
rect 4195 5440 4204 5480
rect 4244 5440 10252 5480
rect 10292 5440 10301 5480
rect 11683 5440 11692 5480
rect 11732 5440 12076 5480
rect 12116 5440 12844 5480
rect 12884 5440 12893 5480
rect 13411 5440 13420 5480
rect 13460 5440 13804 5480
rect 13844 5440 13853 5480
rect 15811 5440 15820 5480
rect 15860 5440 19852 5480
rect 19892 5440 19901 5480
rect 20140 5440 21504 5480
rect 1795 5439 1853 5440
rect 10243 5439 10301 5440
rect 12067 5439 12125 5440
rect 8803 5396 8861 5397
rect 10915 5396 10973 5397
rect 17059 5396 17117 5397
rect 20140 5396 20180 5440
rect 21424 5420 21504 5440
rect 1219 5356 1228 5396
rect 1268 5356 8812 5396
rect 8852 5356 8861 5396
rect 10339 5356 10348 5396
rect 10388 5356 10924 5396
rect 10964 5356 10973 5396
rect 12451 5356 12460 5396
rect 12500 5356 13132 5396
rect 13172 5356 13516 5396
rect 13556 5356 13565 5396
rect 13699 5356 13708 5396
rect 13748 5356 17068 5396
rect 17108 5356 20180 5396
rect 8803 5355 8861 5356
rect 10915 5355 10973 5356
rect 17059 5355 17117 5356
rect 0 5312 80 5332
rect 163 5312 221 5313
rect 18883 5312 18941 5313
rect 0 5272 172 5312
rect 212 5272 221 5312
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 6307 5272 6316 5312
rect 6356 5272 9484 5312
rect 9524 5272 9533 5312
rect 10435 5272 10444 5312
rect 10484 5272 15916 5312
rect 15956 5272 15965 5312
rect 16300 5272 18892 5312
rect 18932 5272 18941 5312
rect 19171 5272 19180 5312
rect 19220 5272 19660 5312
rect 19700 5272 19709 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 0 5252 80 5272
rect 163 5271 221 5272
rect 2179 5228 2237 5229
rect 7459 5228 7517 5229
rect 13891 5228 13949 5229
rect 2083 5188 2092 5228
rect 2132 5188 2188 5228
rect 2228 5188 2237 5228
rect 7363 5188 7372 5228
rect 7412 5188 7468 5228
rect 7508 5188 7517 5228
rect 9667 5188 9676 5228
rect 9716 5188 11308 5228
rect 11348 5188 11357 5228
rect 12355 5188 12364 5228
rect 12404 5188 12652 5228
rect 12692 5188 12701 5228
rect 13806 5188 13900 5228
rect 13940 5188 13949 5228
rect 2179 5187 2237 5188
rect 7459 5187 7517 5188
rect 13891 5187 13949 5188
rect 16300 5144 16340 5272
rect 18883 5271 18941 5272
rect 16579 5188 16588 5228
rect 16628 5188 21004 5228
rect 21044 5188 21053 5228
rect 1411 5104 1420 5144
rect 1460 5104 5836 5144
rect 5876 5104 7180 5144
rect 7220 5104 7229 5144
rect 7939 5104 7948 5144
rect 7988 5104 8236 5144
rect 8276 5104 8285 5144
rect 9379 5104 9388 5144
rect 9428 5104 10924 5144
rect 10964 5104 10973 5144
rect 11212 5104 16340 5144
rect 16483 5144 16541 5145
rect 21424 5144 21504 5164
rect 16483 5104 16492 5144
rect 16532 5104 16626 5144
rect 20140 5104 21504 5144
rect 1411 5060 1469 5061
rect 7459 5060 7517 5061
rect 1411 5020 1420 5060
rect 1460 5020 1996 5060
rect 2036 5020 2045 5060
rect 6883 5020 6892 5060
rect 6932 5020 7468 5060
rect 7508 5020 7517 5060
rect 1411 5019 1469 5020
rect 7459 5019 7517 5020
rect 9676 5020 10484 5060
rect 10531 5020 10540 5060
rect 10580 5020 11116 5060
rect 11156 5020 11165 5060
rect 8419 4976 8477 4977
rect 8707 4976 8765 4977
rect 9571 4976 9629 4977
rect 3139 4936 3148 4976
rect 3188 4936 4492 4976
rect 4532 4936 5932 4976
rect 5972 4936 6124 4976
rect 6164 4936 6173 4976
rect 6787 4936 6796 4976
rect 6836 4936 7756 4976
rect 7796 4936 7805 4976
rect 8419 4936 8428 4976
rect 8468 4936 8716 4976
rect 8756 4936 9004 4976
rect 9044 4936 9053 4976
rect 9486 4936 9580 4976
rect 9620 4936 9629 4976
rect 8419 4935 8477 4936
rect 8707 4935 8765 4936
rect 9571 4935 9629 4936
rect 9676 4892 9716 5020
rect 9955 4976 10013 4977
rect 9870 4936 9964 4976
rect 10004 4936 10013 4976
rect 10444 4976 10484 5020
rect 11212 4976 11252 5104
rect 16483 5103 16541 5104
rect 20140 5060 20180 5104
rect 21424 5084 21504 5104
rect 14179 5020 14188 5060
rect 14228 5020 14860 5060
rect 14900 5020 14909 5060
rect 16291 5020 16300 5060
rect 16340 5020 17452 5060
rect 17492 5020 17501 5060
rect 18508 5020 18796 5060
rect 18836 5020 18845 5060
rect 19267 5020 19276 5060
rect 19316 5020 19756 5060
rect 19796 5020 20180 5060
rect 12163 4976 12221 4977
rect 10444 4936 11252 4976
rect 11875 4936 11884 4976
rect 11924 4936 12172 4976
rect 12212 4936 12221 4976
rect 9955 4935 10013 4936
rect 12163 4935 12221 4936
rect 12355 4976 12413 4977
rect 15235 4976 15293 4977
rect 18508 4976 18548 5020
rect 12355 4936 12364 4976
rect 12404 4936 12498 4976
rect 12643 4936 12652 4976
rect 12692 4936 12844 4976
rect 12884 4936 13324 4976
rect 13364 4936 13373 4976
rect 13987 4936 13996 4976
rect 14036 4936 14476 4976
rect 14516 4936 14525 4976
rect 15235 4936 15244 4976
rect 15284 4936 16108 4976
rect 16148 4936 16492 4976
rect 16532 4936 17660 4976
rect 18307 4936 18316 4976
rect 18356 4936 18508 4976
rect 18548 4936 18557 4976
rect 18691 4936 18700 4976
rect 18740 4936 19084 4976
rect 19124 4936 19948 4976
rect 19988 4936 19997 4976
rect 12355 4935 12413 4936
rect 15235 4935 15293 4936
rect 17620 4892 17660 4936
rect 21283 4892 21341 4893
rect 835 4852 844 4892
rect 884 4852 4972 4892
rect 5012 4852 5644 4892
rect 5684 4852 6508 4892
rect 6548 4852 6557 4892
rect 6979 4852 6988 4892
rect 7028 4852 8332 4892
rect 8372 4852 8381 4892
rect 9187 4852 9196 4892
rect 9236 4852 9484 4892
rect 9524 4852 9716 4892
rect 11299 4852 11308 4892
rect 11348 4852 11500 4892
rect 11540 4852 12460 4892
rect 12500 4852 12509 4892
rect 12739 4852 12748 4892
rect 12788 4852 13612 4892
rect 13652 4852 13661 4892
rect 17620 4852 20716 4892
rect 20756 4852 20765 4892
rect 20812 4852 21292 4892
rect 21332 4852 21341 4892
rect 0 4808 80 4828
rect 18403 4808 18461 4809
rect 20812 4808 20852 4852
rect 21283 4851 21341 4852
rect 21424 4808 21504 4828
rect 0 4768 748 4808
rect 788 4768 797 4808
rect 1219 4768 1228 4808
rect 1268 4768 7756 4808
rect 7796 4768 7805 4808
rect 11971 4768 11980 4808
rect 12020 4768 12556 4808
rect 12596 4768 12605 4808
rect 13507 4768 13516 4808
rect 13556 4768 18412 4808
rect 18452 4768 18461 4808
rect 20035 4768 20044 4808
rect 20084 4768 20852 4808
rect 21100 4768 21504 4808
rect 0 4748 80 4768
rect 18403 4767 18461 4768
rect 2275 4724 2333 4725
rect 4963 4724 5021 4725
rect 17539 4724 17597 4725
rect 21100 4724 21140 4768
rect 21424 4748 21504 4768
rect 2275 4684 2284 4724
rect 2324 4684 2860 4724
rect 2900 4684 3244 4724
rect 3284 4684 3293 4724
rect 4867 4684 4876 4724
rect 4916 4684 4972 4724
rect 5012 4684 5021 4724
rect 2275 4683 2333 4684
rect 4963 4683 5021 4684
rect 6124 4684 12076 4724
rect 12116 4684 12125 4724
rect 12355 4684 12364 4724
rect 12404 4684 13132 4724
rect 13172 4684 13181 4724
rect 13795 4684 13804 4724
rect 13844 4684 17164 4724
rect 17204 4684 17213 4724
rect 17539 4684 17548 4724
rect 17588 4684 21140 4724
rect 5539 4640 5597 4641
rect 6124 4640 6164 4684
rect 17539 4683 17597 4684
rect 9283 4640 9341 4641
rect 10723 4640 10781 4641
rect 1603 4600 1612 4640
rect 1652 4600 5548 4640
rect 5588 4600 6164 4640
rect 9198 4600 9292 4640
rect 9332 4600 9772 4640
rect 9812 4600 10732 4640
rect 10772 4600 10781 4640
rect 5539 4599 5597 4600
rect 9283 4599 9341 4600
rect 10723 4599 10781 4600
rect 10924 4600 18412 4640
rect 18452 4600 18461 4640
rect 10924 4556 10964 4600
rect 12451 4556 12509 4557
rect 17731 4556 17789 4557
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 5347 4516 5356 4556
rect 5396 4516 7948 4556
rect 7988 4516 10196 4556
rect 10915 4516 10924 4556
rect 10964 4516 10973 4556
rect 11395 4516 11404 4556
rect 11444 4516 11692 4556
rect 11732 4516 11741 4556
rect 12366 4516 12460 4556
rect 12500 4516 12509 4556
rect 17539 4516 17548 4556
rect 17588 4516 17740 4556
rect 17780 4516 17789 4556
rect 18211 4516 18220 4556
rect 18260 4516 18269 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 67 4472 125 4473
rect 10156 4472 10196 4516
rect 12451 4515 12509 4516
rect 17731 4515 17789 4516
rect 18220 4472 18260 4516
rect 20131 4472 20189 4473
rect 21424 4472 21504 4492
rect 67 4432 76 4472
rect 116 4432 1804 4472
rect 1844 4432 1853 4472
rect 3427 4432 3436 4472
rect 3476 4432 10060 4472
rect 10100 4432 10109 4472
rect 10156 4432 14092 4472
rect 14132 4432 14141 4472
rect 15907 4432 15916 4472
rect 15956 4432 18836 4472
rect 19555 4432 19564 4472
rect 19604 4432 19613 4472
rect 20131 4432 20140 4472
rect 20180 4432 21504 4472
rect 67 4431 125 4432
rect 17827 4388 17885 4389
rect 18796 4388 18836 4432
rect 19564 4388 19604 4432
rect 20131 4431 20189 4432
rect 21424 4412 21504 4432
rect 1699 4348 1708 4388
rect 1748 4348 4588 4388
rect 4628 4348 4637 4388
rect 4771 4348 4780 4388
rect 4820 4348 6836 4388
rect 6979 4348 6988 4388
rect 7028 4348 13132 4388
rect 13172 4348 13181 4388
rect 17827 4348 17836 4388
rect 17876 4348 18220 4388
rect 18260 4348 18269 4388
rect 18787 4348 18796 4388
rect 18836 4348 18845 4388
rect 19075 4348 19084 4388
rect 19124 4348 19604 4388
rect 0 4304 80 4324
rect 5731 4304 5789 4305
rect 6115 4304 6173 4305
rect 6796 4304 6836 4348
rect 17827 4347 17885 4348
rect 8227 4304 8285 4305
rect 8995 4304 9053 4305
rect 16675 4304 16733 4305
rect 0 4264 268 4304
rect 308 4264 317 4304
rect 5731 4264 5740 4304
rect 5780 4264 5932 4304
rect 5972 4264 6124 4304
rect 6164 4264 6220 4304
rect 6260 4264 6269 4304
rect 6796 4264 7660 4304
rect 7700 4264 8236 4304
rect 8276 4264 8285 4304
rect 8899 4264 8908 4304
rect 8948 4264 9004 4304
rect 9044 4264 9053 4304
rect 9571 4264 9580 4304
rect 9620 4264 9629 4304
rect 10060 4264 10828 4304
rect 10868 4264 11308 4304
rect 11348 4264 12844 4304
rect 12884 4264 12893 4304
rect 15811 4264 15820 4304
rect 15860 4264 16684 4304
rect 16724 4264 17068 4304
rect 17108 4264 17117 4304
rect 17635 4264 17644 4304
rect 17684 4264 18508 4304
rect 18548 4264 19564 4304
rect 19604 4264 19613 4304
rect 0 4244 80 4264
rect 5731 4263 5789 4264
rect 6115 4263 6173 4264
rect 4579 4220 4637 4221
rect 4771 4220 4829 4221
rect 1219 4180 1228 4220
rect 1268 4180 2284 4220
rect 2324 4180 4588 4220
rect 4628 4180 4637 4220
rect 4686 4180 4780 4220
rect 4820 4180 4829 4220
rect 6220 4220 6260 4264
rect 8227 4263 8285 4264
rect 8995 4263 9053 4264
rect 9580 4220 9620 4264
rect 6220 4180 9620 4220
rect 4579 4179 4637 4180
rect 4771 4179 4829 4180
rect 4099 4136 4157 4137
rect 2179 4096 2188 4136
rect 2228 4096 4108 4136
rect 4148 4096 4157 4136
rect 4099 4095 4157 4096
rect 4291 4136 4349 4137
rect 8707 4136 8765 4137
rect 10060 4136 10100 4264
rect 16675 4263 16733 4264
rect 11587 4220 11645 4221
rect 17059 4220 17117 4221
rect 21091 4220 21149 4221
rect 10828 4180 11212 4220
rect 11252 4180 11261 4220
rect 11502 4180 11596 4220
rect 11636 4180 11645 4220
rect 13987 4180 13996 4220
rect 14036 4180 14188 4220
rect 14228 4180 14237 4220
rect 17059 4180 17068 4220
rect 17108 4180 20122 4220
rect 20162 4180 21100 4220
rect 21140 4180 21149 4220
rect 4291 4096 4300 4136
rect 4340 4096 4434 4136
rect 4579 4096 4588 4136
rect 4628 4096 5356 4136
rect 5396 4096 5405 4136
rect 7075 4096 7084 4136
rect 7124 4096 8716 4136
rect 8756 4096 8765 4136
rect 8995 4096 9004 4136
rect 9044 4096 10100 4136
rect 10147 4096 10156 4136
rect 10196 4096 10205 4136
rect 4291 4095 4349 4096
rect 8707 4095 8765 4096
rect 1123 4012 1132 4052
rect 1172 4012 3820 4052
rect 3860 4012 3869 4052
rect 1891 3968 1949 3969
rect 6691 3968 6749 3969
rect 931 3928 940 3968
rect 980 3928 1228 3968
rect 1268 3928 1277 3968
rect 1891 3928 1900 3968
rect 1940 3928 1996 3968
rect 2036 3928 2045 3968
rect 6606 3928 6700 3968
rect 6740 3928 6749 3968
rect 1891 3927 1949 3928
rect 6691 3927 6749 3928
rect 7363 3884 7421 3885
rect 9667 3884 9725 3885
rect 1612 3844 2188 3884
rect 2228 3844 2237 3884
rect 4387 3844 4396 3884
rect 4436 3844 7220 3884
rect 0 3800 80 3820
rect 547 3800 605 3801
rect 1507 3800 1565 3801
rect 0 3760 556 3800
rect 596 3760 605 3800
rect 1422 3760 1516 3800
rect 1556 3760 1565 3800
rect 0 3740 80 3760
rect 547 3759 605 3760
rect 1507 3759 1565 3760
rect 1612 3716 1652 3844
rect 1699 3760 1708 3800
rect 1748 3760 3628 3800
rect 3668 3760 3677 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 5923 3760 5932 3800
rect 5972 3760 6412 3800
rect 6452 3760 6461 3800
rect 2467 3716 2525 3717
rect 7180 3716 7220 3844
rect 7363 3844 7372 3884
rect 7412 3844 7506 3884
rect 8332 3844 8620 3884
rect 8660 3844 8669 3884
rect 9582 3844 9676 3884
rect 9716 3844 9725 3884
rect 7363 3843 7421 3844
rect 8332 3800 8372 3844
rect 9667 3843 9725 3844
rect 10156 3800 10196 4096
rect 10828 4052 10868 4180
rect 11587 4179 11645 4180
rect 17059 4179 17117 4180
rect 21091 4179 21149 4180
rect 15235 4136 15293 4137
rect 19939 4136 19997 4137
rect 21424 4136 21504 4156
rect 10915 4096 10924 4136
rect 10964 4096 10973 4136
rect 11395 4096 11404 4136
rect 11444 4096 11884 4136
rect 11924 4096 11933 4136
rect 12067 4096 12076 4136
rect 12116 4096 15244 4136
rect 15284 4096 15293 4136
rect 15715 4096 15724 4136
rect 15764 4096 16012 4136
rect 16052 4096 16780 4136
rect 16820 4096 16829 4136
rect 17347 4096 17356 4136
rect 17396 4096 17932 4136
rect 17972 4096 17981 4136
rect 19854 4096 19948 4136
rect 19988 4096 19997 4136
rect 10924 4052 10964 4096
rect 15235 4095 15293 4096
rect 19939 4095 19997 4096
rect 20140 4096 21504 4136
rect 20140 4052 20180 4096
rect 21424 4076 21504 4096
rect 10819 4012 10828 4052
rect 10868 4012 10877 4052
rect 10924 4012 11692 4052
rect 11732 4012 17644 4052
rect 17684 4012 17693 4052
rect 19267 4012 19276 4052
rect 19316 4012 20180 4052
rect 11203 3928 11212 3968
rect 11252 3928 11596 3968
rect 11636 3928 11645 3968
rect 11971 3928 11980 3968
rect 12020 3928 15628 3968
rect 15668 3928 15677 3968
rect 19363 3928 19372 3968
rect 19412 3928 20812 3968
rect 20852 3928 20861 3968
rect 19555 3884 19613 3885
rect 10723 3844 10732 3884
rect 10772 3844 19084 3884
rect 19124 3844 19564 3884
rect 19604 3844 19613 3884
rect 19555 3843 19613 3844
rect 21424 3800 21504 3820
rect 7939 3760 7948 3800
rect 7988 3760 8372 3800
rect 8419 3760 8428 3800
rect 8468 3760 10196 3800
rect 10339 3760 10348 3800
rect 10388 3760 11692 3800
rect 11732 3760 12076 3800
rect 12116 3760 12125 3800
rect 13123 3760 13132 3800
rect 13172 3760 13324 3800
rect 13364 3760 14476 3800
rect 14516 3760 16492 3800
rect 16532 3760 16541 3800
rect 17059 3760 17068 3800
rect 17108 3760 17836 3800
rect 17876 3760 17885 3800
rect 18211 3760 18220 3800
rect 18260 3760 18269 3800
rect 18403 3760 18412 3800
rect 18452 3760 19468 3800
rect 19508 3760 19517 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 20707 3760 20716 3800
rect 20756 3760 21504 3800
rect 17155 3716 17213 3717
rect 1603 3676 1612 3716
rect 1652 3676 1661 3716
rect 2467 3676 2476 3716
rect 2516 3676 5452 3716
rect 5492 3676 5501 3716
rect 6307 3676 6316 3716
rect 6356 3676 6836 3716
rect 7180 3676 13612 3716
rect 13652 3676 13661 3716
rect 13891 3676 13900 3716
rect 13940 3676 16396 3716
rect 16436 3676 17164 3716
rect 17204 3676 17213 3716
rect 18220 3716 18260 3760
rect 21424 3740 21504 3760
rect 18220 3676 20084 3716
rect 2467 3675 2525 3676
rect 1411 3632 1469 3633
rect 1326 3592 1420 3632
rect 1460 3592 1469 3632
rect 1411 3591 1469 3592
rect 1603 3632 1661 3633
rect 3235 3632 3293 3633
rect 6796 3632 6836 3676
rect 17155 3675 17213 3676
rect 7555 3632 7613 3633
rect 15715 3632 15773 3633
rect 16387 3632 16445 3633
rect 17251 3632 17309 3633
rect 1603 3592 1612 3632
rect 1652 3592 1900 3632
rect 1940 3592 1949 3632
rect 3235 3592 3244 3632
rect 3284 3592 3340 3632
rect 3380 3592 3389 3632
rect 3523 3592 3532 3632
rect 3572 3592 3724 3632
rect 3764 3592 3773 3632
rect 4483 3592 4492 3632
rect 4532 3592 4972 3632
rect 5012 3592 5021 3632
rect 6787 3592 6796 3632
rect 6836 3592 6845 3632
rect 7555 3592 7564 3632
rect 7604 3592 15148 3632
rect 15188 3592 15197 3632
rect 15523 3592 15532 3632
rect 15572 3592 15724 3632
rect 15764 3592 16204 3632
rect 16244 3592 16253 3632
rect 16387 3592 16396 3632
rect 16436 3592 16588 3632
rect 16628 3592 16637 3632
rect 17166 3592 17260 3632
rect 17300 3592 17309 3632
rect 17539 3592 17548 3632
rect 17588 3592 17597 3632
rect 17731 3592 17740 3632
rect 17780 3592 19948 3632
rect 19988 3592 19997 3632
rect 1603 3591 1661 3592
rect 3235 3591 3293 3592
rect 7555 3591 7613 3592
rect 15715 3591 15773 3592
rect 16387 3591 16445 3592
rect 17251 3591 17309 3592
rect 14947 3548 15005 3549
rect 17548 3548 17588 3592
rect 20044 3548 20084 3676
rect 4099 3508 4108 3548
rect 4148 3508 6316 3548
rect 6356 3508 6365 3548
rect 9196 3508 14956 3548
rect 14996 3508 15005 3548
rect 15619 3508 15628 3548
rect 15668 3508 15820 3548
rect 15860 3508 15869 3548
rect 16675 3508 16684 3548
rect 16724 3508 16972 3548
rect 17012 3508 18356 3548
rect 20035 3508 20044 3548
rect 20084 3508 20093 3548
rect 8035 3464 8093 3465
rect 9196 3464 9236 3508
rect 14947 3507 15005 3508
rect 10147 3464 10205 3465
rect 3715 3424 3724 3464
rect 3764 3424 5740 3464
rect 5780 3424 5789 3464
rect 7950 3424 8044 3464
rect 8084 3424 8093 3464
rect 9187 3424 9196 3464
rect 9236 3424 9245 3464
rect 10062 3424 10156 3464
rect 10196 3424 10205 3464
rect 8035 3423 8093 3424
rect 10147 3423 10205 3424
rect 10339 3464 10397 3465
rect 12643 3464 12701 3465
rect 10339 3424 10348 3464
rect 10388 3424 10482 3464
rect 11779 3424 11788 3464
rect 11828 3424 12076 3464
rect 12116 3424 12125 3464
rect 12643 3424 12652 3464
rect 12692 3424 13516 3464
rect 13556 3424 13565 3464
rect 13987 3424 13996 3464
rect 14036 3424 18220 3464
rect 18260 3424 18269 3464
rect 10339 3423 10397 3424
rect 12643 3423 12701 3424
rect 6691 3380 6749 3381
rect 9763 3380 9821 3381
rect 10723 3380 10781 3381
rect 3427 3340 3436 3380
rect 3476 3340 4012 3380
rect 4052 3340 4492 3380
rect 4532 3340 6124 3380
rect 6164 3340 6700 3380
rect 6740 3340 9004 3380
rect 9044 3340 9053 3380
rect 9678 3340 9772 3380
rect 9812 3340 9821 3380
rect 10638 3340 10732 3380
rect 10772 3340 10781 3380
rect 6691 3339 6749 3340
rect 9763 3339 9821 3340
rect 10723 3339 10781 3340
rect 12163 3380 12221 3381
rect 18316 3380 18356 3508
rect 20515 3464 20573 3465
rect 19267 3424 19276 3464
rect 19316 3424 20524 3464
rect 20564 3424 20573 3464
rect 20515 3423 20573 3424
rect 20803 3464 20861 3465
rect 21424 3464 21504 3484
rect 20803 3424 20812 3464
rect 20852 3424 21504 3464
rect 20803 3423 20861 3424
rect 21424 3404 21504 3424
rect 12163 3340 12172 3380
rect 12212 3340 12268 3380
rect 12308 3340 13228 3380
rect 13268 3340 13277 3380
rect 15043 3340 15052 3380
rect 15092 3340 18028 3380
rect 18068 3340 18077 3380
rect 18316 3340 19796 3380
rect 12163 3339 12221 3340
rect 0 3296 80 3316
rect 6883 3296 6941 3297
rect 14947 3296 15005 3297
rect 15619 3296 15677 3297
rect 18595 3296 18653 3297
rect 19555 3296 19613 3297
rect 19756 3296 19796 3340
rect 19939 3296 19997 3297
rect 0 3256 172 3296
rect 212 3256 221 3296
rect 3043 3256 3052 3296
rect 3092 3256 6412 3296
rect 6452 3256 6461 3296
rect 6883 3256 6892 3296
rect 6932 3256 14956 3296
rect 14996 3256 15005 3296
rect 15139 3256 15148 3296
rect 15188 3256 15436 3296
rect 15476 3256 15485 3296
rect 15619 3256 15628 3296
rect 15668 3256 16436 3296
rect 16483 3256 16492 3296
rect 16532 3256 17260 3296
rect 17300 3256 17309 3296
rect 17731 3256 17740 3296
rect 17780 3256 18412 3296
rect 18452 3256 18461 3296
rect 18595 3256 18604 3296
rect 18644 3256 18796 3296
rect 18836 3256 18845 3296
rect 19470 3256 19564 3296
rect 19604 3256 19613 3296
rect 19747 3256 19756 3296
rect 19796 3256 19948 3296
rect 19988 3256 19997 3296
rect 0 3236 80 3256
rect 6883 3255 6941 3256
rect 14947 3255 15005 3256
rect 15619 3255 15677 3256
rect 2179 3212 2237 3213
rect 12547 3212 12605 3213
rect 16396 3212 16436 3256
rect 18595 3255 18653 3256
rect 19555 3255 19613 3256
rect 19939 3255 19997 3256
rect 17443 3212 17501 3213
rect 2083 3172 2092 3212
rect 2132 3172 2188 3212
rect 2228 3172 2237 3212
rect 3331 3172 3340 3212
rect 3380 3172 4684 3212
rect 4724 3172 4733 3212
rect 4963 3172 4972 3212
rect 5012 3172 7948 3212
rect 7988 3172 7997 3212
rect 11779 3172 11788 3212
rect 11828 3172 12172 3212
rect 12212 3172 12221 3212
rect 12547 3172 12556 3212
rect 12596 3172 15724 3212
rect 15764 3172 15773 3212
rect 16396 3172 17452 3212
rect 17492 3172 18068 3212
rect 18115 3172 18124 3212
rect 18164 3172 20129 3212
rect 20169 3172 20178 3212
rect 2179 3171 2237 3172
rect 12547 3171 12605 3172
rect 17443 3171 17501 3172
rect 15235 3128 15293 3129
rect 18028 3128 18068 3172
rect 19747 3128 19805 3129
rect 21424 3128 21504 3148
rect 2467 3088 2476 3128
rect 2516 3088 4204 3128
rect 4244 3088 4253 3128
rect 4300 3088 7852 3128
rect 7892 3088 7901 3128
rect 15235 3088 15244 3128
rect 15284 3088 16876 3128
rect 16916 3088 16925 3128
rect 18028 3088 19316 3128
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 4300 2960 4340 3088
rect 7852 3044 7892 3088
rect 15235 3087 15293 3088
rect 19276 3044 19316 3088
rect 19747 3088 19756 3128
rect 19796 3088 21504 3128
rect 19747 3087 19805 3088
rect 21424 3068 21504 3088
rect 6211 3004 6220 3044
rect 6260 3004 7468 3044
rect 7508 3004 7796 3044
rect 7852 3004 13460 3044
rect 13507 3004 13516 3044
rect 13556 3004 17548 3044
rect 17588 3004 17597 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 19276 3004 20180 3044
rect 7651 2960 7709 2961
rect 3235 2920 3244 2960
rect 3284 2920 3436 2960
rect 3476 2920 4340 2960
rect 7363 2920 7372 2960
rect 7412 2920 7660 2960
rect 7700 2920 7709 2960
rect 7756 2960 7796 3004
rect 13420 2960 13460 3004
rect 7756 2920 12748 2960
rect 12788 2920 12797 2960
rect 13420 2920 14284 2960
rect 14324 2920 15340 2960
rect 15380 2920 15916 2960
rect 15956 2920 15965 2960
rect 18019 2920 18028 2960
rect 18068 2920 19660 2960
rect 19700 2920 19709 2960
rect 7651 2919 7709 2920
rect 10915 2876 10973 2877
rect 17251 2876 17309 2877
rect 1228 2836 1516 2876
rect 1556 2836 1565 2876
rect 3532 2836 4972 2876
rect 5012 2836 5021 2876
rect 5068 2836 10636 2876
rect 10676 2836 10685 2876
rect 10915 2836 10924 2876
rect 10964 2836 11596 2876
rect 11636 2836 16300 2876
rect 16340 2836 16349 2876
rect 17251 2836 17260 2876
rect 17300 2836 19852 2876
rect 19892 2836 19901 2876
rect 0 2792 80 2812
rect 1228 2792 1268 2836
rect 0 2752 1268 2792
rect 1315 2752 1324 2792
rect 1364 2752 1612 2792
rect 1652 2752 1661 2792
rect 0 2732 80 2752
rect 3532 2708 3572 2836
rect 5068 2792 5108 2836
rect 10915 2835 10973 2836
rect 17251 2835 17309 2836
rect 5923 2792 5981 2793
rect 9091 2792 9149 2793
rect 11779 2792 11837 2793
rect 20140 2792 20180 3004
rect 21424 2792 21504 2812
rect 5059 2752 5068 2792
rect 5108 2752 5117 2792
rect 5635 2752 5644 2792
rect 5684 2752 5932 2792
rect 5972 2752 5981 2792
rect 6115 2752 6124 2792
rect 6164 2752 7756 2792
rect 7796 2752 7805 2792
rect 9091 2752 9100 2792
rect 9140 2752 9292 2792
rect 9332 2752 10732 2792
rect 10772 2752 11212 2792
rect 11252 2752 11261 2792
rect 11779 2752 11788 2792
rect 11828 2752 13900 2792
rect 13940 2752 14956 2792
rect 14996 2752 15005 2792
rect 15139 2752 15148 2792
rect 15188 2752 17548 2792
rect 17588 2752 17932 2792
rect 17972 2752 17981 2792
rect 20140 2752 21504 2792
rect 5923 2751 5981 2752
rect 9091 2751 9149 2752
rect 11779 2751 11837 2752
rect 21424 2732 21504 2752
rect 16195 2708 16253 2709
rect 3523 2668 3532 2708
rect 3572 2668 3581 2708
rect 4771 2668 4780 2708
rect 4820 2668 8428 2708
rect 8468 2668 8477 2708
rect 9868 2668 12116 2708
rect 12163 2668 12172 2708
rect 12212 2668 12460 2708
rect 12500 2668 12509 2708
rect 13699 2668 13708 2708
rect 13748 2668 16204 2708
rect 16244 2668 16780 2708
rect 16820 2668 16829 2708
rect 9868 2625 9908 2668
rect 2659 2624 2717 2625
rect 6307 2624 6365 2625
rect 2179 2584 2188 2624
rect 2228 2584 2668 2624
rect 2708 2584 2717 2624
rect 3619 2584 3628 2624
rect 3668 2584 5548 2624
rect 5588 2584 5932 2624
rect 5972 2584 5981 2624
rect 6222 2584 6316 2624
rect 6356 2584 6365 2624
rect 2659 2583 2717 2584
rect 6307 2583 6365 2584
rect 6883 2624 6941 2625
rect 9859 2624 9917 2625
rect 12076 2624 12116 2668
rect 16195 2667 16253 2668
rect 17059 2624 17117 2625
rect 17539 2624 17597 2625
rect 6883 2584 6892 2624
rect 6932 2584 6988 2624
rect 7028 2584 7037 2624
rect 8131 2584 8140 2624
rect 8180 2584 8756 2624
rect 9763 2584 9772 2624
rect 9812 2584 9868 2624
rect 9908 2584 9917 2624
rect 6883 2583 6941 2584
rect 5827 2540 5885 2541
rect 6499 2540 6557 2541
rect 7555 2540 7613 2541
rect 8716 2540 8756 2584
rect 9859 2583 9917 2584
rect 11212 2584 11500 2624
rect 11540 2584 11549 2624
rect 12076 2584 12652 2624
rect 12692 2584 16012 2624
rect 16052 2584 16061 2624
rect 17059 2584 17068 2624
rect 17108 2584 17492 2624
rect 11212 2540 11252 2584
rect 17059 2583 17117 2584
rect 17452 2540 17492 2584
rect 17539 2584 17548 2624
rect 17588 2584 18028 2624
rect 18068 2584 18077 2624
rect 17539 2583 17597 2584
rect 20131 2540 20189 2541
rect 5220 2500 5260 2540
rect 5300 2500 5309 2540
rect 5742 2500 5836 2540
rect 5876 2500 5885 2540
rect 6019 2500 6028 2540
rect 6068 2500 6508 2540
rect 6548 2500 6557 2540
rect 7470 2500 7564 2540
rect 7604 2500 7613 2540
rect 8580 2500 8620 2540
rect 8660 2500 8669 2540
rect 8712 2500 8721 2540
rect 8761 2500 8770 2540
rect 9924 2500 9964 2540
rect 10004 2500 10013 2540
rect 10819 2500 10828 2540
rect 10868 2500 11020 2540
rect 11060 2500 11069 2540
rect 11203 2500 11212 2540
rect 11252 2500 11261 2540
rect 11320 2500 11444 2540
rect 16099 2500 16108 2540
rect 16148 2500 16300 2540
rect 16340 2500 16349 2540
rect 17124 2500 17164 2540
rect 17204 2500 17213 2540
rect 17452 2500 17548 2540
rect 17588 2500 17597 2540
rect 18084 2500 18124 2540
rect 18164 2500 18173 2540
rect 20131 2500 20140 2540
rect 20180 2500 20274 2540
rect 5260 2456 5300 2500
rect 5827 2499 5885 2500
rect 6499 2499 6557 2500
rect 7555 2499 7613 2500
rect 5923 2456 5981 2457
rect 8620 2456 8660 2500
rect 9964 2456 10004 2500
rect 3139 2416 3148 2456
rect 3188 2416 3436 2456
rect 3476 2416 3485 2456
rect 4579 2416 4588 2456
rect 4628 2416 5164 2456
rect 5204 2416 5213 2456
rect 5260 2416 5452 2456
rect 5492 2416 5501 2456
rect 5923 2416 5932 2456
rect 5972 2416 7852 2456
rect 7892 2416 7901 2456
rect 8620 2416 10004 2456
rect 10243 2456 10301 2457
rect 11320 2456 11360 2500
rect 10243 2416 10252 2456
rect 10292 2416 11360 2456
rect 11404 2456 11444 2500
rect 16771 2456 16829 2457
rect 11404 2416 13420 2456
rect 13460 2416 16780 2456
rect 16820 2416 16829 2456
rect 17164 2456 17204 2500
rect 18124 2456 18164 2500
rect 20131 2499 20189 2500
rect 17164 2416 18164 2456
rect 18403 2456 18461 2457
rect 21424 2456 21504 2476
rect 18403 2416 18412 2456
rect 18452 2416 19948 2456
rect 19988 2416 19997 2456
rect 20803 2416 20812 2456
rect 20852 2416 21504 2456
rect 5923 2415 5981 2416
rect 10243 2415 10301 2416
rect 16771 2415 16829 2416
rect 18403 2415 18461 2416
rect 21424 2396 21504 2416
rect 5731 2372 5789 2373
rect 4483 2332 4492 2372
rect 4532 2332 5740 2372
rect 5780 2332 5789 2372
rect 5731 2331 5789 2332
rect 7267 2372 7325 2373
rect 17731 2372 17789 2373
rect 7267 2332 7276 2372
rect 7316 2332 7468 2372
rect 7508 2332 7517 2372
rect 10339 2332 10348 2372
rect 10388 2332 12172 2372
rect 12212 2332 12221 2372
rect 12547 2332 12556 2372
rect 12596 2332 15572 2372
rect 7267 2331 7325 2332
rect 4387 2288 4445 2289
rect 8419 2288 8477 2289
rect 1699 2248 1708 2288
rect 1748 2248 2956 2288
rect 2996 2248 4108 2288
rect 4148 2248 4396 2288
rect 4436 2248 4445 2288
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 5731 2248 5740 2288
rect 5780 2248 8428 2288
rect 8468 2248 8477 2288
rect 4387 2247 4445 2248
rect 8419 2247 8477 2248
rect 8707 2288 8765 2289
rect 15532 2288 15572 2332
rect 17731 2332 17740 2372
rect 17780 2332 19276 2372
rect 19316 2332 19325 2372
rect 17731 2331 17789 2332
rect 8707 2248 8716 2288
rect 8756 2248 11980 2288
rect 12020 2248 15244 2288
rect 15284 2248 15293 2288
rect 15532 2248 19372 2288
rect 19412 2248 19852 2288
rect 19892 2248 19901 2288
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 8707 2247 8765 2248
rect 5635 2204 5693 2205
rect 8803 2204 8861 2205
rect 4003 2164 4012 2204
rect 4052 2164 4204 2204
rect 4244 2164 4396 2204
rect 4436 2164 5644 2204
rect 5684 2164 5693 2204
rect 5923 2164 5932 2204
rect 5972 2164 7660 2204
rect 7700 2164 7709 2204
rect 8803 2164 8812 2204
rect 8852 2164 8946 2204
rect 9667 2164 9676 2204
rect 9716 2164 11020 2204
rect 11060 2164 11069 2204
rect 11980 2164 12460 2204
rect 12500 2164 12509 2204
rect 13027 2164 13036 2204
rect 13076 2164 18220 2204
rect 18260 2164 18269 2204
rect 5068 2120 5108 2164
rect 5635 2163 5693 2164
rect 8803 2163 8861 2164
rect 11020 2120 11060 2164
rect 5059 2080 5068 2120
rect 5108 2080 5148 2120
rect 5539 2080 5548 2120
rect 5588 2080 9580 2120
rect 9620 2080 9629 2120
rect 9955 2080 9964 2120
rect 10004 2080 10252 2120
rect 10292 2080 10301 2120
rect 11020 2080 11404 2120
rect 11444 2080 11453 2120
rect 11980 2036 12020 2164
rect 20611 2120 20669 2121
rect 21424 2120 21504 2140
rect 12163 2080 12172 2120
rect 12212 2080 12556 2120
rect 12596 2080 12605 2120
rect 13123 2080 13132 2120
rect 13172 2080 13612 2120
rect 13652 2080 18028 2120
rect 18068 2080 18077 2120
rect 18595 2080 18604 2120
rect 18644 2080 19660 2120
rect 19700 2080 19709 2120
rect 20611 2080 20620 2120
rect 20660 2080 21504 2120
rect 20611 2079 20669 2080
rect 21424 2060 21504 2080
rect 1987 1996 1996 2036
rect 2036 1996 12020 2036
rect 15523 1996 15532 2036
rect 15572 1996 17740 2036
rect 17780 1996 17789 2036
rect 2083 1952 2141 1953
rect 6499 1952 6557 1953
rect 7171 1952 7229 1953
rect 9571 1952 9629 1953
rect 16771 1952 16829 1953
rect 2083 1912 2092 1952
rect 2132 1912 4012 1952
rect 4052 1912 4061 1952
rect 6414 1912 6508 1952
rect 6548 1912 6557 1952
rect 6979 1912 6988 1952
rect 7028 1912 7180 1952
rect 7220 1912 7229 1952
rect 7843 1912 7852 1952
rect 7892 1912 8524 1952
rect 8564 1912 8573 1952
rect 9571 1912 9580 1952
rect 9620 1912 9772 1952
rect 9812 1912 9821 1952
rect 10531 1912 10540 1952
rect 10580 1912 15916 1952
rect 15956 1912 15965 1952
rect 16771 1912 16780 1952
rect 16820 1912 17932 1952
rect 17972 1912 17981 1952
rect 18499 1912 18508 1952
rect 18548 1912 20127 1952
rect 20167 1912 20176 1952
rect 2083 1911 2141 1912
rect 6499 1911 6557 1912
rect 7171 1911 7229 1912
rect 6883 1868 6941 1869
rect 6798 1828 6892 1868
rect 6932 1828 6941 1868
rect 8524 1868 8564 1912
rect 9571 1911 9629 1912
rect 16771 1911 16829 1912
rect 17731 1868 17789 1869
rect 8524 1828 12692 1868
rect 6883 1827 6941 1828
rect 3619 1744 3628 1784
rect 3668 1744 6796 1784
rect 6836 1744 6845 1784
rect 9763 1744 9772 1784
rect 9812 1744 11360 1784
rect 11491 1744 11500 1784
rect 11540 1744 12172 1784
rect 12212 1744 12221 1784
rect 11320 1700 11360 1744
rect 12652 1700 12692 1828
rect 15436 1828 17452 1868
rect 17492 1828 17501 1868
rect 17646 1828 17740 1868
rect 17780 1828 17789 1868
rect 15436 1784 15476 1828
rect 17731 1827 17789 1828
rect 18595 1784 18653 1785
rect 20707 1784 20765 1785
rect 21424 1784 21504 1804
rect 12739 1744 12748 1784
rect 12788 1744 13804 1784
rect 13844 1744 15436 1784
rect 15476 1744 15485 1784
rect 16195 1744 16204 1784
rect 16244 1744 17164 1784
rect 17204 1744 17213 1784
rect 18595 1744 18604 1784
rect 18644 1744 19852 1784
rect 19892 1744 19901 1784
rect 20707 1744 20716 1784
rect 20756 1744 21504 1784
rect 18595 1743 18653 1744
rect 20707 1743 20765 1744
rect 21424 1724 21504 1744
rect 2851 1660 2860 1700
rect 2900 1660 2996 1700
rect 6115 1660 6124 1700
rect 6164 1660 10252 1700
rect 10292 1660 10301 1700
rect 11320 1660 11732 1700
rect 12652 1660 14132 1700
rect 14179 1660 14188 1700
rect 14228 1660 15052 1700
rect 15092 1660 17452 1700
rect 17492 1660 17501 1700
rect 2851 1616 2909 1617
rect 2179 1576 2188 1616
rect 2228 1576 2860 1616
rect 2900 1576 2909 1616
rect 2956 1616 2996 1660
rect 11692 1616 11732 1660
rect 2956 1576 10540 1616
rect 10580 1576 10589 1616
rect 10915 1576 10924 1616
rect 10964 1576 11596 1616
rect 11636 1576 11645 1616
rect 11692 1576 13132 1616
rect 13172 1576 13181 1616
rect 13315 1576 13324 1616
rect 13364 1576 13708 1616
rect 13748 1576 13757 1616
rect 2851 1575 2909 1576
rect 11203 1532 11261 1533
rect 14092 1532 14132 1660
rect 15427 1616 15485 1617
rect 15427 1576 15436 1616
rect 15476 1576 20180 1616
rect 15427 1575 15485 1576
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 4291 1492 4300 1532
rect 4340 1492 11212 1532
rect 11252 1492 11261 1532
rect 11779 1492 11788 1532
rect 11828 1492 12364 1532
rect 12404 1492 12413 1532
rect 14092 1492 16876 1532
rect 16916 1492 16925 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 11203 1491 11261 1492
rect 20140 1448 20180 1576
rect 21424 1448 21504 1468
rect 1411 1408 1420 1448
rect 1460 1408 8812 1448
rect 8852 1408 8861 1448
rect 11299 1408 11308 1448
rect 11348 1408 15436 1448
rect 15476 1408 15485 1448
rect 16387 1408 16396 1448
rect 16436 1408 19276 1448
rect 19316 1408 19325 1448
rect 20140 1408 21504 1448
rect 21424 1388 21504 1408
rect 5347 1364 5405 1365
rect 8035 1364 8093 1365
rect 1699 1324 1708 1364
rect 1748 1324 3052 1364
rect 3092 1324 3101 1364
rect 4003 1324 4012 1364
rect 4052 1324 5356 1364
rect 5396 1324 5405 1364
rect 7267 1324 7276 1364
rect 7316 1324 8044 1364
rect 8084 1324 8236 1364
rect 8276 1324 8285 1364
rect 9763 1324 9772 1364
rect 9812 1324 17548 1364
rect 17588 1324 17597 1364
rect 5347 1323 5405 1324
rect 8035 1323 8093 1324
rect 2755 1280 2813 1281
rect 3331 1280 3389 1281
rect 6211 1280 6269 1281
rect 6595 1280 6653 1281
rect 2275 1240 2284 1280
rect 2324 1240 2476 1280
rect 2516 1240 2525 1280
rect 2670 1240 2764 1280
rect 2804 1240 2813 1280
rect 3246 1240 3340 1280
rect 3380 1240 3389 1280
rect 3907 1240 3916 1280
rect 3956 1240 4204 1280
rect 4244 1240 4253 1280
rect 4771 1240 4780 1280
rect 4820 1240 5644 1280
rect 5684 1240 5693 1280
rect 6126 1240 6220 1280
rect 6260 1240 6269 1280
rect 6510 1240 6604 1280
rect 6644 1240 6653 1280
rect 2755 1239 2813 1240
rect 3331 1239 3389 1240
rect 6211 1239 6269 1240
rect 6595 1239 6653 1240
rect 6787 1280 6845 1281
rect 6979 1280 7037 1281
rect 7171 1280 7229 1281
rect 7747 1280 7805 1281
rect 8131 1280 8189 1281
rect 6787 1240 6796 1280
rect 6836 1240 6930 1280
rect 6979 1240 6988 1280
rect 7028 1240 7122 1280
rect 7171 1240 7180 1280
rect 7220 1240 7314 1280
rect 7662 1240 7756 1280
rect 7796 1240 7805 1280
rect 8046 1240 8140 1280
rect 8180 1240 8189 1280
rect 6787 1239 6845 1240
rect 6979 1239 7037 1240
rect 7171 1239 7229 1240
rect 7747 1239 7805 1240
rect 8131 1239 8189 1240
rect 8323 1280 8381 1281
rect 8899 1280 8957 1281
rect 13315 1280 13373 1281
rect 14275 1280 14333 1281
rect 14467 1280 14525 1281
rect 8323 1240 8332 1280
rect 8372 1240 8466 1280
rect 8515 1240 8524 1280
rect 8564 1240 8908 1280
rect 8948 1240 8957 1280
rect 11011 1240 11020 1280
rect 11060 1240 12940 1280
rect 12980 1240 12989 1280
rect 13230 1240 13324 1280
rect 13364 1240 13373 1280
rect 14190 1240 14284 1280
rect 14324 1240 14333 1280
rect 14382 1240 14476 1280
rect 14516 1240 14525 1280
rect 8323 1239 8381 1240
rect 8899 1239 8957 1240
rect 13315 1239 13373 1240
rect 14275 1239 14333 1240
rect 14467 1239 14525 1240
rect 14659 1280 14717 1281
rect 16963 1280 17021 1281
rect 14659 1240 14668 1280
rect 14708 1240 14802 1280
rect 16878 1240 16972 1280
rect 17012 1240 17021 1280
rect 14659 1239 14717 1240
rect 16963 1239 17021 1240
rect 17155 1280 17213 1281
rect 17923 1280 17981 1281
rect 18499 1280 18557 1281
rect 17155 1240 17164 1280
rect 17204 1240 17492 1280
rect 17838 1240 17932 1280
rect 17972 1240 17981 1280
rect 18414 1240 18508 1280
rect 18548 1240 18557 1280
rect 17155 1239 17213 1240
rect 1507 1196 1565 1197
rect 5251 1196 5309 1197
rect 9379 1196 9437 1197
rect 15139 1196 15197 1197
rect 16291 1196 16349 1197
rect 17452 1196 17492 1240
rect 17923 1239 17981 1240
rect 18499 1239 18557 1240
rect 18691 1280 18749 1281
rect 18691 1240 18700 1280
rect 18740 1240 18834 1280
rect 18691 1239 18749 1240
rect 1422 1156 1516 1196
rect 1556 1156 1565 1196
rect 2563 1156 2572 1196
rect 2612 1156 4724 1196
rect 5166 1156 5260 1196
rect 5300 1156 5309 1196
rect 5443 1156 5452 1196
rect 5492 1156 6124 1196
rect 6164 1156 6173 1196
rect 7459 1156 7468 1196
rect 7508 1156 8428 1196
rect 8468 1156 8477 1196
rect 9283 1156 9292 1196
rect 9332 1156 9388 1196
rect 9428 1156 9437 1196
rect 10723 1156 10732 1196
rect 10772 1156 13900 1196
rect 13940 1156 13949 1196
rect 14371 1156 14380 1196
rect 14420 1156 14860 1196
rect 14900 1156 14909 1196
rect 15139 1156 15148 1196
rect 15188 1156 16300 1196
rect 16340 1156 16349 1196
rect 16483 1156 16492 1196
rect 16532 1156 17356 1196
rect 17396 1156 17405 1196
rect 17452 1156 20180 1196
rect 1507 1155 1565 1156
rect 4291 1112 4349 1113
rect 4684 1112 4724 1156
rect 5251 1155 5309 1156
rect 9379 1155 9437 1156
rect 15139 1155 15197 1156
rect 16291 1155 16349 1156
rect 20140 1112 20180 1156
rect 21424 1112 21504 1132
rect 2083 1072 2092 1112
rect 2132 1072 3148 1112
rect 3188 1072 3197 1112
rect 4099 1072 4108 1112
rect 4148 1072 4300 1112
rect 4340 1072 4349 1112
rect 4675 1072 4684 1112
rect 4724 1072 5356 1112
rect 5396 1072 5405 1112
rect 7075 1072 7084 1112
rect 7124 1072 9964 1112
rect 10004 1072 10013 1112
rect 13123 1072 13132 1112
rect 13172 1072 13420 1112
rect 13460 1072 13469 1112
rect 14947 1072 14956 1112
rect 14996 1072 15628 1112
rect 15668 1072 15677 1112
rect 16291 1072 16300 1112
rect 16340 1072 17740 1112
rect 17780 1072 17789 1112
rect 20140 1072 21504 1112
rect 4291 1071 4349 1072
rect 21424 1052 21504 1072
rect 4867 988 4876 1028
rect 4916 988 8044 1028
rect 8084 988 8093 1028
rect 8227 988 8236 1028
rect 8276 988 8908 1028
rect 8948 988 10156 1028
rect 10196 988 10205 1028
rect 13219 988 13228 1028
rect 13268 988 17548 1028
rect 17588 988 17597 1028
rect 3523 944 3581 945
rect 6019 944 6077 945
rect 835 904 844 944
rect 884 904 1996 944
rect 2036 904 2045 944
rect 3438 904 3532 944
rect 3572 904 3581 944
rect 5934 904 6028 944
rect 6068 904 6077 944
rect 3523 903 3581 904
rect 6019 903 6077 904
rect 6403 944 6461 945
rect 8611 944 8669 945
rect 12547 944 12605 945
rect 12931 944 12989 945
rect 13507 944 13565 945
rect 6403 904 6412 944
rect 6452 904 7372 944
rect 7412 904 7421 944
rect 7555 904 7564 944
rect 7604 904 8620 944
rect 8660 904 8669 944
rect 9475 904 9484 944
rect 9524 904 11212 944
rect 11252 904 11261 944
rect 12462 904 12556 944
rect 12596 904 12605 944
rect 12846 904 12940 944
rect 12980 904 12989 944
rect 13422 904 13516 944
rect 13556 904 13565 944
rect 6403 903 6461 904
rect 8611 903 8669 904
rect 12547 903 12605 904
rect 12931 903 12989 904
rect 13507 903 13565 904
rect 13699 944 13757 945
rect 17635 944 17693 945
rect 18211 944 18269 945
rect 13699 904 13708 944
rect 13748 904 13842 944
rect 17635 904 17644 944
rect 17684 904 17740 944
rect 17780 904 17789 944
rect 18211 904 18220 944
rect 18260 904 19084 944
rect 19124 904 19133 944
rect 20035 904 20044 944
rect 20084 904 20093 944
rect 13699 903 13757 904
rect 17635 903 17693 904
rect 18211 903 18269 904
rect 7939 860 7997 861
rect 13123 860 13181 861
rect 20044 860 20084 904
rect 3427 820 3436 860
rect 3476 820 7508 860
rect 7854 820 7948 860
rect 7988 820 7997 860
rect 13038 820 13132 860
rect 13172 820 13181 860
rect 15235 820 15244 860
rect 15284 820 20084 860
rect 7468 776 7508 820
rect 7939 819 7997 820
rect 13123 819 13181 820
rect 16003 776 16061 777
rect 20515 776 20573 777
rect 21424 776 21504 796
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 7468 736 15820 776
rect 15860 736 15869 776
rect 16003 736 16012 776
rect 16052 736 19468 776
rect 19508 736 19517 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 20515 736 20524 776
rect 20564 736 21504 776
rect 16003 735 16061 736
rect 20515 735 20573 736
rect 21424 716 21504 736
rect 5443 692 5501 693
rect 7075 692 7133 693
rect 13891 692 13949 693
rect 5358 652 5452 692
rect 5492 652 5501 692
rect 5827 652 5836 692
rect 5876 652 7084 692
rect 7124 652 7133 692
rect 8803 652 8812 692
rect 8852 652 9292 692
rect 9332 652 9341 692
rect 13806 652 13900 692
rect 13940 652 13949 692
rect 5443 651 5501 652
rect 7075 651 7133 652
rect 13891 651 13949 652
rect 15331 692 15389 693
rect 15331 652 15340 692
rect 15380 652 18316 692
rect 18356 652 18365 692
rect 15331 651 15389 652
rect 4675 608 4733 609
rect 5539 608 5597 609
rect 7459 608 7517 609
rect 15139 608 15197 609
rect 4675 568 4684 608
rect 4724 568 4876 608
rect 4916 568 4925 608
rect 5251 568 5260 608
rect 5300 568 5548 608
rect 5588 568 5597 608
rect 6403 568 6412 608
rect 6452 568 7468 608
rect 7508 568 7517 608
rect 7843 568 7852 608
rect 7892 568 14188 608
rect 14228 568 14237 608
rect 14284 568 15148 608
rect 15188 568 15197 608
rect 4675 567 4733 568
rect 5539 567 5597 568
rect 7459 567 7517 568
rect 14284 524 14324 568
rect 15139 567 15197 568
rect 15715 608 15773 609
rect 15715 568 15724 608
rect 15764 568 19276 608
rect 19316 568 19325 608
rect 15715 567 15773 568
rect 1699 484 1708 524
rect 1748 484 2540 524
rect 5923 484 5932 524
rect 5972 484 11020 524
rect 11060 484 11069 524
rect 12739 484 12748 524
rect 12788 484 14324 524
rect 14851 484 14860 524
rect 14900 484 19660 524
rect 19700 484 19709 524
rect 2500 356 2540 484
rect 18883 440 18941 441
rect 5539 400 5548 440
rect 5588 400 15052 440
rect 15092 400 15101 440
rect 15811 400 15820 440
rect 15860 400 16108 440
rect 16148 400 16157 440
rect 16867 400 16876 440
rect 16916 400 17548 440
rect 17588 400 17597 440
rect 18798 400 18892 440
rect 18932 400 18941 440
rect 18883 399 18941 400
rect 19651 440 19709 441
rect 21424 440 21504 460
rect 19651 400 19660 440
rect 19700 400 21504 440
rect 19651 399 19709 400
rect 21424 380 21504 400
rect 12163 356 12221 357
rect 2500 316 8908 356
rect 8948 316 8957 356
rect 10915 316 10924 356
rect 10964 316 12172 356
rect 12212 316 16780 356
rect 16820 316 16829 356
rect 12163 315 12221 316
rect 15619 272 15677 273
rect 5347 232 5356 272
rect 5396 232 10636 272
rect 10676 232 10685 272
rect 11491 232 11500 272
rect 11540 232 11549 272
rect 15534 232 15628 272
rect 15668 232 15677 272
rect 6115 148 6124 188
rect 6164 148 6173 188
rect 9763 148 9772 188
rect 9812 148 11404 188
rect 11444 148 11453 188
rect 5059 104 5117 105
rect 4974 64 5068 104
rect 5108 64 5117 104
rect 6124 104 6164 148
rect 11500 104 11540 232
rect 15619 231 15677 232
rect 12451 148 12460 188
rect 12500 148 14380 188
rect 14420 148 17164 188
rect 17204 148 17213 188
rect 17539 104 17597 105
rect 18115 104 18173 105
rect 21424 104 21504 124
rect 6124 64 10828 104
rect 10868 64 10877 104
rect 11500 64 17548 104
rect 17588 64 17597 104
rect 18030 64 18124 104
rect 18164 64 18173 104
rect 21187 64 21196 104
rect 21236 64 21504 104
rect 5059 63 5117 64
rect 17539 63 17597 64
rect 18115 63 18173 64
rect 21424 44 21504 64
<< via3 >>
rect 15532 42904 15572 42944
rect 1420 42820 1460 42860
rect 21100 42736 21140 42776
rect 7564 42652 7604 42692
rect 18316 42652 18356 42692
rect 9484 42568 9524 42608
rect 18028 42568 18068 42608
rect 460 42484 500 42524
rect 1036 42400 1076 42440
rect 21292 42064 21332 42104
rect 6412 41980 6452 42020
rect 16300 41980 16340 42020
rect 5452 41896 5492 41936
rect 17932 41896 17972 41936
rect 5548 41812 5588 41852
rect 7852 41812 7892 41852
rect 18220 41812 18260 41852
rect 16396 41728 16436 41768
rect 3148 41560 3188 41600
rect 5836 41644 5876 41684
rect 11404 41644 11444 41684
rect 19468 41644 19508 41684
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 6604 41560 6644 41600
rect 6796 41560 6836 41600
rect 7180 41560 7220 41600
rect 7372 41560 7412 41600
rect 7948 41560 7988 41600
rect 9292 41560 9332 41600
rect 9868 41560 9908 41600
rect 10252 41560 10292 41600
rect 11020 41560 11060 41600
rect 11500 41560 11540 41600
rect 11788 41560 11828 41600
rect 12268 41560 12308 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 1132 41476 1172 41516
rect 15724 41476 15764 41516
rect 17164 41476 17204 41516
rect 17260 41392 17300 41432
rect 18316 41308 18356 41348
rect 3052 41224 3092 41264
rect 7468 41140 7508 41180
rect 15628 41140 15668 41180
rect 16396 41140 16436 41180
rect 19660 41140 19700 41180
rect 19852 41140 19892 41180
rect 20140 41056 20180 41096
rect 10828 40972 10868 41012
rect 15436 40972 15476 41012
rect 16396 40972 16436 41012
rect 16588 40972 16628 41012
rect 17068 40972 17108 41012
rect 17548 40972 17588 41012
rect 18316 40972 18356 41012
rect 19084 40972 19124 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 12940 40720 12980 40760
rect 17740 40720 17780 40760
rect 16588 40636 16628 40676
rect 12844 40552 12884 40592
rect 18124 40552 18164 40592
rect 19276 40552 19316 40592
rect 268 40468 308 40508
rect 1324 40384 1364 40424
rect 2284 40468 2324 40508
rect 5740 40468 5780 40508
rect 6508 40468 6548 40508
rect 8812 40468 8852 40508
rect 2956 40384 2996 40424
rect 12652 40384 12692 40424
rect 16108 40384 16148 40424
rect 16396 40384 16436 40424
rect 16972 40384 17012 40424
rect 17452 40384 17492 40424
rect 4204 40300 4244 40340
rect 6796 40300 6836 40340
rect 10156 40300 10196 40340
rect 16300 40300 16340 40340
rect 18412 40300 18452 40340
rect 18604 40300 18644 40340
rect 6988 40216 7028 40256
rect 15148 40216 15188 40256
rect 18508 40216 18548 40256
rect 15052 40132 15092 40172
rect 15628 40132 15668 40172
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 8044 39964 8084 40004
rect 15724 40048 15764 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 15244 39964 15284 40004
rect 16108 39964 16148 40004
rect 16972 39880 17012 39920
rect 18700 39880 18740 39920
rect 6796 39796 6836 39836
rect 19372 39796 19412 39836
rect 2188 39712 2228 39752
rect 2860 39712 2900 39752
rect 16396 39712 16436 39752
rect 5356 39628 5396 39668
rect 7084 39628 7124 39668
rect 8524 39628 8564 39668
rect 8908 39628 8948 39668
rect 17836 39628 17876 39668
rect 19948 39628 19988 39668
rect 2380 39544 2420 39584
rect 12556 39544 12596 39584
rect 8908 39460 8948 39500
rect 15820 39460 15860 39500
rect 16492 39460 16532 39500
rect 14572 39376 14612 39416
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 17644 39292 17684 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 2092 39208 2132 39248
rect 16396 39208 16436 39248
rect 17164 39124 17204 39164
rect 1324 39040 1364 39080
rect 1900 39040 1940 39080
rect 10636 39040 10676 39080
rect 12172 39040 12212 39080
rect 20140 39040 20180 39080
rect 1804 38956 1844 38996
rect 8812 38956 8852 38996
rect 3052 38872 3092 38912
rect 14956 38872 14996 38912
rect 15628 38956 15668 38996
rect 19564 38956 19604 38996
rect 15148 38872 15188 38912
rect 1996 38704 2036 38744
rect 3532 38704 3572 38744
rect 4300 38704 4340 38744
rect 4588 38704 4628 38744
rect 6316 38704 6356 38744
rect 6988 38704 7028 38744
rect 15148 38704 15188 38744
rect 16972 38704 17012 38744
rect 18412 38704 18452 38744
rect 20524 38704 20564 38744
rect 20812 38704 20852 38744
rect 18700 38620 18740 38660
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 18604 38536 18644 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 18508 38452 18548 38492
rect 2764 38284 2804 38324
rect 13324 38368 13364 38408
rect 15244 38368 15284 38408
rect 5836 38284 5876 38324
rect 5356 38200 5396 38240
rect 1516 38116 1556 38156
rect 1708 38116 1748 38156
rect 2572 38116 2612 38156
rect 3340 38116 3380 38156
rect 20140 38368 20180 38408
rect 13708 38284 13748 38324
rect 16588 38284 16628 38324
rect 16972 38284 17012 38324
rect 19276 38284 19316 38324
rect 6700 38200 6740 38240
rect 16108 38200 16148 38240
rect 7468 38116 7508 38156
rect 17260 38116 17300 38156
rect 6220 38032 6260 38072
rect 14188 38032 14228 38072
rect 15628 38032 15668 38072
rect 18700 38032 18740 38072
rect 15052 37948 15092 37988
rect 17548 37948 17588 37988
rect 2476 37864 2516 37904
rect 2764 37864 2804 37904
rect 6988 37864 7028 37904
rect 12460 37864 12500 37904
rect 20140 38032 20180 38072
rect 12652 37864 12692 37904
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 6316 37780 6356 37820
rect 13900 37780 13940 37820
rect 14476 37864 14516 37904
rect 17836 37864 17876 37904
rect 15724 37780 15764 37820
rect 1420 37612 1460 37652
rect 6988 37696 7028 37736
rect 15340 37696 15380 37736
rect 1708 37612 1748 37652
rect 2572 37528 2612 37568
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 20140 37696 20180 37736
rect 9964 37612 10004 37652
rect 13900 37612 13940 37652
rect 17836 37612 17876 37652
rect 21196 37612 21236 37652
rect 16396 37528 16436 37568
rect 16780 37528 16820 37568
rect 18412 37528 18452 37568
rect 19372 37528 19412 37568
rect 3532 37444 3572 37484
rect 6028 37444 6068 37484
rect 9388 37444 9428 37484
rect 20044 37444 20084 37484
rect 9004 37360 9044 37400
rect 20332 37360 20372 37400
rect 12364 37276 12404 37316
rect 3052 37192 3092 37232
rect 3820 37192 3860 37232
rect 4492 37192 4532 37232
rect 8908 37192 8948 37232
rect 13900 37192 13940 37232
rect 19276 37192 19316 37232
rect 3244 37108 3284 37148
rect 5644 37108 5684 37148
rect 13996 37108 14036 37148
rect 17452 37108 17492 37148
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 15244 37024 15284 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20620 37024 20660 37064
rect 15340 36940 15380 36980
rect 18604 36940 18644 36980
rect 2572 36856 2612 36896
rect 14476 36856 14516 36896
rect 17932 36856 17972 36896
rect 2668 36772 2708 36812
rect 12652 36772 12692 36812
rect 10348 36688 10388 36728
rect 17068 36772 17108 36812
rect 15340 36688 15380 36728
rect 6988 36604 7028 36644
rect 9580 36604 9620 36644
rect 16012 36604 16052 36644
rect 19468 36604 19508 36644
rect 3052 36520 3092 36560
rect 12460 36520 12500 36560
rect 20140 36520 20180 36560
rect 2572 36436 2612 36476
rect 15244 36352 15284 36392
rect 15724 36352 15764 36392
rect 17356 36352 17396 36392
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 3052 36184 3092 36224
rect 4588 36184 4628 36224
rect 2860 36100 2900 36140
rect 11308 36184 11348 36224
rect 19372 36184 19412 36224
rect 1228 36016 1268 36056
rect 13708 36016 13748 36056
rect 364 35932 404 35972
rect 1900 35932 1940 35972
rect 16300 36100 16340 36140
rect 17836 36100 17876 36140
rect 17068 36016 17108 36056
rect 18508 36016 18548 36056
rect 19948 36016 19988 36056
rect 20140 36016 20180 36056
rect 1612 35848 1652 35888
rect 2668 35848 2708 35888
rect 4780 35848 4820 35888
rect 8044 35848 8084 35888
rect 2764 35764 2804 35804
rect 6028 35764 6068 35804
rect 11308 35764 11348 35804
rect 2188 35680 2228 35720
rect 12748 35764 12788 35804
rect 16108 35764 16148 35804
rect 16396 35764 16436 35804
rect 3628 35680 3668 35720
rect 10828 35680 10868 35720
rect 12940 35680 12980 35720
rect 20716 35680 20756 35720
rect 20908 35680 20948 35720
rect 1420 35596 1460 35636
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 7660 35428 7700 35468
rect 13228 35428 13268 35468
rect 16684 35428 16724 35468
rect 17164 35344 17204 35384
rect 4108 35260 4148 35300
rect 2188 35176 2228 35216
rect 4780 35176 4820 35216
rect 5260 35176 5300 35216
rect 844 35092 884 35132
rect 4396 35092 4436 35132
rect 1900 34924 1940 34964
rect 6892 35176 6932 35216
rect 9964 35260 10004 35300
rect 10444 35260 10484 35300
rect 10828 35260 10868 35300
rect 17644 35344 17684 35384
rect 16012 35260 16052 35300
rect 18796 35260 18836 35300
rect 7756 35176 7796 35216
rect 14092 35176 14132 35216
rect 7084 35092 7124 35132
rect 14572 35092 14612 35132
rect 17836 35092 17876 35132
rect 3532 35008 3572 35048
rect 6316 35008 6356 35048
rect 9388 35008 9428 35048
rect 10060 35008 10100 35048
rect 13516 35008 13556 35048
rect 17740 35008 17780 35048
rect 3052 34924 3092 34964
rect 16396 34924 16436 34964
rect 5644 34840 5684 34880
rect 10060 34840 10100 34880
rect 2188 34756 2228 34796
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 11116 34756 11156 34796
rect 11884 34756 11924 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 2956 34672 2996 34712
rect 20140 34672 20180 34712
rect 1612 34588 1652 34628
rect 4684 34588 4724 34628
rect 6700 34588 6740 34628
rect 13420 34588 13460 34628
rect 4492 34504 4532 34544
rect 17644 34504 17684 34544
rect 19948 34504 19988 34544
rect 4876 34420 4916 34460
rect 6796 34420 6836 34460
rect 7564 34420 7604 34460
rect 8428 34420 8468 34460
rect 4780 34336 4820 34376
rect 5644 34336 5684 34376
rect 7276 34336 7316 34376
rect 8044 34336 8084 34376
rect 9964 34336 10004 34376
rect 11692 34336 11732 34376
rect 17452 34336 17492 34376
rect 20524 34336 20564 34376
rect 3628 34252 3668 34292
rect 13036 34252 13076 34292
rect 16492 34252 16532 34292
rect 1900 34168 1940 34208
rect 6124 34168 6164 34208
rect 10060 34168 10100 34208
rect 10732 34168 10772 34208
rect 15148 34168 15188 34208
rect 10636 34084 10676 34124
rect 12076 34084 12116 34124
rect 15724 34084 15764 34124
rect 3532 34000 3572 34040
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 5932 34000 5972 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 6892 33832 6932 33872
rect 7660 33832 7700 33872
rect 7564 33748 7604 33788
rect 16204 33916 16244 33956
rect 16588 33832 16628 33872
rect 21388 33832 21428 33872
rect 13324 33748 13364 33788
rect 19564 33748 19604 33788
rect 10540 33664 10580 33704
rect 17932 33664 17972 33704
rect 4588 33580 4628 33620
rect 13324 33580 13364 33620
rect 19468 33580 19508 33620
rect 6700 33496 6740 33536
rect 10540 33496 10580 33536
rect 19852 33496 19892 33536
rect 2572 33412 2612 33452
rect 15436 33412 15476 33452
rect 10924 33328 10964 33368
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 6796 33244 6836 33284
rect 16300 33244 16340 33284
rect 17740 33244 17780 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 12460 33160 12500 33200
rect 15916 33160 15956 33200
rect 2284 33076 2324 33116
rect 6124 33076 6164 33116
rect 7756 33076 7796 33116
rect 13804 33076 13844 33116
rect 18508 33076 18548 33116
rect 19660 33076 19700 33116
rect 6508 32992 6548 33032
rect 11980 32992 12020 33032
rect 2188 32908 2228 32948
rect 2284 32824 2324 32864
rect 2764 32824 2804 32864
rect 6700 32908 6740 32948
rect 14284 32908 14324 32948
rect 3244 32824 3284 32864
rect 3532 32824 3572 32864
rect 8236 32824 8276 32864
rect 8428 32824 8468 32864
rect 11596 32824 11636 32864
rect 4684 32740 4724 32780
rect 6220 32740 6260 32780
rect 14092 32740 14132 32780
rect 21196 32656 21236 32696
rect 6220 32572 6260 32612
rect 11116 32572 11156 32612
rect 16012 32572 16052 32612
rect 16300 32572 16340 32612
rect 17068 32572 17108 32612
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 6316 32488 6356 32528
rect 6988 32488 7028 32528
rect 7756 32488 7796 32528
rect 11308 32488 11348 32528
rect 13900 32488 13940 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 14284 32404 14324 32444
rect 1324 32236 1364 32276
rect 3340 32320 3380 32360
rect 7564 32320 7604 32360
rect 16012 32320 16052 32360
rect 11980 32236 12020 32276
rect 18220 32236 18260 32276
rect 18700 32236 18740 32276
rect 1420 32068 1460 32108
rect 4204 32152 4244 32192
rect 8620 32152 8660 32192
rect 11116 32152 11156 32192
rect 1612 32068 1652 32108
rect 7180 31984 7220 32024
rect 3052 31900 3092 31940
rect 3532 31900 3572 31940
rect 7564 31900 7604 31940
rect 11596 31900 11636 31940
rect 14572 31900 14612 31940
rect 16684 31900 16724 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 9964 31732 10004 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 20140 31648 20180 31688
rect 13804 31564 13844 31604
rect 16396 31564 16436 31604
rect 18700 31564 18740 31604
rect 5452 31480 5492 31520
rect 7564 31480 7604 31520
rect 8812 31480 8852 31520
rect 9100 31480 9140 31520
rect 10444 31480 10484 31520
rect 15724 31480 15764 31520
rect 20908 31480 20948 31520
rect 8428 31396 8468 31436
rect 11980 31396 12020 31436
rect 12844 31396 12884 31436
rect 17068 31396 17108 31436
rect 18508 31396 18548 31436
rect 21196 31396 21236 31436
rect 5644 31312 5684 31352
rect 10060 31312 10100 31352
rect 10348 31312 10388 31352
rect 10732 31312 10772 31352
rect 13804 31312 13844 31352
rect 20716 31312 20756 31352
rect 7660 31228 7700 31268
rect 10924 31228 10964 31268
rect 13708 31228 13748 31268
rect 16204 31228 16244 31268
rect 12076 31144 12116 31184
rect 14284 31144 14324 31184
rect 17740 31144 17780 31184
rect 19564 31144 19604 31184
rect 19660 31060 19700 31100
rect 3436 30976 3476 31016
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 5932 30976 5972 31016
rect 11884 30976 11924 31016
rect 16204 30976 16244 31016
rect 17932 30976 17972 31016
rect 19852 30976 19892 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 2572 30892 2612 30932
rect 11116 30892 11156 30932
rect 12172 30892 12212 30932
rect 3436 30808 3476 30848
rect 14092 30892 14132 30932
rect 16876 30808 16916 30848
rect 5548 30724 5588 30764
rect 11884 30724 11924 30764
rect 12844 30724 12884 30764
rect 7660 30640 7700 30680
rect 16012 30640 16052 30680
rect 17740 30724 17780 30764
rect 6124 30556 6164 30596
rect 5932 30472 5972 30512
rect 11116 30472 11156 30512
rect 9004 30388 9044 30428
rect 652 30304 692 30344
rect 5644 30304 5684 30344
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 4780 30220 4820 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 12076 30136 12116 30176
rect 12844 30136 12884 30176
rect 4780 30052 4820 30092
rect 16588 30052 16628 30092
rect 8140 29968 8180 30008
rect 15052 29968 15092 30008
rect 12364 29884 12404 29924
rect 12748 29884 12788 29924
rect 16684 29884 16724 29924
rect 2860 29800 2900 29840
rect 1996 29716 2036 29756
rect 2476 29716 2516 29756
rect 8716 29716 8756 29756
rect 9196 29716 9236 29756
rect 16492 29716 16532 29756
rect 19852 29800 19892 29840
rect 3244 29632 3284 29672
rect 7180 29632 7220 29672
rect 11884 29632 11924 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 9676 29464 9716 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 6124 29380 6164 29420
rect 9004 29380 9044 29420
rect 13900 29380 13940 29420
rect 18220 29380 18260 29420
rect 2956 29296 2996 29336
rect 8428 29296 8468 29336
rect 9196 29296 9236 29336
rect 3244 29212 3284 29252
rect 7564 29212 7604 29252
rect 12268 29212 12308 29252
rect 13324 29212 13364 29252
rect 15436 29212 15476 29252
rect 3340 29128 3380 29168
rect 4204 29128 4244 29168
rect 4780 29128 4820 29168
rect 8428 29128 8468 29168
rect 10732 29128 10772 29168
rect 13420 29128 13460 29168
rect 17548 29128 17588 29168
rect 5452 29044 5492 29084
rect 13900 29044 13940 29084
rect 15820 29044 15860 29084
rect 19372 29044 19412 29084
rect 6700 28876 6740 28916
rect 9964 28876 10004 28916
rect 13708 28876 13748 28916
rect 17740 28876 17780 28916
rect 20524 28876 20564 28916
rect 3244 28792 3284 28832
rect 12076 28792 12116 28832
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 6988 28708 7028 28748
rect 9964 28708 10004 28748
rect 18220 28708 18260 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 5548 28624 5588 28664
rect 10060 28624 10100 28664
rect 10348 28624 10388 28664
rect 11884 28624 11924 28664
rect 18604 28624 18644 28664
rect 19276 28624 19316 28664
rect 5740 28540 5780 28580
rect 16012 28540 16052 28580
rect 16876 28540 16916 28580
rect 20812 28540 20852 28580
rect 7948 28456 7988 28496
rect 17260 28456 17300 28496
rect 3628 28372 3668 28412
rect 4108 28372 4148 28412
rect 7468 28372 7508 28412
rect 8140 28372 8180 28412
rect 5548 28204 5588 28244
rect 8428 28204 8468 28244
rect 16012 28288 16052 28328
rect 16204 28288 16244 28328
rect 21100 28204 21140 28244
rect 3436 28120 3476 28160
rect 1996 27952 2036 27992
rect 11596 28036 11636 28076
rect 12748 28036 12788 28076
rect 18220 28036 18260 28076
rect 4588 27952 4628 27992
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 3244 27868 3284 27908
rect 4108 27868 4148 27908
rect 5452 27868 5492 27908
rect 11020 27868 11060 27908
rect 12364 27784 12404 27824
rect 4492 27700 4532 27740
rect 11884 27700 11924 27740
rect 6220 27616 6260 27656
rect 8524 27616 8564 27656
rect 9388 27616 9428 27656
rect 11980 27616 12020 27656
rect 4300 27532 4340 27572
rect 3436 27448 3476 27488
rect 7372 27448 7412 27488
rect 9292 27448 9332 27488
rect 1324 27364 1364 27404
rect 3532 27364 3572 27404
rect 6700 27364 6740 27404
rect 6988 27364 7028 27404
rect 20524 27364 20564 27404
rect 5644 27280 5684 27320
rect 12076 27280 12116 27320
rect 17260 27280 17300 27320
rect 21292 27280 21332 27320
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 19372 27196 19412 27236
rect 11308 27112 11348 27152
rect 4108 27028 4148 27068
rect 15532 27028 15572 27068
rect 19372 27028 19412 27068
rect 1420 26944 1460 26984
rect 1804 26944 1844 26984
rect 15532 26860 15572 26900
rect 11980 26776 12020 26816
rect 17452 26776 17492 26816
rect 20812 26776 20852 26816
rect 2284 26692 2324 26732
rect 1324 26524 1364 26564
rect 2284 26524 2324 26564
rect 6700 26608 6740 26648
rect 10924 26608 10964 26648
rect 11308 26524 11348 26564
rect 12844 26524 12884 26564
rect 17740 26524 17780 26564
rect 19468 26524 19508 26564
rect 20908 26524 20948 26564
rect 3532 26440 3572 26480
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 6508 26440 6548 26480
rect 8620 26440 8660 26480
rect 8812 26440 8852 26480
rect 9004 26440 9044 26480
rect 9580 26440 9620 26480
rect 13900 26440 13940 26480
rect 15244 26440 15284 26480
rect 16492 26440 16532 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 1900 26356 1940 26396
rect 1228 26188 1268 26228
rect 4300 26188 4340 26228
rect 2860 26104 2900 26144
rect 12268 26020 12308 26060
rect 76 25936 116 25976
rect 1420 25936 1460 25976
rect 7948 25852 7988 25892
rect 11020 25852 11060 25892
rect 5740 25768 5780 25808
rect 17452 25768 17492 25808
rect 17644 25768 17684 25808
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 13996 25684 14036 25724
rect 16012 25684 16052 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 5836 25600 5876 25640
rect 17548 25600 17588 25640
rect 20908 25600 20948 25640
rect 6412 25516 6452 25556
rect 10540 25516 10580 25556
rect 12556 25516 12596 25556
rect 14764 25516 14804 25556
rect 12268 25432 12308 25472
rect 18028 25432 18068 25472
rect 3532 25348 3572 25388
rect 4588 25348 4628 25388
rect 7468 25348 7508 25388
rect 9676 25348 9716 25388
rect 10732 25348 10772 25388
rect 11116 25348 11156 25388
rect 12844 25348 12884 25388
rect 14572 25348 14612 25388
rect 2668 25264 2708 25304
rect 5068 25264 5108 25304
rect 19372 25264 19412 25304
rect 2380 25012 2420 25052
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 6892 24928 6932 24968
rect 18700 24928 18740 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 748 24760 788 24800
rect 6412 24760 6452 24800
rect 6700 24760 6740 24800
rect 8524 24760 8564 24800
rect 14956 24760 14996 24800
rect 17260 24760 17300 24800
rect 19852 24760 19892 24800
rect 2476 24592 2516 24632
rect 4204 24592 4244 24632
rect 10348 24592 10388 24632
rect 15244 24592 15284 24632
rect 20812 24928 20852 24968
rect 18028 24592 18068 24632
rect 8140 24508 8180 24548
rect 10924 24508 10964 24548
rect 15436 24424 15476 24464
rect 2476 24340 2516 24380
rect 4204 24340 4244 24380
rect 13036 24340 13076 24380
rect 14764 24256 14804 24296
rect 1804 24172 1844 24212
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 11788 24172 11828 24212
rect 16492 24172 16532 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 1516 24088 1556 24128
rect 7276 24088 7316 24128
rect 7372 24004 7412 24044
rect 15340 24088 15380 24128
rect 10060 24004 10100 24044
rect 13228 24004 13268 24044
rect 19276 24004 19316 24044
rect 20908 24004 20948 24044
rect 76 23920 116 23960
rect 556 23920 596 23960
rect 8140 23920 8180 23960
rect 12652 23920 12692 23960
rect 13036 23920 13076 23960
rect 13612 23920 13652 23960
rect 16780 23920 16820 23960
rect 6700 23836 6740 23876
rect 11788 23752 11828 23792
rect 12652 23752 12692 23792
rect 6412 23668 6452 23708
rect 7372 23668 7412 23708
rect 13996 23668 14036 23708
rect 18700 23668 18740 23708
rect 1900 23584 1940 23624
rect 8812 23584 8852 23624
rect 11308 23584 11348 23624
rect 19852 23584 19892 23624
rect 9196 23500 9236 23540
rect 10252 23500 10292 23540
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 7468 23416 7508 23456
rect 14764 23416 14804 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 9292 23332 9332 23372
rect 6316 23248 6356 23288
rect 7852 23248 7892 23288
rect 8524 23248 8564 23288
rect 16876 23248 16916 23288
rect 19948 23248 19988 23288
rect 2476 23164 2516 23204
rect 5932 23164 5972 23204
rect 1228 23080 1268 23120
rect 2188 22996 2228 23036
rect 3340 22996 3380 23036
rect 4588 22996 4628 23036
rect 5932 22996 5972 23036
rect 6412 22996 6452 23036
rect 10732 22996 10772 23036
rect 6220 22828 6260 22868
rect 6700 22828 6740 22868
rect 12076 22828 12116 22868
rect 13036 22828 13076 22868
rect 2764 22744 2804 22784
rect 7180 22744 7220 22784
rect 19468 22744 19508 22784
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 16300 22660 16340 22700
rect 16780 22660 16820 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 19372 22660 19412 22700
rect 268 22576 308 22616
rect 940 22492 980 22532
rect 6604 22492 6644 22532
rect 13612 22492 13652 22532
rect 1228 22408 1268 22448
rect 4684 22408 4724 22448
rect 13996 22408 14036 22448
rect 2668 22324 2708 22364
rect 7852 22324 7892 22364
rect 13420 22324 13460 22364
rect 19660 22240 19700 22280
rect 4492 22156 4532 22196
rect 15916 22156 15956 22196
rect 12652 22072 12692 22112
rect 16588 22072 16628 22112
rect 17548 22072 17588 22112
rect 460 21988 500 22028
rect 9196 21988 9236 22028
rect 12748 21988 12788 22028
rect 1036 21904 1076 21944
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 6892 21904 6932 21944
rect 15916 21904 15956 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 1132 21736 1172 21776
rect 1900 21736 1940 21776
rect 3532 21736 3572 21776
rect 3724 21736 3764 21776
rect 4492 21736 4532 21776
rect 6988 21736 7028 21776
rect 3052 21568 3092 21608
rect 9580 21568 9620 21608
rect 20620 21568 20660 21608
rect 460 21484 500 21524
rect 1420 21484 1460 21524
rect 2092 21484 2132 21524
rect 3244 21484 3284 21524
rect 16204 21484 16244 21524
rect 5356 21316 5396 21356
rect 9676 21316 9716 21356
rect 13228 21316 13268 21356
rect 19372 21316 19412 21356
rect 1900 21232 1940 21272
rect 7276 21232 7316 21272
rect 17644 21232 17684 21272
rect 21292 21232 21332 21272
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 12844 21064 12884 21104
rect 15628 21064 15668 21104
rect 17452 21064 17492 21104
rect 1516 20980 1556 21020
rect 11596 20980 11636 21020
rect 19948 20896 19988 20936
rect 1420 20812 1460 20852
rect 4300 20812 4340 20852
rect 12172 20812 12212 20852
rect 5548 20728 5588 20768
rect 5932 20728 5972 20768
rect 11596 20728 11636 20768
rect 9868 20644 9908 20684
rect 14188 20560 14228 20600
rect 15436 20560 15476 20600
rect 2380 20476 2420 20516
rect 268 20392 308 20432
rect 16396 20644 16436 20684
rect 19756 20560 19796 20600
rect 19852 20476 19892 20516
rect 2572 20392 2612 20432
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 3148 20308 3188 20348
rect 14188 20308 14228 20348
rect 12364 20224 12404 20264
rect 12652 20224 12692 20264
rect 13612 20140 13652 20180
rect 14764 20140 14804 20180
rect 12268 20056 12308 20096
rect 17548 20140 17588 20180
rect 18700 20140 18740 20180
rect 16396 20056 16436 20096
rect 1228 19888 1268 19928
rect 2956 19888 2996 19928
rect 3148 19888 3188 19928
rect 7372 19888 7412 19928
rect 8236 19972 8276 20012
rect 15340 19972 15380 20012
rect 10828 19888 10868 19928
rect 15628 19972 15668 20012
rect 19660 19972 19700 20012
rect 2572 19804 2612 19844
rect 3436 19804 3476 19844
rect 6604 19804 6644 19844
rect 15340 19720 15380 19760
rect 16204 19720 16244 19760
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 13612 19636 13652 19676
rect 14956 19636 14996 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 844 19552 884 19592
rect 10060 19552 10100 19592
rect 21004 19552 21044 19592
rect 10828 19468 10868 19508
rect 11020 19468 11060 19508
rect 1324 19384 1364 19424
rect 8236 19384 8276 19424
rect 2860 19216 2900 19256
rect 10732 19216 10772 19256
rect 12844 19216 12884 19256
rect 14188 19216 14228 19256
rect 14956 19216 14996 19256
rect 20524 19216 20564 19256
rect 4396 19132 4436 19172
rect 5356 19132 5396 19172
rect 16684 19132 16724 19172
rect 172 19048 212 19088
rect 6412 19048 6452 19088
rect 12076 19048 12116 19088
rect 19468 19132 19508 19172
rect 18700 19048 18740 19088
rect 2092 18964 2132 19004
rect 11884 18964 11924 19004
rect 12172 18964 12212 19004
rect 16876 18964 16916 19004
rect 3148 18880 3188 18920
rect 4396 18880 4436 18920
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 6124 18880 6164 18920
rect 11500 18880 11540 18920
rect 13900 18880 13940 18920
rect 14092 18880 14132 18920
rect 17164 18880 17204 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 6412 18796 6452 18836
rect 9964 18796 10004 18836
rect 16396 18796 16436 18836
rect 5644 18712 5684 18752
rect 14380 18712 14420 18752
rect 10156 18628 10196 18668
rect 12460 18544 12500 18584
rect 16492 18628 16532 18668
rect 21004 18628 21044 18668
rect 12652 18544 12692 18584
rect 17164 18544 17204 18584
rect 12268 18460 12308 18500
rect 1228 18376 1268 18416
rect 5740 18376 5780 18416
rect 13420 18376 13460 18416
rect 1708 18292 1748 18332
rect 4780 18292 4820 18332
rect 11692 18292 11732 18332
rect 14956 18292 14996 18332
rect 18508 18544 18548 18584
rect 19468 18544 19508 18584
rect 20620 18376 20660 18416
rect 19372 18292 19412 18332
rect 21196 18208 21236 18248
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 11596 18124 11636 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 844 18040 884 18080
rect 4396 18040 4436 18080
rect 19660 18040 19700 18080
rect 16396 17956 16436 17996
rect 19948 17956 19988 17996
rect 556 17872 596 17912
rect 1324 17872 1364 17912
rect 14380 17872 14420 17912
rect 19564 17872 19604 17912
rect 2476 17788 2516 17828
rect 1804 17704 1844 17744
rect 4108 17788 4148 17828
rect 5452 17788 5492 17828
rect 17644 17788 17684 17828
rect 19756 17788 19796 17828
rect 2380 17704 2420 17744
rect 2668 17704 2708 17744
rect 4492 17704 4532 17744
rect 4780 17704 4820 17744
rect 9004 17704 9044 17744
rect 9196 17704 9236 17744
rect 9580 17704 9620 17744
rect 14188 17704 14228 17744
rect 556 17620 596 17660
rect 844 17620 884 17660
rect 9964 17620 10004 17660
rect 10156 17620 10196 17660
rect 10348 17620 10388 17660
rect 13708 17620 13748 17660
rect 13900 17620 13940 17660
rect 14956 17704 14996 17744
rect 2764 17536 2804 17576
rect 4588 17452 4628 17492
rect 6988 17452 7028 17492
rect 13612 17452 13652 17492
rect 16876 17620 16916 17660
rect 19852 17620 19892 17660
rect 20620 17536 20660 17576
rect 14092 17452 14132 17492
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 6892 17368 6932 17408
rect 9196 17368 9236 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 1036 17284 1076 17324
rect 5644 17284 5684 17324
rect 6412 17284 6452 17324
rect 2284 17200 2324 17240
rect 5740 17200 5780 17240
rect 17452 17200 17492 17240
rect 4108 17116 4148 17156
rect 5548 17116 5588 17156
rect 15916 17116 15956 17156
rect 1324 17032 1364 17072
rect 6412 17032 6452 17072
rect 16972 16948 17012 16988
rect 1228 16864 1268 16904
rect 13900 16864 13940 16904
rect 1132 16780 1172 16820
rect 16012 16780 16052 16820
rect 4396 16696 4436 16736
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 12844 16612 12884 16652
rect 14188 16612 14228 16652
rect 15340 16612 15380 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 1804 16528 1844 16568
rect 4300 16528 4340 16568
rect 17644 16528 17684 16568
rect 1324 16444 1364 16484
rect 940 16360 980 16400
rect 4108 16360 4148 16400
rect 4492 16360 4532 16400
rect 6412 16360 6452 16400
rect 8716 16360 8756 16400
rect 11500 16360 11540 16400
rect 12556 16360 12596 16400
rect 19564 16360 19604 16400
rect 1516 16276 1556 16316
rect 3436 16276 3476 16316
rect 13324 16192 13364 16232
rect 13900 16192 13940 16232
rect 14956 16192 14996 16232
rect 16588 16192 16628 16232
rect 15628 16108 15668 16148
rect 9580 16024 9620 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 10540 15856 10580 15896
rect 13420 15856 13460 15896
rect 844 15772 884 15812
rect 14572 15856 14612 15896
rect 16012 15856 16052 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20716 15856 20756 15896
rect 12556 15772 12596 15812
rect 17356 15772 17396 15812
rect 4108 15688 4148 15728
rect 6988 15520 7028 15560
rect 7180 15520 7220 15560
rect 1804 15436 1844 15476
rect 7564 15352 7604 15392
rect 8908 15604 8948 15644
rect 10924 15604 10964 15644
rect 19660 15604 19700 15644
rect 20524 15604 20564 15644
rect 11596 15520 11636 15560
rect 15820 15520 15860 15560
rect 19372 15520 19412 15560
rect 19756 15520 19796 15560
rect 14188 15436 14228 15476
rect 15052 15436 15092 15476
rect 15916 15436 15956 15476
rect 9484 15352 9524 15392
rect 19276 15352 19316 15392
rect 19564 15352 19604 15392
rect 3628 15268 3668 15308
rect 5548 15268 5588 15308
rect 7660 15184 7700 15224
rect 8044 15184 8084 15224
rect 15820 15184 15860 15224
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 13420 15100 13460 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 11308 15016 11348 15056
rect 19852 15016 19892 15056
rect 10156 14932 10196 14972
rect 13900 14932 13940 14972
rect 1516 14848 1556 14888
rect 4300 14848 4340 14888
rect 11020 14848 11060 14888
rect 14668 14848 14708 14888
rect 15436 14848 15476 14888
rect 16588 14848 16628 14888
rect 20812 14848 20852 14888
rect 3724 14764 3764 14804
rect 11116 14764 11156 14804
rect 1900 14680 1940 14720
rect 13708 14680 13748 14720
rect 14380 14680 14420 14720
rect 19756 14680 19796 14720
rect 4780 14596 4820 14636
rect 8908 14596 8948 14636
rect 13324 14596 13364 14636
rect 13612 14596 13652 14636
rect 19468 14596 19508 14636
rect 5740 14512 5780 14552
rect 6412 14512 6452 14552
rect 16108 14512 16148 14552
rect 21100 14512 21140 14552
rect 3148 14428 3188 14468
rect 12172 14428 12212 14468
rect 17164 14428 17204 14468
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 9196 14344 9236 14384
rect 16300 14344 16340 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 3148 14260 3188 14300
rect 20908 14260 20948 14300
rect 4204 14176 4244 14216
rect 5452 14176 5492 14216
rect 6988 14176 7028 14216
rect 8908 14092 8948 14132
rect 17164 14092 17204 14132
rect 16108 14008 16148 14048
rect 1324 13924 1364 13964
rect 2380 13924 2420 13964
rect 3436 13924 3476 13964
rect 10156 13924 10196 13964
rect 17644 13924 17684 13964
rect 1132 13840 1172 13880
rect 10060 13840 10100 13880
rect 18316 13840 18356 13880
rect 18700 13840 18740 13880
rect 19852 13840 19892 13880
rect 1996 13756 2036 13796
rect 2476 13756 2516 13796
rect 5836 13756 5876 13796
rect 11308 13756 11348 13796
rect 14092 13756 14132 13796
rect 15436 13756 15476 13796
rect 17068 13756 17108 13796
rect 18604 13756 18644 13796
rect 1996 13588 2036 13628
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 10348 13588 10388 13628
rect 11020 13588 11060 13628
rect 1804 13504 1844 13544
rect 12364 13504 12404 13544
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 9676 13420 9716 13460
rect 10540 13420 10580 13460
rect 19564 13420 19604 13460
rect 1708 13336 1748 13376
rect 18700 13336 18740 13376
rect 19276 13336 19316 13376
rect 11596 13252 11636 13292
rect 16684 13252 16724 13292
rect 1516 13168 1556 13208
rect 4492 13168 4532 13208
rect 5740 13168 5780 13208
rect 8236 13168 8276 13208
rect 8524 13168 8564 13208
rect 4588 13084 4628 13124
rect 10444 13168 10484 13208
rect 11116 13084 11156 13124
rect 16300 13084 16340 13124
rect 2476 13000 2516 13040
rect 4492 13000 4532 13040
rect 19372 13000 19412 13040
rect 2188 12916 2228 12956
rect 20524 13168 20564 13208
rect 7948 12916 7988 12956
rect 17164 12916 17204 12956
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 17548 12832 17588 12872
rect 19468 12832 19508 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 9580 12748 9620 12788
rect 16396 12748 16436 12788
rect 2092 12664 2132 12704
rect 9676 12664 9716 12704
rect 8428 12580 8468 12620
rect 8908 12580 8948 12620
rect 12172 12580 12212 12620
rect 17836 12580 17876 12620
rect 2956 12496 2996 12536
rect 18412 12580 18452 12620
rect 20620 12580 20660 12620
rect 4108 12412 4148 12452
rect 6508 12412 6548 12452
rect 3148 12244 3188 12284
rect 3436 12244 3476 12284
rect 4108 12244 4148 12284
rect 9676 12412 9716 12452
rect 15916 12412 15956 12452
rect 19756 12412 19796 12452
rect 9580 12328 9620 12368
rect 5548 12244 5588 12284
rect 7852 12244 7892 12284
rect 10444 12244 10484 12284
rect 11500 12244 11540 12284
rect 10348 12160 10388 12200
rect 16972 12160 17012 12200
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 9196 12076 9236 12116
rect 13996 12076 14036 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 7372 11992 7412 12032
rect 11308 11992 11348 12032
rect 17356 11992 17396 12032
rect 8044 11908 8084 11948
rect 7564 11824 7604 11864
rect 8428 11824 8468 11864
rect 9196 11824 9236 11864
rect 13900 11824 13940 11864
rect 16684 11824 16724 11864
rect 1228 11656 1268 11696
rect 5740 11740 5780 11780
rect 10444 11740 10484 11780
rect 4204 11656 4244 11696
rect 2092 11488 2132 11528
rect 7948 11656 7988 11696
rect 10732 11656 10772 11696
rect 9292 11572 9332 11612
rect 1420 11404 1460 11444
rect 7276 11488 7316 11528
rect 9580 11488 9620 11528
rect 8428 11404 8468 11444
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 5932 11320 5972 11360
rect 15436 11572 15476 11612
rect 16108 11488 16148 11528
rect 17452 11404 17492 11444
rect 6700 11320 6740 11360
rect 7660 11320 7700 11360
rect 11308 11320 11348 11360
rect 16108 11320 16148 11360
rect 5740 11236 5780 11276
rect 7276 11236 7316 11276
rect 7564 11236 7604 11276
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 11980 11152 12020 11192
rect 18124 11152 18164 11192
rect 3052 11068 3092 11108
rect 5740 11068 5780 11108
rect 15340 11068 15380 11108
rect 7852 10984 7892 11024
rect 13036 10984 13076 11024
rect 5548 10900 5588 10940
rect 11500 10900 11540 10940
rect 8812 10816 8852 10856
rect 9580 10816 9620 10856
rect 11596 10816 11636 10856
rect 11788 10648 11828 10688
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 10540 10564 10580 10604
rect 16300 10564 16340 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 11116 10480 11156 10520
rect 15244 10480 15284 10520
rect 15436 10480 15476 10520
rect 20620 10480 20660 10520
rect 5740 10396 5780 10436
rect 7660 10396 7700 10436
rect 17164 10396 17204 10436
rect 8812 10228 8852 10268
rect 11020 10312 11060 10352
rect 11884 10312 11924 10352
rect 12364 10312 12404 10352
rect 13036 10312 13076 10352
rect 19468 10312 19508 10352
rect 12748 10228 12788 10268
rect 3436 10144 3476 10184
rect 10348 10144 10388 10184
rect 19468 10144 19508 10184
rect 20716 10144 20756 10184
rect 4108 10060 4148 10100
rect 7948 10060 7988 10100
rect 11116 10060 11156 10100
rect 12076 10060 12116 10100
rect 13324 10060 13364 10100
rect 9196 9976 9236 10016
rect 11308 9976 11348 10016
rect 4588 9892 4628 9932
rect 18508 9892 18548 9932
rect 1228 9808 1268 9848
rect 3436 9808 3476 9848
rect 4300 9808 4340 9848
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 11116 9808 11156 9848
rect 19564 9892 19604 9932
rect 11788 9808 11828 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 1516 9724 1556 9764
rect 3148 9640 3188 9680
rect 4396 9640 4436 9680
rect 9580 9640 9620 9680
rect 10348 9724 10388 9764
rect 13900 9724 13940 9764
rect 10540 9640 10580 9680
rect 1900 9556 1940 9596
rect 2188 9556 2228 9596
rect 3052 9556 3092 9596
rect 10636 9556 10676 9596
rect 11020 9640 11060 9680
rect 12556 9640 12596 9680
rect 13708 9640 13748 9680
rect 3820 9472 3860 9512
rect 9580 9472 9620 9512
rect 15436 9304 15476 9344
rect 16396 9304 16436 9344
rect 1036 9220 1076 9260
rect 9676 9220 9716 9260
rect 9868 9220 9908 9260
rect 15244 9220 15284 9260
rect 18700 9388 18740 9428
rect 16204 9136 16244 9176
rect 18124 9136 18164 9176
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 4204 9052 4244 9092
rect 12364 9052 12404 9092
rect 12556 9052 12596 9092
rect 13324 9052 13364 9092
rect 18028 9052 18068 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 6316 8968 6356 9008
rect 5740 8884 5780 8924
rect 6124 8884 6164 8924
rect 12652 8968 12692 9008
rect 17068 8968 17108 9008
rect 10540 8884 10580 8924
rect 20812 8884 20852 8924
rect 6700 8800 6740 8840
rect 9196 8800 9236 8840
rect 17548 8800 17588 8840
rect 18796 8800 18836 8840
rect 21388 8800 21428 8840
rect 652 8716 692 8756
rect 12076 8716 12116 8756
rect 12364 8716 12404 8756
rect 12652 8716 12692 8756
rect 1228 8632 1268 8672
rect 2188 8632 2228 8672
rect 15340 8632 15380 8672
rect 17452 8632 17492 8672
rect 748 8548 788 8588
rect 12268 8548 12308 8588
rect 18124 8548 18164 8588
rect 6892 8464 6932 8504
rect 11980 8464 12020 8504
rect 12748 8464 12788 8504
rect 18700 8464 18740 8504
rect 19948 8464 19988 8504
rect 2380 8380 2420 8420
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 5740 8296 5780 8336
rect 10540 8296 10580 8336
rect 5644 8212 5684 8252
rect 13900 8296 13940 8336
rect 14092 8296 14132 8336
rect 15820 8296 15860 8336
rect 16204 8296 16244 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 15244 8212 15284 8252
rect 18124 8128 18164 8168
rect 19948 8128 19988 8168
rect 12844 8044 12884 8084
rect 18412 8044 18452 8084
rect 19564 8044 19604 8084
rect 4108 7876 4148 7916
rect 4396 7876 4436 7916
rect 8044 7960 8084 8000
rect 8236 7960 8276 8000
rect 17260 7960 17300 8000
rect 9868 7876 9908 7916
rect 13900 7876 13940 7916
rect 1132 7792 1172 7832
rect 4204 7792 4244 7832
rect 11788 7792 11828 7832
rect 2188 7708 2228 7748
rect 12172 7708 12212 7748
rect 9484 7624 9524 7664
rect 11596 7624 11636 7664
rect 16300 7624 16340 7664
rect 18124 7624 18164 7664
rect 18700 7624 18740 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 9196 7540 9236 7580
rect 11980 7540 12020 7580
rect 12844 7540 12884 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 9292 7456 9332 7496
rect 21004 7456 21044 7496
rect 2956 7372 2996 7412
rect 5644 7372 5684 7412
rect 8044 7372 8084 7412
rect 18700 7372 18740 7412
rect 15340 7288 15380 7328
rect 15628 7288 15668 7328
rect 7372 7204 7412 7244
rect 4300 7120 4340 7160
rect 1516 6952 1556 6992
rect 364 6868 404 6908
rect 8524 7204 8564 7244
rect 12652 7204 12692 7244
rect 6508 7120 6548 7160
rect 9004 7120 9044 7160
rect 14572 7120 14612 7160
rect 19468 7120 19508 7160
rect 7564 7036 7604 7076
rect 11404 7036 11444 7076
rect 8044 6952 8084 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 16396 6784 16436 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 1996 6616 2036 6656
rect 11596 6616 11636 6656
rect 12364 6616 12404 6656
rect 15340 6616 15380 6656
rect 16684 6700 16724 6740
rect 16588 6616 16628 6656
rect 14572 6532 14612 6572
rect 16492 6532 16532 6572
rect 3820 6448 3860 6488
rect 7564 6448 7604 6488
rect 13036 6448 13076 6488
rect 15052 6448 15092 6488
rect 20620 6448 20660 6488
rect 7660 6364 7700 6404
rect 8812 6364 8852 6404
rect 11788 6364 11828 6404
rect 8524 6280 8564 6320
rect 14860 6280 14900 6320
rect 16588 6280 16628 6320
rect 19564 6280 19604 6320
rect 2572 6196 2612 6236
rect 10348 6196 10388 6236
rect 14188 6196 14228 6236
rect 15724 6196 15764 6236
rect 16108 6196 16148 6236
rect 15916 6112 15956 6152
rect 2380 6028 2420 6068
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 10156 5860 10196 5900
rect 11980 6028 12020 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 460 5776 500 5816
rect 18892 5776 18932 5816
rect 19276 5776 19316 5816
rect 10444 5608 10484 5648
rect 11788 5608 11828 5648
rect 7468 5524 7508 5564
rect 12460 5524 12500 5564
rect 1804 5440 1844 5480
rect 10252 5440 10292 5480
rect 12076 5440 12116 5480
rect 8812 5356 8852 5396
rect 10924 5356 10964 5396
rect 17068 5356 17108 5396
rect 172 5272 212 5312
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 18892 5272 18932 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 2188 5188 2228 5228
rect 7468 5188 7508 5228
rect 13900 5188 13940 5228
rect 16492 5104 16532 5144
rect 1420 5020 1460 5060
rect 7468 5020 7508 5060
rect 8428 4936 8468 4976
rect 8716 4936 8756 4976
rect 9580 4936 9620 4976
rect 9964 4936 10004 4976
rect 12172 4936 12212 4976
rect 12364 4936 12404 4976
rect 15244 4936 15284 4976
rect 21292 4852 21332 4892
rect 18412 4768 18452 4808
rect 2284 4684 2324 4724
rect 4972 4684 5012 4724
rect 17548 4684 17588 4724
rect 5548 4600 5588 4640
rect 9292 4600 9332 4640
rect 10732 4600 10772 4640
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 12460 4516 12500 4556
rect 17740 4516 17780 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 76 4432 116 4472
rect 20140 4432 20180 4472
rect 17836 4348 17876 4388
rect 5740 4264 5780 4304
rect 6124 4264 6164 4304
rect 8236 4264 8276 4304
rect 9004 4264 9044 4304
rect 16684 4264 16724 4304
rect 4588 4180 4628 4220
rect 4780 4180 4820 4220
rect 4108 4096 4148 4136
rect 11596 4180 11636 4220
rect 17068 4180 17108 4220
rect 21100 4180 21140 4220
rect 4300 4096 4340 4136
rect 8716 4096 8756 4136
rect 1900 3928 1940 3968
rect 6700 3928 6740 3968
rect 556 3760 596 3800
rect 1516 3760 1556 3800
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 7372 3844 7412 3884
rect 9676 3844 9716 3884
rect 15244 4096 15284 4136
rect 19948 4096 19988 4136
rect 19564 3844 19604 3884
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 2476 3676 2516 3716
rect 17164 3676 17204 3716
rect 1420 3592 1460 3632
rect 1612 3592 1652 3632
rect 3244 3592 3284 3632
rect 7564 3592 7604 3632
rect 15724 3592 15764 3632
rect 16396 3592 16436 3632
rect 17260 3592 17300 3632
rect 14956 3508 14996 3548
rect 8044 3424 8084 3464
rect 10156 3424 10196 3464
rect 10348 3424 10388 3464
rect 12652 3424 12692 3464
rect 6700 3340 6740 3380
rect 9772 3340 9812 3380
rect 10732 3340 10772 3380
rect 20524 3424 20564 3464
rect 20812 3424 20852 3464
rect 12172 3340 12212 3380
rect 6892 3256 6932 3296
rect 14956 3256 14996 3296
rect 15628 3256 15668 3296
rect 18604 3256 18644 3296
rect 19564 3256 19604 3296
rect 19948 3256 19988 3296
rect 2188 3172 2228 3212
rect 12556 3172 12596 3212
rect 17452 3172 17492 3212
rect 15244 3088 15284 3128
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 19756 3088 19796 3128
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 7660 2920 7700 2960
rect 10924 2836 10964 2876
rect 17260 2836 17300 2876
rect 5932 2752 5972 2792
rect 9100 2752 9140 2792
rect 11788 2752 11828 2792
rect 16204 2668 16244 2708
rect 2668 2584 2708 2624
rect 6316 2584 6356 2624
rect 6892 2584 6932 2624
rect 9868 2584 9908 2624
rect 17068 2584 17108 2624
rect 17548 2584 17588 2624
rect 5836 2500 5876 2540
rect 6508 2500 6548 2540
rect 7564 2500 7604 2540
rect 20140 2500 20180 2540
rect 5932 2416 5972 2456
rect 10252 2416 10292 2456
rect 16780 2416 16820 2456
rect 18412 2416 18452 2456
rect 5740 2332 5780 2372
rect 7276 2332 7316 2372
rect 4396 2248 4436 2288
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 8428 2248 8468 2288
rect 17740 2332 17780 2372
rect 8716 2248 8756 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 5644 2164 5684 2204
rect 8812 2164 8852 2204
rect 20620 2080 20660 2120
rect 2092 1912 2132 1952
rect 6508 1912 6548 1952
rect 7180 1912 7220 1952
rect 9580 1912 9620 1952
rect 16780 1912 16820 1952
rect 6892 1828 6932 1868
rect 17740 1828 17780 1868
rect 18604 1744 18644 1784
rect 20716 1744 20756 1784
rect 2860 1576 2900 1616
rect 15436 1576 15476 1616
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 11212 1492 11252 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 5356 1324 5396 1364
rect 8044 1324 8084 1364
rect 2764 1240 2804 1280
rect 3340 1240 3380 1280
rect 6220 1240 6260 1280
rect 6604 1240 6644 1280
rect 6796 1240 6836 1280
rect 6988 1240 7028 1280
rect 7180 1240 7220 1280
rect 7756 1240 7796 1280
rect 8140 1240 8180 1280
rect 8332 1240 8372 1280
rect 8908 1240 8948 1280
rect 13324 1240 13364 1280
rect 14284 1240 14324 1280
rect 14476 1240 14516 1280
rect 14668 1240 14708 1280
rect 16972 1240 17012 1280
rect 17164 1240 17204 1280
rect 17932 1240 17972 1280
rect 18508 1240 18548 1280
rect 18700 1240 18740 1280
rect 1516 1156 1556 1196
rect 5260 1156 5300 1196
rect 9388 1156 9428 1196
rect 15148 1156 15188 1196
rect 16300 1156 16340 1196
rect 4300 1072 4340 1112
rect 3532 904 3572 944
rect 6028 904 6068 944
rect 6412 904 6452 944
rect 8620 904 8660 944
rect 12556 904 12596 944
rect 12940 904 12980 944
rect 13516 904 13556 944
rect 13708 904 13748 944
rect 17644 904 17684 944
rect 18220 904 18260 944
rect 7948 820 7988 860
rect 13132 820 13172 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 16012 736 16052 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 20524 736 20564 776
rect 5452 652 5492 692
rect 7084 652 7124 692
rect 13900 652 13940 692
rect 15340 652 15380 692
rect 4684 568 4724 608
rect 5548 568 5588 608
rect 7468 568 7508 608
rect 15148 568 15188 608
rect 15724 568 15764 608
rect 18892 400 18932 440
rect 19660 400 19700 440
rect 12172 316 12212 356
rect 15628 232 15668 272
rect 5068 64 5108 104
rect 17548 64 17588 104
rect 18124 64 18164 104
<< metal4 >>
rect 15532 42944 15572 42953
rect 1420 42860 1460 42869
rect 460 42524 500 42533
rect 268 40508 308 40517
rect 76 25976 116 25987
rect 76 25901 116 25936
rect 75 25892 117 25901
rect 75 25852 76 25892
rect 116 25852 117 25892
rect 75 25843 117 25852
rect 76 23960 116 23969
rect 76 4472 116 23920
rect 268 22616 308 40468
rect 268 22567 308 22576
rect 364 35972 404 35981
rect 268 20432 308 20441
rect 172 19088 212 19097
rect 172 5312 212 19048
rect 268 18509 308 20392
rect 267 18500 309 18509
rect 267 18460 268 18500
rect 308 18460 309 18500
rect 267 18451 309 18460
rect 364 6908 404 35932
rect 460 22028 500 42484
rect 1036 42440 1076 42449
rect 555 35888 597 35897
rect 555 35848 556 35888
rect 596 35848 597 35888
rect 555 35839 597 35848
rect 556 23960 596 35839
rect 844 35132 884 35141
rect 556 23911 596 23920
rect 652 30344 692 30353
rect 460 21979 500 21988
rect 364 6859 404 6868
rect 460 21524 500 21533
rect 460 5816 500 21484
rect 555 17912 597 17921
rect 555 17872 556 17912
rect 596 17872 597 17912
rect 555 17863 597 17872
rect 556 17778 596 17863
rect 460 5767 500 5776
rect 556 17660 596 17669
rect 172 5263 212 5272
rect 76 4423 116 4432
rect 556 3800 596 17620
rect 652 8756 692 30304
rect 652 8707 692 8716
rect 748 24800 788 24809
rect 748 8588 788 24760
rect 844 19592 884 35092
rect 1036 29000 1076 42400
rect 940 28960 1076 29000
rect 1132 41516 1172 41525
rect 940 22532 980 28960
rect 1035 23288 1077 23297
rect 1035 23248 1036 23288
rect 1076 23248 1077 23288
rect 1035 23239 1077 23248
rect 940 22483 980 22492
rect 1036 21944 1076 23239
rect 1036 21895 1076 21904
rect 1132 21776 1172 41476
rect 1324 40424 1364 40433
rect 1324 39080 1364 40384
rect 1228 36056 1268 36065
rect 1228 30017 1268 36016
rect 1324 35636 1364 39040
rect 1420 37652 1460 42820
rect 7564 42692 7604 42701
rect 6795 42272 6837 42281
rect 6795 42232 6796 42272
rect 6836 42232 6837 42272
rect 6795 42223 6837 42232
rect 6412 42020 6452 42029
rect 5452 41936 5492 41945
rect 3148 41600 3188 41609
rect 3052 41264 3092 41273
rect 2284 40508 2324 40517
rect 2188 39752 2228 39761
rect 2092 39248 2132 39257
rect 1900 39080 1940 39089
rect 1804 38996 1844 39005
rect 1420 37603 1460 37612
rect 1516 38156 1556 38165
rect 1420 35636 1460 35645
rect 1324 35596 1420 35636
rect 1323 34544 1365 34553
rect 1323 34504 1324 34544
rect 1364 34504 1365 34544
rect 1323 34495 1365 34504
rect 1324 32276 1364 34495
rect 1227 30008 1269 30017
rect 1227 29968 1228 30008
rect 1268 29968 1269 30008
rect 1227 29959 1269 29968
rect 1324 27404 1364 32236
rect 1420 32108 1460 35596
rect 1420 32059 1460 32068
rect 1516 30773 1556 38116
rect 1708 38156 1748 38165
rect 1708 37652 1748 38116
rect 1612 35888 1652 35897
rect 1612 34628 1652 35848
rect 1612 32108 1652 34588
rect 1612 32059 1652 32068
rect 1708 31940 1748 37612
rect 1612 31900 1748 31940
rect 1515 30764 1557 30773
rect 1515 30724 1516 30764
rect 1556 30724 1557 30764
rect 1515 30715 1557 30724
rect 1324 26564 1364 27364
rect 1324 26515 1364 26524
rect 1420 26984 1460 26993
rect 1228 26228 1268 26237
rect 1228 25901 1268 26188
rect 1420 25976 1460 26944
rect 1227 25892 1269 25901
rect 1227 25852 1228 25892
rect 1268 25852 1269 25892
rect 1227 25843 1269 25852
rect 1228 23120 1268 25843
rect 1228 23071 1268 23080
rect 1227 22448 1269 22457
rect 1227 22408 1228 22448
rect 1268 22408 1269 22448
rect 1227 22399 1269 22408
rect 1228 22314 1268 22399
rect 1132 21727 1172 21736
rect 1420 21524 1460 25936
rect 1420 21475 1460 21484
rect 1516 24128 1556 24137
rect 1516 21020 1556 24088
rect 1516 20971 1556 20980
rect 1420 20852 1460 20861
rect 1227 19928 1269 19937
rect 1227 19888 1228 19928
rect 1268 19888 1269 19928
rect 1227 19879 1269 19888
rect 1228 19794 1268 19879
rect 844 19543 884 19552
rect 1324 19424 1364 19433
rect 1227 18416 1269 18425
rect 1227 18376 1228 18416
rect 1268 18376 1269 18416
rect 1227 18367 1269 18376
rect 1228 18282 1268 18367
rect 844 18080 884 18089
rect 844 17660 884 18040
rect 1324 17912 1364 19384
rect 1324 17863 1364 17872
rect 844 17611 884 17620
rect 1420 17585 1460 20812
rect 1419 17576 1461 17585
rect 1419 17536 1420 17576
rect 1460 17536 1461 17576
rect 1419 17527 1461 17536
rect 1036 17324 1076 17333
rect 939 16400 981 16409
rect 939 16360 940 16400
rect 980 16360 981 16400
rect 939 16351 981 16360
rect 940 16266 980 16351
rect 843 15812 885 15821
rect 843 15772 844 15812
rect 884 15772 885 15812
rect 843 15763 885 15772
rect 844 15678 884 15763
rect 1036 9260 1076 17284
rect 1324 17072 1364 17081
rect 1227 16904 1269 16913
rect 1227 16864 1228 16904
rect 1268 16864 1269 16904
rect 1227 16855 1269 16864
rect 1132 16820 1172 16829
rect 1132 13880 1172 16780
rect 1228 16770 1268 16855
rect 1324 16652 1364 17032
rect 1132 13831 1172 13840
rect 1228 16612 1364 16652
rect 1131 11948 1173 11957
rect 1131 11908 1132 11948
rect 1172 11908 1173 11948
rect 1131 11899 1173 11908
rect 1036 9211 1076 9220
rect 748 8539 788 8548
rect 1132 7832 1172 11899
rect 1228 11696 1268 16612
rect 1324 16484 1364 16493
rect 1324 13964 1364 16444
rect 1516 16316 1556 16325
rect 1324 13915 1364 13924
rect 1420 16276 1516 16316
rect 1228 11647 1268 11656
rect 1420 11444 1460 16276
rect 1516 16267 1556 16276
rect 1515 14888 1557 14897
rect 1515 14848 1516 14888
rect 1556 14848 1557 14888
rect 1515 14839 1557 14848
rect 1516 14754 1556 14839
rect 1420 11395 1460 11404
rect 1516 13208 1556 13217
rect 1227 10016 1269 10025
rect 1227 9976 1228 10016
rect 1268 9976 1269 10016
rect 1227 9967 1269 9976
rect 1228 9848 1268 9967
rect 1516 9932 1556 13168
rect 1228 9799 1268 9808
rect 1420 9892 1556 9932
rect 1420 9521 1460 9892
rect 1516 9764 1556 9773
rect 1419 9512 1461 9521
rect 1419 9472 1420 9512
rect 1460 9472 1461 9512
rect 1419 9463 1461 9472
rect 1228 8672 1268 8683
rect 1228 8597 1268 8632
rect 1227 8588 1269 8597
rect 1227 8548 1228 8588
rect 1268 8548 1269 8588
rect 1227 8539 1269 8548
rect 1132 7783 1172 7792
rect 1420 5060 1460 9463
rect 1420 5011 1460 5020
rect 1516 6992 1556 9724
rect 556 3751 596 3760
rect 1516 3800 1556 6952
rect 1516 3751 1556 3760
rect 1419 3632 1461 3641
rect 1419 3592 1420 3632
rect 1460 3592 1461 3632
rect 1419 3583 1461 3592
rect 1612 3632 1652 31900
rect 1707 31772 1749 31781
rect 1707 31732 1708 31772
rect 1748 31732 1749 31772
rect 1707 31723 1749 31732
rect 1708 18593 1748 31723
rect 1804 26984 1844 38956
rect 1900 35972 1940 39040
rect 1996 38744 2036 38753
rect 1996 38081 2036 38704
rect 1995 38072 2037 38081
rect 1995 38032 1996 38072
rect 2036 38032 2037 38072
rect 1995 38023 2037 38032
rect 1995 36812 2037 36821
rect 1995 36772 1996 36812
rect 2036 36772 2037 36812
rect 1995 36763 2037 36772
rect 1900 35923 1940 35932
rect 1996 35804 2036 36763
rect 1900 35764 2036 35804
rect 1900 34964 1940 35764
rect 1900 34208 1940 34924
rect 1900 31781 1940 34168
rect 1899 31772 1941 31781
rect 1899 31732 1900 31772
rect 1940 31732 1941 31772
rect 1899 31723 1941 31732
rect 1804 26935 1844 26944
rect 1996 29756 2036 29765
rect 1996 27992 2036 29716
rect 1900 26396 1940 26405
rect 1804 24212 1844 24221
rect 1804 21272 1844 24172
rect 1900 23624 1940 26356
rect 1900 23575 1940 23584
rect 1899 21776 1941 21785
rect 1899 21736 1900 21776
rect 1940 21736 1941 21776
rect 1899 21727 1941 21736
rect 1900 21642 1940 21727
rect 1900 21272 1940 21281
rect 1804 21232 1900 21272
rect 1707 18584 1749 18593
rect 1707 18544 1708 18584
rect 1748 18544 1749 18584
rect 1707 18535 1749 18544
rect 1708 18332 1748 18341
rect 1708 13376 1748 18292
rect 1803 17744 1845 17753
rect 1803 17704 1804 17744
rect 1844 17704 1845 17744
rect 1803 17695 1845 17704
rect 1804 17610 1844 17695
rect 1804 16568 1844 16577
rect 1804 15476 1844 16528
rect 1804 15427 1844 15436
rect 1900 14720 1940 21232
rect 1708 13327 1748 13336
rect 1804 13544 1844 13553
rect 1804 5480 1844 13504
rect 1900 9773 1940 14680
rect 1996 13796 2036 27952
rect 2092 21524 2132 39208
rect 2188 36653 2228 39712
rect 2187 36644 2229 36653
rect 2187 36604 2188 36644
rect 2228 36604 2229 36644
rect 2187 36595 2229 36604
rect 2187 35720 2229 35729
rect 2187 35680 2188 35720
rect 2228 35680 2229 35720
rect 2187 35671 2229 35680
rect 2188 35586 2228 35671
rect 2188 35216 2228 35225
rect 2188 34796 2228 35176
rect 2188 34747 2228 34756
rect 2284 33116 2324 40468
rect 2956 40424 2996 40433
rect 2860 39752 2900 39761
rect 2380 39584 2420 39593
rect 2380 36821 2420 39544
rect 2764 38324 2804 38333
rect 2572 38156 2612 38165
rect 2476 37904 2516 37913
rect 2379 36812 2421 36821
rect 2379 36772 2380 36812
rect 2420 36772 2421 36812
rect 2379 36763 2421 36772
rect 2379 36644 2421 36653
rect 2379 36604 2380 36644
rect 2420 36604 2421 36644
rect 2379 36595 2421 36604
rect 2284 33067 2324 33076
rect 2188 32948 2228 32957
rect 2188 23036 2228 32908
rect 2284 32864 2324 32873
rect 2284 28841 2324 32824
rect 2380 29000 2420 36595
rect 2476 29756 2516 37864
rect 2572 37568 2612 38116
rect 2764 37904 2804 38284
rect 2764 37855 2804 37864
rect 2860 37736 2900 39712
rect 2572 37519 2612 37528
rect 2764 37696 2900 37736
rect 2572 36896 2612 36905
rect 2572 36476 2612 36856
rect 2572 36427 2612 36436
rect 2668 36812 2708 36821
rect 2668 35888 2708 36772
rect 2476 29707 2516 29716
rect 2572 33452 2612 33461
rect 2572 30932 2612 33412
rect 2572 29168 2612 30892
rect 2668 29429 2708 35848
rect 2764 35804 2804 37696
rect 2764 35755 2804 35764
rect 2860 36140 2900 36149
rect 2763 33032 2805 33041
rect 2763 32992 2764 33032
rect 2804 32992 2805 33032
rect 2763 32983 2805 32992
rect 2764 32864 2804 32983
rect 2764 32815 2804 32824
rect 2860 29840 2900 36100
rect 2956 34889 2996 40384
rect 3052 38912 3092 41224
rect 3052 38863 3092 38872
rect 3052 37232 3092 37241
rect 3052 36737 3092 37192
rect 3051 36728 3093 36737
rect 3051 36688 3052 36728
rect 3092 36688 3093 36728
rect 3051 36679 3093 36688
rect 3052 36560 3092 36569
rect 3052 36224 3092 36520
rect 3052 36175 3092 36184
rect 3052 34964 3092 34973
rect 2955 34880 2997 34889
rect 2955 34840 2956 34880
rect 2996 34840 2997 34880
rect 2955 34831 2997 34840
rect 2956 34712 2996 34721
rect 2956 31268 2996 34672
rect 3052 31940 3092 34924
rect 3052 31891 3092 31900
rect 2956 31228 3092 31268
rect 2955 30008 2997 30017
rect 2955 29968 2956 30008
rect 2996 29968 2997 30008
rect 2955 29959 2997 29968
rect 2667 29420 2709 29429
rect 2667 29380 2668 29420
rect 2708 29380 2709 29420
rect 2667 29371 2709 29380
rect 2860 29345 2900 29800
rect 2859 29336 2901 29345
rect 2859 29296 2860 29336
rect 2900 29296 2901 29336
rect 2859 29287 2901 29296
rect 2956 29336 2996 29959
rect 2572 29128 2708 29168
rect 2571 29000 2613 29009
rect 2380 28960 2516 29000
rect 2283 28832 2325 28841
rect 2283 28792 2284 28832
rect 2324 28792 2325 28832
rect 2283 28783 2325 28792
rect 2284 26741 2324 26826
rect 2283 26732 2325 26741
rect 2283 26692 2284 26732
rect 2324 26692 2325 26732
rect 2283 26683 2325 26692
rect 2188 22987 2228 22996
rect 2284 26564 2324 26573
rect 2092 21475 2132 21484
rect 2284 20180 2324 26524
rect 2380 25052 2420 25061
rect 2380 20516 2420 25012
rect 2476 24632 2516 28960
rect 2571 28960 2572 29000
rect 2612 28960 2613 29000
rect 2571 28951 2613 28960
rect 2476 24380 2516 24592
rect 2476 24331 2516 24340
rect 2380 20467 2420 20476
rect 2476 23204 2516 23213
rect 2284 20140 2420 20180
rect 1996 13747 2036 13756
rect 2092 19004 2132 19013
rect 1996 13628 2036 13637
rect 1899 9764 1941 9773
rect 1899 9724 1900 9764
rect 1940 9724 1941 9764
rect 1899 9715 1941 9724
rect 1804 5431 1844 5440
rect 1900 9596 1940 9605
rect 1900 3968 1940 9556
rect 1996 6656 2036 13588
rect 2092 12704 2132 18964
rect 2187 18584 2229 18593
rect 2187 18544 2188 18584
rect 2228 18544 2229 18584
rect 2187 18535 2229 18544
rect 2188 12956 2228 18535
rect 2380 17744 2420 20140
rect 2476 17828 2516 23164
rect 2572 20432 2612 28951
rect 2668 25304 2708 29128
rect 2859 28916 2901 28925
rect 2859 28876 2860 28916
rect 2900 28876 2901 28916
rect 2859 28867 2901 28876
rect 2763 28832 2805 28841
rect 2763 28792 2764 28832
rect 2804 28792 2805 28832
rect 2763 28783 2805 28792
rect 2668 25255 2708 25264
rect 2764 22784 2804 28783
rect 2764 22735 2804 22744
rect 2860 26144 2900 28867
rect 2667 22364 2709 22373
rect 2667 22324 2668 22364
rect 2708 22324 2709 22364
rect 2667 22315 2709 22324
rect 2668 22230 2708 22315
rect 2572 20383 2612 20392
rect 2476 17779 2516 17788
rect 2572 19844 2612 19853
rect 2380 17695 2420 17704
rect 2284 17240 2324 17249
rect 2284 12965 2324 17200
rect 2380 13964 2420 13973
rect 2188 12907 2228 12916
rect 2283 12956 2325 12965
rect 2283 12916 2284 12956
rect 2324 12916 2325 12956
rect 2283 12907 2325 12916
rect 2092 12655 2132 12664
rect 2380 12620 2420 13924
rect 2476 13796 2516 13805
rect 2476 13040 2516 13756
rect 2476 12991 2516 13000
rect 2475 12872 2517 12881
rect 2475 12832 2476 12872
rect 2516 12832 2517 12872
rect 2475 12823 2517 12832
rect 2188 12580 2420 12620
rect 1996 6607 2036 6616
rect 2092 11528 2132 11537
rect 1900 3919 1940 3928
rect 1612 3583 1652 3592
rect 1420 3498 1460 3583
rect 2092 1952 2132 11488
rect 2188 9596 2228 12580
rect 2283 9764 2325 9773
rect 2283 9724 2284 9764
rect 2324 9724 2325 9764
rect 2283 9715 2325 9724
rect 2188 9547 2228 9556
rect 2187 8672 2229 8681
rect 2187 8632 2188 8672
rect 2228 8632 2229 8672
rect 2187 8623 2229 8632
rect 2188 8538 2228 8623
rect 2188 7748 2228 7757
rect 2188 5228 2228 7708
rect 2188 5179 2228 5188
rect 2284 4724 2324 9715
rect 2380 8420 2420 8429
rect 2380 6068 2420 8380
rect 2380 6019 2420 6028
rect 2284 4675 2324 4684
rect 2476 3716 2516 12823
rect 2572 6236 2612 19804
rect 2860 19256 2900 26104
rect 2572 6187 2612 6196
rect 2668 17744 2708 17753
rect 2476 3667 2516 3676
rect 2187 3212 2229 3221
rect 2187 3172 2188 3212
rect 2228 3172 2229 3212
rect 2187 3163 2229 3172
rect 2188 3078 2228 3163
rect 2668 2717 2708 17704
rect 2764 17576 2804 17585
rect 2667 2708 2709 2717
rect 2667 2668 2668 2708
rect 2708 2668 2709 2708
rect 2667 2659 2709 2668
rect 2668 2624 2708 2659
rect 2668 2574 2708 2584
rect 2092 1903 2132 1912
rect 2764 1280 2804 17536
rect 2860 1616 2900 19216
rect 2956 19928 2996 29296
rect 3052 21608 3092 31228
rect 3148 27749 3188 41560
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 4204 40340 4244 40349
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 3532 38744 3572 38753
rect 3532 38417 3572 38704
rect 3531 38408 3573 38417
rect 3531 38368 3532 38408
rect 3572 38368 3573 38408
rect 3531 38359 3573 38368
rect 3340 38156 3380 38165
rect 3244 37148 3284 37157
rect 3244 32864 3284 37108
rect 3244 32815 3284 32824
rect 3340 32360 3380 38116
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3532 37484 3572 37493
rect 3532 35981 3572 37444
rect 3819 37232 3861 37241
rect 3819 37192 3820 37232
rect 3860 37192 3861 37232
rect 3819 37183 3861 37192
rect 3820 37098 3860 37183
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3531 35972 3573 35981
rect 3531 35932 3532 35972
rect 3572 35932 3573 35972
rect 3531 35923 3573 35932
rect 3628 35720 3668 35729
rect 3628 35225 3668 35680
rect 4108 35300 4148 35309
rect 3627 35216 3669 35225
rect 3627 35176 3628 35216
rect 3668 35176 3669 35216
rect 3627 35167 3669 35176
rect 3532 35048 3572 35057
rect 3435 34880 3477 34889
rect 3435 34840 3436 34880
rect 3476 34840 3477 34880
rect 3435 34831 3477 34840
rect 3340 32311 3380 32320
rect 3436 31016 3476 34831
rect 3532 34040 3572 35008
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3532 33991 3572 34000
rect 3628 34292 3668 34301
rect 3628 33452 3668 34252
rect 3532 33412 3668 33452
rect 3532 32864 3572 33412
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 3532 32815 3572 32824
rect 3436 30967 3476 30976
rect 3532 31940 3572 31949
rect 3436 30848 3476 30857
rect 3244 29672 3284 29681
rect 3244 29261 3284 29632
rect 3243 29252 3285 29261
rect 3243 29212 3244 29252
rect 3284 29212 3285 29252
rect 3243 29203 3285 29212
rect 3244 29118 3284 29203
rect 3339 29168 3381 29177
rect 3339 29128 3340 29168
rect 3380 29128 3381 29168
rect 3339 29119 3381 29128
rect 3340 29034 3380 29119
rect 3244 28832 3284 28841
rect 3244 27908 3284 28792
rect 3244 27859 3284 27868
rect 3436 28160 3476 30808
rect 3147 27740 3189 27749
rect 3147 27700 3148 27740
rect 3188 27700 3189 27740
rect 3147 27691 3189 27700
rect 3436 27488 3476 28120
rect 3052 21559 3092 21568
rect 3340 23036 3380 23045
rect 3244 21524 3284 21533
rect 2956 18341 2996 19888
rect 3148 20348 3188 20357
rect 3148 19928 3188 20308
rect 3148 19879 3188 19888
rect 3148 18920 3188 18929
rect 2955 18332 2997 18341
rect 2955 18292 2956 18332
rect 2996 18292 2997 18332
rect 2955 18283 2997 18292
rect 3148 14468 3188 18880
rect 3148 14419 3188 14428
rect 3148 14300 3188 14309
rect 2956 12536 2996 12545
rect 2956 7412 2996 12496
rect 3148 12284 3188 14260
rect 3052 11108 3092 11117
rect 3052 9596 3092 11068
rect 3148 9689 3188 12244
rect 3147 9680 3189 9689
rect 3147 9640 3148 9680
rect 3188 9640 3189 9680
rect 3147 9631 3189 9640
rect 3052 9547 3092 9556
rect 3148 9546 3188 9631
rect 2956 7363 2996 7372
rect 3244 3632 3284 21484
rect 3244 3583 3284 3592
rect 2860 1567 2900 1576
rect 2764 1231 2804 1240
rect 3340 1280 3380 22996
rect 3436 19844 3476 27448
rect 3532 27404 3572 31900
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3628 28412 3668 28421
rect 3628 28253 3668 28372
rect 4108 28412 4148 35260
rect 4204 32192 4244 40300
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 5356 39668 5396 39677
rect 5356 39509 5396 39628
rect 5355 39500 5397 39509
rect 5355 39460 5356 39500
rect 5396 39460 5397 39500
rect 5355 39451 5397 39460
rect 4204 32143 4244 32152
rect 4300 38744 4340 38753
rect 4300 29177 4340 38704
rect 4587 38744 4629 38753
rect 4587 38704 4588 38744
rect 4628 38704 4629 38744
rect 4587 38695 4629 38704
rect 4588 38610 4628 38695
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5356 38240 5396 38249
rect 4492 37232 4532 37241
rect 4492 36485 4532 37192
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4491 36476 4533 36485
rect 4491 36436 4492 36476
rect 4532 36436 4533 36476
rect 4491 36427 4533 36436
rect 4588 36224 4628 36233
rect 4396 35132 4436 35141
rect 3627 28244 3669 28253
rect 3627 28204 3628 28244
rect 3668 28204 3669 28244
rect 3627 28195 3669 28204
rect 4108 27908 4148 28372
rect 4108 27859 4148 27868
rect 4204 29168 4244 29177
rect 4107 27656 4149 27665
rect 4107 27616 4108 27656
rect 4148 27616 4149 27656
rect 4107 27607 4149 27616
rect 3532 27355 3572 27364
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 4108 27068 4148 27607
rect 3532 26480 3572 26489
rect 3532 25388 3572 26440
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3532 25339 3572 25348
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 4108 22541 4148 27028
rect 4204 24632 4244 29128
rect 4299 29168 4341 29177
rect 4299 29128 4300 29168
rect 4340 29128 4341 29168
rect 4299 29119 4341 29128
rect 4300 27572 4340 27581
rect 4300 26657 4340 27532
rect 4299 26648 4341 26657
rect 4299 26608 4300 26648
rect 4340 26608 4341 26648
rect 4299 26599 4341 26608
rect 4204 24583 4244 24592
rect 4300 26228 4340 26237
rect 4204 24380 4244 24389
rect 4107 22532 4149 22541
rect 4107 22492 4108 22532
rect 4148 22492 4149 22532
rect 4107 22483 4149 22492
rect 4107 22280 4149 22289
rect 4107 22240 4108 22280
rect 4148 22240 4149 22280
rect 4107 22231 4149 22240
rect 3436 19795 3476 19804
rect 3532 21776 3572 21785
rect 3436 16316 3476 16325
rect 3436 13964 3476 16276
rect 3436 13915 3476 13924
rect 3436 12284 3476 12293
rect 3436 10361 3476 12244
rect 3435 10352 3477 10361
rect 3435 10312 3436 10352
rect 3476 10312 3477 10352
rect 3435 10303 3477 10312
rect 3436 10184 3476 10193
rect 3436 9848 3476 10144
rect 3436 9799 3476 9808
rect 3340 1231 3380 1240
rect 1515 1196 1557 1205
rect 1515 1156 1516 1196
rect 1556 1156 1557 1196
rect 1515 1147 1557 1156
rect 1516 1062 1556 1147
rect 3532 944 3572 21736
rect 3723 21776 3765 21785
rect 3723 21736 3724 21776
rect 3764 21736 3765 21776
rect 3723 21727 3765 21736
rect 3724 21642 3764 21727
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 4108 17828 4148 22231
rect 4108 17779 4148 17788
rect 4108 17156 4148 17165
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 4108 16400 4148 17116
rect 4108 16351 4148 16360
rect 4108 15728 4148 15737
rect 3628 15317 3668 15402
rect 3627 15308 3669 15317
rect 3627 15268 3628 15308
rect 3668 15268 3669 15308
rect 3627 15259 3669 15268
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3723 14804 3765 14813
rect 3723 14764 3724 14804
rect 3764 14764 3765 14804
rect 3723 14755 3765 14764
rect 3724 14670 3764 14755
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 4108 12452 4148 15688
rect 4204 14216 4244 24340
rect 4300 22961 4340 26188
rect 4396 24716 4436 35092
rect 4492 34544 4532 34555
rect 4492 34469 4532 34504
rect 4491 34460 4533 34469
rect 4491 34420 4492 34460
rect 4532 34420 4533 34460
rect 4491 34411 4533 34420
rect 4588 33620 4628 36184
rect 4780 35888 4820 35897
rect 4780 35216 4820 35848
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4780 35167 4820 35176
rect 5260 35216 5300 35225
rect 5260 34973 5300 35176
rect 5259 34964 5301 34973
rect 5259 34924 5260 34964
rect 5300 34924 5301 34964
rect 5259 34915 5301 34924
rect 4683 34628 4725 34637
rect 4683 34588 4684 34628
rect 4724 34588 4725 34628
rect 4683 34579 4725 34588
rect 4684 34494 4724 34579
rect 4875 34460 4917 34469
rect 4875 34420 4876 34460
rect 4916 34420 4917 34460
rect 4875 34411 4917 34420
rect 4780 34376 4820 34385
rect 4780 34217 4820 34336
rect 4876 34326 4916 34411
rect 4779 34208 4821 34217
rect 4779 34168 4780 34208
rect 4820 34168 4821 34208
rect 4779 34159 4821 34168
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4588 27992 4628 33580
rect 4588 27943 4628 27952
rect 4684 32780 4724 32789
rect 4491 27740 4533 27749
rect 4491 27700 4492 27740
rect 4532 27700 4533 27740
rect 4491 27691 4533 27700
rect 4492 27606 4532 27691
rect 4588 25388 4628 25397
rect 4396 24676 4532 24716
rect 4395 24548 4437 24557
rect 4395 24508 4396 24548
rect 4436 24508 4437 24548
rect 4395 24499 4437 24508
rect 4299 22952 4341 22961
rect 4299 22912 4300 22952
rect 4340 22912 4341 22952
rect 4299 22903 4341 22912
rect 4300 22289 4340 22903
rect 4299 22280 4341 22289
rect 4299 22240 4300 22280
rect 4340 22240 4341 22280
rect 4299 22231 4341 22240
rect 4300 20852 4340 20861
rect 4300 19097 4340 20812
rect 4396 19172 4436 24499
rect 4492 22196 4532 24676
rect 4588 23633 4628 25348
rect 4587 23624 4629 23633
rect 4587 23584 4588 23624
rect 4628 23584 4629 23624
rect 4587 23575 4629 23584
rect 4587 23036 4629 23045
rect 4587 22996 4588 23036
rect 4628 22996 4629 23036
rect 4587 22987 4629 22996
rect 4588 22902 4628 22987
rect 4587 22532 4629 22541
rect 4587 22492 4588 22532
rect 4628 22492 4629 22532
rect 4587 22483 4629 22492
rect 4492 22147 4532 22156
rect 4396 19123 4436 19132
rect 4492 21776 4532 21785
rect 4299 19088 4341 19097
rect 4299 19048 4300 19088
rect 4340 19048 4341 19088
rect 4299 19039 4341 19048
rect 4396 18920 4436 18929
rect 4396 18080 4436 18880
rect 4396 18031 4436 18040
rect 4492 17744 4532 21736
rect 4492 17695 4532 17704
rect 4588 17492 4628 22483
rect 4588 17443 4628 17452
rect 4684 22448 4724 32740
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4780 30260 4820 30269
rect 4780 30092 4820 30220
rect 4780 29168 4820 30052
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 4780 24557 4820 29128
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 5067 25304 5109 25313
rect 5067 25264 5068 25304
rect 5108 25264 5109 25304
rect 5067 25255 5109 25264
rect 5068 25170 5108 25255
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 4779 24548 4821 24557
rect 4779 24508 4780 24548
rect 4820 24508 4821 24548
rect 4779 24499 4821 24508
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 4396 16736 4436 16745
rect 4300 16568 4340 16577
rect 4300 14888 4340 16528
rect 4300 14839 4340 14848
rect 4204 14167 4244 14176
rect 4108 12403 4148 12412
rect 4108 12284 4148 12293
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 3819 10352 3861 10361
rect 3819 10312 3820 10352
rect 3860 10312 3861 10352
rect 3819 10303 3861 10312
rect 3820 9512 3860 10303
rect 4108 10100 4148 12244
rect 4108 10051 4148 10060
rect 4204 11696 4244 11705
rect 3820 9463 3860 9472
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 4204 9092 4244 11656
rect 4300 9848 4340 9857
rect 4300 9512 4340 9808
rect 4396 9680 4436 16696
rect 4492 16400 4532 16409
rect 4492 13208 4532 16360
rect 4492 13159 4532 13168
rect 4588 13124 4628 13133
rect 4396 9631 4436 9640
rect 4492 13040 4532 13049
rect 4300 9472 4436 9512
rect 4204 9043 4244 9052
rect 4108 7916 4148 7925
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3819 6992 3861 7001
rect 3819 6952 3820 6992
rect 3860 6952 3861 6992
rect 3819 6943 3861 6952
rect 3820 6488 3860 6943
rect 4108 6497 4148 7876
rect 4396 7916 4436 9472
rect 4396 7867 4436 7876
rect 4204 7832 4244 7841
rect 3820 6439 3860 6448
rect 4107 6488 4149 6497
rect 4107 6448 4108 6488
rect 4148 6448 4149 6488
rect 4107 6439 4149 6448
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4204 4397 4244 7792
rect 4299 7160 4341 7169
rect 4299 7120 4300 7160
rect 4340 7120 4341 7160
rect 4299 7111 4341 7120
rect 4300 7026 4340 7111
rect 4203 4388 4245 4397
rect 4203 4348 4204 4388
rect 4244 4348 4245 4388
rect 4203 4339 4245 4348
rect 4107 4136 4149 4145
rect 4107 4096 4108 4136
rect 4148 4096 4149 4136
rect 4107 4087 4149 4096
rect 4300 4136 4340 4145
rect 4108 4002 4148 4087
rect 4300 3977 4340 4096
rect 4299 3968 4341 3977
rect 4299 3928 4300 3968
rect 4340 3928 4341 3968
rect 4299 3919 4341 3928
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 4492 2540 4532 13000
rect 4588 9932 4628 13084
rect 4588 9883 4628 9892
rect 4684 6572 4724 22408
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 5356 21356 5396 38200
rect 5452 31520 5492 41896
rect 5452 31471 5492 31480
rect 5548 41852 5588 41861
rect 5548 30932 5588 41812
rect 5836 41684 5876 41693
rect 5740 40508 5780 40517
rect 5644 37148 5684 37157
rect 5644 35309 5684 37108
rect 5643 35300 5685 35309
rect 5643 35260 5644 35300
rect 5684 35260 5685 35300
rect 5643 35251 5685 35260
rect 5644 34880 5684 34889
rect 5644 34376 5684 34840
rect 5644 31352 5684 34336
rect 5644 31303 5684 31312
rect 5452 30892 5588 30932
rect 5452 29084 5492 30892
rect 5547 30764 5589 30773
rect 5547 30724 5548 30764
rect 5588 30724 5589 30764
rect 5547 30715 5589 30724
rect 5548 30630 5588 30715
rect 5452 29035 5492 29044
rect 5644 30344 5684 30353
rect 5548 28664 5588 28673
rect 5548 28244 5588 28624
rect 5452 27908 5492 27917
rect 5452 27581 5492 27868
rect 5451 27572 5493 27581
rect 5451 27532 5452 27572
rect 5492 27532 5493 27572
rect 5451 27523 5493 27532
rect 5451 24716 5493 24725
rect 5451 24676 5452 24716
rect 5492 24676 5493 24716
rect 5451 24667 5493 24676
rect 5452 21785 5492 24667
rect 5451 21776 5493 21785
rect 5451 21736 5452 21776
rect 5492 21736 5493 21776
rect 5451 21727 5493 21736
rect 5548 21608 5588 28204
rect 5644 27320 5684 30304
rect 5740 28580 5780 40468
rect 5836 40349 5876 41644
rect 5835 40340 5877 40349
rect 5835 40300 5836 40340
rect 5876 40300 5877 40340
rect 5835 40291 5877 40300
rect 6316 38744 6356 38753
rect 5740 28531 5780 28540
rect 5836 38324 5876 38333
rect 5644 27271 5684 27280
rect 5643 25892 5685 25901
rect 5643 25852 5644 25892
rect 5684 25852 5685 25892
rect 5643 25843 5685 25852
rect 5356 21307 5396 21316
rect 5452 21568 5588 21608
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 5356 19172 5396 19181
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 4779 18332 4821 18341
rect 4779 18292 4780 18332
rect 4820 18292 4821 18332
rect 4779 18283 4821 18292
rect 4780 18198 4820 18283
rect 4780 17744 4820 17753
rect 4780 14636 4820 17704
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 4780 8597 4820 14596
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4779 8588 4821 8597
rect 4779 8548 4780 8588
rect 4820 8548 4821 8588
rect 4779 8539 4821 8548
rect 4780 7169 4820 8539
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4779 7160 4821 7169
rect 4779 7120 4780 7160
rect 4820 7120 4821 7160
rect 4779 7111 4821 7120
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 4684 6532 4820 6572
rect 4683 6236 4725 6245
rect 4683 6196 4684 6236
rect 4724 6196 4725 6236
rect 4683 6187 4725 6196
rect 4587 4640 4629 4649
rect 4587 4600 4588 4640
rect 4628 4600 4629 4640
rect 4587 4591 4629 4600
rect 4588 4220 4628 4591
rect 4588 4171 4628 4180
rect 4396 2500 4532 2540
rect 4396 2288 4436 2500
rect 4396 2239 4436 2248
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 4299 1448 4341 1457
rect 4299 1408 4300 1448
rect 4340 1408 4341 1448
rect 4299 1399 4341 1408
rect 4300 1112 4340 1399
rect 4300 1063 4340 1072
rect 3532 895 3572 904
rect 4684 608 4724 6187
rect 4780 5144 4820 6532
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4780 5104 4916 5144
rect 4779 4220 4821 4229
rect 4779 4180 4780 4220
rect 4820 4180 4821 4220
rect 4779 4171 4821 4180
rect 4780 4086 4820 4171
rect 4876 4145 4916 5104
rect 4971 4724 5013 4733
rect 4971 4684 4972 4724
rect 5012 4684 5013 4724
rect 4971 4675 5013 4684
rect 4972 4590 5012 4675
rect 4875 4136 4917 4145
rect 4875 4096 4876 4136
rect 4916 4096 4917 4136
rect 4875 4087 4917 4096
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5356 1364 5396 19132
rect 5452 17828 5492 21568
rect 5452 17779 5492 17788
rect 5548 20768 5588 20777
rect 5548 17156 5588 20728
rect 5644 18752 5684 25843
rect 5644 18703 5684 18712
rect 5740 25808 5780 25817
rect 5740 18416 5780 25768
rect 5836 25640 5876 38284
rect 6220 38072 6260 38081
rect 6220 37913 6260 38032
rect 6219 37904 6261 37913
rect 6219 37864 6220 37904
rect 6260 37864 6261 37904
rect 6219 37855 6261 37864
rect 6028 37484 6068 37493
rect 6028 35804 6068 37444
rect 5931 34964 5973 34973
rect 5931 34924 5932 34964
rect 5972 34924 5973 34964
rect 5931 34915 5973 34924
rect 5932 34040 5972 34915
rect 5932 33991 5972 34000
rect 5836 25591 5876 25600
rect 5932 31016 5972 31025
rect 5932 30512 5972 30976
rect 5932 23204 5972 30472
rect 5932 23036 5972 23164
rect 5932 22987 5972 22996
rect 5931 22364 5973 22373
rect 5931 22324 5932 22364
rect 5972 22324 5973 22364
rect 5931 22315 5973 22324
rect 5740 17660 5780 18376
rect 5932 20768 5972 22315
rect 5740 17620 5876 17660
rect 5548 17107 5588 17116
rect 5644 17324 5684 17333
rect 5548 15308 5588 15317
rect 5356 1315 5396 1324
rect 5452 14216 5492 14225
rect 5259 1196 5301 1205
rect 5259 1156 5260 1196
rect 5300 1156 5301 1196
rect 5259 1147 5301 1156
rect 5260 1062 5300 1147
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5452 692 5492 14176
rect 5548 12284 5588 15268
rect 5548 12235 5588 12244
rect 5644 11360 5684 17284
rect 5740 17240 5780 17249
rect 5740 14552 5780 17200
rect 5740 14503 5780 14512
rect 5836 13964 5876 17620
rect 5548 11320 5684 11360
rect 5740 13924 5876 13964
rect 5740 13208 5780 13924
rect 5740 11780 5780 13168
rect 5548 10940 5588 11320
rect 5740 11276 5780 11740
rect 5740 11108 5780 11236
rect 5740 11059 5780 11068
rect 5836 13796 5876 13805
rect 5548 4640 5588 10900
rect 5739 10772 5781 10781
rect 5739 10732 5740 10772
rect 5780 10732 5781 10772
rect 5739 10723 5781 10732
rect 5740 10436 5780 10723
rect 5740 10387 5780 10396
rect 5740 8924 5780 8933
rect 5740 8336 5780 8884
rect 5740 8287 5780 8296
rect 5644 8252 5684 8261
rect 5644 7412 5684 8212
rect 5644 7363 5684 7372
rect 5548 4591 5588 4600
rect 5740 4304 5780 4313
rect 5643 2624 5685 2633
rect 5643 2584 5644 2624
rect 5684 2584 5685 2624
rect 5643 2575 5685 2584
rect 5644 2204 5684 2575
rect 5740 2372 5780 4264
rect 5836 2540 5876 13756
rect 5932 11360 5972 20728
rect 5932 11311 5972 11320
rect 5836 2491 5876 2500
rect 5932 2792 5972 2801
rect 5932 2456 5972 2752
rect 5932 2407 5972 2416
rect 5740 2323 5780 2332
rect 5644 2155 5684 2164
rect 5547 2036 5589 2045
rect 5547 1996 5548 2036
rect 5588 1996 5589 2036
rect 5547 1987 5589 1996
rect 5452 643 5492 652
rect 4684 559 4724 568
rect 5548 608 5588 1987
rect 6028 944 6068 35764
rect 6123 35216 6165 35225
rect 6123 35176 6124 35216
rect 6164 35176 6165 35216
rect 6123 35167 6165 35176
rect 6124 34208 6164 35167
rect 6124 34159 6164 34168
rect 6124 33116 6164 33125
rect 6124 30596 6164 33076
rect 6220 32780 6260 37855
rect 6316 37820 6356 38704
rect 6316 37771 6356 37780
rect 6315 35048 6357 35057
rect 6315 35008 6316 35048
rect 6356 35008 6357 35048
rect 6315 34999 6357 35008
rect 6316 34914 6356 34999
rect 6220 32731 6260 32740
rect 6124 29420 6164 30556
rect 6124 29371 6164 29380
rect 6220 32612 6260 32621
rect 6220 27656 6260 32572
rect 6220 27607 6260 27616
rect 6316 32528 6356 32537
rect 6123 26732 6165 26741
rect 6123 26692 6124 26732
rect 6164 26692 6165 26732
rect 6123 26683 6165 26692
rect 6124 20180 6164 26683
rect 6219 25136 6261 25145
rect 6219 25096 6220 25136
rect 6260 25096 6261 25136
rect 6219 25087 6261 25096
rect 6220 23036 6260 25087
rect 6316 23288 6356 32488
rect 6412 25556 6452 41980
rect 6604 41600 6644 41609
rect 6508 40508 6548 40517
rect 6508 34301 6548 40468
rect 6507 34292 6549 34301
rect 6507 34252 6508 34292
rect 6548 34252 6549 34292
rect 6507 34243 6549 34252
rect 6508 33032 6548 34243
rect 6508 32983 6548 32992
rect 6412 25507 6452 25516
rect 6508 26480 6548 26489
rect 6412 24800 6452 24809
rect 6412 23708 6452 24760
rect 6412 23659 6452 23668
rect 6316 23239 6356 23248
rect 6412 23036 6452 23045
rect 6220 22996 6356 23036
rect 6219 22868 6261 22877
rect 6219 22828 6220 22868
rect 6260 22828 6261 22868
rect 6219 22819 6261 22828
rect 6220 22734 6260 22819
rect 6316 22037 6356 22996
rect 6315 22028 6357 22037
rect 6315 21988 6316 22028
rect 6356 21988 6357 22028
rect 6315 21979 6357 21988
rect 6124 20140 6260 20180
rect 6124 18920 6164 18929
rect 6124 8924 6164 18880
rect 6124 4304 6164 8884
rect 6124 4255 6164 4264
rect 6220 1280 6260 20140
rect 6412 19088 6452 22996
rect 6412 19039 6452 19048
rect 6412 18836 6452 18845
rect 6412 17660 6452 18796
rect 6508 17837 6548 26440
rect 6604 22532 6644 41560
rect 6796 41600 6836 42223
rect 6796 41551 6836 41560
rect 7180 41600 7220 41609
rect 6796 40340 6836 40349
rect 6796 39836 6836 40300
rect 6699 38240 6741 38249
rect 6699 38200 6700 38240
rect 6740 38200 6741 38240
rect 6699 38191 6741 38200
rect 6700 38106 6740 38191
rect 6700 34628 6740 34637
rect 6700 33536 6740 34588
rect 6700 33487 6740 33496
rect 6796 34460 6836 39796
rect 6988 40256 7028 40265
rect 6988 38744 7028 40216
rect 7083 39668 7125 39677
rect 7083 39628 7084 39668
rect 7124 39628 7125 39668
rect 7083 39619 7125 39628
rect 7084 39534 7124 39619
rect 6988 38695 7028 38704
rect 6988 37904 7028 37913
rect 6988 37736 7028 37864
rect 6988 37687 7028 37696
rect 6988 36644 7028 36653
rect 6892 35216 6932 35225
rect 6892 34469 6932 35176
rect 6796 33284 6836 34420
rect 6891 34460 6933 34469
rect 6891 34420 6892 34460
rect 6932 34420 6933 34460
rect 6891 34411 6933 34420
rect 6796 33235 6836 33244
rect 6892 33872 6932 33881
rect 6699 32948 6741 32957
rect 6699 32908 6700 32948
rect 6740 32908 6741 32948
rect 6699 32899 6741 32908
rect 6700 32814 6740 32899
rect 6700 28916 6740 28925
rect 6700 27404 6740 28876
rect 6795 27572 6837 27581
rect 6795 27532 6796 27572
rect 6836 27532 6837 27572
rect 6795 27523 6837 27532
rect 6700 27355 6740 27364
rect 6699 26732 6741 26741
rect 6699 26692 6700 26732
rect 6740 26692 6741 26732
rect 6699 26683 6741 26692
rect 6700 26648 6740 26683
rect 6700 26597 6740 26608
rect 6700 24800 6740 24809
rect 6700 23876 6740 24760
rect 6700 23827 6740 23836
rect 6699 22952 6741 22961
rect 6699 22912 6700 22952
rect 6740 22912 6741 22952
rect 6699 22903 6741 22912
rect 6700 22868 6740 22903
rect 6700 22817 6740 22828
rect 6604 22483 6644 22492
rect 6699 22028 6741 22037
rect 6699 21988 6700 22028
rect 6740 21988 6741 22028
rect 6699 21979 6741 21988
rect 6604 19844 6644 19853
rect 6507 17828 6549 17837
rect 6507 17788 6508 17828
rect 6548 17788 6549 17828
rect 6507 17779 6549 17788
rect 6412 17620 6548 17660
rect 6412 17324 6452 17333
rect 6412 17072 6452 17284
rect 6412 17023 6452 17032
rect 6412 16400 6452 16409
rect 6315 15728 6357 15737
rect 6315 15688 6316 15728
rect 6356 15688 6357 15728
rect 6315 15679 6357 15688
rect 6316 9008 6356 15679
rect 6412 14552 6452 16360
rect 6412 14503 6452 14512
rect 6411 12620 6453 12629
rect 6411 12580 6412 12620
rect 6452 12580 6453 12620
rect 6411 12571 6453 12580
rect 6316 8959 6356 8968
rect 6315 3632 6357 3641
rect 6315 3592 6316 3632
rect 6356 3592 6357 3632
rect 6315 3583 6357 3592
rect 6316 2624 6356 3583
rect 6316 2575 6356 2584
rect 6220 1231 6260 1240
rect 6028 895 6068 904
rect 6412 944 6452 12571
rect 6508 12452 6548 17620
rect 6508 12403 6548 12412
rect 6508 7160 6548 7169
rect 6508 2540 6548 7120
rect 6508 2491 6548 2500
rect 6507 1952 6549 1961
rect 6507 1912 6508 1952
rect 6548 1912 6549 1952
rect 6507 1903 6549 1912
rect 6508 1818 6548 1903
rect 6604 1280 6644 19804
rect 6700 11360 6740 21979
rect 6700 11311 6740 11320
rect 6700 8840 6740 8849
rect 6700 4565 6740 8800
rect 6699 4556 6741 4565
rect 6699 4516 6700 4556
rect 6740 4516 6741 4556
rect 6699 4507 6741 4516
rect 6700 3968 6740 3977
rect 6700 3380 6740 3928
rect 6700 3331 6740 3340
rect 6604 1231 6644 1240
rect 6796 1280 6836 27523
rect 6892 25145 6932 33832
rect 6988 32528 7028 36604
rect 6988 32479 7028 32488
rect 7084 35132 7124 35141
rect 6988 28748 7028 28757
rect 6988 27404 7028 28708
rect 6891 25136 6933 25145
rect 6891 25096 6892 25136
rect 6932 25096 6933 25136
rect 6891 25087 6933 25096
rect 6892 24968 6932 24977
rect 6892 21944 6932 24928
rect 6892 21895 6932 21904
rect 6988 21776 7028 27364
rect 6988 21727 7028 21736
rect 6988 17492 7028 17501
rect 6892 17408 6932 17417
rect 6892 11360 6932 17368
rect 6988 15560 7028 17452
rect 6988 14216 7028 15520
rect 6988 14167 7028 14176
rect 6892 11320 7028 11360
rect 6892 8504 6932 8513
rect 6892 3296 6932 8464
rect 6892 2624 6932 3256
rect 6892 2575 6932 2584
rect 6891 1868 6933 1877
rect 6891 1828 6892 1868
rect 6932 1828 6933 1868
rect 6891 1819 6933 1828
rect 6892 1734 6932 1819
rect 6796 1231 6836 1240
rect 6988 1280 7028 11320
rect 6988 1231 7028 1240
rect 6412 895 6452 904
rect 7084 692 7124 35092
rect 7180 32024 7220 41560
rect 7372 41600 7412 41609
rect 7275 36728 7317 36737
rect 7275 36688 7276 36728
rect 7316 36688 7317 36728
rect 7275 36679 7317 36688
rect 7276 34376 7316 36679
rect 7276 34327 7316 34336
rect 7180 31975 7220 31984
rect 7180 29672 7220 29681
rect 7180 23372 7220 29632
rect 7372 29000 7412 41560
rect 7468 41180 7508 41189
rect 7468 41021 7508 41140
rect 7467 41012 7509 41021
rect 7467 40972 7468 41012
rect 7508 40972 7509 41012
rect 7467 40963 7509 40972
rect 7276 28960 7412 29000
rect 7468 38156 7508 38165
rect 7276 24128 7316 28960
rect 7468 28580 7508 38116
rect 7564 35729 7604 42652
rect 9484 42608 9524 42617
rect 7852 41852 7892 41861
rect 7563 35720 7605 35729
rect 7563 35680 7564 35720
rect 7604 35680 7605 35720
rect 7563 35671 7605 35680
rect 7660 35468 7700 35477
rect 7563 34460 7605 34469
rect 7563 34420 7564 34460
rect 7604 34420 7605 34460
rect 7563 34411 7605 34420
rect 7564 33788 7604 34411
rect 7660 33872 7700 35428
rect 7660 33823 7700 33832
rect 7756 35216 7796 35225
rect 7564 32360 7604 33748
rect 7756 33116 7796 35176
rect 7756 33067 7796 33076
rect 7564 31940 7604 32320
rect 7564 31891 7604 31900
rect 7756 32528 7796 32537
rect 7564 31520 7604 31529
rect 7564 29252 7604 31480
rect 7660 31268 7700 31277
rect 7660 30680 7700 31228
rect 7660 30631 7700 30640
rect 7564 29203 7604 29212
rect 7372 28540 7508 28580
rect 7372 27488 7412 28540
rect 7467 28412 7509 28421
rect 7467 28372 7468 28412
rect 7508 28372 7509 28412
rect 7467 28363 7509 28372
rect 7468 28278 7508 28363
rect 7372 27439 7412 27448
rect 7276 24079 7316 24088
rect 7468 25388 7508 25397
rect 7371 24044 7413 24053
rect 7371 24004 7372 24044
rect 7412 24004 7413 24044
rect 7371 23995 7413 24004
rect 7372 23910 7412 23995
rect 7468 23960 7508 25348
rect 7468 23920 7604 23960
rect 7372 23708 7412 23717
rect 7180 23332 7316 23372
rect 7180 22784 7220 22793
rect 7180 15560 7220 22744
rect 7276 21272 7316 23332
rect 7276 15737 7316 21232
rect 7372 19928 7412 23668
rect 7372 19879 7412 19888
rect 7468 23456 7508 23465
rect 7275 15728 7317 15737
rect 7275 15688 7276 15728
rect 7316 15688 7317 15728
rect 7275 15679 7317 15688
rect 7180 6740 7220 15520
rect 7371 12452 7413 12461
rect 7371 12412 7372 12452
rect 7412 12412 7413 12452
rect 7371 12403 7413 12412
rect 7372 12032 7412 12403
rect 7276 11528 7316 11537
rect 7276 11276 7316 11488
rect 7276 11227 7316 11236
rect 7372 7244 7412 11992
rect 7372 7195 7412 7204
rect 7180 6700 7316 6740
rect 7179 4808 7221 4817
rect 7179 4768 7180 4808
rect 7220 4768 7221 4808
rect 7179 4759 7221 4768
rect 7180 4229 7220 4759
rect 7276 4733 7316 6700
rect 7468 5564 7508 23416
rect 7564 15821 7604 23920
rect 7563 15812 7605 15821
rect 7563 15772 7564 15812
rect 7604 15772 7605 15812
rect 7563 15763 7605 15772
rect 7564 15392 7604 15401
rect 7564 15233 7604 15352
rect 7563 15224 7605 15233
rect 7563 15184 7564 15224
rect 7604 15184 7605 15224
rect 7563 15175 7605 15184
rect 7660 15224 7700 15233
rect 7660 12041 7700 15184
rect 7659 12032 7701 12041
rect 7659 11992 7660 12032
rect 7700 11992 7701 12032
rect 7659 11983 7701 11992
rect 7564 11864 7604 11873
rect 7564 11276 7604 11824
rect 7564 11227 7604 11236
rect 7660 11360 7700 11369
rect 7660 10436 7700 11320
rect 7660 10387 7700 10396
rect 7563 9680 7605 9689
rect 7563 9640 7564 9680
rect 7604 9640 7605 9680
rect 7563 9631 7605 9640
rect 7564 7076 7604 9631
rect 7564 7027 7604 7036
rect 7563 6488 7605 6497
rect 7563 6448 7564 6488
rect 7604 6448 7605 6488
rect 7563 6439 7605 6448
rect 7564 6354 7604 6439
rect 7660 6404 7700 6415
rect 7660 6329 7700 6364
rect 7659 6320 7701 6329
rect 7659 6280 7660 6320
rect 7700 6280 7701 6320
rect 7659 6271 7701 6280
rect 7371 5228 7413 5237
rect 7371 5188 7372 5228
rect 7412 5188 7413 5228
rect 7371 5179 7413 5188
rect 7468 5228 7508 5524
rect 7468 5179 7508 5188
rect 7275 4724 7317 4733
rect 7275 4684 7276 4724
rect 7316 4684 7317 4724
rect 7275 4675 7317 4684
rect 7275 4556 7317 4565
rect 7275 4516 7276 4556
rect 7316 4516 7317 4556
rect 7275 4507 7317 4516
rect 7179 4220 7221 4229
rect 7179 4180 7180 4220
rect 7220 4180 7221 4220
rect 7179 4171 7221 4180
rect 7180 1952 7220 4171
rect 7276 2372 7316 4507
rect 7372 3884 7412 5179
rect 7372 3835 7412 3844
rect 7468 5060 7508 5069
rect 7276 2323 7316 2332
rect 7180 1903 7220 1912
rect 7179 1280 7221 1289
rect 7179 1240 7180 1280
rect 7220 1240 7221 1280
rect 7179 1231 7221 1240
rect 7180 1146 7220 1231
rect 7084 643 7124 652
rect 5548 559 5588 568
rect 7468 608 7508 5020
rect 7564 3632 7604 3641
rect 7564 2717 7604 3592
rect 7660 2960 7700 6271
rect 7660 2911 7700 2920
rect 7563 2708 7605 2717
rect 7563 2668 7564 2708
rect 7604 2668 7605 2708
rect 7563 2659 7605 2668
rect 7564 2540 7604 2659
rect 7564 2491 7604 2500
rect 7756 1280 7796 32488
rect 7852 23288 7892 41812
rect 7948 41600 7988 41609
rect 7948 28496 7988 41560
rect 9292 41600 9332 41609
rect 8812 40508 8852 40517
rect 8044 40004 8084 40013
rect 8044 35888 8084 39964
rect 8044 35839 8084 35848
rect 8524 39668 8564 39677
rect 8427 34460 8469 34469
rect 8427 34420 8428 34460
rect 8468 34420 8469 34460
rect 8427 34411 8469 34420
rect 8043 34376 8085 34385
rect 8043 34336 8044 34376
rect 8084 34336 8085 34376
rect 8043 34327 8085 34336
rect 8044 34242 8084 34327
rect 8428 34326 8468 34411
rect 8043 32948 8085 32957
rect 8043 32908 8044 32948
rect 8084 32908 8085 32948
rect 8043 32899 8085 32908
rect 7948 28447 7988 28456
rect 7947 25892 7989 25901
rect 7947 25852 7948 25892
rect 7988 25852 7989 25892
rect 7947 25843 7989 25852
rect 7948 25758 7988 25843
rect 7852 23239 7892 23248
rect 7852 22364 7892 22373
rect 7852 12629 7892 22324
rect 8044 15224 8084 32899
rect 8236 32864 8276 32873
rect 8140 30008 8180 30017
rect 8140 28673 8180 29968
rect 8139 28664 8181 28673
rect 8139 28624 8140 28664
rect 8180 28624 8181 28664
rect 8139 28615 8181 28624
rect 8140 28412 8180 28421
rect 8140 24548 8180 28372
rect 8140 23960 8180 24508
rect 8140 23911 8180 23920
rect 8236 20012 8276 32824
rect 8428 32864 8468 32873
rect 8428 31436 8468 32824
rect 8428 31387 8468 31396
rect 8428 29336 8468 29345
rect 8331 29168 8373 29177
rect 8331 29128 8332 29168
rect 8372 29128 8373 29168
rect 8331 29119 8373 29128
rect 8428 29168 8468 29296
rect 8428 29119 8468 29128
rect 8236 19424 8276 19972
rect 8236 19375 8276 19384
rect 8139 17576 8181 17585
rect 8139 17536 8140 17576
rect 8180 17536 8181 17576
rect 8139 17527 8181 17536
rect 8044 15175 8084 15184
rect 7948 12956 7988 12965
rect 7851 12620 7893 12629
rect 7851 12580 7852 12620
rect 7892 12580 7893 12620
rect 7851 12571 7893 12580
rect 7852 12284 7892 12293
rect 7852 11024 7892 12244
rect 7852 10975 7892 10984
rect 7948 11696 7988 12916
rect 7948 10100 7988 11656
rect 8044 11948 8084 11957
rect 8044 11453 8084 11908
rect 8043 11444 8085 11453
rect 8043 11404 8044 11444
rect 8084 11404 8085 11444
rect 8043 11395 8085 11404
rect 7948 10051 7988 10060
rect 8044 8000 8084 11395
rect 8044 7951 8084 7960
rect 8044 7412 8084 7421
rect 8044 6992 8084 7372
rect 8044 6943 8084 6952
rect 8044 3464 8084 3473
rect 8044 1364 8084 3424
rect 8044 1315 8084 1324
rect 7756 1231 7796 1240
rect 8140 1280 8180 17527
rect 8236 13208 8276 13217
rect 8236 8000 8276 13168
rect 8236 4304 8276 7960
rect 8236 4255 8276 4264
rect 8140 1231 8180 1240
rect 8332 1280 8372 29119
rect 8524 29000 8564 39628
rect 8812 38996 8852 40468
rect 8812 38947 8852 38956
rect 8908 39668 8948 39677
rect 8908 39500 8948 39628
rect 8908 37820 8948 39460
rect 8812 37780 8948 37820
rect 8620 32192 8660 32201
rect 8620 29597 8660 32152
rect 8812 31520 8852 37780
rect 9004 37400 9044 37409
rect 8908 37232 8948 37241
rect 8908 35309 8948 37192
rect 8907 35300 8949 35309
rect 8907 35260 8908 35300
rect 8948 35260 8949 35300
rect 8907 35251 8949 35260
rect 8812 31471 8852 31480
rect 9004 30596 9044 37360
rect 9099 37232 9141 37241
rect 9099 37192 9100 37232
rect 9140 37192 9141 37232
rect 9099 37183 9141 37192
rect 9100 31949 9140 37183
rect 9099 31940 9141 31949
rect 9099 31900 9100 31940
rect 9140 31900 9141 31940
rect 9099 31891 9141 31900
rect 8908 30556 9044 30596
rect 9100 31520 9140 31529
rect 8716 29756 8756 29765
rect 8619 29588 8661 29597
rect 8619 29548 8620 29588
rect 8660 29548 8661 29588
rect 8619 29539 8661 29548
rect 8619 29252 8661 29261
rect 8619 29212 8620 29252
rect 8660 29212 8661 29252
rect 8619 29203 8661 29212
rect 8428 28960 8564 29000
rect 8428 28244 8468 28960
rect 8523 28664 8565 28673
rect 8523 28624 8524 28664
rect 8564 28624 8565 28664
rect 8523 28615 8565 28624
rect 8428 12620 8468 28204
rect 8524 27656 8564 28615
rect 8524 27607 8564 27616
rect 8620 26480 8660 29203
rect 8716 29093 8756 29716
rect 8715 29084 8757 29093
rect 8715 29044 8716 29084
rect 8756 29044 8757 29084
rect 8715 29035 8757 29044
rect 8811 27572 8853 27581
rect 8811 27532 8812 27572
rect 8852 27532 8853 27572
rect 8811 27523 8853 27532
rect 8620 26431 8660 26440
rect 8812 26480 8852 27523
rect 8812 26431 8852 26440
rect 8524 24800 8564 24809
rect 8524 23288 8564 24760
rect 8908 23717 8948 30556
rect 9004 30428 9044 30437
rect 9004 29420 9044 30388
rect 9004 29371 9044 29380
rect 9003 26480 9045 26489
rect 9003 26440 9004 26480
rect 9044 26440 9045 26480
rect 9003 26431 9045 26440
rect 9004 26346 9044 26431
rect 8907 23708 8949 23717
rect 8907 23668 8908 23708
rect 8948 23668 8949 23708
rect 8907 23659 8949 23668
rect 8524 13208 8564 23248
rect 8812 23624 8852 23633
rect 8716 16400 8756 16409
rect 8619 15812 8661 15821
rect 8619 15772 8620 15812
rect 8660 15772 8661 15812
rect 8619 15763 8661 15772
rect 8524 13159 8564 13168
rect 8428 12571 8468 12580
rect 8428 11864 8468 11873
rect 8428 11444 8468 11824
rect 8428 11395 8468 11404
rect 8524 7244 8564 7253
rect 8524 6320 8564 7204
rect 8524 6271 8564 6280
rect 8428 4976 8468 4985
rect 8428 2288 8468 4936
rect 8428 2239 8468 2248
rect 8332 1231 8372 1240
rect 8620 944 8660 15763
rect 8716 4976 8756 16360
rect 8812 10856 8852 23584
rect 9004 17744 9044 17753
rect 8907 15644 8949 15653
rect 8907 15604 8908 15644
rect 8948 15604 8949 15644
rect 8907 15595 8949 15604
rect 8908 15510 8948 15595
rect 8908 14636 8948 14645
rect 8908 14132 8948 14596
rect 8908 14083 8948 14092
rect 8812 10807 8852 10816
rect 8908 12620 8948 12629
rect 8812 10268 8852 10277
rect 8812 6404 8852 10228
rect 8812 6355 8852 6364
rect 8716 4927 8756 4936
rect 8812 5396 8852 5405
rect 8716 4136 8756 4145
rect 8716 2288 8756 4096
rect 8716 2239 8756 2248
rect 8812 2204 8852 5356
rect 8812 2155 8852 2164
rect 8908 1280 8948 12580
rect 9004 7160 9044 17704
rect 9004 7111 9044 7120
rect 9003 4304 9045 4313
rect 9003 4264 9004 4304
rect 9044 4264 9045 4304
rect 9003 4255 9045 4264
rect 9004 4170 9044 4255
rect 9100 2792 9140 31480
rect 9196 29756 9236 29765
rect 9196 29336 9236 29716
rect 9196 23540 9236 29296
rect 9292 27488 9332 41560
rect 9387 37484 9429 37493
rect 9387 37444 9388 37484
rect 9428 37444 9429 37484
rect 9387 37435 9429 37444
rect 9388 37350 9428 37435
rect 9387 35048 9429 35057
rect 9387 35008 9388 35048
rect 9428 35008 9429 35048
rect 9387 34999 9429 35008
rect 9388 34914 9428 34999
rect 9484 34637 9524 42568
rect 11404 41684 11444 41693
rect 9868 41600 9908 41609
rect 9580 36644 9620 36653
rect 9483 34628 9525 34637
rect 9483 34588 9484 34628
rect 9524 34588 9525 34628
rect 9483 34579 9525 34588
rect 9387 27656 9429 27665
rect 9387 27616 9388 27656
rect 9428 27616 9429 27656
rect 9387 27607 9429 27616
rect 9388 27522 9428 27607
rect 9292 27439 9332 27448
rect 9196 23491 9236 23500
rect 9292 23372 9332 23381
rect 9196 22028 9236 22037
rect 9196 17744 9236 21988
rect 9196 17695 9236 17704
rect 9196 17408 9236 17417
rect 9196 14384 9236 17368
rect 9196 14335 9236 14344
rect 9196 12116 9236 12125
rect 9196 11864 9236 12076
rect 9292 11957 9332 23332
rect 9484 20180 9524 34579
rect 9580 26480 9620 36604
rect 9580 26431 9620 26440
rect 9676 29504 9716 29513
rect 9676 25388 9716 29464
rect 9771 29084 9813 29093
rect 9771 29044 9772 29084
rect 9812 29044 9813 29084
rect 9771 29035 9813 29044
rect 9676 25339 9716 25348
rect 9388 20140 9524 20180
rect 9580 21608 9620 21617
rect 9291 11948 9333 11957
rect 9291 11908 9292 11948
rect 9332 11908 9333 11948
rect 9291 11899 9333 11908
rect 9196 10016 9236 11824
rect 9196 9967 9236 9976
rect 9292 11612 9332 11621
rect 9196 8840 9236 8849
rect 9196 7580 9236 8800
rect 9196 7531 9236 7540
rect 9292 7496 9332 11572
rect 9292 7447 9332 7456
rect 9291 4640 9333 4649
rect 9291 4600 9292 4640
rect 9332 4600 9333 4640
rect 9291 4591 9333 4600
rect 9292 4506 9332 4591
rect 9100 2743 9140 2752
rect 9388 2465 9428 20140
rect 9580 17744 9620 21568
rect 9676 21356 9716 21365
rect 9676 18929 9716 21316
rect 9675 18920 9717 18929
rect 9675 18880 9676 18920
rect 9716 18880 9717 18920
rect 9675 18871 9717 18880
rect 9580 16325 9620 17704
rect 9579 16316 9621 16325
rect 9579 16276 9580 16316
rect 9620 16276 9621 16316
rect 9579 16267 9621 16276
rect 9580 16064 9620 16267
rect 9580 16015 9620 16024
rect 9484 15392 9524 15401
rect 9484 7664 9524 15352
rect 9676 13460 9716 13469
rect 9580 12788 9620 12797
rect 9580 12368 9620 12748
rect 9676 12704 9716 13420
rect 9676 12655 9716 12664
rect 9580 11528 9620 12328
rect 9580 11479 9620 11488
rect 9676 12452 9716 12461
rect 9580 10856 9620 10865
rect 9580 9680 9620 10816
rect 9580 9631 9620 9640
rect 9579 9512 9621 9521
rect 9579 9472 9580 9512
rect 9620 9472 9621 9512
rect 9579 9463 9621 9472
rect 9580 9378 9620 9463
rect 9676 9260 9716 12412
rect 9676 9211 9716 9220
rect 9484 7615 9524 7624
rect 9579 5060 9621 5069
rect 9579 5020 9580 5060
rect 9620 5020 9621 5060
rect 9579 5011 9621 5020
rect 9580 4976 9620 5011
rect 9580 4925 9620 4936
rect 9772 4220 9812 29035
rect 9868 20684 9908 41560
rect 9963 41600 10005 41609
rect 9963 41560 9964 41600
rect 10004 41560 10005 41600
rect 9963 41551 10005 41560
rect 10252 41600 10292 41609
rect 9964 37652 10004 41551
rect 10156 40340 10196 40349
rect 10059 38744 10101 38753
rect 10059 38704 10060 38744
rect 10100 38704 10101 38744
rect 10059 38695 10101 38704
rect 9964 37603 10004 37612
rect 9964 35300 10004 35309
rect 9964 34376 10004 35260
rect 10060 35048 10100 38695
rect 10060 34999 10100 35008
rect 9964 34327 10004 34336
rect 10060 34880 10100 34889
rect 10060 34208 10100 34840
rect 10060 34159 10100 34168
rect 9964 31772 10004 31781
rect 9964 28916 10004 31732
rect 9964 28867 10004 28876
rect 10060 31352 10100 31361
rect 9868 20635 9908 20644
rect 9964 28748 10004 28757
rect 9964 18836 10004 28708
rect 10060 28664 10100 31312
rect 10060 28615 10100 28624
rect 10059 25304 10101 25313
rect 10059 25264 10060 25304
rect 10100 25264 10101 25304
rect 10059 25255 10101 25264
rect 10060 24044 10100 25255
rect 10060 23995 10100 24004
rect 9964 18787 10004 18796
rect 10060 19592 10100 19601
rect 9964 17660 10004 17669
rect 9867 14804 9909 14813
rect 9867 14764 9868 14804
rect 9908 14764 9909 14804
rect 9867 14755 9909 14764
rect 9868 9260 9908 14755
rect 9868 9211 9908 9220
rect 9964 8177 10004 17620
rect 10060 13880 10100 19552
rect 10156 18668 10196 40300
rect 10252 23540 10292 41560
rect 11020 41600 11060 41609
rect 10828 41012 10868 41021
rect 10636 39080 10676 39089
rect 10636 37913 10676 39040
rect 10731 38408 10773 38417
rect 10731 38368 10732 38408
rect 10772 38368 10773 38408
rect 10731 38359 10773 38368
rect 10635 37904 10677 37913
rect 10635 37864 10636 37904
rect 10676 37864 10677 37904
rect 10635 37855 10677 37864
rect 10348 36728 10388 36737
rect 10348 31352 10388 36688
rect 10636 36569 10676 37855
rect 10635 36560 10677 36569
rect 10635 36520 10636 36560
rect 10676 36520 10677 36560
rect 10635 36511 10677 36520
rect 10444 35300 10484 35309
rect 10444 35057 10484 35260
rect 10443 35048 10485 35057
rect 10443 35008 10444 35048
rect 10484 35008 10485 35048
rect 10443 34999 10485 35008
rect 10732 34973 10772 38359
rect 10828 35720 10868 40972
rect 10828 35671 10868 35680
rect 10828 35300 10868 35309
rect 10731 34964 10773 34973
rect 10731 34924 10732 34964
rect 10772 34924 10773 34964
rect 10731 34915 10773 34924
rect 10732 34208 10772 34217
rect 10636 34124 10676 34133
rect 10540 33704 10580 33713
rect 10540 33536 10580 33664
rect 10348 31303 10388 31312
rect 10444 31520 10484 31529
rect 10348 28664 10388 28673
rect 10348 24632 10388 28624
rect 10348 24583 10388 24592
rect 10252 23491 10292 23500
rect 10251 23036 10293 23045
rect 10251 22996 10252 23036
rect 10292 22996 10293 23036
rect 10251 22987 10293 22996
rect 10156 17660 10196 18628
rect 10156 17611 10196 17620
rect 10156 14972 10196 14981
rect 10156 13964 10196 14932
rect 10156 13915 10196 13924
rect 10060 13831 10100 13840
rect 10155 13796 10197 13805
rect 10155 13756 10156 13796
rect 10196 13756 10197 13796
rect 10155 13747 10197 13756
rect 10059 10688 10101 10697
rect 10059 10648 10060 10688
rect 10100 10648 10101 10688
rect 10059 10639 10101 10648
rect 9963 8168 10005 8177
rect 9963 8128 9964 8168
rect 10004 8128 10005 8168
rect 9963 8119 10005 8128
rect 9580 4180 9812 4220
rect 9868 7916 9908 7925
rect 9387 2456 9429 2465
rect 9387 2416 9388 2456
rect 9428 2416 9429 2456
rect 9387 2407 9429 2416
rect 8908 1231 8948 1240
rect 9388 1196 9428 2407
rect 9580 1952 9620 4180
rect 9675 3968 9717 3977
rect 9675 3928 9676 3968
rect 9716 3928 9717 3968
rect 9675 3919 9717 3928
rect 9676 3884 9716 3919
rect 9676 3833 9716 3844
rect 9771 3380 9813 3389
rect 9771 3340 9772 3380
rect 9812 3340 9813 3380
rect 9771 3331 9813 3340
rect 9772 3246 9812 3331
rect 9868 2624 9908 7876
rect 9964 4976 10004 8119
rect 9964 4927 10004 4936
rect 10060 2633 10100 10639
rect 10156 5900 10196 13747
rect 10252 6245 10292 22987
rect 10348 17660 10388 17669
rect 10348 13805 10388 17620
rect 10347 13796 10389 13805
rect 10347 13756 10348 13796
rect 10388 13756 10389 13796
rect 10347 13747 10389 13756
rect 10348 13628 10388 13637
rect 10348 12200 10388 13588
rect 10444 13208 10484 31480
rect 10540 30353 10580 33496
rect 10539 30344 10581 30353
rect 10539 30304 10540 30344
rect 10580 30304 10581 30344
rect 10539 30295 10581 30304
rect 10539 27740 10581 27749
rect 10539 27700 10540 27740
rect 10580 27700 10581 27740
rect 10539 27691 10581 27700
rect 10540 25556 10580 27691
rect 10636 27665 10676 34084
rect 10732 31352 10772 34168
rect 10732 31303 10772 31312
rect 10731 29168 10773 29177
rect 10731 29128 10732 29168
rect 10772 29128 10773 29168
rect 10731 29119 10773 29128
rect 10732 29034 10772 29119
rect 10635 27656 10677 27665
rect 10635 27616 10636 27656
rect 10676 27616 10677 27656
rect 10635 27607 10677 27616
rect 10540 25507 10580 25516
rect 10732 25388 10772 25397
rect 10732 23036 10772 25348
rect 10732 20180 10772 22996
rect 10636 20140 10772 20180
rect 10444 13159 10484 13168
rect 10540 15896 10580 15905
rect 10540 13460 10580 15856
rect 10348 12151 10388 12160
rect 10444 12284 10484 12293
rect 10444 11780 10484 12244
rect 10348 10184 10388 10193
rect 10348 9764 10388 10144
rect 10348 9715 10388 9724
rect 10251 6236 10293 6245
rect 10251 6196 10252 6236
rect 10292 6196 10293 6236
rect 10251 6187 10293 6196
rect 10348 6236 10388 6245
rect 10156 5851 10196 5860
rect 10252 5480 10292 5489
rect 10155 3464 10197 3473
rect 10155 3424 10156 3464
rect 10196 3424 10197 3464
rect 10155 3415 10197 3424
rect 10156 3330 10196 3415
rect 9868 2575 9908 2584
rect 10059 2624 10101 2633
rect 10059 2584 10060 2624
rect 10100 2584 10101 2624
rect 10059 2575 10101 2584
rect 10252 2456 10292 5440
rect 10348 3464 10388 6196
rect 10444 5648 10484 11740
rect 10540 10604 10580 13420
rect 10540 10109 10580 10564
rect 10539 10100 10581 10109
rect 10539 10060 10540 10100
rect 10580 10060 10581 10100
rect 10539 10051 10581 10060
rect 10540 9680 10580 9689
rect 10540 8924 10580 9640
rect 10636 9596 10676 20140
rect 10828 19928 10868 35260
rect 10924 33368 10964 33377
rect 10924 31268 10964 33328
rect 10924 27497 10964 31228
rect 11020 27908 11060 41560
rect 11308 36224 11348 36233
rect 11308 35804 11348 36184
rect 11308 35755 11348 35764
rect 11116 34796 11156 34805
rect 11116 32612 11156 34756
rect 11211 34208 11253 34217
rect 11211 34168 11212 34208
rect 11252 34168 11253 34208
rect 11211 34159 11253 34168
rect 11116 32192 11156 32572
rect 11116 32143 11156 32152
rect 11116 30932 11156 30941
rect 11116 30512 11156 30892
rect 11116 30463 11156 30472
rect 11115 30344 11157 30353
rect 11115 30304 11116 30344
rect 11156 30304 11157 30344
rect 11115 30295 11157 30304
rect 11020 27859 11060 27868
rect 11019 27656 11061 27665
rect 11019 27616 11020 27656
rect 11060 27616 11061 27656
rect 11019 27607 11061 27616
rect 10923 27488 10965 27497
rect 10923 27448 10924 27488
rect 10964 27448 10965 27488
rect 10923 27439 10965 27448
rect 11020 26825 11060 27607
rect 11019 26816 11061 26825
rect 11019 26776 11020 26816
rect 11060 26776 11061 26816
rect 11019 26767 11061 26776
rect 10828 19508 10868 19888
rect 10828 19459 10868 19468
rect 10924 26648 10964 26657
rect 10924 24548 10964 26608
rect 11020 25892 11060 26767
rect 11020 25843 11060 25852
rect 11116 25388 11156 30295
rect 11116 25339 11156 25348
rect 10732 19256 10772 19265
rect 10732 14057 10772 19216
rect 10827 15644 10869 15653
rect 10827 15604 10828 15644
rect 10868 15604 10869 15644
rect 10827 15595 10869 15604
rect 10924 15644 10964 24508
rect 10924 15595 10964 15604
rect 11020 19508 11060 19517
rect 10731 14048 10773 14057
rect 10731 14008 10732 14048
rect 10772 14008 10773 14048
rect 10731 13999 10773 14008
rect 10732 11696 10772 13999
rect 10732 11647 10772 11656
rect 10636 9547 10676 9556
rect 10540 8875 10580 8884
rect 10539 8756 10581 8765
rect 10539 8716 10540 8756
rect 10580 8716 10581 8756
rect 10539 8707 10581 8716
rect 10540 8336 10580 8707
rect 10540 8287 10580 8296
rect 10444 5599 10484 5608
rect 10348 3415 10388 3424
rect 10732 4640 10772 4649
rect 10732 3380 10772 4600
rect 10732 3331 10772 3340
rect 10252 2407 10292 2416
rect 9580 1903 9620 1912
rect 10828 1877 10868 15595
rect 11020 15476 11060 19468
rect 10924 15436 11060 15476
rect 10924 5396 10964 15436
rect 11020 14888 11060 14897
rect 11020 13628 11060 14848
rect 11020 13579 11060 13588
rect 11116 14804 11156 14813
rect 11116 13124 11156 14764
rect 11116 13075 11156 13084
rect 11115 10520 11157 10529
rect 11115 10480 11116 10520
rect 11156 10480 11157 10520
rect 11115 10471 11157 10480
rect 11116 10386 11156 10471
rect 11020 10352 11060 10361
rect 11020 9680 11060 10312
rect 11115 10100 11157 10109
rect 11115 10060 11116 10100
rect 11156 10060 11157 10100
rect 11115 10051 11157 10060
rect 11116 9966 11156 10051
rect 11115 9848 11157 9857
rect 11115 9808 11116 9848
rect 11156 9808 11157 9848
rect 11115 9799 11157 9808
rect 11116 9714 11156 9799
rect 11020 9631 11060 9640
rect 10924 2876 10964 5356
rect 10924 2827 10964 2836
rect 10827 1868 10869 1877
rect 10827 1828 10828 1868
rect 10868 1828 10869 1868
rect 10827 1819 10869 1828
rect 11212 1532 11252 34159
rect 11308 32528 11348 32537
rect 11308 27152 11348 32488
rect 11308 27103 11348 27112
rect 11308 26573 11348 26658
rect 11307 26564 11349 26573
rect 11307 26524 11308 26564
rect 11348 26524 11349 26564
rect 11307 26515 11349 26524
rect 11308 23624 11348 23633
rect 11308 15056 11348 23584
rect 11308 15007 11348 15016
rect 11308 13796 11348 13805
rect 11308 12032 11348 13756
rect 11308 11983 11348 11992
rect 11308 11360 11348 11369
rect 11308 10529 11348 11320
rect 11404 10697 11444 41644
rect 14763 41684 14805 41693
rect 14763 41644 14764 41684
rect 14804 41644 14805 41684
rect 14763 41635 14805 41644
rect 11500 41600 11540 41609
rect 11500 23120 11540 41560
rect 11788 41600 11828 41609
rect 11692 34376 11732 34385
rect 11595 32864 11637 32873
rect 11595 32824 11596 32864
rect 11636 32824 11637 32864
rect 11595 32815 11637 32824
rect 11596 32730 11636 32815
rect 11596 31940 11636 31949
rect 11596 28076 11636 31900
rect 11596 28027 11636 28036
rect 11500 23080 11636 23120
rect 11499 22448 11541 22457
rect 11499 22408 11500 22448
rect 11540 22408 11541 22448
rect 11499 22399 11541 22408
rect 11500 18920 11540 22399
rect 11596 21020 11636 23080
rect 11596 20971 11636 20980
rect 11500 18871 11540 18880
rect 11596 20768 11636 20777
rect 11596 18164 11636 20728
rect 11692 18332 11732 34336
rect 11788 24212 11828 41560
rect 12268 41600 12308 41609
rect 12172 39080 12212 39089
rect 11884 34796 11924 34805
rect 11884 31016 11924 34756
rect 12075 34628 12117 34637
rect 12075 34588 12076 34628
rect 12116 34588 12117 34628
rect 12075 34579 12117 34588
rect 12076 34124 12116 34579
rect 12076 34075 12116 34084
rect 11980 33032 12020 33041
rect 11980 32276 12020 32992
rect 11980 32227 12020 32236
rect 11884 30764 11924 30976
rect 11884 30715 11924 30724
rect 11980 31436 12020 31445
rect 11884 29672 11924 29681
rect 11884 28664 11924 29632
rect 11884 27740 11924 28624
rect 11884 27691 11924 27700
rect 11980 27656 12020 31396
rect 12076 31184 12116 31193
rect 12076 30176 12116 31144
rect 12172 30932 12212 39040
rect 12172 30883 12212 30892
rect 12268 30764 12308 41560
rect 12843 41348 12885 41357
rect 12843 41308 12844 41348
rect 12884 41308 12885 41348
rect 12843 41299 12885 41308
rect 12459 41096 12501 41105
rect 12459 41056 12460 41096
rect 12500 41056 12501 41096
rect 12459 41047 12501 41056
rect 12460 37904 12500 41047
rect 12844 40592 12884 41299
rect 12844 40543 12884 40552
rect 12940 40760 12980 40769
rect 12652 40424 12692 40433
rect 12555 39584 12597 39593
rect 12555 39544 12556 39584
rect 12596 39544 12597 39584
rect 12555 39535 12597 39544
rect 12556 39450 12596 39535
rect 12460 37855 12500 37864
rect 12652 37904 12692 40384
rect 12843 39668 12885 39677
rect 12843 39628 12844 39668
rect 12884 39628 12885 39668
rect 12843 39619 12885 39628
rect 12747 38072 12789 38081
rect 12747 38032 12748 38072
rect 12788 38032 12789 38072
rect 12747 38023 12789 38032
rect 12652 37855 12692 37864
rect 12076 30127 12116 30136
rect 12172 30724 12308 30764
rect 12364 37316 12404 37325
rect 11980 27607 12020 27616
rect 12076 28832 12116 28841
rect 12076 27320 12116 28792
rect 12076 27271 12116 27280
rect 11979 26816 12021 26825
rect 11979 26776 11980 26816
rect 12020 26776 12021 26816
rect 11979 26767 12021 26776
rect 11980 26682 12020 26767
rect 11788 24163 11828 24172
rect 11692 18283 11732 18292
rect 11788 23792 11828 23801
rect 11596 18115 11636 18124
rect 11691 17828 11733 17837
rect 11691 17788 11692 17828
rect 11732 17788 11733 17828
rect 11691 17779 11733 17788
rect 11500 16400 11540 16409
rect 11500 12284 11540 16360
rect 11596 15560 11636 15569
rect 11596 13292 11636 15520
rect 11596 13243 11636 13252
rect 11500 12235 11540 12244
rect 11500 10940 11540 10949
rect 11403 10688 11445 10697
rect 11403 10648 11404 10688
rect 11444 10648 11445 10688
rect 11403 10639 11445 10648
rect 11307 10520 11349 10529
rect 11307 10480 11308 10520
rect 11348 10480 11444 10520
rect 11307 10471 11349 10480
rect 11308 10386 11348 10471
rect 11212 1483 11252 1492
rect 11308 10016 11348 10025
rect 9388 1147 9428 1156
rect 8620 895 8660 904
rect 7947 860 7989 869
rect 7947 820 7948 860
rect 7988 820 7989 860
rect 7947 811 7989 820
rect 7948 726 7988 811
rect 7468 559 7508 568
rect 11308 449 11348 9976
rect 11404 7076 11444 10480
rect 11404 7027 11444 7036
rect 11500 6656 11540 10900
rect 11596 10856 11636 10865
rect 11596 7664 11636 10816
rect 11596 7615 11636 7624
rect 11596 6656 11636 6665
rect 11500 6616 11596 6656
rect 11596 6607 11636 6616
rect 11595 4220 11637 4229
rect 11595 4180 11596 4220
rect 11636 4180 11637 4220
rect 11595 4171 11637 4180
rect 11596 4086 11636 4171
rect 11307 440 11349 449
rect 11307 400 11308 440
rect 11348 400 11349 440
rect 11307 391 11349 400
rect 5068 113 5108 198
rect 11692 113 11732 17779
rect 11788 10865 11828 23752
rect 12076 22868 12116 22877
rect 12076 19256 12116 22828
rect 12172 20852 12212 30724
rect 12364 30092 12404 37276
rect 12652 36812 12692 36821
rect 12460 36560 12500 36569
rect 12460 33368 12500 36520
rect 12555 36560 12597 36569
rect 12555 36520 12556 36560
rect 12596 36520 12597 36560
rect 12555 36511 12597 36520
rect 12556 33629 12596 36511
rect 12555 33620 12597 33629
rect 12555 33580 12556 33620
rect 12596 33580 12597 33620
rect 12555 33571 12597 33580
rect 12460 33328 12596 33368
rect 12268 30052 12404 30092
rect 12460 33200 12500 33209
rect 12268 29252 12308 30052
rect 12268 29203 12308 29212
rect 12364 29924 12404 29933
rect 12364 27824 12404 29884
rect 12364 27775 12404 27784
rect 12460 27665 12500 33160
rect 12267 27656 12309 27665
rect 12267 27616 12268 27656
rect 12308 27616 12309 27656
rect 12267 27607 12309 27616
rect 12459 27656 12501 27665
rect 12459 27616 12460 27656
rect 12500 27616 12501 27656
rect 12459 27607 12501 27616
rect 12268 26060 12308 27607
rect 12459 27488 12501 27497
rect 12459 27448 12460 27488
rect 12500 27448 12501 27488
rect 12459 27439 12501 27448
rect 12268 26011 12308 26020
rect 12172 20803 12212 20812
rect 12268 25472 12308 25481
rect 12268 20096 12308 25432
rect 12268 20047 12308 20056
rect 12364 20264 12404 20273
rect 12076 19216 12212 19256
rect 12076 19088 12116 19097
rect 11884 19004 11924 19013
rect 11787 10856 11829 10865
rect 11787 10816 11788 10856
rect 11828 10816 11829 10856
rect 11787 10807 11829 10816
rect 11788 10688 11828 10697
rect 11788 9848 11828 10648
rect 11884 10352 11924 18964
rect 12076 11201 12116 19048
rect 12172 19004 12212 19216
rect 12172 18955 12212 18964
rect 12268 18500 12308 18509
rect 12172 14468 12212 14477
rect 12172 12620 12212 14428
rect 12172 12571 12212 12580
rect 11980 11192 12020 11201
rect 11980 10781 12020 11152
rect 12075 11192 12117 11201
rect 12075 11152 12076 11192
rect 12116 11152 12117 11192
rect 12075 11143 12117 11152
rect 12171 10856 12213 10865
rect 12171 10816 12172 10856
rect 12212 10816 12213 10856
rect 12171 10807 12213 10816
rect 11979 10772 12021 10781
rect 11979 10732 11980 10772
rect 12020 10732 12021 10772
rect 11979 10723 12021 10732
rect 11884 10303 11924 10312
rect 11788 9799 11828 9808
rect 12076 10100 12116 10109
rect 12076 8756 12116 10060
rect 12076 8707 12116 8716
rect 11980 8504 12020 8513
rect 11788 7832 11828 7841
rect 11788 6404 11828 7792
rect 11883 7832 11925 7841
rect 11883 7792 11884 7832
rect 11924 7792 11925 7832
rect 11883 7783 11925 7792
rect 11788 6355 11828 6364
rect 11788 5648 11828 5657
rect 11788 2792 11828 5608
rect 11788 2743 11828 2752
rect 11884 113 11924 7783
rect 11980 7580 12020 8464
rect 11980 6068 12020 7540
rect 11980 6019 12020 6028
rect 12172 7748 12212 10807
rect 12268 8588 12308 18460
rect 12364 13544 12404 20224
rect 12364 13495 12404 13504
rect 12460 18584 12500 27439
rect 12556 25556 12596 33328
rect 12556 25507 12596 25516
rect 12652 23960 12692 36772
rect 12748 35804 12788 38023
rect 12748 35755 12788 35764
rect 12844 33461 12884 39619
rect 12940 36989 12980 40720
rect 14667 39920 14709 39929
rect 14667 39880 14668 39920
rect 14708 39880 14709 39920
rect 14667 39871 14709 39880
rect 13131 39500 13173 39509
rect 13131 39460 13132 39500
rect 13172 39460 13173 39500
rect 13131 39451 13173 39460
rect 14571 39500 14613 39509
rect 14571 39460 14572 39500
rect 14612 39460 14613 39500
rect 14571 39451 14613 39460
rect 12939 36980 12981 36989
rect 12939 36940 12940 36980
rect 12980 36940 12981 36980
rect 12939 36931 12981 36940
rect 12940 35720 12980 35729
rect 12843 33452 12885 33461
rect 12843 33412 12844 33452
rect 12884 33412 12885 33452
rect 12843 33403 12885 33412
rect 12844 31436 12884 31445
rect 12844 30764 12884 31396
rect 12844 30715 12884 30724
rect 12844 30176 12884 30185
rect 12748 29924 12788 29933
rect 12748 28076 12788 29884
rect 12748 28027 12788 28036
rect 12844 27749 12884 30136
rect 12843 27740 12885 27749
rect 12843 27700 12844 27740
rect 12884 27700 12885 27740
rect 12843 27691 12885 27700
rect 12844 26573 12884 26658
rect 12843 26564 12885 26573
rect 12843 26524 12844 26564
rect 12884 26524 12885 26564
rect 12843 26515 12885 26524
rect 12652 23911 12692 23920
rect 12844 25388 12884 25397
rect 12652 23792 12692 23801
rect 12652 22112 12692 23752
rect 12652 22063 12692 22072
rect 12748 22028 12788 22037
rect 12460 12461 12500 18544
rect 12652 20264 12692 20273
rect 12652 18584 12692 20224
rect 12652 18535 12692 18544
rect 12556 16400 12596 16409
rect 12556 15812 12596 16360
rect 12556 15763 12596 15772
rect 12459 12452 12501 12461
rect 12459 12412 12460 12452
rect 12500 12412 12501 12452
rect 12459 12403 12501 12412
rect 12748 10445 12788 21988
rect 12844 21104 12884 25348
rect 12844 21055 12884 21064
rect 12844 19256 12884 19265
rect 12844 16652 12884 19216
rect 12844 16603 12884 16612
rect 12843 16316 12885 16325
rect 12843 16276 12844 16316
rect 12884 16276 12885 16316
rect 12843 16267 12885 16276
rect 12555 10436 12597 10445
rect 12555 10396 12556 10436
rect 12596 10396 12597 10436
rect 12555 10387 12597 10396
rect 12747 10436 12789 10445
rect 12747 10396 12748 10436
rect 12788 10396 12789 10436
rect 12747 10387 12789 10396
rect 12364 10352 12404 10361
rect 12364 9092 12404 10312
rect 12556 9848 12596 10387
rect 12748 10268 12788 10277
rect 12556 9808 12692 9848
rect 12364 9043 12404 9052
rect 12556 9680 12596 9689
rect 12556 9092 12596 9640
rect 12556 9043 12596 9052
rect 12652 9008 12692 9808
rect 12652 8959 12692 8968
rect 12364 8756 12404 8765
rect 12364 8597 12404 8716
rect 12651 8756 12693 8765
rect 12651 8716 12652 8756
rect 12692 8716 12693 8756
rect 12651 8707 12693 8716
rect 12652 8622 12692 8707
rect 12268 8539 12308 8548
rect 12363 8588 12405 8597
rect 12363 8548 12364 8588
rect 12404 8548 12405 8588
rect 12363 8539 12405 8548
rect 12748 8504 12788 10228
rect 12748 8455 12788 8464
rect 12076 5480 12116 5489
rect 12076 4313 12116 5440
rect 12172 4976 12212 7708
rect 12844 8084 12884 16267
rect 12267 7664 12309 7673
rect 12267 7624 12268 7664
rect 12308 7624 12309 7664
rect 12267 7615 12309 7624
rect 12172 4927 12212 4936
rect 12075 4304 12117 4313
rect 12075 4264 12076 4304
rect 12116 4264 12117 4304
rect 12075 4255 12117 4264
rect 12076 3380 12116 4255
rect 12172 3380 12212 3389
rect 12076 3340 12172 3380
rect 12172 356 12212 3340
rect 12268 2540 12308 7615
rect 12555 7580 12597 7589
rect 12555 7540 12556 7580
rect 12596 7540 12597 7580
rect 12555 7531 12597 7540
rect 12844 7580 12884 8044
rect 12844 7531 12884 7540
rect 12364 6656 12404 6665
rect 12364 4976 12404 6616
rect 12364 4927 12404 4936
rect 12460 5564 12500 5573
rect 12460 4556 12500 5524
rect 12460 4507 12500 4516
rect 12556 3380 12596 7531
rect 12652 7244 12692 7253
rect 12652 3464 12692 7204
rect 12652 3415 12692 3424
rect 12460 3340 12596 3380
rect 12460 2540 12500 3340
rect 12555 3212 12597 3221
rect 12555 3172 12556 3212
rect 12596 3172 12597 3212
rect 12555 3163 12597 3172
rect 12556 3078 12596 3163
rect 12268 2500 12404 2540
rect 12460 2500 12596 2540
rect 12364 1121 12404 2500
rect 12363 1112 12405 1121
rect 12363 1072 12364 1112
rect 12404 1072 12405 1112
rect 12363 1063 12405 1072
rect 12556 944 12596 2500
rect 12556 895 12596 904
rect 12940 944 12980 35680
rect 13035 34544 13077 34553
rect 13035 34504 13036 34544
rect 13076 34504 13077 34544
rect 13035 34495 13077 34504
rect 13036 34292 13076 34495
rect 13036 34243 13076 34252
rect 13035 33452 13077 33461
rect 13035 33412 13036 33452
rect 13076 33412 13077 33452
rect 13035 33403 13077 33412
rect 13036 24380 13076 33403
rect 13036 24331 13076 24340
rect 13036 23960 13076 23969
rect 13036 22868 13076 23920
rect 13036 22819 13076 22828
rect 13035 16316 13077 16325
rect 13035 16276 13036 16316
rect 13076 16276 13077 16316
rect 13035 16267 13077 16276
rect 13036 11024 13076 16267
rect 13036 10975 13076 10984
rect 13036 10352 13076 10361
rect 13036 6488 13076 10312
rect 13036 6439 13076 6448
rect 13132 2045 13172 39451
rect 14572 39416 14612 39451
rect 14572 39365 14612 39376
rect 13899 39248 13941 39257
rect 13899 39208 13900 39248
rect 13940 39208 13941 39248
rect 13899 39199 13941 39208
rect 13324 38408 13364 38417
rect 13228 35468 13268 35477
rect 13228 24044 13268 35428
rect 13324 33788 13364 38368
rect 13708 38324 13748 38333
rect 13611 38072 13653 38081
rect 13611 38032 13612 38072
rect 13652 38032 13653 38072
rect 13611 38023 13653 38032
rect 13516 35048 13556 35057
rect 13324 33620 13364 33748
rect 13324 33571 13364 33580
rect 13420 34628 13460 34637
rect 13228 23995 13268 24004
rect 13324 29252 13364 29261
rect 13228 21356 13268 21365
rect 13228 10025 13268 21316
rect 13324 16232 13364 29212
rect 13420 29177 13460 34588
rect 13419 29168 13461 29177
rect 13419 29128 13420 29168
rect 13460 29128 13461 29168
rect 13419 29119 13461 29128
rect 13420 29034 13460 29119
rect 13420 22364 13460 22373
rect 13420 18416 13460 22324
rect 13420 18367 13460 18376
rect 13324 15140 13364 16192
rect 13419 15896 13461 15905
rect 13419 15856 13420 15896
rect 13460 15856 13461 15896
rect 13419 15847 13461 15856
rect 13420 15762 13460 15847
rect 13420 15140 13460 15149
rect 13324 15100 13420 15140
rect 13324 14636 13364 14645
rect 13324 10100 13364 14596
rect 13324 10051 13364 10060
rect 13227 10016 13269 10025
rect 13227 9976 13228 10016
rect 13268 9976 13269 10016
rect 13227 9967 13269 9976
rect 13420 9857 13460 15100
rect 13419 9848 13461 9857
rect 13419 9808 13420 9848
rect 13460 9808 13461 9848
rect 13419 9799 13461 9808
rect 13324 9092 13364 9101
rect 13131 2036 13173 2045
rect 13131 1996 13132 2036
rect 13172 1996 13173 2036
rect 13131 1987 13173 1996
rect 13324 1280 13364 9052
rect 13324 1231 13364 1240
rect 12940 895 12980 904
rect 13516 944 13556 35008
rect 13612 23960 13652 38023
rect 13708 36056 13748 38284
rect 13900 37820 13940 39199
rect 14187 38912 14229 38921
rect 14187 38872 14188 38912
rect 14228 38872 14229 38912
rect 14187 38863 14229 38872
rect 14188 38072 14228 38863
rect 14379 38492 14421 38501
rect 14379 38452 14380 38492
rect 14420 38452 14421 38492
rect 14379 38443 14421 38452
rect 14188 38023 14228 38032
rect 13900 37771 13940 37780
rect 13900 37652 13940 37661
rect 13900 37232 13940 37612
rect 13900 37183 13940 37192
rect 13708 36007 13748 36016
rect 13996 37148 14036 37157
rect 13996 34469 14036 37108
rect 14187 35300 14229 35309
rect 14187 35260 14188 35300
rect 14228 35260 14229 35300
rect 14187 35251 14229 35260
rect 14092 35216 14132 35225
rect 13995 34460 14037 34469
rect 13995 34420 13996 34460
rect 14036 34420 14037 34460
rect 13995 34411 14037 34420
rect 13803 33116 13845 33125
rect 13803 33076 13804 33116
rect 13844 33076 13845 33116
rect 13803 33067 13845 33076
rect 13804 32957 13844 33067
rect 13803 32948 13845 32957
rect 13803 32908 13804 32948
rect 13844 32908 13845 32948
rect 13803 32899 13845 32908
rect 13899 32528 13941 32537
rect 13899 32488 13900 32528
rect 13940 32488 13941 32528
rect 13899 32479 13941 32488
rect 13900 32394 13940 32479
rect 13804 31604 13844 31613
rect 13804 31352 13844 31564
rect 13804 31303 13844 31312
rect 13707 31268 13749 31277
rect 13707 31228 13708 31268
rect 13748 31228 13749 31268
rect 13707 31219 13749 31228
rect 13708 31134 13748 31219
rect 13900 29420 13940 29429
rect 13900 29084 13940 29380
rect 13612 23911 13652 23920
rect 13708 28916 13748 28925
rect 13611 22532 13653 22541
rect 13611 22492 13612 22532
rect 13652 22492 13653 22532
rect 13611 22483 13653 22492
rect 13612 22398 13652 22483
rect 13612 20180 13652 20189
rect 13612 19676 13652 20140
rect 13612 19627 13652 19636
rect 13708 17660 13748 28876
rect 13900 26480 13940 29044
rect 13996 29000 14036 34411
rect 14092 33041 14132 35176
rect 14091 33032 14133 33041
rect 14091 32992 14092 33032
rect 14132 32992 14133 33032
rect 14091 32983 14133 32992
rect 14092 32780 14132 32789
rect 14092 30932 14132 32740
rect 14092 30883 14132 30892
rect 14188 29000 14228 35251
rect 14283 33032 14325 33041
rect 14283 32992 14284 33032
rect 14324 32992 14325 33032
rect 14283 32983 14325 32992
rect 14284 32948 14324 32983
rect 14284 32897 14324 32908
rect 14284 32444 14324 32453
rect 14284 31184 14324 32404
rect 14284 31135 14324 31144
rect 13996 28960 14132 29000
rect 14188 28960 14324 29000
rect 13900 26431 13940 26440
rect 13996 25724 14036 25733
rect 13996 23708 14036 25684
rect 13996 23659 14036 23668
rect 13996 22448 14036 22457
rect 13900 18920 13940 18929
rect 13612 17492 13652 17501
rect 13612 14636 13652 17452
rect 13708 14720 13748 17620
rect 13804 18880 13900 18920
rect 13804 15737 13844 18880
rect 13900 18871 13940 18880
rect 13900 17753 13940 17755
rect 13899 17744 13941 17753
rect 13899 17704 13900 17744
rect 13940 17704 13941 17744
rect 13899 17695 13941 17704
rect 13900 17660 13940 17695
rect 13900 17611 13940 17620
rect 13900 16904 13940 16913
rect 13900 16232 13940 16864
rect 13803 15728 13845 15737
rect 13803 15688 13804 15728
rect 13844 15688 13845 15728
rect 13803 15679 13845 15688
rect 13708 14671 13748 14680
rect 13612 14587 13652 14596
rect 13516 895 13556 904
rect 13708 9680 13748 9689
rect 13708 944 13748 9640
rect 13804 5069 13844 15679
rect 13900 14972 13940 16192
rect 13900 11864 13940 14932
rect 13900 11815 13940 11824
rect 13996 12116 14036 22408
rect 14092 18920 14132 28960
rect 14092 18871 14132 18880
rect 14188 20600 14228 20609
rect 14188 20348 14228 20560
rect 14188 19256 14228 20308
rect 14188 17744 14228 19216
rect 14188 17695 14228 17704
rect 14092 17492 14132 17501
rect 14092 13796 14132 17452
rect 14092 13747 14132 13756
rect 14188 16652 14228 16661
rect 14188 15476 14228 16612
rect 13996 11453 14036 12076
rect 13995 11444 14037 11453
rect 13995 11404 13996 11444
rect 14036 11404 14037 11444
rect 13995 11395 14037 11404
rect 13899 10100 13941 10109
rect 13899 10060 13900 10100
rect 13940 10060 13941 10100
rect 13899 10051 13941 10060
rect 13900 9764 13940 10051
rect 13900 9715 13940 9724
rect 14188 9680 14228 15436
rect 13996 9640 14228 9680
rect 13900 8336 13940 8345
rect 13900 7916 13940 8296
rect 13900 7867 13940 7876
rect 13899 6488 13941 6497
rect 13899 6448 13900 6488
rect 13940 6448 13941 6488
rect 13899 6439 13941 6448
rect 13900 5228 13940 6439
rect 13900 5179 13940 5188
rect 13803 5060 13845 5069
rect 13803 5020 13804 5060
rect 13844 5020 13845 5060
rect 13803 5011 13845 5020
rect 13996 4817 14036 9640
rect 14187 9512 14229 9521
rect 14187 9472 14188 9512
rect 14228 9472 14229 9512
rect 14187 9463 14229 9472
rect 14092 8336 14132 8345
rect 14092 6497 14132 8296
rect 14091 6488 14133 6497
rect 14091 6448 14092 6488
rect 14132 6448 14133 6488
rect 14091 6439 14133 6448
rect 14188 6236 14228 9463
rect 14188 6187 14228 6196
rect 13995 4808 14037 4817
rect 13995 4768 13996 4808
rect 14036 4768 14037 4808
rect 13995 4759 14037 4768
rect 14284 1280 14324 28960
rect 14380 23297 14420 38443
rect 14476 37904 14516 37913
rect 14476 36896 14516 37864
rect 14476 36847 14516 36856
rect 14572 35132 14612 35141
rect 14475 34124 14517 34133
rect 14475 34084 14476 34124
rect 14516 34084 14517 34124
rect 14475 34075 14517 34084
rect 14379 23288 14421 23297
rect 14379 23248 14380 23288
rect 14420 23248 14421 23288
rect 14379 23239 14421 23248
rect 14380 18752 14420 18761
rect 14380 17912 14420 18712
rect 14380 17863 14420 17872
rect 14380 14720 14420 14729
rect 14380 1793 14420 14680
rect 14379 1784 14421 1793
rect 14379 1744 14380 1784
rect 14420 1744 14421 1784
rect 14379 1735 14421 1744
rect 14284 1231 14324 1240
rect 14476 1280 14516 34075
rect 14572 31940 14612 35092
rect 14572 31891 14612 31900
rect 14572 25388 14612 25397
rect 14572 15896 14612 25348
rect 14572 15847 14612 15856
rect 14668 15728 14708 39871
rect 14764 25556 14804 41635
rect 15436 41012 15476 41021
rect 15147 40424 15189 40433
rect 15147 40384 15148 40424
rect 15188 40384 15189 40424
rect 15147 40375 15189 40384
rect 15148 40256 15188 40375
rect 15148 40207 15188 40216
rect 15052 40172 15092 40181
rect 14859 38996 14901 39005
rect 14859 38956 14860 38996
rect 14900 38956 14901 38996
rect 14859 38947 14901 38956
rect 14764 25507 14804 25516
rect 14764 24296 14804 24305
rect 14764 23456 14804 24256
rect 14764 23407 14804 23416
rect 14763 22700 14805 22709
rect 14763 22660 14764 22700
rect 14804 22660 14805 22700
rect 14763 22651 14805 22660
rect 14764 20180 14804 22651
rect 14764 20131 14804 20140
rect 14763 18920 14805 18929
rect 14763 18880 14764 18920
rect 14804 18880 14805 18920
rect 14763 18871 14805 18880
rect 14572 15688 14708 15728
rect 14572 11360 14612 15688
rect 14667 15224 14709 15233
rect 14667 15184 14668 15224
rect 14708 15184 14709 15224
rect 14667 15175 14709 15184
rect 14668 14888 14708 15175
rect 14668 14839 14708 14848
rect 14572 11320 14708 11360
rect 14571 7160 14613 7169
rect 14571 7120 14572 7160
rect 14612 7120 14613 7160
rect 14571 7111 14613 7120
rect 14572 6572 14612 7111
rect 14572 6523 14612 6532
rect 14476 1231 14516 1240
rect 14668 1280 14708 11320
rect 14764 1289 14804 18871
rect 14860 6320 14900 38947
rect 14955 38912 14997 38921
rect 14955 38872 14956 38912
rect 14996 38872 14997 38912
rect 14955 38863 14997 38872
rect 14956 38778 14996 38863
rect 15052 37988 15092 40132
rect 15244 40004 15284 40013
rect 15244 39761 15284 39964
rect 15243 39752 15285 39761
rect 15243 39712 15244 39752
rect 15284 39712 15285 39752
rect 15243 39703 15285 39712
rect 15148 38912 15188 38921
rect 15148 38744 15188 38872
rect 15148 38695 15188 38704
rect 15052 37939 15092 37948
rect 15244 38408 15284 38417
rect 15244 37064 15284 38368
rect 15244 37015 15284 37024
rect 15340 37736 15380 37745
rect 15340 36980 15380 37696
rect 15340 36728 15380 36940
rect 15244 36392 15284 36401
rect 15147 34208 15189 34217
rect 15147 34168 15148 34208
rect 15188 34168 15189 34208
rect 15147 34159 15189 34168
rect 14955 34040 14997 34049
rect 14955 34000 14956 34040
rect 14996 34000 14997 34040
rect 14955 33991 14997 34000
rect 14956 24800 14996 33991
rect 14956 24751 14996 24760
rect 15052 30008 15092 30017
rect 14955 19928 14997 19937
rect 14955 19888 14956 19928
rect 14996 19888 14997 19928
rect 14955 19879 14997 19888
rect 14956 19676 14996 19879
rect 14956 19627 14996 19636
rect 14956 19256 14996 19265
rect 14956 18332 14996 19216
rect 14956 18283 14996 18292
rect 14956 17753 14996 17838
rect 14955 17744 14997 17753
rect 14955 17704 14956 17744
rect 14996 17704 14997 17744
rect 14955 17695 14997 17704
rect 14860 6271 14900 6280
rect 14956 16232 14996 16241
rect 14956 3548 14996 16192
rect 15052 15476 15092 29968
rect 15052 15427 15092 15436
rect 15051 6488 15093 6497
rect 15051 6448 15052 6488
rect 15092 6448 15093 6488
rect 15051 6439 15093 6448
rect 15052 6354 15092 6439
rect 14956 3499 14996 3508
rect 14955 3296 14997 3305
rect 14955 3256 14956 3296
rect 14996 3256 14997 3296
rect 14955 3247 14997 3256
rect 14956 3162 14996 3247
rect 15148 2540 15188 34159
rect 15244 26480 15284 36352
rect 15244 26431 15284 26440
rect 15244 24632 15284 24641
rect 15244 10688 15284 24592
rect 15340 24128 15380 36688
rect 15436 35225 15476 40972
rect 15435 35216 15477 35225
rect 15435 35176 15436 35216
rect 15476 35176 15477 35216
rect 15435 35167 15477 35176
rect 15436 33452 15476 33461
rect 15436 29252 15476 33412
rect 15436 29203 15476 29212
rect 15532 27068 15572 42904
rect 21100 42776 21140 42785
rect 18316 42692 18356 42701
rect 18028 42608 18068 42617
rect 16395 42272 16437 42281
rect 16395 42232 16396 42272
rect 16436 42232 16437 42272
rect 16395 42223 16437 42232
rect 16300 42020 16340 42029
rect 16300 41600 16340 41980
rect 16396 41768 16436 42223
rect 16396 41719 16436 41728
rect 17932 41936 17972 41945
rect 16300 41560 16436 41600
rect 15724 41516 15764 41525
rect 15628 41180 15668 41189
rect 15628 40172 15668 41140
rect 15628 40123 15668 40132
rect 15724 40088 15764 41476
rect 16396 41180 16436 41560
rect 16396 41131 16436 41140
rect 17164 41516 17204 41525
rect 16396 41012 16436 41021
rect 16011 40928 16053 40937
rect 16011 40888 16012 40928
rect 16052 40888 16053 40928
rect 16011 40879 16053 40888
rect 15724 40039 15764 40048
rect 15820 39500 15860 39509
rect 15628 38996 15668 39005
rect 15628 38072 15668 38956
rect 15628 38023 15668 38032
rect 15724 37820 15764 37829
rect 15724 36392 15764 37780
rect 15724 36343 15764 36352
rect 15627 34376 15669 34385
rect 15627 34336 15628 34376
rect 15668 34336 15669 34376
rect 15627 34327 15669 34336
rect 15628 31352 15668 34327
rect 15724 34124 15764 34133
rect 15724 31520 15764 34084
rect 15724 31471 15764 31480
rect 15628 31312 15764 31352
rect 15627 29588 15669 29597
rect 15627 29548 15628 29588
rect 15668 29548 15669 29588
rect 15627 29539 15669 29548
rect 15532 27019 15572 27028
rect 15532 26900 15572 26909
rect 15340 24079 15380 24088
rect 15436 24464 15476 24473
rect 15436 20600 15476 24424
rect 15436 20551 15476 20560
rect 15340 20012 15380 20021
rect 15340 19760 15380 19972
rect 15340 19711 15380 19720
rect 15435 16904 15477 16913
rect 15435 16864 15436 16904
rect 15476 16864 15477 16904
rect 15435 16855 15477 16864
rect 15340 16652 15380 16661
rect 15340 11108 15380 16612
rect 15436 14888 15476 16855
rect 15436 14839 15476 14848
rect 15436 13796 15476 13805
rect 15436 11612 15476 13756
rect 15436 11563 15476 11572
rect 15340 11059 15380 11068
rect 15244 10648 15380 10688
rect 15244 10520 15284 10529
rect 15244 9260 15284 10480
rect 15244 9211 15284 9220
rect 15340 8681 15380 10648
rect 15436 10520 15476 10529
rect 15436 9344 15476 10480
rect 15436 9295 15476 9304
rect 15435 8756 15477 8765
rect 15435 8716 15436 8756
rect 15476 8716 15477 8756
rect 15435 8707 15477 8716
rect 15339 8672 15381 8681
rect 15339 8632 15340 8672
rect 15380 8632 15381 8672
rect 15339 8623 15381 8632
rect 15340 8538 15380 8623
rect 15244 8252 15284 8261
rect 15244 4976 15284 8212
rect 15340 7328 15380 7337
rect 15340 6656 15380 7288
rect 15340 6607 15380 6616
rect 15244 4927 15284 4936
rect 15244 4136 15284 4145
rect 15244 3128 15284 4096
rect 15244 3079 15284 3088
rect 15148 2500 15380 2540
rect 14668 1231 14708 1240
rect 14763 1280 14805 1289
rect 14763 1240 14764 1280
rect 14804 1240 14805 1280
rect 14763 1231 14805 1240
rect 13708 895 13748 904
rect 15148 1196 15188 1205
rect 13131 860 13173 869
rect 13131 820 13132 860
rect 13172 820 13173 860
rect 13131 811 13173 820
rect 13132 726 13172 811
rect 13899 692 13941 701
rect 13899 652 13900 692
rect 13940 652 13941 692
rect 13899 643 13941 652
rect 13900 558 13940 643
rect 15148 608 15188 1156
rect 15340 692 15380 2500
rect 15436 1616 15476 8707
rect 15532 2540 15572 26860
rect 15628 24641 15668 29539
rect 15627 24632 15669 24641
rect 15627 24592 15628 24632
rect 15668 24592 15669 24632
rect 15627 24583 15669 24592
rect 15628 21104 15668 21113
rect 15628 20012 15668 21064
rect 15628 19963 15668 19972
rect 15628 16148 15668 16157
rect 15628 7328 15668 16108
rect 15724 7664 15764 31312
rect 15820 29084 15860 39460
rect 16012 39341 16052 40879
rect 16108 40424 16148 40433
rect 16108 40004 16148 40384
rect 16396 40424 16436 40972
rect 16588 41012 16628 41021
rect 16588 40676 16628 40972
rect 17067 41012 17109 41021
rect 17067 40972 17068 41012
rect 17108 40972 17109 41012
rect 17067 40963 17109 40972
rect 17068 40878 17108 40963
rect 16588 40627 16628 40636
rect 16396 40375 16436 40384
rect 16971 40424 17013 40433
rect 16971 40384 16972 40424
rect 17012 40384 17013 40424
rect 16971 40375 17013 40384
rect 16108 39955 16148 39964
rect 16300 40340 16340 40349
rect 16011 39332 16053 39341
rect 16011 39292 16012 39332
rect 16052 39292 16053 39332
rect 16011 39283 16053 39292
rect 16203 39332 16245 39341
rect 16203 39292 16204 39332
rect 16244 39292 16245 39332
rect 16203 39283 16245 39292
rect 15915 39080 15957 39089
rect 15915 39040 15916 39080
rect 15956 39040 15957 39080
rect 15915 39031 15957 39040
rect 15916 34049 15956 39031
rect 16011 38744 16053 38753
rect 16011 38704 16012 38744
rect 16052 38704 16053 38744
rect 16011 38695 16053 38704
rect 16012 36644 16052 38695
rect 16012 36595 16052 36604
rect 16108 38240 16148 38249
rect 16108 35804 16148 38200
rect 16012 35300 16052 35309
rect 15915 34040 15957 34049
rect 15915 34000 15916 34040
rect 15956 34000 15957 34040
rect 15915 33991 15957 34000
rect 15820 29035 15860 29044
rect 15916 33200 15956 33209
rect 15819 24632 15861 24641
rect 15819 24592 15820 24632
rect 15860 24592 15861 24632
rect 15819 24583 15861 24592
rect 15820 15560 15860 24583
rect 15916 22196 15956 33160
rect 16012 33125 16052 35260
rect 16011 33116 16053 33125
rect 16011 33076 16012 33116
rect 16052 33076 16053 33116
rect 16011 33067 16053 33076
rect 16012 32612 16052 32621
rect 16012 32360 16052 32572
rect 16012 32311 16052 32320
rect 16012 30680 16052 30689
rect 16012 28580 16052 30640
rect 16012 28531 16052 28540
rect 15916 22147 15956 22156
rect 16012 28328 16052 28337
rect 16012 25724 16052 28288
rect 15916 21944 15956 21953
rect 15916 17156 15956 21904
rect 15916 16325 15956 17116
rect 16012 16820 16052 25684
rect 16012 16771 16052 16780
rect 15915 16316 15957 16325
rect 15915 16276 15916 16316
rect 15956 16276 15957 16316
rect 15915 16267 15957 16276
rect 15820 15511 15860 15520
rect 16012 15896 16052 15905
rect 15916 15476 15956 15485
rect 15820 15224 15860 15233
rect 15820 8336 15860 15184
rect 15916 12452 15956 15436
rect 15916 12403 15956 12412
rect 15915 12032 15957 12041
rect 15915 11992 15916 12032
rect 15956 11992 15957 12032
rect 15915 11983 15957 11992
rect 15820 8287 15860 8296
rect 15724 7624 15860 7664
rect 15628 7279 15668 7288
rect 15724 6236 15764 6245
rect 15724 3632 15764 6196
rect 15724 3583 15764 3592
rect 15627 3296 15669 3305
rect 15627 3256 15628 3296
rect 15668 3256 15669 3296
rect 15627 3247 15669 3256
rect 15628 3162 15668 3247
rect 15532 2500 15764 2540
rect 15436 1567 15476 1576
rect 15340 643 15380 652
rect 15148 559 15188 568
rect 15724 608 15764 2500
rect 15820 1961 15860 7624
rect 15916 6152 15956 11983
rect 15916 6103 15956 6112
rect 15819 1952 15861 1961
rect 15819 1912 15820 1952
rect 15860 1912 15861 1952
rect 15819 1903 15861 1912
rect 16012 776 16052 15856
rect 16108 14552 16148 35764
rect 16204 34133 16244 39283
rect 16300 36140 16340 40300
rect 16972 40290 17012 40375
rect 16972 39920 17012 39929
rect 16395 39752 16437 39761
rect 16395 39712 16396 39752
rect 16436 39712 16437 39752
rect 16395 39703 16437 39712
rect 16396 39618 16436 39703
rect 16491 39500 16533 39509
rect 16491 39460 16492 39500
rect 16532 39460 16533 39500
rect 16491 39451 16533 39460
rect 16492 39366 16532 39451
rect 16395 39248 16437 39257
rect 16395 39208 16396 39248
rect 16436 39208 16437 39248
rect 16395 39199 16437 39208
rect 16396 39114 16436 39199
rect 16875 39164 16917 39173
rect 16875 39124 16876 39164
rect 16916 39124 16917 39164
rect 16875 39115 16917 39124
rect 16683 38408 16725 38417
rect 16683 38368 16684 38408
rect 16724 38368 16725 38408
rect 16683 38359 16725 38368
rect 16588 38324 16628 38333
rect 16300 36091 16340 36100
rect 16396 37568 16436 37577
rect 16396 35804 16436 37528
rect 16396 35755 16436 35764
rect 16396 34964 16436 34973
rect 16203 34124 16245 34133
rect 16203 34084 16204 34124
rect 16244 34084 16245 34124
rect 16203 34075 16245 34084
rect 16204 33956 16244 33965
rect 16204 31268 16244 33916
rect 16300 33284 16340 33293
rect 16300 32612 16340 33244
rect 16300 32563 16340 32572
rect 16396 31604 16436 34924
rect 16396 31555 16436 31564
rect 16492 34292 16532 34301
rect 16204 31219 16244 31228
rect 16204 31016 16244 31025
rect 16204 28328 16244 30976
rect 16204 28279 16244 28288
rect 16492 29756 16532 34252
rect 16588 33872 16628 38284
rect 16684 35468 16724 38359
rect 16684 35419 16724 35428
rect 16780 37568 16820 37577
rect 16588 30092 16628 33832
rect 16588 30043 16628 30052
rect 16684 31940 16724 31949
rect 16684 29924 16724 31900
rect 16684 29875 16724 29884
rect 16492 26480 16532 29716
rect 16492 26431 16532 26440
rect 16492 24212 16532 24221
rect 16300 22700 16340 22709
rect 16204 21524 16244 21533
rect 16204 19760 16244 21484
rect 16204 19711 16244 19720
rect 16300 15056 16340 22660
rect 16396 20684 16436 20693
rect 16396 20096 16436 20644
rect 16396 20047 16436 20056
rect 16396 18836 16436 18845
rect 16396 17996 16436 18796
rect 16492 18668 16532 24172
rect 16780 23960 16820 37528
rect 16876 30848 16916 39115
rect 16972 38744 17012 39880
rect 17164 39164 17204 41476
rect 17164 39115 17204 39124
rect 17260 41432 17300 41441
rect 16972 38324 17012 38704
rect 16972 38275 17012 38284
rect 17260 38156 17300 41392
rect 17548 41012 17588 41021
rect 17452 40424 17492 40433
rect 17452 39173 17492 40384
rect 17548 40349 17588 40972
rect 17740 40760 17780 40769
rect 17547 40340 17589 40349
rect 17547 40300 17548 40340
rect 17588 40300 17589 40340
rect 17547 40291 17589 40300
rect 17643 39332 17685 39341
rect 17643 39292 17644 39332
rect 17684 39292 17685 39332
rect 17643 39283 17685 39292
rect 17644 39198 17684 39283
rect 17451 39164 17493 39173
rect 17451 39124 17452 39164
rect 17492 39124 17493 39164
rect 17451 39115 17493 39124
rect 16971 37400 17013 37409
rect 16971 37360 16972 37400
rect 17012 37360 17013 37400
rect 16971 37351 17013 37360
rect 16876 30799 16916 30808
rect 16780 23911 16820 23920
rect 16876 28580 16916 28589
rect 16683 23624 16725 23633
rect 16683 23584 16684 23624
rect 16724 23584 16725 23624
rect 16683 23575 16725 23584
rect 16492 18619 16532 18628
rect 16588 22112 16628 22121
rect 16396 17947 16436 17956
rect 16588 16232 16628 22072
rect 16588 16183 16628 16192
rect 16684 19172 16724 23575
rect 16876 23288 16916 28540
rect 16876 23239 16916 23248
rect 16395 15308 16437 15317
rect 16395 15268 16396 15308
rect 16436 15268 16437 15308
rect 16395 15259 16437 15268
rect 16108 14503 16148 14512
rect 16204 15016 16340 15056
rect 16107 14048 16149 14057
rect 16107 14008 16108 14048
rect 16148 14008 16149 14048
rect 16107 13999 16149 14008
rect 16108 13914 16148 13999
rect 16108 11528 16148 11537
rect 16108 11360 16148 11488
rect 16108 11311 16148 11320
rect 16107 9848 16149 9857
rect 16107 9808 16108 9848
rect 16148 9808 16149 9848
rect 16107 9799 16149 9808
rect 16108 6236 16148 9799
rect 16204 9176 16244 15016
rect 16299 14384 16341 14393
rect 16299 14344 16300 14384
rect 16340 14344 16341 14384
rect 16299 14335 16341 14344
rect 16300 14250 16340 14335
rect 16300 13124 16340 13133
rect 16300 10604 16340 13084
rect 16396 12788 16436 15259
rect 16491 15140 16533 15149
rect 16491 15100 16492 15140
rect 16532 15100 16533 15140
rect 16491 15091 16533 15100
rect 16396 12739 16436 12748
rect 16395 12620 16437 12629
rect 16395 12580 16396 12620
rect 16436 12580 16437 12620
rect 16395 12571 16437 12580
rect 16300 10555 16340 10564
rect 16396 9344 16436 12571
rect 16396 9295 16436 9304
rect 16204 9127 16244 9136
rect 16108 6187 16148 6196
rect 16204 8336 16244 8345
rect 16204 2708 16244 8296
rect 16204 2659 16244 2668
rect 16300 7664 16340 7673
rect 16300 1196 16340 7624
rect 16492 7589 16532 15091
rect 16588 14888 16628 14897
rect 16588 12629 16628 14848
rect 16684 13292 16724 19132
rect 16684 13243 16724 13252
rect 16780 22700 16820 22709
rect 16587 12620 16629 12629
rect 16587 12580 16588 12620
rect 16628 12580 16629 12620
rect 16587 12571 16629 12580
rect 16684 11864 16724 11873
rect 16491 7580 16533 7589
rect 16491 7540 16492 7580
rect 16532 7540 16533 7580
rect 16491 7531 16533 7540
rect 16396 6824 16436 6833
rect 16396 3632 16436 6784
rect 16684 6740 16724 11824
rect 16588 6656 16628 6665
rect 16396 3583 16436 3592
rect 16492 6572 16532 6581
rect 16492 5144 16532 6532
rect 16588 6320 16628 6616
rect 16588 6271 16628 6280
rect 16492 3473 16532 5104
rect 16684 4304 16724 6700
rect 16684 4255 16724 4264
rect 16491 3464 16533 3473
rect 16491 3424 16492 3464
rect 16532 3424 16533 3464
rect 16491 3415 16533 3424
rect 16780 2456 16820 22660
rect 16972 22541 17012 37351
rect 17068 36812 17108 36821
rect 17068 36056 17108 36772
rect 17068 36007 17108 36016
rect 17164 35384 17204 35393
rect 17068 32612 17108 32623
rect 17068 32537 17108 32572
rect 17067 32528 17109 32537
rect 17067 32488 17068 32528
rect 17108 32488 17109 32528
rect 17067 32479 17109 32488
rect 17068 31436 17108 32479
rect 17068 31387 17108 31396
rect 16971 22532 17013 22541
rect 16971 22492 16972 22532
rect 17012 22492 17013 22532
rect 16971 22483 17013 22492
rect 16876 19004 16916 19013
rect 16876 17660 16916 18964
rect 17164 18920 17204 35344
rect 17260 28496 17300 38116
rect 17548 37988 17588 37997
rect 17452 37148 17492 37157
rect 17260 28447 17300 28456
rect 17356 36392 17396 36401
rect 17260 27320 17300 27329
rect 17260 24800 17300 27280
rect 17260 24751 17300 24760
rect 17356 22877 17396 36352
rect 17452 34637 17492 37108
rect 17451 34628 17493 34637
rect 17451 34588 17452 34628
rect 17492 34588 17493 34628
rect 17451 34579 17493 34588
rect 17452 34376 17492 34385
rect 17452 33041 17492 34336
rect 17451 33032 17493 33041
rect 17451 32992 17452 33032
rect 17492 32992 17493 33032
rect 17451 32983 17493 32992
rect 17452 26816 17492 32983
rect 17548 29168 17588 37948
rect 17643 36476 17685 36485
rect 17643 36436 17644 36476
rect 17684 36436 17685 36476
rect 17643 36427 17685 36436
rect 17644 35384 17684 36427
rect 17644 35335 17684 35344
rect 17740 35048 17780 40720
rect 17836 39668 17876 39677
rect 17836 37904 17876 39628
rect 17836 37855 17876 37864
rect 17836 37652 17876 37661
rect 17836 36140 17876 37612
rect 17932 36896 17972 41896
rect 17932 36847 17972 36856
rect 17836 36091 17876 36100
rect 17740 34999 17780 35008
rect 17836 35132 17876 35141
rect 17548 29119 17588 29128
rect 17644 34544 17684 34553
rect 17452 26767 17492 26776
rect 17452 25808 17492 25817
rect 17355 22868 17397 22877
rect 17355 22828 17356 22868
rect 17396 22828 17397 22868
rect 17355 22819 17397 22828
rect 17452 21104 17492 25768
rect 17644 25808 17684 34504
rect 17740 33284 17780 33293
rect 17740 31184 17780 33244
rect 17740 31135 17780 31144
rect 17740 30764 17780 30773
rect 17740 28916 17780 30724
rect 17740 28867 17780 28876
rect 17644 25759 17684 25768
rect 17740 26564 17780 26573
rect 17548 25640 17588 25649
rect 17548 22112 17588 25600
rect 17548 22063 17588 22072
rect 17452 21055 17492 21064
rect 17644 21272 17684 21281
rect 17164 18584 17204 18880
rect 17164 18535 17204 18544
rect 17548 20180 17588 20189
rect 17259 18500 17301 18509
rect 17259 18460 17260 18500
rect 17300 18460 17301 18500
rect 17259 18451 17301 18460
rect 17163 18416 17205 18425
rect 17163 18376 17164 18416
rect 17204 18376 17205 18416
rect 17163 18367 17205 18376
rect 16876 4061 16916 17620
rect 16972 16988 17012 16997
rect 16972 15905 17012 16948
rect 17067 16400 17109 16409
rect 17067 16360 17068 16400
rect 17108 16360 17109 16400
rect 17067 16351 17109 16360
rect 16971 15896 17013 15905
rect 16971 15856 16972 15896
rect 17012 15856 17013 15896
rect 16971 15847 17013 15856
rect 16972 13628 17012 15847
rect 17068 13796 17108 16351
rect 17164 14468 17204 18367
rect 17164 14419 17204 14428
rect 17163 14300 17205 14309
rect 17163 14260 17164 14300
rect 17204 14260 17205 14300
rect 17163 14251 17205 14260
rect 17164 14132 17204 14251
rect 17164 14083 17204 14092
rect 17068 13747 17108 13756
rect 16972 13588 17108 13628
rect 16972 12200 17012 12209
rect 16875 4052 16917 4061
rect 16875 4012 16876 4052
rect 16916 4012 16917 4052
rect 16875 4003 16917 4012
rect 16780 1952 16820 2416
rect 16780 1903 16820 1912
rect 16972 1280 17012 12160
rect 17068 11873 17108 13588
rect 17164 12956 17204 12965
rect 17067 11864 17109 11873
rect 17067 11824 17068 11864
rect 17108 11824 17109 11864
rect 17067 11815 17109 11824
rect 17164 10436 17204 12916
rect 17068 9008 17108 9017
rect 17068 5396 17108 8968
rect 17068 5347 17108 5356
rect 17067 4388 17109 4397
rect 17067 4348 17068 4388
rect 17108 4348 17109 4388
rect 17067 4339 17109 4348
rect 17068 4220 17108 4339
rect 17068 2624 17108 4180
rect 17164 3716 17204 10396
rect 17260 8000 17300 18451
rect 17452 17240 17492 17249
rect 17356 15812 17396 15821
rect 17356 12032 17396 15772
rect 17452 14897 17492 17200
rect 17451 14888 17493 14897
rect 17451 14848 17452 14888
rect 17492 14848 17493 14888
rect 17451 14839 17493 14848
rect 17451 14720 17493 14729
rect 17451 14680 17452 14720
rect 17492 14680 17493 14720
rect 17451 14671 17493 14680
rect 17356 11983 17396 11992
rect 17355 11864 17397 11873
rect 17355 11824 17356 11864
rect 17396 11824 17397 11864
rect 17355 11815 17397 11824
rect 17260 7951 17300 7960
rect 17164 3667 17204 3676
rect 17260 3632 17300 3641
rect 17163 3464 17205 3473
rect 17163 3424 17164 3464
rect 17204 3424 17205 3464
rect 17163 3415 17205 3424
rect 17068 2575 17108 2584
rect 16972 1231 17012 1240
rect 17164 1280 17204 3415
rect 17260 2876 17300 3592
rect 17260 2827 17300 2836
rect 17356 2540 17396 11815
rect 17452 11444 17492 14671
rect 17548 12872 17588 20140
rect 17644 17828 17684 21232
rect 17644 17779 17684 17788
rect 17644 16568 17684 16577
rect 17644 13964 17684 16528
rect 17644 13915 17684 13924
rect 17548 12823 17588 12832
rect 17452 11395 17492 11404
rect 17740 11360 17780 26524
rect 17836 22709 17876 35092
rect 17932 33704 17972 33713
rect 17932 31193 17972 33664
rect 17931 31184 17973 31193
rect 17931 31144 17932 31184
rect 17972 31144 17973 31184
rect 17931 31135 17973 31144
rect 17932 31016 17972 31025
rect 17835 22700 17877 22709
rect 17835 22660 17836 22700
rect 17876 22660 17877 22700
rect 17835 22651 17877 22660
rect 17644 11320 17780 11360
rect 17836 12620 17876 12629
rect 17548 8840 17588 8849
rect 17452 8672 17492 8681
rect 17452 3212 17492 8632
rect 17548 8597 17588 8800
rect 17547 8588 17589 8597
rect 17547 8548 17548 8588
rect 17588 8548 17589 8588
rect 17547 8539 17589 8548
rect 17548 4724 17588 4733
rect 17548 4061 17588 4684
rect 17547 4052 17589 4061
rect 17547 4012 17548 4052
rect 17588 4012 17589 4052
rect 17547 4003 17589 4012
rect 17452 3163 17492 3172
rect 17548 2624 17588 2633
rect 17548 2540 17588 2584
rect 17356 2500 17588 2540
rect 17164 1231 17204 1240
rect 16300 1147 16340 1156
rect 16012 727 16052 736
rect 15724 559 15764 568
rect 12172 307 12212 316
rect 15627 272 15669 281
rect 15627 232 15628 272
rect 15668 232 15669 272
rect 15627 223 15669 232
rect 15628 138 15668 223
rect 5067 104 5109 113
rect 5067 64 5068 104
rect 5108 64 5109 104
rect 5067 55 5109 64
rect 11691 104 11733 113
rect 11691 64 11692 104
rect 11732 64 11733 104
rect 11691 55 11733 64
rect 11883 104 11925 113
rect 11883 64 11884 104
rect 11924 64 11925 104
rect 11883 55 11925 64
rect 17548 104 17588 2500
rect 17644 944 17684 11320
rect 17740 4556 17780 4565
rect 17740 2372 17780 4516
rect 17836 4388 17876 12580
rect 17836 4339 17876 4348
rect 17740 2323 17780 2332
rect 17739 1868 17781 1877
rect 17739 1828 17740 1868
rect 17780 1828 17781 1868
rect 17739 1819 17781 1828
rect 17740 1734 17780 1819
rect 17932 1280 17972 30976
rect 18028 27581 18068 42568
rect 18220 41852 18260 41861
rect 18124 40592 18164 40601
rect 18027 27572 18069 27581
rect 18027 27532 18028 27572
rect 18068 27532 18069 27572
rect 18027 27523 18069 27532
rect 18028 25472 18068 25481
rect 18028 24632 18068 25432
rect 18028 24583 18068 24592
rect 18124 11360 18164 40552
rect 18220 32276 18260 41812
rect 18316 41609 18356 42652
rect 19467 41684 19509 41693
rect 19467 41644 19468 41684
rect 19508 41644 19509 41684
rect 19467 41635 19509 41644
rect 18315 41600 18357 41609
rect 18315 41560 18316 41600
rect 18356 41560 18357 41600
rect 18315 41551 18357 41560
rect 19468 41550 19508 41635
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 18315 41348 18357 41357
rect 18315 41308 18316 41348
rect 18356 41308 18357 41348
rect 18315 41299 18357 41308
rect 18316 41214 18356 41299
rect 19660 41180 19700 41189
rect 19084 41021 19124 41106
rect 18220 32227 18260 32236
rect 18316 41012 18356 41021
rect 18219 31184 18261 31193
rect 18219 31144 18220 31184
rect 18260 31144 18261 31184
rect 18219 31135 18261 31144
rect 18220 29420 18260 31135
rect 18220 28748 18260 29380
rect 18220 28699 18260 28708
rect 18028 11320 18164 11360
rect 18220 28076 18260 28085
rect 18028 9092 18068 11320
rect 18123 11192 18165 11201
rect 18123 11152 18124 11192
rect 18164 11152 18165 11192
rect 18123 11143 18165 11152
rect 18124 11058 18164 11143
rect 18028 9043 18068 9052
rect 18124 9176 18164 9185
rect 18124 8588 18164 9136
rect 18124 8539 18164 8548
rect 18124 8168 18164 8177
rect 18124 7664 18164 8128
rect 18124 7615 18164 7624
rect 17932 1231 17972 1240
rect 17644 895 17684 904
rect 18220 944 18260 28036
rect 18316 13880 18356 40972
rect 19083 41012 19125 41021
rect 19083 40972 19084 41012
rect 19124 40972 19125 41012
rect 19083 40963 19125 40972
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 19276 40592 19316 40601
rect 18412 40340 18452 40349
rect 18412 39593 18452 40300
rect 18604 40340 18644 40349
rect 18508 40256 18548 40265
rect 18411 39584 18453 39593
rect 18411 39544 18412 39584
rect 18452 39544 18453 39584
rect 18411 39535 18453 39544
rect 18412 38744 18452 38753
rect 18412 38501 18452 38704
rect 18411 38492 18453 38501
rect 18411 38452 18412 38492
rect 18452 38452 18453 38492
rect 18411 38443 18453 38452
rect 18508 38492 18548 40216
rect 18604 38921 18644 40300
rect 18699 39920 18741 39929
rect 18699 39880 18700 39920
rect 18740 39880 18741 39920
rect 18699 39871 18741 39880
rect 18700 39786 18740 39871
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19276 39005 19316 40552
rect 19372 39836 19412 39845
rect 19275 38996 19317 39005
rect 19275 38956 19276 38996
rect 19316 38956 19317 38996
rect 19275 38947 19317 38956
rect 18603 38912 18645 38921
rect 18603 38872 18604 38912
rect 18644 38872 18645 38912
rect 18603 38863 18645 38872
rect 18700 38660 18740 38669
rect 18508 38443 18548 38452
rect 18604 38576 18644 38585
rect 18316 13831 18356 13840
rect 18412 37568 18452 37577
rect 18412 12620 18452 37528
rect 18604 37148 18644 38536
rect 18700 38072 18740 38620
rect 18700 38023 18740 38032
rect 19276 38324 19316 38333
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 19276 37400 19316 38284
rect 19372 37568 19412 39796
rect 19372 37519 19412 37528
rect 19564 38996 19604 39005
rect 19276 37360 19412 37400
rect 18508 37108 18644 37148
rect 19276 37232 19316 37241
rect 18508 36056 18548 37108
rect 18508 36007 18548 36016
rect 18604 36980 18644 36989
rect 18508 33116 18548 33125
rect 18508 31436 18548 33076
rect 18508 31277 18548 31396
rect 18507 31268 18549 31277
rect 18507 31228 18508 31268
rect 18548 31228 18549 31268
rect 18507 31219 18549 31228
rect 18604 28664 18644 36940
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 18795 35972 18837 35981
rect 18795 35932 18796 35972
rect 18836 35932 18837 35972
rect 18795 35923 18837 35932
rect 18796 35300 18836 35923
rect 18796 35251 18836 35260
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 19276 34385 19316 37192
rect 19372 36224 19412 37360
rect 19467 36644 19509 36653
rect 19467 36604 19468 36644
rect 19508 36604 19509 36644
rect 19467 36595 19509 36604
rect 19468 36510 19508 36595
rect 19372 36175 19412 36184
rect 19275 34376 19317 34385
rect 19275 34336 19276 34376
rect 19316 34336 19317 34376
rect 19275 34327 19317 34336
rect 19564 33788 19604 38956
rect 19564 33739 19604 33748
rect 19467 33620 19509 33629
rect 19467 33580 19468 33620
rect 19508 33580 19509 33620
rect 19467 33571 19509 33580
rect 19468 33486 19508 33571
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 19660 33116 19700 41140
rect 19468 33076 19660 33116
rect 18700 32276 18740 32285
rect 18700 31604 18740 32236
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18700 31555 18740 31564
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 19372 29084 19412 29093
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18604 28615 18644 28624
rect 19276 28664 19316 28673
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18700 24968 18740 24977
rect 18700 23708 18740 24928
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 19276 24044 19316 28624
rect 19372 27236 19412 29044
rect 19372 27187 19412 27196
rect 19372 27068 19412 27077
rect 19372 25304 19412 27028
rect 19468 26564 19508 33076
rect 19660 33067 19700 33076
rect 19852 41180 19892 41189
rect 19852 33536 19892 41140
rect 20139 41096 20181 41105
rect 20139 41056 20140 41096
rect 20180 41056 20181 41096
rect 20139 41047 20181 41056
rect 20140 40962 20180 41047
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 19948 39668 19988 39677
rect 19948 36056 19988 39628
rect 20139 39080 20181 39089
rect 20139 39040 20140 39080
rect 20180 39040 20181 39080
rect 20139 39031 20181 39040
rect 20140 38946 20180 39031
rect 20524 38744 20564 38753
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 20139 38408 20181 38417
rect 20139 38368 20140 38408
rect 20180 38368 20181 38408
rect 20139 38359 20181 38368
rect 20140 38274 20180 38359
rect 20139 38072 20181 38081
rect 20139 38032 20140 38072
rect 20180 38032 20181 38072
rect 20139 38023 20181 38032
rect 20140 37938 20180 38023
rect 20140 37736 20180 37745
rect 20044 37696 20140 37736
rect 20044 37484 20084 37696
rect 20140 37687 20180 37696
rect 20044 37435 20084 37444
rect 20331 37400 20373 37409
rect 20331 37360 20332 37400
rect 20372 37360 20373 37400
rect 20331 37351 20373 37360
rect 20332 37266 20372 37351
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 19948 36007 19988 36016
rect 20140 36560 20180 36569
rect 20140 36056 20180 36520
rect 20140 36007 20180 36016
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 20139 34712 20181 34721
rect 20139 34672 20140 34712
rect 20180 34672 20181 34712
rect 20139 34663 20181 34672
rect 20140 34578 20180 34663
rect 19468 26515 19508 26524
rect 19564 31184 19604 31193
rect 19372 25255 19412 25264
rect 19276 23995 19316 24004
rect 18700 20180 18740 23668
rect 19468 22784 19508 22793
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 19372 22700 19412 22709
rect 19372 21356 19412 22660
rect 19372 21307 19412 21316
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 19468 20273 19508 22744
rect 19467 20264 19509 20273
rect 19467 20224 19468 20264
rect 19508 20224 19509 20264
rect 19467 20215 19509 20224
rect 18700 19088 18740 20140
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 18700 19039 18740 19048
rect 19468 19172 19508 19181
rect 18412 12571 18452 12580
rect 18508 18584 18548 18593
rect 18508 11360 18548 18544
rect 19468 18584 19508 19132
rect 19468 18535 19508 18544
rect 19372 18332 19412 18341
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 19372 15737 19412 18292
rect 19564 17912 19604 31144
rect 19660 31100 19700 31109
rect 19660 22280 19700 31060
rect 19852 31016 19892 33496
rect 19852 30967 19892 30976
rect 19948 34544 19988 34553
rect 19852 29840 19892 29849
rect 19755 26648 19797 26657
rect 19755 26608 19756 26648
rect 19796 26608 19797 26648
rect 19755 26599 19797 26608
rect 19756 23456 19796 26599
rect 19852 26480 19892 29800
rect 19948 26657 19988 34504
rect 20524 34376 20564 38704
rect 20811 38744 20853 38753
rect 20811 38704 20812 38744
rect 20852 38704 20853 38744
rect 20811 38695 20853 38704
rect 20812 38610 20852 38695
rect 20620 37064 20660 37073
rect 20620 35897 20660 37024
rect 20619 35888 20661 35897
rect 20619 35848 20620 35888
rect 20660 35848 20661 35888
rect 20619 35839 20661 35848
rect 20524 34327 20564 34336
rect 20716 35720 20756 35729
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 20139 31688 20181 31697
rect 20139 31648 20140 31688
rect 20180 31648 20181 31688
rect 20139 31639 20181 31648
rect 20140 31554 20180 31639
rect 20716 31352 20756 35680
rect 20908 35720 20948 35729
rect 20908 32780 20948 35680
rect 20716 31303 20756 31312
rect 20812 32740 20948 32780
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 20524 28916 20564 28925
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 20524 27404 20564 28876
rect 20812 28580 20852 32740
rect 20908 31520 20948 31529
rect 20908 29000 20948 31480
rect 20908 28960 21044 29000
rect 20812 28531 20852 28540
rect 20524 27355 20564 27364
rect 20812 26816 20852 26825
rect 19947 26648 19989 26657
rect 19947 26608 19948 26648
rect 19988 26608 19989 26648
rect 19947 26599 19989 26608
rect 20048 26480 20416 26489
rect 19852 26440 19988 26480
rect 19852 24800 19892 24809
rect 19852 23624 19892 24760
rect 19852 23575 19892 23584
rect 19756 23416 19892 23456
rect 19660 22231 19700 22240
rect 19756 20600 19796 20609
rect 19660 20012 19700 20021
rect 19660 18080 19700 19972
rect 19660 18031 19700 18040
rect 19564 17863 19604 17872
rect 19756 17828 19796 20560
rect 19852 20516 19892 23416
rect 19948 23288 19988 26440
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20812 24968 20852 26776
rect 20908 26564 20948 26573
rect 20908 25640 20948 26524
rect 20908 25591 20948 25600
rect 20812 24919 20852 24928
rect 20908 24044 20948 24053
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 19948 23239 19988 23248
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20620 21608 20660 21617
rect 19852 20467 19892 20476
rect 19948 20936 19988 20945
rect 19851 20264 19893 20273
rect 19851 20224 19852 20264
rect 19892 20224 19893 20264
rect 19851 20215 19893 20224
rect 19756 17779 19796 17788
rect 19852 17660 19892 20215
rect 19948 17996 19988 20896
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 20524 19256 20564 19265
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 19948 17947 19988 17956
rect 19852 17611 19892 17620
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 19564 16400 19604 16409
rect 19371 15728 19413 15737
rect 19371 15688 19372 15728
rect 19412 15688 19413 15728
rect 19371 15679 19413 15688
rect 19372 15560 19412 15569
rect 19276 15392 19316 15401
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 18700 13880 18740 13889
rect 18316 11320 18548 11360
rect 18604 13796 18644 13805
rect 18316 3389 18356 11320
rect 18508 9932 18548 9941
rect 18412 8084 18452 8093
rect 18412 4808 18452 8044
rect 18315 3380 18357 3389
rect 18315 3340 18316 3380
rect 18356 3340 18357 3380
rect 18315 3331 18357 3340
rect 18412 2456 18452 4768
rect 18412 2407 18452 2416
rect 18508 1280 18548 9892
rect 18604 3296 18644 13756
rect 18700 13376 18740 13840
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18700 13327 18740 13336
rect 19276 13376 19316 15352
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18700 9428 18740 9437
rect 18700 8840 18740 9388
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18796 8840 18836 8849
rect 18700 8800 18796 8840
rect 18796 8791 18836 8800
rect 18700 8504 18740 8513
rect 18700 7664 18740 8464
rect 18700 7615 18740 7624
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 18604 3247 18644 3256
rect 18700 7412 18740 7421
rect 18700 2540 18740 7372
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18892 5816 18932 5825
rect 18892 5312 18932 5776
rect 19276 5816 19316 13336
rect 19372 13040 19412 15520
rect 19564 15392 19604 16360
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 19755 15728 19797 15737
rect 19755 15688 19756 15728
rect 19796 15688 19797 15728
rect 19755 15679 19797 15688
rect 19564 15343 19604 15352
rect 19660 15644 19700 15653
rect 19372 12991 19412 13000
rect 19468 14636 19508 14645
rect 19468 12872 19508 14596
rect 19468 12823 19508 12832
rect 19564 13460 19604 13469
rect 19468 10352 19508 10361
rect 19468 10184 19508 10312
rect 19468 7160 19508 10144
rect 19564 9932 19604 13420
rect 19564 9883 19604 9892
rect 19468 6329 19508 7120
rect 19564 8084 19604 8093
rect 19467 6320 19509 6329
rect 19467 6280 19468 6320
rect 19508 6280 19509 6320
rect 19467 6271 19509 6280
rect 19564 6320 19604 8044
rect 19564 6271 19604 6280
rect 19276 5767 19316 5776
rect 18892 5263 18932 5272
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 19564 3884 19604 3893
rect 19564 3296 19604 3844
rect 19660 3557 19700 15604
rect 19756 15560 19796 15679
rect 20524 15644 20564 19216
rect 20620 18416 20660 21568
rect 20620 18367 20660 18376
rect 20524 15595 20564 15604
rect 20620 17576 20660 17585
rect 19756 15511 19796 15520
rect 19852 15056 19892 15065
rect 19756 14720 19796 14729
rect 19756 12452 19796 14680
rect 19852 13880 19892 15016
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 19852 13831 19892 13840
rect 20524 13208 20564 13217
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 19756 8177 19796 12412
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 19948 8504 19988 8513
rect 19755 8168 19797 8177
rect 19755 8128 19756 8168
rect 19796 8128 19797 8168
rect 19755 8119 19797 8128
rect 19948 8168 19988 8464
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19948 8119 19988 8128
rect 19659 3548 19701 3557
rect 19659 3508 19660 3548
rect 19700 3508 19701 3548
rect 19659 3499 19701 3508
rect 19564 3247 19604 3256
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18604 2500 18740 2540
rect 18604 1784 18644 2500
rect 18604 1735 18644 1744
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18508 1231 18548 1240
rect 18699 1280 18741 1289
rect 18699 1240 18700 1280
rect 18740 1240 18741 1280
rect 18699 1231 18741 1240
rect 18700 1146 18740 1231
rect 18220 895 18260 904
rect 18891 440 18933 449
rect 18891 400 18892 440
rect 18932 400 18933 440
rect 18891 391 18933 400
rect 19660 440 19700 3499
rect 19756 3128 19796 8119
rect 20524 7001 20564 13168
rect 20620 12620 20660 17536
rect 20620 12571 20660 12580
rect 20716 15896 20756 15905
rect 20620 10520 20660 10529
rect 20523 6992 20565 7001
rect 20523 6952 20524 6992
rect 20564 6952 20565 6992
rect 20523 6943 20565 6952
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 20043 4808 20085 4817
rect 20043 4768 20044 4808
rect 20084 4768 20085 4808
rect 20043 4759 20085 4768
rect 20044 4472 20084 4759
rect 20140 4472 20180 4481
rect 20044 4432 20140 4472
rect 20140 4404 20180 4432
rect 19948 4136 19988 4145
rect 19948 3296 19988 4096
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20524 3464 20564 6943
rect 20620 6488 20660 10480
rect 20716 10184 20756 15856
rect 20716 10135 20756 10144
rect 20812 14888 20852 14897
rect 20812 8924 20852 14848
rect 20908 14300 20948 24004
rect 21004 19592 21044 28960
rect 21100 28244 21140 42736
rect 21292 42104 21332 42113
rect 21196 37652 21236 37661
rect 21196 32696 21236 37612
rect 21196 32647 21236 32656
rect 21100 28195 21140 28204
rect 21196 31436 21236 31445
rect 21004 19543 21044 19552
rect 20908 14251 20948 14260
rect 21004 18668 21044 18677
rect 20812 8875 20852 8884
rect 21004 7496 21044 18628
rect 21196 18248 21236 31396
rect 21292 27320 21332 42064
rect 21292 27271 21332 27280
rect 21388 33872 21428 33881
rect 21196 18199 21236 18208
rect 21292 21272 21332 21281
rect 21004 7447 21044 7456
rect 21100 14552 21140 14561
rect 20620 6439 20660 6448
rect 20811 4724 20853 4733
rect 20811 4684 20812 4724
rect 20852 4684 20853 4724
rect 20811 4675 20853 4684
rect 20524 3415 20564 3424
rect 20812 3464 20852 4675
rect 21100 4220 21140 14512
rect 21292 4892 21332 21232
rect 21388 8840 21428 33832
rect 21388 8791 21428 8800
rect 21292 4843 21332 4852
rect 21100 4171 21140 4180
rect 20812 3415 20852 3424
rect 20619 3380 20661 3389
rect 20619 3340 20620 3380
rect 20660 3340 20661 3380
rect 20619 3331 20661 3340
rect 19948 3247 19988 3256
rect 19756 3079 19796 3088
rect 20140 2549 20180 2634
rect 20139 2540 20181 2549
rect 20139 2500 20140 2540
rect 20180 2500 20181 2540
rect 20139 2491 20181 2500
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 20620 2120 20660 3331
rect 20620 2071 20660 2080
rect 20523 1952 20565 1961
rect 20523 1912 20524 1952
rect 20564 1912 20565 1952
rect 20523 1903 20565 1912
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 20524 776 20564 1903
rect 20715 1784 20757 1793
rect 20715 1744 20716 1784
rect 20756 1744 20757 1784
rect 20715 1735 20757 1744
rect 20716 1650 20756 1735
rect 20524 727 20564 736
rect 19660 391 19700 400
rect 18892 306 18932 391
rect 18124 113 18164 198
rect 17548 55 17588 64
rect 18123 104 18165 113
rect 18123 64 18124 104
rect 18164 64 18165 104
rect 18123 55 18165 64
<< via4 >>
rect 76 25852 116 25892
rect 268 18460 308 18500
rect 556 35848 596 35888
rect 556 17872 596 17912
rect 1036 23248 1076 23288
rect 6796 42232 6836 42272
rect 1324 34504 1364 34544
rect 1228 29968 1268 30008
rect 1516 30724 1556 30764
rect 1228 25852 1268 25892
rect 1228 22408 1268 22448
rect 1228 19888 1268 19928
rect 1228 18376 1268 18416
rect 1420 17536 1460 17576
rect 940 16360 980 16400
rect 844 15772 884 15812
rect 1228 16864 1268 16904
rect 1132 11908 1172 11948
rect 1516 14848 1556 14888
rect 1228 9976 1268 10016
rect 1420 9472 1460 9512
rect 1228 8548 1268 8588
rect 1420 3592 1460 3632
rect 1708 31732 1748 31772
rect 1996 38032 2036 38072
rect 1996 36772 2036 36812
rect 1900 31732 1940 31772
rect 1900 21736 1940 21776
rect 1708 18544 1748 18584
rect 1804 17704 1844 17744
rect 2188 36604 2228 36644
rect 2188 35680 2228 35720
rect 2380 36772 2420 36812
rect 2380 36604 2420 36644
rect 2764 32992 2804 33032
rect 3052 36688 3092 36728
rect 2956 34840 2996 34880
rect 2956 29968 2996 30008
rect 2668 29380 2708 29420
rect 2860 29296 2900 29336
rect 2284 28792 2324 28832
rect 2284 26692 2324 26732
rect 2572 28960 2612 29000
rect 1900 9724 1940 9764
rect 2188 18544 2228 18584
rect 2860 28876 2900 28916
rect 2764 28792 2804 28832
rect 2668 22324 2708 22364
rect 2284 12916 2324 12956
rect 2476 12832 2516 12872
rect 2284 9724 2324 9764
rect 2188 8632 2228 8672
rect 2188 3172 2228 3212
rect 2668 2668 2708 2708
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 3532 38368 3572 38408
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3820 37192 3860 37232
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 3532 35932 3572 35972
rect 3628 35176 3668 35216
rect 3436 34840 3476 34880
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 3244 29212 3284 29252
rect 3340 29128 3380 29168
rect 3148 27700 3188 27740
rect 2956 18292 2996 18332
rect 3148 9640 3188 9680
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 5356 39460 5396 39500
rect 4588 38704 4628 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 4492 36436 4532 36476
rect 3628 28204 3668 28244
rect 4108 27616 4148 27656
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 4300 29128 4340 29168
rect 4300 26608 4340 26648
rect 4108 22492 4148 22532
rect 4108 22240 4148 22280
rect 3436 10312 3476 10352
rect 1516 1156 1556 1196
rect 3724 21736 3764 21776
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3628 15268 3668 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3724 14764 3764 14804
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 4492 34420 4532 34460
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 5260 34924 5300 34964
rect 4684 34588 4724 34628
rect 4876 34420 4916 34460
rect 4780 34168 4820 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4492 27700 4532 27740
rect 4396 24508 4436 24548
rect 4300 22912 4340 22952
rect 4300 22240 4340 22280
rect 4588 23584 4628 23624
rect 4588 22996 4628 23036
rect 4588 22492 4628 22532
rect 4300 19048 4340 19088
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 5068 25264 5108 25304
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4780 24508 4820 24548
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3820 10312 3860 10352
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3820 6952 3860 6992
rect 4108 6448 4148 6488
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4300 7120 4340 7160
rect 4204 4348 4244 4388
rect 4108 4096 4148 4136
rect 4300 3928 4340 3968
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 5644 35260 5684 35300
rect 5548 30724 5588 30764
rect 5452 27532 5492 27572
rect 5452 24676 5492 24716
rect 5452 21736 5492 21776
rect 5836 40300 5876 40340
rect 5644 25852 5684 25892
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4780 18292 4820 18332
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4780 8548 4820 8588
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4780 7120 4820 7160
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4684 6196 4724 6236
rect 4588 4600 4628 4640
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4300 1408 4340 1448
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 4780 4180 4820 4220
rect 4972 4684 5012 4724
rect 4876 4096 4916 4136
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 6220 37864 6260 37904
rect 5932 34924 5972 34964
rect 5932 22324 5972 22364
rect 5260 1156 5300 1196
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5740 10732 5780 10772
rect 5644 2584 5684 2624
rect 5548 1996 5588 2036
rect 6124 35176 6164 35216
rect 6316 35008 6356 35048
rect 6124 26692 6164 26732
rect 6220 25096 6260 25136
rect 6508 34252 6548 34292
rect 6220 22828 6260 22868
rect 6316 21988 6356 22028
rect 6700 38200 6740 38240
rect 7084 39628 7124 39668
rect 6892 34420 6932 34460
rect 6700 32908 6740 32948
rect 6796 27532 6836 27572
rect 6700 26692 6740 26732
rect 6700 22912 6740 22952
rect 6700 21988 6740 22028
rect 6508 17788 6548 17828
rect 6316 15688 6356 15728
rect 6412 12580 6452 12620
rect 6316 3592 6356 3632
rect 6508 1912 6548 1952
rect 6700 4516 6740 4556
rect 6892 25096 6932 25136
rect 6892 1828 6932 1868
rect 7276 36688 7316 36728
rect 7468 40972 7508 41012
rect 7564 35680 7604 35720
rect 7564 34420 7604 34460
rect 7468 28372 7508 28412
rect 7372 24004 7412 24044
rect 7276 15688 7316 15728
rect 7372 12412 7412 12452
rect 7180 4768 7220 4808
rect 7564 15772 7604 15812
rect 7564 15184 7604 15224
rect 7660 11992 7700 12032
rect 7564 9640 7604 9680
rect 7564 6448 7604 6488
rect 7660 6280 7700 6320
rect 7372 5188 7412 5228
rect 7276 4684 7316 4724
rect 7276 4516 7316 4556
rect 7180 4180 7220 4220
rect 7180 1240 7220 1280
rect 7564 2668 7604 2708
rect 8428 34420 8468 34460
rect 8044 34336 8084 34376
rect 8044 32908 8084 32948
rect 7948 25852 7988 25892
rect 8140 28624 8180 28664
rect 8332 29128 8372 29168
rect 8140 17536 8180 17576
rect 7852 12580 7892 12620
rect 8044 11404 8084 11444
rect 8908 35260 8948 35300
rect 9100 37192 9140 37232
rect 9100 31900 9140 31940
rect 8620 29548 8660 29588
rect 8620 29212 8660 29252
rect 8524 28624 8564 28664
rect 8716 29044 8756 29084
rect 8812 27532 8852 27572
rect 9004 26440 9044 26480
rect 8908 23668 8948 23708
rect 8620 15772 8660 15812
rect 8908 15604 8948 15644
rect 9004 4264 9044 4304
rect 9388 37444 9428 37484
rect 9388 35008 9428 35048
rect 9484 34588 9524 34628
rect 9388 27616 9428 27656
rect 9772 29044 9812 29084
rect 9292 11908 9332 11948
rect 9292 4600 9332 4640
rect 9676 18880 9716 18920
rect 9580 16276 9620 16316
rect 9580 9472 9620 9512
rect 9580 5020 9620 5060
rect 9964 41560 10004 41600
rect 10060 38704 10100 38744
rect 10060 25264 10100 25304
rect 9868 14764 9908 14804
rect 10732 38368 10772 38408
rect 10636 37864 10676 37904
rect 10636 36520 10676 36560
rect 10444 35008 10484 35048
rect 10732 34924 10772 34964
rect 10252 22996 10292 23036
rect 10156 13756 10196 13796
rect 10060 10648 10100 10688
rect 9964 8128 10004 8168
rect 9388 2416 9428 2456
rect 9676 3928 9716 3968
rect 9772 3340 9812 3380
rect 10348 13756 10388 13796
rect 10540 30304 10580 30344
rect 10540 27700 10580 27740
rect 10732 29128 10772 29168
rect 10636 27616 10676 27656
rect 10252 6196 10292 6236
rect 10156 3424 10196 3464
rect 10060 2584 10100 2624
rect 10540 10060 10580 10100
rect 11212 34168 11252 34208
rect 11116 30304 11156 30344
rect 11020 27616 11060 27656
rect 10924 27448 10964 27488
rect 11020 26776 11060 26816
rect 10828 15604 10868 15644
rect 10732 14008 10772 14048
rect 10540 8716 10580 8756
rect 11116 10480 11156 10520
rect 11116 10060 11156 10100
rect 11116 9808 11156 9848
rect 10828 1828 10868 1868
rect 11308 26524 11348 26564
rect 14764 41644 14804 41684
rect 11596 32824 11636 32864
rect 11500 22408 11540 22448
rect 12076 34588 12116 34628
rect 12844 41308 12884 41348
rect 12460 41056 12500 41096
rect 12556 39544 12596 39584
rect 12844 39628 12884 39668
rect 12748 38032 12788 38072
rect 11980 26776 12020 26816
rect 11692 17788 11732 17828
rect 11404 10648 11444 10688
rect 11308 10480 11348 10520
rect 7948 820 7988 860
rect 11596 4180 11636 4220
rect 11308 400 11348 440
rect 12556 36520 12596 36560
rect 12556 33580 12596 33620
rect 12268 27616 12308 27656
rect 12460 27616 12500 27656
rect 12460 27448 12500 27488
rect 11788 10816 11828 10856
rect 12076 11152 12116 11192
rect 12172 10816 12212 10856
rect 11980 10732 12020 10772
rect 11884 7792 11924 7832
rect 14668 39880 14708 39920
rect 13132 39460 13172 39500
rect 14572 39460 14612 39500
rect 12940 36940 12980 36980
rect 12844 33412 12884 33452
rect 12844 27700 12884 27740
rect 12844 26524 12884 26564
rect 12460 12412 12500 12452
rect 12844 16276 12884 16316
rect 12556 10396 12596 10436
rect 12748 10396 12788 10436
rect 12652 8716 12692 8756
rect 12364 8548 12404 8588
rect 12268 7624 12308 7664
rect 12076 4264 12116 4304
rect 12556 7540 12596 7580
rect 12556 3172 12596 3212
rect 12364 1072 12404 1112
rect 13036 34504 13076 34544
rect 13036 33412 13076 33452
rect 13036 16276 13076 16316
rect 13900 39208 13940 39248
rect 13612 38032 13652 38072
rect 13420 29128 13460 29168
rect 13420 15856 13460 15896
rect 13228 9976 13268 10016
rect 13420 9808 13460 9848
rect 13132 1996 13172 2036
rect 14188 38872 14228 38912
rect 14380 38452 14420 38492
rect 14188 35260 14228 35300
rect 13996 34420 14036 34460
rect 13804 33076 13844 33116
rect 13804 32908 13844 32948
rect 13900 32488 13940 32528
rect 13708 31228 13748 31268
rect 13612 22492 13652 22532
rect 14092 32992 14132 33032
rect 14284 32992 14324 33032
rect 13900 17704 13940 17744
rect 13804 15688 13844 15728
rect 13996 11404 14036 11444
rect 13900 10060 13940 10100
rect 13900 6448 13940 6488
rect 13804 5020 13844 5060
rect 14188 9472 14228 9512
rect 14092 6448 14132 6488
rect 13996 4768 14036 4808
rect 14476 34084 14516 34124
rect 14380 23248 14420 23288
rect 14380 1744 14420 1784
rect 15148 40384 15188 40424
rect 14860 38956 14900 38996
rect 14764 22660 14804 22700
rect 14764 18880 14804 18920
rect 14668 15184 14708 15224
rect 14572 7120 14612 7160
rect 14956 38872 14996 38912
rect 15244 39712 15284 39752
rect 15148 34168 15188 34208
rect 14956 34000 14996 34040
rect 14956 19888 14996 19928
rect 14956 17704 14996 17744
rect 15052 6448 15092 6488
rect 14956 3256 14996 3296
rect 15436 35176 15476 35216
rect 16396 42232 16436 42272
rect 16012 40888 16052 40928
rect 15628 34336 15668 34376
rect 15628 29548 15668 29588
rect 15436 16864 15476 16904
rect 15436 8716 15476 8756
rect 15340 8632 15380 8672
rect 14764 1240 14804 1280
rect 13132 820 13172 860
rect 13900 652 13940 692
rect 15628 24592 15668 24632
rect 17068 40972 17108 41012
rect 16972 40384 17012 40424
rect 16012 39292 16052 39332
rect 16204 39292 16244 39332
rect 15916 39040 15956 39080
rect 16012 38704 16052 38744
rect 15916 34000 15956 34040
rect 15820 24592 15860 24632
rect 16012 33076 16052 33116
rect 15916 16276 15956 16316
rect 15916 11992 15956 12032
rect 15628 3256 15668 3296
rect 15820 1912 15860 1952
rect 16396 39712 16436 39752
rect 16492 39460 16532 39500
rect 16396 39208 16436 39248
rect 16876 39124 16916 39164
rect 16684 38368 16724 38408
rect 16204 34084 16244 34124
rect 17548 40300 17588 40340
rect 17644 39292 17684 39332
rect 17452 39124 17492 39164
rect 16972 37360 17012 37400
rect 16684 23584 16724 23624
rect 16396 15268 16436 15308
rect 16108 14008 16148 14048
rect 16108 9808 16148 9848
rect 16300 14344 16340 14384
rect 16492 15100 16532 15140
rect 16396 12580 16436 12620
rect 16588 12580 16628 12620
rect 16492 7540 16532 7580
rect 16492 3424 16532 3464
rect 17068 32488 17108 32528
rect 16972 22492 17012 22532
rect 17452 34588 17492 34628
rect 17452 32992 17492 33032
rect 17644 36436 17684 36476
rect 17356 22828 17396 22868
rect 17260 18460 17300 18500
rect 17164 18376 17204 18416
rect 17068 16360 17108 16400
rect 16972 15856 17012 15896
rect 17164 14260 17204 14300
rect 16876 4012 16916 4052
rect 17068 11824 17108 11864
rect 17068 4348 17108 4388
rect 17452 14848 17492 14888
rect 17452 14680 17492 14720
rect 17356 11824 17396 11864
rect 17164 3424 17204 3464
rect 17932 31144 17972 31184
rect 17836 22660 17876 22700
rect 17548 8548 17588 8588
rect 17548 4012 17588 4052
rect 15628 232 15668 272
rect 5068 64 5108 104
rect 11692 64 11732 104
rect 11884 64 11924 104
rect 17740 1828 17780 1868
rect 18028 27532 18068 27572
rect 19468 41644 19508 41684
rect 18316 41560 18356 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 18316 41308 18356 41348
rect 18220 31144 18260 31184
rect 18124 11152 18164 11192
rect 19084 40972 19124 41012
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 18412 39544 18452 39584
rect 18412 38452 18452 38492
rect 18700 39880 18740 39920
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 19276 38956 19316 38996
rect 18604 38872 18644 38912
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18508 31228 18548 31268
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 18796 35932 18836 35972
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 19468 36604 19508 36644
rect 19276 34336 19316 34376
rect 19468 33580 19508 33620
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 20140 41056 20180 41096
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 20140 39040 20180 39080
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20140 38368 20180 38408
rect 20140 38032 20180 38072
rect 20332 37360 20372 37400
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20140 34672 20180 34712
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 19468 20224 19508 20264
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 19756 26608 19796 26648
rect 20812 38704 20852 38744
rect 20620 35848 20660 35888
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20140 31648 20180 31688
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 19948 26608 19988 26648
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 19852 20224 19892 20264
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 19372 15688 19412 15728
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18316 3340 18356 3380
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 19756 15688 19796 15728
rect 19468 6280 19508 6320
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19756 8128 19796 8168
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19660 3508 19700 3548
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 18700 1240 18740 1280
rect 18892 400 18932 440
rect 20524 6952 20564 6992
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 20044 4768 20084 4808
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20812 4684 20852 4724
rect 20620 3340 20660 3380
rect 20140 2500 20180 2540
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 20524 1912 20564 1952
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 20716 1744 20756 1784
rect 18124 64 18164 104
<< metal5 >>
rect 6787 42232 6796 42272
rect 6836 42232 16396 42272
rect 16436 42232 16445 42272
rect 14755 41644 14764 41684
rect 14804 41644 19468 41684
rect 19508 41644 19517 41684
rect 4919 41623 5305 41642
rect 4919 41600 4985 41623
rect 5071 41600 5153 41623
rect 5239 41600 5305 41623
rect 20039 41623 20425 41642
rect 20039 41600 20105 41623
rect 20191 41600 20273 41623
rect 20359 41600 20425 41623
rect 4919 41560 4928 41600
rect 4968 41560 4985 41600
rect 5071 41560 5092 41600
rect 5132 41560 5153 41600
rect 5239 41560 5256 41600
rect 5296 41560 5305 41600
rect 9955 41560 9964 41600
rect 10004 41560 18316 41600
rect 18356 41560 18365 41600
rect 20039 41560 20048 41600
rect 20088 41560 20105 41600
rect 20191 41560 20212 41600
rect 20252 41560 20273 41600
rect 20359 41560 20376 41600
rect 20416 41560 20425 41600
rect 4919 41537 4985 41560
rect 5071 41537 5153 41560
rect 5239 41537 5305 41560
rect 4919 41518 5305 41537
rect 20039 41537 20105 41560
rect 20191 41537 20273 41560
rect 20359 41537 20425 41560
rect 20039 41518 20425 41537
rect 12835 41308 12844 41348
rect 12884 41308 18316 41348
rect 18356 41308 18365 41348
rect 12451 41056 12460 41096
rect 12500 41056 20140 41096
rect 20180 41056 20189 41096
rect 7459 40972 7468 41012
rect 7508 40972 17068 41012
rect 17108 40972 17117 41012
rect 17180 40972 19084 41012
rect 19124 40972 19133 41012
rect 17180 40928 17220 40972
rect 16003 40888 16012 40928
rect 16052 40888 17220 40928
rect 3679 40867 4065 40886
rect 3679 40844 3745 40867
rect 3831 40844 3913 40867
rect 3999 40844 4065 40867
rect 3679 40804 3688 40844
rect 3728 40804 3745 40844
rect 3831 40804 3852 40844
rect 3892 40804 3913 40844
rect 3999 40804 4016 40844
rect 4056 40804 4065 40844
rect 3679 40781 3745 40804
rect 3831 40781 3913 40804
rect 3999 40781 4065 40804
rect 3679 40762 4065 40781
rect 18799 40867 19185 40886
rect 18799 40844 18865 40867
rect 18951 40844 19033 40867
rect 19119 40844 19185 40867
rect 18799 40804 18808 40844
rect 18848 40804 18865 40844
rect 18951 40804 18972 40844
rect 19012 40804 19033 40844
rect 19119 40804 19136 40844
rect 19176 40804 19185 40844
rect 18799 40781 18865 40804
rect 18951 40781 19033 40804
rect 19119 40781 19185 40804
rect 18799 40762 19185 40781
rect 15139 40384 15148 40424
rect 15188 40384 16972 40424
rect 17012 40384 17021 40424
rect 2090 40363 2214 40382
rect 2090 40277 2109 40363
rect 2195 40340 2214 40363
rect 17138 40363 17262 40382
rect 2195 40300 5836 40340
rect 5876 40300 5885 40340
rect 2195 40277 2214 40300
rect 2090 40258 2214 40277
rect 17138 40277 17157 40363
rect 17243 40340 17262 40363
rect 17243 40300 17548 40340
rect 17588 40300 17597 40340
rect 17243 40277 17262 40300
rect 17138 40258 17262 40277
rect 4919 40111 5305 40130
rect 4919 40088 4985 40111
rect 5071 40088 5153 40111
rect 5239 40088 5305 40111
rect 4919 40048 4928 40088
rect 4968 40048 4985 40088
rect 5071 40048 5092 40088
rect 5132 40048 5153 40088
rect 5239 40048 5256 40088
rect 5296 40048 5305 40088
rect 4919 40025 4985 40048
rect 5071 40025 5153 40048
rect 5239 40025 5305 40048
rect 4919 40006 5305 40025
rect 20039 40111 20425 40130
rect 20039 40088 20105 40111
rect 20191 40088 20273 40111
rect 20359 40088 20425 40111
rect 20039 40048 20048 40088
rect 20088 40048 20105 40088
rect 20191 40048 20212 40088
rect 20252 40048 20273 40088
rect 20359 40048 20376 40088
rect 20416 40048 20425 40088
rect 20039 40025 20105 40048
rect 20191 40025 20273 40048
rect 20359 40025 20425 40048
rect 20039 40006 20425 40025
rect 14659 39880 14668 39920
rect 14708 39880 18700 39920
rect 18740 39880 18749 39920
rect 15235 39712 15244 39752
rect 15284 39712 16396 39752
rect 16436 39712 16445 39752
rect 7075 39628 7084 39668
rect 7124 39628 12844 39668
rect 12884 39628 12893 39668
rect 12547 39544 12556 39584
rect 12596 39544 18412 39584
rect 18452 39544 18461 39584
rect 5347 39460 5356 39500
rect 5396 39460 13132 39500
rect 13172 39460 13181 39500
rect 14563 39460 14572 39500
rect 14612 39460 16492 39500
rect 16532 39460 16541 39500
rect 3679 39355 4065 39374
rect 3679 39332 3745 39355
rect 3831 39332 3913 39355
rect 3999 39332 4065 39355
rect 3679 39292 3688 39332
rect 3728 39292 3745 39332
rect 3831 39292 3852 39332
rect 3892 39292 3913 39332
rect 3999 39292 4016 39332
rect 4056 39292 4065 39332
rect 3679 39269 3745 39292
rect 3831 39269 3913 39292
rect 3999 39269 4065 39292
rect 3679 39250 4065 39269
rect 13034 39355 13158 39374
rect 13034 39269 13053 39355
rect 13139 39332 13158 39355
rect 18799 39355 19185 39374
rect 18799 39332 18865 39355
rect 18951 39332 19033 39355
rect 19119 39332 19185 39355
rect 13139 39292 16012 39332
rect 16052 39292 16061 39332
rect 16195 39292 16204 39332
rect 16244 39292 17644 39332
rect 17684 39292 17693 39332
rect 18799 39292 18808 39332
rect 18848 39292 18865 39332
rect 18951 39292 18972 39332
rect 19012 39292 19033 39332
rect 19119 39292 19136 39332
rect 19176 39292 19185 39332
rect 13139 39269 13158 39292
rect 13034 39250 13158 39269
rect 18799 39269 18865 39292
rect 18951 39269 19033 39292
rect 19119 39269 19185 39292
rect 18799 39250 19185 39269
rect 13891 39208 13900 39248
rect 13940 39208 16396 39248
rect 16436 39208 16445 39248
rect 16867 39124 16876 39164
rect 16916 39124 17452 39164
rect 17492 39124 17501 39164
rect 15907 39040 15916 39080
rect 15956 39040 20140 39080
rect 20180 39040 20189 39080
rect 14851 38956 14860 38996
rect 14900 38956 19276 38996
rect 19316 38956 19325 38996
rect 14179 38872 14188 38912
rect 14228 38872 14956 38912
rect 14996 38872 18604 38912
rect 18644 38872 18653 38912
rect 4579 38704 4588 38744
rect 4628 38704 10060 38744
rect 10100 38704 10109 38744
rect 16003 38704 16012 38744
rect 16052 38704 20812 38744
rect 20852 38704 20861 38744
rect 4919 38599 5305 38618
rect 4919 38576 4985 38599
rect 5071 38576 5153 38599
rect 5239 38576 5305 38599
rect 4919 38536 4928 38576
rect 4968 38536 4985 38576
rect 5071 38536 5092 38576
rect 5132 38536 5153 38576
rect 5239 38536 5256 38576
rect 5296 38536 5305 38576
rect 4919 38513 4985 38536
rect 5071 38513 5153 38536
rect 5239 38513 5305 38536
rect 4919 38494 5305 38513
rect 20039 38599 20425 38618
rect 20039 38576 20105 38599
rect 20191 38576 20273 38599
rect 20359 38576 20425 38599
rect 20039 38536 20048 38576
rect 20088 38536 20105 38576
rect 20191 38536 20212 38576
rect 20252 38536 20273 38576
rect 20359 38536 20376 38576
rect 20416 38536 20425 38576
rect 20039 38513 20105 38536
rect 20191 38513 20273 38536
rect 20359 38513 20425 38536
rect 20039 38494 20425 38513
rect 14371 38452 14380 38492
rect 14420 38452 18412 38492
rect 18452 38452 18461 38492
rect 3523 38368 3532 38408
rect 3572 38368 10732 38408
rect 10772 38368 10781 38408
rect 16675 38368 16684 38408
rect 16724 38368 20140 38408
rect 20180 38368 20189 38408
rect 7106 38263 7230 38282
rect 7106 38240 7125 38263
rect 6691 38200 6700 38240
rect 6740 38200 7125 38240
rect 7106 38177 7125 38200
rect 7211 38177 7230 38263
rect 7106 38158 7230 38177
rect 1987 38032 1996 38072
rect 2036 38032 12748 38072
rect 12788 38032 12797 38072
rect 13603 38032 13612 38072
rect 13652 38032 20140 38072
rect 20180 38032 20189 38072
rect 6211 37864 6220 37904
rect 6260 37864 10636 37904
rect 10676 37864 10685 37904
rect 3679 37843 4065 37862
rect 3679 37820 3745 37843
rect 3831 37820 3913 37843
rect 3999 37820 4065 37843
rect 3679 37780 3688 37820
rect 3728 37780 3745 37820
rect 3831 37780 3852 37820
rect 3892 37780 3913 37820
rect 3999 37780 4016 37820
rect 4056 37780 4065 37820
rect 3679 37757 3745 37780
rect 3831 37757 3913 37780
rect 3999 37757 4065 37780
rect 3679 37738 4065 37757
rect 18799 37843 19185 37862
rect 18799 37820 18865 37843
rect 18951 37820 19033 37843
rect 19119 37820 19185 37843
rect 18799 37780 18808 37820
rect 18848 37780 18865 37820
rect 18951 37780 18972 37820
rect 19012 37780 19033 37820
rect 19119 37780 19136 37820
rect 19176 37780 19185 37820
rect 18799 37757 18865 37780
rect 18951 37757 19033 37780
rect 19119 37757 19185 37780
rect 18799 37738 19185 37757
rect 8930 37507 9054 37526
rect 8930 37421 8949 37507
rect 9035 37484 9054 37507
rect 9035 37444 9388 37484
rect 9428 37444 9437 37484
rect 9035 37421 9054 37444
rect 8930 37402 9054 37421
rect 16963 37360 16972 37400
rect 17012 37360 20332 37400
rect 20372 37360 20381 37400
rect 3811 37192 3820 37232
rect 3860 37192 9100 37232
rect 9140 37192 9149 37232
rect 4919 37087 5305 37106
rect 4919 37064 4985 37087
rect 5071 37064 5153 37087
rect 5239 37064 5305 37087
rect 4919 37024 4928 37064
rect 4968 37024 4985 37064
rect 5071 37024 5092 37064
rect 5132 37024 5153 37064
rect 5239 37024 5256 37064
rect 5296 37024 5305 37064
rect 4919 37001 4985 37024
rect 5071 37001 5153 37024
rect 5239 37001 5305 37024
rect 20039 37087 20425 37106
rect 20039 37064 20105 37087
rect 20191 37064 20273 37087
rect 20359 37064 20425 37087
rect 20039 37024 20048 37064
rect 20088 37024 20105 37064
rect 20191 37024 20212 37064
rect 20252 37024 20273 37064
rect 20359 37024 20376 37064
rect 20416 37024 20425 37064
rect 4919 36982 5305 37001
rect 13946 37003 14070 37022
rect 13946 36980 13965 37003
rect 12931 36940 12940 36980
rect 12980 36940 13965 36980
rect 13946 36917 13965 36940
rect 14051 36917 14070 37003
rect 20039 37001 20105 37024
rect 20191 37001 20273 37024
rect 20359 37001 20425 37024
rect 20039 36982 20425 37001
rect 13946 36898 14070 36917
rect 1987 36772 1996 36812
rect 2036 36772 2380 36812
rect 2420 36772 2429 36812
rect 3043 36688 3052 36728
rect 3092 36688 7276 36728
rect 7316 36688 7325 36728
rect 2179 36604 2188 36644
rect 2228 36604 2380 36644
rect 2420 36604 19468 36644
rect 19508 36604 19517 36644
rect 10627 36520 10636 36560
rect 10676 36520 12556 36560
rect 12596 36520 12605 36560
rect 4483 36436 4492 36476
rect 4532 36436 17644 36476
rect 17684 36436 17693 36476
rect 3679 36331 4065 36350
rect 3679 36308 3745 36331
rect 3831 36308 3913 36331
rect 3999 36308 4065 36331
rect 3679 36268 3688 36308
rect 3728 36268 3745 36308
rect 3831 36268 3852 36308
rect 3892 36268 3913 36308
rect 3999 36268 4016 36308
rect 4056 36268 4065 36308
rect 3679 36245 3745 36268
rect 3831 36245 3913 36268
rect 3999 36245 4065 36268
rect 3679 36226 4065 36245
rect 18799 36331 19185 36350
rect 18799 36308 18865 36331
rect 18951 36308 19033 36331
rect 19119 36308 19185 36331
rect 18799 36268 18808 36308
rect 18848 36268 18865 36308
rect 18951 36268 18972 36308
rect 19012 36268 19033 36308
rect 19119 36268 19136 36308
rect 19176 36268 19185 36308
rect 18799 36245 18865 36268
rect 18951 36245 19033 36268
rect 19119 36245 19185 36268
rect 18799 36226 19185 36245
rect 3523 35932 3532 35972
rect 3572 35932 18796 35972
rect 18836 35932 18845 35972
rect 547 35848 556 35888
rect 596 35848 20620 35888
rect 20660 35848 20669 35888
rect 2179 35680 2188 35720
rect 2228 35680 7564 35720
rect 7604 35680 7613 35720
rect 4919 35575 5305 35594
rect 4919 35552 4985 35575
rect 5071 35552 5153 35575
rect 5239 35552 5305 35575
rect 4919 35512 4928 35552
rect 4968 35512 4985 35552
rect 5071 35512 5092 35552
rect 5132 35512 5153 35552
rect 5239 35512 5256 35552
rect 5296 35512 5305 35552
rect 4919 35489 4985 35512
rect 5071 35489 5153 35512
rect 5239 35489 5305 35512
rect 4919 35470 5305 35489
rect 20039 35575 20425 35594
rect 20039 35552 20105 35575
rect 20191 35552 20273 35575
rect 20359 35552 20425 35575
rect 20039 35512 20048 35552
rect 20088 35512 20105 35552
rect 20191 35512 20212 35552
rect 20252 35512 20273 35552
rect 20359 35512 20376 35552
rect 20416 35512 20425 35552
rect 20039 35489 20105 35512
rect 20191 35489 20273 35512
rect 20359 35489 20425 35512
rect 20039 35470 20425 35489
rect 5635 35260 5644 35300
rect 5684 35260 5820 35300
rect 8899 35260 8908 35300
rect 8948 35260 14188 35300
rect 14228 35260 14237 35300
rect 5780 35216 5820 35260
rect 3619 35176 3628 35216
rect 3668 35176 5820 35216
rect 6115 35176 6124 35216
rect 6164 35176 15436 35216
rect 15476 35176 15485 35216
rect 5780 35048 5820 35176
rect 5780 35008 6316 35048
rect 6356 35008 6365 35048
rect 9379 35008 9388 35048
rect 9428 35008 10444 35048
rect 10484 35008 10493 35048
rect 5251 34924 5260 34964
rect 5300 34924 5932 34964
rect 5972 34924 5981 34964
rect 10723 34924 10732 34964
rect 10772 34924 20180 34964
rect 2947 34840 2956 34880
rect 2996 34840 3436 34880
rect 3476 34840 3485 34880
rect 3679 34819 4065 34838
rect 3679 34796 3745 34819
rect 3831 34796 3913 34819
rect 3999 34796 4065 34819
rect 3679 34756 3688 34796
rect 3728 34756 3745 34796
rect 3831 34756 3852 34796
rect 3892 34756 3913 34796
rect 3999 34756 4016 34796
rect 4056 34756 4065 34796
rect 3679 34733 3745 34756
rect 3831 34733 3913 34756
rect 3999 34733 4065 34756
rect 3679 34714 4065 34733
rect 18799 34819 19185 34838
rect 18799 34796 18865 34819
rect 18951 34796 19033 34819
rect 19119 34796 19185 34819
rect 18799 34756 18808 34796
rect 18848 34756 18865 34796
rect 18951 34756 18972 34796
rect 19012 34756 19033 34796
rect 19119 34756 19136 34796
rect 19176 34756 19185 34796
rect 18799 34733 18865 34756
rect 18951 34733 19033 34756
rect 19119 34733 19185 34756
rect 18799 34714 19185 34733
rect 20140 34712 20180 34924
rect 20131 34672 20140 34712
rect 20180 34672 20189 34712
rect 4675 34588 4684 34628
rect 4724 34588 9484 34628
rect 9524 34588 9533 34628
rect 12067 34588 12076 34628
rect 12116 34588 17452 34628
rect 17492 34588 17501 34628
rect 1315 34504 1324 34544
rect 1364 34504 13036 34544
rect 13076 34504 13085 34544
rect 4483 34420 4492 34460
rect 4532 34420 4876 34460
rect 4916 34420 4925 34460
rect 6883 34420 6892 34460
rect 6932 34420 7564 34460
rect 7604 34420 7613 34460
rect 8419 34420 8428 34460
rect 8468 34420 13996 34460
rect 14036 34420 14045 34460
rect 8035 34336 8044 34376
rect 8084 34336 15628 34376
rect 15668 34336 19276 34376
rect 19316 34336 19325 34376
rect 6499 34252 6508 34292
rect 6548 34252 11360 34292
rect 11320 34208 11360 34252
rect 4771 34168 4780 34208
rect 4820 34168 11212 34208
rect 11252 34168 11261 34208
rect 11320 34168 15148 34208
rect 15188 34168 15197 34208
rect 14467 34084 14476 34124
rect 14516 34084 16204 34124
rect 16244 34084 16253 34124
rect 4919 34063 5305 34082
rect 4919 34040 4985 34063
rect 5071 34040 5153 34063
rect 5239 34040 5305 34063
rect 20039 34063 20425 34082
rect 20039 34040 20105 34063
rect 20191 34040 20273 34063
rect 20359 34040 20425 34063
rect 4919 34000 4928 34040
rect 4968 34000 4985 34040
rect 5071 34000 5092 34040
rect 5132 34000 5153 34040
rect 5239 34000 5256 34040
rect 5296 34000 5305 34040
rect 14947 34000 14956 34040
rect 14996 34000 15916 34040
rect 15956 34000 15965 34040
rect 20039 34000 20048 34040
rect 20088 34000 20105 34040
rect 20191 34000 20212 34040
rect 20252 34000 20273 34040
rect 20359 34000 20376 34040
rect 20416 34000 20425 34040
rect 4919 33977 4985 34000
rect 5071 33977 5153 34000
rect 5239 33977 5305 34000
rect 4919 33958 5305 33977
rect 20039 33977 20105 34000
rect 20191 33977 20273 34000
rect 20359 33977 20425 34000
rect 20039 33958 20425 33977
rect 12547 33580 12556 33620
rect 12596 33580 19468 33620
rect 19508 33580 19517 33620
rect 12835 33412 12844 33452
rect 12884 33412 13036 33452
rect 13076 33412 13085 33452
rect 3679 33307 4065 33326
rect 3679 33284 3745 33307
rect 3831 33284 3913 33307
rect 3999 33284 4065 33307
rect 3679 33244 3688 33284
rect 3728 33244 3745 33284
rect 3831 33244 3852 33284
rect 3892 33244 3913 33284
rect 3999 33244 4016 33284
rect 4056 33244 4065 33284
rect 3679 33221 3745 33244
rect 3831 33221 3913 33244
rect 3999 33221 4065 33244
rect 3679 33202 4065 33221
rect 18799 33307 19185 33326
rect 18799 33284 18865 33307
rect 18951 33284 19033 33307
rect 19119 33284 19185 33307
rect 18799 33244 18808 33284
rect 18848 33244 18865 33284
rect 18951 33244 18972 33284
rect 19012 33244 19033 33284
rect 19119 33244 19136 33284
rect 19176 33244 19185 33284
rect 18799 33221 18865 33244
rect 18951 33221 19033 33244
rect 19119 33221 19185 33244
rect 18799 33202 19185 33221
rect 13795 33076 13804 33116
rect 13844 33076 16012 33116
rect 16052 33076 16061 33116
rect 2755 32992 2764 33032
rect 2804 32992 14092 33032
rect 14132 32992 14141 33032
rect 14275 32992 14284 33032
rect 14324 32992 17452 33032
rect 17492 32992 17501 33032
rect 6691 32908 6700 32948
rect 6740 32908 8044 32948
rect 8084 32908 13804 32948
rect 13844 32908 13853 32948
rect 15770 32887 15894 32906
rect 15770 32864 15789 32887
rect 11587 32824 11596 32864
rect 11636 32824 15789 32864
rect 15770 32801 15789 32824
rect 15875 32801 15894 32887
rect 15770 32782 15894 32801
rect 4919 32551 5305 32570
rect 4919 32528 4985 32551
rect 5071 32528 5153 32551
rect 5239 32528 5305 32551
rect 20039 32551 20425 32570
rect 20039 32528 20105 32551
rect 20191 32528 20273 32551
rect 20359 32528 20425 32551
rect 4919 32488 4928 32528
rect 4968 32488 4985 32528
rect 5071 32488 5092 32528
rect 5132 32488 5153 32528
rect 5239 32488 5256 32528
rect 5296 32488 5305 32528
rect 13891 32488 13900 32528
rect 13940 32488 17068 32528
rect 17108 32488 17117 32528
rect 20039 32488 20048 32528
rect 20088 32488 20105 32528
rect 20191 32488 20212 32528
rect 20252 32488 20273 32528
rect 20359 32488 20376 32528
rect 20416 32488 20425 32528
rect 4919 32465 4985 32488
rect 5071 32465 5153 32488
rect 5239 32465 5305 32488
rect 4919 32446 5305 32465
rect 20039 32465 20105 32488
rect 20191 32465 20273 32488
rect 20359 32465 20425 32488
rect 20039 32446 20425 32465
rect 9091 31900 9100 31940
rect 9140 31900 20180 31940
rect 3679 31795 4065 31814
rect 3679 31772 3745 31795
rect 3831 31772 3913 31795
rect 3999 31772 4065 31795
rect 1699 31732 1708 31772
rect 1748 31732 1900 31772
rect 1940 31732 1949 31772
rect 3679 31732 3688 31772
rect 3728 31732 3745 31772
rect 3831 31732 3852 31772
rect 3892 31732 3913 31772
rect 3999 31732 4016 31772
rect 4056 31732 4065 31772
rect 3679 31709 3745 31732
rect 3831 31709 3913 31732
rect 3999 31709 4065 31732
rect 3679 31690 4065 31709
rect 18799 31795 19185 31814
rect 18799 31772 18865 31795
rect 18951 31772 19033 31795
rect 19119 31772 19185 31795
rect 18799 31732 18808 31772
rect 18848 31732 18865 31772
rect 18951 31732 18972 31772
rect 19012 31732 19033 31772
rect 19119 31732 19136 31772
rect 19176 31732 19185 31772
rect 18799 31709 18865 31732
rect 18951 31709 19033 31732
rect 19119 31709 19185 31732
rect 18799 31690 19185 31709
rect 20140 31688 20180 31900
rect 20131 31648 20140 31688
rect 20180 31648 20189 31688
rect 13699 31228 13708 31268
rect 13748 31228 18508 31268
rect 18548 31228 18557 31268
rect 17923 31144 17932 31184
rect 17972 31144 18220 31184
rect 18260 31144 18269 31184
rect 4919 31039 5305 31058
rect 4919 31016 4985 31039
rect 5071 31016 5153 31039
rect 5239 31016 5305 31039
rect 4919 30976 4928 31016
rect 4968 30976 4985 31016
rect 5071 30976 5092 31016
rect 5132 30976 5153 31016
rect 5239 30976 5256 31016
rect 5296 30976 5305 31016
rect 4919 30953 4985 30976
rect 5071 30953 5153 30976
rect 5239 30953 5305 30976
rect 4919 30934 5305 30953
rect 20039 31039 20425 31058
rect 20039 31016 20105 31039
rect 20191 31016 20273 31039
rect 20359 31016 20425 31039
rect 20039 30976 20048 31016
rect 20088 30976 20105 31016
rect 20191 30976 20212 31016
rect 20252 30976 20273 31016
rect 20359 30976 20376 31016
rect 20416 30976 20425 31016
rect 20039 30953 20105 30976
rect 20191 30953 20273 30976
rect 20359 30953 20425 30976
rect 20039 30934 20425 30953
rect 1507 30724 1516 30764
rect 1556 30724 5548 30764
rect 5588 30724 5597 30764
rect 10531 30304 10540 30344
rect 10580 30304 11116 30344
rect 11156 30304 11165 30344
rect 3679 30283 4065 30302
rect 3679 30260 3745 30283
rect 3831 30260 3913 30283
rect 3999 30260 4065 30283
rect 3679 30220 3688 30260
rect 3728 30220 3745 30260
rect 3831 30220 3852 30260
rect 3892 30220 3913 30260
rect 3999 30220 4016 30260
rect 4056 30220 4065 30260
rect 3679 30197 3745 30220
rect 3831 30197 3913 30220
rect 3999 30197 4065 30220
rect 3679 30178 4065 30197
rect 18799 30283 19185 30302
rect 18799 30260 18865 30283
rect 18951 30260 19033 30283
rect 19119 30260 19185 30283
rect 18799 30220 18808 30260
rect 18848 30220 18865 30260
rect 18951 30220 18972 30260
rect 19012 30220 19033 30260
rect 19119 30220 19136 30260
rect 19176 30220 19185 30260
rect 18799 30197 18865 30220
rect 18951 30197 19033 30220
rect 19119 30197 19185 30220
rect 18799 30178 19185 30197
rect 1219 29968 1228 30008
rect 1268 29968 2956 30008
rect 2996 29968 3005 30008
rect 8611 29548 8620 29588
rect 8660 29548 15628 29588
rect 15668 29548 15677 29588
rect 4919 29527 5305 29546
rect 4919 29504 4985 29527
rect 5071 29504 5153 29527
rect 5239 29504 5305 29527
rect 4919 29464 4928 29504
rect 4968 29464 4985 29504
rect 5071 29464 5092 29504
rect 5132 29464 5153 29504
rect 5239 29464 5256 29504
rect 5296 29464 5305 29504
rect 4919 29441 4985 29464
rect 5071 29441 5153 29464
rect 5239 29441 5305 29464
rect 4919 29422 5305 29441
rect 20039 29527 20425 29546
rect 20039 29504 20105 29527
rect 20191 29504 20273 29527
rect 20359 29504 20425 29527
rect 20039 29464 20048 29504
rect 20088 29464 20105 29504
rect 20191 29464 20212 29504
rect 20252 29464 20273 29504
rect 20359 29464 20376 29504
rect 20416 29464 20425 29504
rect 20039 29441 20105 29464
rect 20191 29441 20273 29464
rect 20359 29441 20425 29464
rect 20039 29422 20425 29441
rect 2659 29380 2668 29420
rect 2708 29380 2996 29420
rect 2588 29296 2860 29336
rect 2900 29296 2909 29336
rect 2588 29000 2628 29296
rect 2956 29252 2996 29380
rect 2563 28960 2572 29000
rect 2612 28960 2628 29000
rect 2860 29212 2996 29252
rect 3235 29212 3244 29252
rect 3284 29212 8620 29252
rect 8660 29212 8669 29252
rect 2860 28916 2900 29212
rect 3331 29128 3340 29168
rect 3380 29128 4300 29168
rect 4340 29128 8332 29168
rect 8372 29128 8381 29168
rect 10723 29128 10732 29168
rect 10772 29128 13420 29168
rect 13460 29128 13469 29168
rect 8707 29044 8716 29084
rect 8756 29044 9772 29084
rect 9812 29044 9821 29084
rect 2851 28876 2860 28916
rect 2900 28876 2909 28916
rect 2275 28792 2284 28832
rect 2324 28792 2764 28832
rect 2804 28792 2813 28832
rect 3679 28771 4065 28790
rect 3679 28748 3745 28771
rect 3831 28748 3913 28771
rect 3999 28748 4065 28771
rect 3679 28708 3688 28748
rect 3728 28708 3745 28748
rect 3831 28708 3852 28748
rect 3892 28708 3913 28748
rect 3999 28708 4016 28748
rect 4056 28708 4065 28748
rect 3679 28685 3745 28708
rect 3831 28685 3913 28708
rect 3999 28685 4065 28708
rect 3679 28666 4065 28685
rect 18799 28771 19185 28790
rect 18799 28748 18865 28771
rect 18951 28748 19033 28771
rect 19119 28748 19185 28771
rect 18799 28708 18808 28748
rect 18848 28708 18865 28748
rect 18951 28708 18972 28748
rect 19012 28708 19033 28748
rect 19119 28708 19136 28748
rect 19176 28708 19185 28748
rect 18799 28685 18865 28708
rect 18951 28685 19033 28708
rect 19119 28685 19185 28708
rect 18799 28666 19185 28685
rect 8131 28624 8140 28664
rect 8180 28624 8524 28664
rect 8564 28624 8573 28664
rect 8018 28435 8142 28454
rect 8018 28412 8037 28435
rect 7459 28372 7468 28412
rect 7508 28372 8037 28412
rect 8018 28349 8037 28372
rect 8123 28349 8142 28435
rect 8018 28330 8142 28349
rect 11666 28267 11790 28286
rect 11666 28244 11685 28267
rect 3619 28204 3628 28244
rect 3668 28204 11685 28244
rect 11666 28181 11685 28204
rect 11771 28181 11790 28267
rect 11666 28162 11790 28181
rect 4919 28015 5305 28034
rect 4919 27992 4985 28015
rect 5071 27992 5153 28015
rect 5239 27992 5305 28015
rect 4919 27952 4928 27992
rect 4968 27952 4985 27992
rect 5071 27952 5092 27992
rect 5132 27952 5153 27992
rect 5239 27952 5256 27992
rect 5296 27952 5305 27992
rect 4919 27929 4985 27952
rect 5071 27929 5153 27952
rect 5239 27929 5305 27952
rect 4919 27910 5305 27929
rect 20039 28015 20425 28034
rect 20039 27992 20105 28015
rect 20191 27992 20273 28015
rect 20359 27992 20425 28015
rect 20039 27952 20048 27992
rect 20088 27952 20105 27992
rect 20191 27952 20212 27992
rect 20252 27952 20273 27992
rect 20359 27952 20376 27992
rect 20416 27952 20425 27992
rect 20039 27929 20105 27952
rect 20191 27929 20273 27952
rect 20359 27929 20425 27952
rect 20039 27910 20425 27929
rect 3139 27700 3148 27740
rect 3188 27700 4492 27740
rect 4532 27700 4541 27740
rect 10531 27700 10540 27740
rect 10580 27700 12844 27740
rect 12884 27700 12893 27740
rect 4099 27616 4108 27656
rect 4148 27616 9388 27656
rect 9428 27616 9437 27656
rect 10627 27616 10636 27656
rect 10676 27616 11020 27656
rect 11060 27616 11069 27656
rect 12259 27616 12268 27656
rect 12308 27616 12460 27656
rect 12500 27616 12509 27656
rect 5443 27532 5452 27572
rect 5492 27532 6796 27572
rect 6836 27532 6845 27572
rect 8803 27532 8812 27572
rect 8852 27532 18028 27572
rect 18068 27532 18077 27572
rect 10915 27448 10924 27488
rect 10964 27448 12460 27488
rect 12500 27448 12509 27488
rect 3679 27259 4065 27278
rect 3679 27236 3745 27259
rect 3831 27236 3913 27259
rect 3999 27236 4065 27259
rect 3679 27196 3688 27236
rect 3728 27196 3745 27236
rect 3831 27196 3852 27236
rect 3892 27196 3913 27236
rect 3999 27196 4016 27236
rect 4056 27196 4065 27236
rect 3679 27173 3745 27196
rect 3831 27173 3913 27196
rect 3999 27173 4065 27196
rect 3679 27154 4065 27173
rect 18799 27259 19185 27278
rect 18799 27236 18865 27259
rect 18951 27236 19033 27259
rect 19119 27236 19185 27259
rect 18799 27196 18808 27236
rect 18848 27196 18865 27236
rect 18951 27196 18972 27236
rect 19012 27196 19033 27236
rect 19119 27196 19136 27236
rect 19176 27196 19185 27236
rect 18799 27173 18865 27196
rect 18951 27173 19033 27196
rect 19119 27173 19185 27196
rect 18799 27154 19185 27173
rect 11011 26776 11020 26816
rect 11060 26776 11980 26816
rect 12020 26776 12029 26816
rect 2275 26692 2284 26732
rect 2324 26692 6124 26732
rect 6164 26692 6700 26732
rect 6740 26692 6749 26732
rect 9842 26671 9966 26690
rect 9842 26648 9861 26671
rect 4291 26608 4300 26648
rect 4340 26608 9861 26648
rect 9842 26585 9861 26608
rect 9947 26585 9966 26671
rect 19747 26608 19756 26648
rect 19796 26608 19948 26648
rect 19988 26608 19997 26648
rect 9842 26566 9966 26585
rect 11299 26524 11308 26564
rect 11348 26524 12844 26564
rect 12884 26524 12893 26564
rect 4919 26503 5305 26522
rect 4919 26480 4985 26503
rect 5071 26480 5153 26503
rect 5239 26480 5305 26503
rect 4919 26440 4928 26480
rect 4968 26440 4985 26480
rect 5071 26440 5092 26480
rect 5132 26440 5153 26480
rect 5239 26440 5256 26480
rect 5296 26440 5305 26480
rect 4919 26417 4985 26440
rect 5071 26417 5153 26440
rect 5239 26417 5305 26440
rect 4919 26398 5305 26417
rect 8930 26503 9054 26522
rect 8930 26417 8949 26503
rect 9035 26480 9054 26503
rect 9044 26440 9054 26480
rect 9035 26417 9054 26440
rect 8930 26398 9054 26417
rect 20039 26503 20425 26522
rect 20039 26480 20105 26503
rect 20191 26480 20273 26503
rect 20359 26480 20425 26503
rect 20039 26440 20048 26480
rect 20088 26440 20105 26480
rect 20191 26440 20212 26480
rect 20252 26440 20273 26480
rect 20359 26440 20376 26480
rect 20416 26440 20425 26480
rect 20039 26417 20105 26440
rect 20191 26417 20273 26440
rect 20359 26417 20425 26440
rect 20039 26398 20425 26417
rect 67 25852 76 25892
rect 116 25852 1228 25892
rect 1268 25852 5644 25892
rect 5684 25852 7948 25892
rect 7988 25852 7997 25892
rect 3679 25747 4065 25766
rect 3679 25724 3745 25747
rect 3831 25724 3913 25747
rect 3999 25724 4065 25747
rect 3679 25684 3688 25724
rect 3728 25684 3745 25724
rect 3831 25684 3852 25724
rect 3892 25684 3913 25724
rect 3999 25684 4016 25724
rect 4056 25684 4065 25724
rect 3679 25661 3745 25684
rect 3831 25661 3913 25684
rect 3999 25661 4065 25684
rect 3679 25642 4065 25661
rect 18799 25747 19185 25766
rect 18799 25724 18865 25747
rect 18951 25724 19033 25747
rect 19119 25724 19185 25747
rect 18799 25684 18808 25724
rect 18848 25684 18865 25724
rect 18951 25684 18972 25724
rect 19012 25684 19033 25724
rect 19119 25684 19136 25724
rect 19176 25684 19185 25724
rect 18799 25661 18865 25684
rect 18951 25661 19033 25684
rect 19119 25661 19185 25684
rect 18799 25642 19185 25661
rect 5059 25264 5068 25304
rect 5108 25264 10060 25304
rect 10100 25264 10109 25304
rect 6211 25096 6220 25136
rect 6260 25096 6892 25136
rect 6932 25096 6941 25136
rect 4919 24991 5305 25010
rect 4919 24968 4985 24991
rect 5071 24968 5153 24991
rect 5239 24968 5305 24991
rect 4919 24928 4928 24968
rect 4968 24928 4985 24968
rect 5071 24928 5092 24968
rect 5132 24928 5153 24968
rect 5239 24928 5256 24968
rect 5296 24928 5305 24968
rect 4919 24905 4985 24928
rect 5071 24905 5153 24928
rect 5239 24905 5305 24928
rect 4919 24886 5305 24905
rect 20039 24991 20425 25010
rect 20039 24968 20105 24991
rect 20191 24968 20273 24991
rect 20359 24968 20425 24991
rect 20039 24928 20048 24968
rect 20088 24928 20105 24968
rect 20191 24928 20212 24968
rect 20252 24928 20273 24968
rect 20359 24928 20376 24968
rect 20416 24928 20425 24968
rect 20039 24905 20105 24928
rect 20191 24905 20273 24928
rect 20359 24905 20425 24928
rect 20039 24886 20425 24905
rect 7106 24739 7230 24758
rect 7106 24716 7125 24739
rect 5443 24676 5452 24716
rect 5492 24676 7125 24716
rect 7106 24653 7125 24676
rect 7211 24653 7230 24739
rect 7106 24634 7230 24653
rect 15619 24592 15628 24632
rect 15668 24592 15820 24632
rect 15860 24592 15869 24632
rect 4387 24508 4396 24548
rect 4436 24508 4780 24548
rect 4820 24508 4829 24548
rect 3679 24235 4065 24254
rect 3679 24212 3745 24235
rect 3831 24212 3913 24235
rect 3999 24212 4065 24235
rect 3679 24172 3688 24212
rect 3728 24172 3745 24212
rect 3831 24172 3852 24212
rect 3892 24172 3913 24212
rect 3999 24172 4016 24212
rect 4056 24172 4065 24212
rect 3679 24149 3745 24172
rect 3831 24149 3913 24172
rect 3999 24149 4065 24172
rect 3679 24130 4065 24149
rect 18799 24235 19185 24254
rect 18799 24212 18865 24235
rect 18951 24212 19033 24235
rect 19119 24212 19185 24235
rect 18799 24172 18808 24212
rect 18848 24172 18865 24212
rect 18951 24172 18972 24212
rect 19012 24172 19033 24212
rect 19119 24172 19136 24212
rect 19176 24172 19185 24212
rect 18799 24149 18865 24172
rect 18951 24149 19033 24172
rect 19119 24149 19185 24172
rect 18799 24130 19185 24149
rect 7106 24067 7230 24086
rect 7106 23981 7125 24067
rect 7211 24044 7230 24067
rect 7211 24004 7372 24044
rect 7412 24004 7421 24044
rect 7211 23981 7230 24004
rect 7106 23962 7230 23981
rect 1178 23731 1302 23750
rect 1178 23645 1197 23731
rect 1283 23708 1302 23731
rect 1283 23668 8908 23708
rect 8948 23668 8957 23708
rect 1283 23645 1302 23668
rect 1178 23626 1302 23645
rect 4579 23584 4588 23624
rect 4628 23584 16684 23624
rect 16724 23584 16733 23624
rect 4919 23479 5305 23498
rect 4919 23456 4985 23479
rect 5071 23456 5153 23479
rect 5239 23456 5305 23479
rect 4919 23416 4928 23456
rect 4968 23416 4985 23456
rect 5071 23416 5092 23456
rect 5132 23416 5153 23456
rect 5239 23416 5256 23456
rect 5296 23416 5305 23456
rect 4919 23393 4985 23416
rect 5071 23393 5153 23416
rect 5239 23393 5305 23416
rect 4919 23374 5305 23393
rect 20039 23479 20425 23498
rect 20039 23456 20105 23479
rect 20191 23456 20273 23479
rect 20359 23456 20425 23479
rect 20039 23416 20048 23456
rect 20088 23416 20105 23456
rect 20191 23416 20212 23456
rect 20252 23416 20273 23456
rect 20359 23416 20376 23456
rect 20416 23416 20425 23456
rect 20039 23393 20105 23416
rect 20191 23393 20273 23416
rect 20359 23393 20425 23416
rect 20039 23374 20425 23393
rect 1027 23248 1036 23288
rect 1076 23248 14380 23288
rect 14420 23248 14429 23288
rect 4579 22996 4588 23036
rect 4628 22996 10252 23036
rect 10292 22996 10301 23036
rect 4291 22912 4300 22952
rect 4340 22912 6700 22952
rect 6740 22912 6749 22952
rect 6211 22828 6220 22868
rect 6260 22828 17356 22868
rect 17396 22828 17405 22868
rect 3679 22723 4065 22742
rect 3679 22700 3745 22723
rect 3831 22700 3913 22723
rect 3999 22700 4065 22723
rect 18799 22723 19185 22742
rect 18799 22700 18865 22723
rect 18951 22700 19033 22723
rect 19119 22700 19185 22723
rect 3679 22660 3688 22700
rect 3728 22660 3745 22700
rect 3831 22660 3852 22700
rect 3892 22660 3913 22700
rect 3999 22660 4016 22700
rect 4056 22660 4065 22700
rect 14755 22660 14764 22700
rect 14804 22660 17836 22700
rect 17876 22660 17885 22700
rect 18799 22660 18808 22700
rect 18848 22660 18865 22700
rect 18951 22660 18972 22700
rect 19012 22660 19033 22700
rect 19119 22660 19136 22700
rect 19176 22660 19185 22700
rect 3679 22637 3745 22660
rect 3831 22637 3913 22660
rect 3999 22637 4065 22660
rect 3679 22618 4065 22637
rect 18799 22637 18865 22660
rect 18951 22637 19033 22660
rect 19119 22637 19185 22660
rect 18799 22618 19185 22637
rect 4099 22492 4108 22532
rect 4148 22492 4588 22532
rect 4628 22492 4637 22532
rect 13603 22492 13612 22532
rect 13652 22492 16972 22532
rect 17012 22492 17021 22532
rect 1219 22408 1228 22448
rect 1268 22408 11500 22448
rect 11540 22408 11549 22448
rect 2659 22324 2668 22364
rect 2708 22324 5932 22364
rect 5972 22324 5981 22364
rect 4099 22240 4108 22280
rect 4148 22240 4300 22280
rect 4340 22240 4349 22280
rect 6307 21988 6316 22028
rect 6356 21988 6700 22028
rect 6740 21988 6749 22028
rect 4919 21967 5305 21986
rect 4919 21944 4985 21967
rect 5071 21944 5153 21967
rect 5239 21944 5305 21967
rect 4919 21904 4928 21944
rect 4968 21904 4985 21944
rect 5071 21904 5092 21944
rect 5132 21904 5153 21944
rect 5239 21904 5256 21944
rect 5296 21904 5305 21944
rect 4919 21881 4985 21904
rect 5071 21881 5153 21904
rect 5239 21881 5305 21904
rect 4919 21862 5305 21881
rect 20039 21967 20425 21986
rect 20039 21944 20105 21967
rect 20191 21944 20273 21967
rect 20359 21944 20425 21967
rect 20039 21904 20048 21944
rect 20088 21904 20105 21944
rect 20191 21904 20212 21944
rect 20252 21904 20273 21944
rect 20359 21904 20376 21944
rect 20416 21904 20425 21944
rect 20039 21881 20105 21904
rect 20191 21881 20273 21904
rect 20359 21881 20425 21904
rect 20039 21862 20425 21881
rect 2090 21799 2214 21818
rect 2090 21776 2109 21799
rect 1891 21736 1900 21776
rect 1940 21736 2109 21776
rect 2090 21713 2109 21736
rect 2195 21713 2214 21799
rect 3715 21736 3724 21776
rect 3764 21736 5452 21776
rect 5492 21736 5501 21776
rect 2090 21694 2214 21713
rect 3679 21211 4065 21230
rect 3679 21188 3745 21211
rect 3831 21188 3913 21211
rect 3999 21188 4065 21211
rect 3679 21148 3688 21188
rect 3728 21148 3745 21188
rect 3831 21148 3852 21188
rect 3892 21148 3913 21188
rect 3999 21148 4016 21188
rect 4056 21148 4065 21188
rect 3679 21125 3745 21148
rect 3831 21125 3913 21148
rect 3999 21125 4065 21148
rect 3679 21106 4065 21125
rect 18799 21211 19185 21230
rect 18799 21188 18865 21211
rect 18951 21188 19033 21211
rect 19119 21188 19185 21211
rect 18799 21148 18808 21188
rect 18848 21148 18865 21188
rect 18951 21148 18972 21188
rect 19012 21148 19033 21188
rect 19119 21148 19136 21188
rect 19176 21148 19185 21188
rect 18799 21125 18865 21148
rect 18951 21125 19033 21148
rect 19119 21125 19185 21148
rect 18799 21106 19185 21125
rect 4919 20455 5305 20474
rect 4919 20432 4985 20455
rect 5071 20432 5153 20455
rect 5239 20432 5305 20455
rect 4919 20392 4928 20432
rect 4968 20392 4985 20432
rect 5071 20392 5092 20432
rect 5132 20392 5153 20432
rect 5239 20392 5256 20432
rect 5296 20392 5305 20432
rect 4919 20369 4985 20392
rect 5071 20369 5153 20392
rect 5239 20369 5305 20392
rect 4919 20350 5305 20369
rect 20039 20455 20425 20474
rect 20039 20432 20105 20455
rect 20191 20432 20273 20455
rect 20359 20432 20425 20455
rect 20039 20392 20048 20432
rect 20088 20392 20105 20432
rect 20191 20392 20212 20432
rect 20252 20392 20273 20432
rect 20359 20392 20376 20432
rect 20416 20392 20425 20432
rect 20039 20369 20105 20392
rect 20191 20369 20273 20392
rect 20359 20369 20425 20392
rect 20039 20350 20425 20369
rect 19459 20224 19468 20264
rect 19508 20224 19852 20264
rect 19892 20224 19901 20264
rect 1219 19888 1228 19928
rect 1268 19888 14956 19928
rect 14996 19888 15005 19928
rect 3679 19699 4065 19718
rect 3679 19676 3745 19699
rect 3831 19676 3913 19699
rect 3999 19676 4065 19699
rect 3679 19636 3688 19676
rect 3728 19636 3745 19676
rect 3831 19636 3852 19676
rect 3892 19636 3913 19676
rect 3999 19636 4016 19676
rect 4056 19636 4065 19676
rect 3679 19613 3745 19636
rect 3831 19613 3913 19636
rect 3999 19613 4065 19636
rect 3679 19594 4065 19613
rect 18799 19699 19185 19718
rect 18799 19676 18865 19699
rect 18951 19676 19033 19699
rect 19119 19676 19185 19699
rect 18799 19636 18808 19676
rect 18848 19636 18865 19676
rect 18951 19636 18972 19676
rect 19012 19636 19033 19676
rect 19119 19636 19136 19676
rect 19176 19636 19185 19676
rect 18799 19613 18865 19636
rect 18951 19613 19033 19636
rect 19119 19613 19185 19636
rect 18799 19594 19185 19613
rect 10754 19111 10878 19130
rect 10754 19088 10773 19111
rect 4291 19048 4300 19088
rect 4340 19048 10773 19088
rect 10754 19025 10773 19048
rect 10859 19025 10878 19111
rect 10754 19006 10878 19025
rect 4919 18943 5305 18962
rect 4919 18920 4985 18943
rect 5071 18920 5153 18943
rect 5239 18920 5305 18943
rect 20039 18943 20425 18962
rect 20039 18920 20105 18943
rect 20191 18920 20273 18943
rect 20359 18920 20425 18943
rect 4919 18880 4928 18920
rect 4968 18880 4985 18920
rect 5071 18880 5092 18920
rect 5132 18880 5153 18920
rect 5239 18880 5256 18920
rect 5296 18880 5305 18920
rect 9667 18880 9676 18920
rect 9716 18880 14764 18920
rect 14804 18880 14813 18920
rect 20039 18880 20048 18920
rect 20088 18880 20105 18920
rect 20191 18880 20212 18920
rect 20252 18880 20273 18920
rect 20359 18880 20376 18920
rect 20416 18880 20425 18920
rect 4919 18857 4985 18880
rect 5071 18857 5153 18880
rect 5239 18857 5305 18880
rect 4919 18838 5305 18857
rect 20039 18857 20105 18880
rect 20191 18857 20273 18880
rect 20359 18857 20425 18880
rect 20039 18838 20425 18857
rect 1699 18544 1708 18584
rect 1748 18544 2188 18584
rect 2228 18544 2237 18584
rect 259 18460 268 18500
rect 308 18460 17260 18500
rect 17300 18460 17309 18500
rect 1219 18376 1228 18416
rect 1268 18376 17164 18416
rect 17204 18376 17213 18416
rect 2947 18292 2956 18332
rect 2996 18292 4780 18332
rect 4820 18292 4829 18332
rect 3679 18187 4065 18206
rect 3679 18164 3745 18187
rect 3831 18164 3913 18187
rect 3999 18164 4065 18187
rect 3679 18124 3688 18164
rect 3728 18124 3745 18164
rect 3831 18124 3852 18164
rect 3892 18124 3913 18164
rect 3999 18124 4016 18164
rect 4056 18124 4065 18164
rect 3679 18101 3745 18124
rect 3831 18101 3913 18124
rect 3999 18101 4065 18124
rect 3679 18082 4065 18101
rect 18799 18187 19185 18206
rect 18799 18164 18865 18187
rect 18951 18164 19033 18187
rect 19119 18164 19185 18187
rect 18799 18124 18808 18164
rect 18848 18124 18865 18164
rect 18951 18124 18972 18164
rect 19012 18124 19033 18164
rect 19119 18124 19136 18164
rect 19176 18124 19185 18164
rect 18799 18101 18865 18124
rect 18951 18101 19033 18124
rect 19119 18101 19185 18124
rect 18799 18082 19185 18101
rect 1178 17935 1302 17954
rect 1178 17912 1197 17935
rect 547 17872 556 17912
rect 596 17872 1197 17912
rect 1178 17849 1197 17872
rect 1283 17849 1302 17935
rect 1178 17830 1302 17849
rect 6499 17788 6508 17828
rect 6548 17788 11692 17828
rect 11732 17788 11741 17828
rect 2090 17767 2214 17786
rect 2090 17744 2109 17767
rect 1795 17704 1804 17744
rect 1844 17704 2109 17744
rect 2090 17681 2109 17704
rect 2195 17681 2214 17767
rect 13891 17704 13900 17744
rect 13940 17704 14956 17744
rect 14996 17704 15005 17744
rect 2090 17662 2214 17681
rect 1411 17536 1420 17576
rect 1460 17536 8140 17576
rect 8180 17536 8189 17576
rect 4919 17431 5305 17450
rect 4919 17408 4985 17431
rect 5071 17408 5153 17431
rect 5239 17408 5305 17431
rect 4919 17368 4928 17408
rect 4968 17368 4985 17408
rect 5071 17368 5092 17408
rect 5132 17368 5153 17408
rect 5239 17368 5256 17408
rect 5296 17368 5305 17408
rect 4919 17345 4985 17368
rect 5071 17345 5153 17368
rect 5239 17345 5305 17368
rect 4919 17326 5305 17345
rect 20039 17431 20425 17450
rect 20039 17408 20105 17431
rect 20191 17408 20273 17431
rect 20359 17408 20425 17431
rect 20039 17368 20048 17408
rect 20088 17368 20105 17408
rect 20191 17368 20212 17408
rect 20252 17368 20273 17408
rect 20359 17368 20376 17408
rect 20416 17368 20425 17408
rect 20039 17345 20105 17368
rect 20191 17345 20273 17368
rect 20359 17345 20425 17368
rect 20039 17326 20425 17345
rect 1219 16864 1228 16904
rect 1268 16864 15436 16904
rect 15476 16864 15485 16904
rect 3679 16675 4065 16694
rect 3679 16652 3745 16675
rect 3831 16652 3913 16675
rect 3999 16652 4065 16675
rect 3679 16612 3688 16652
rect 3728 16612 3745 16652
rect 3831 16612 3852 16652
rect 3892 16612 3913 16652
rect 3999 16612 4016 16652
rect 4056 16612 4065 16652
rect 3679 16589 3745 16612
rect 3831 16589 3913 16612
rect 3999 16589 4065 16612
rect 3679 16570 4065 16589
rect 18799 16675 19185 16694
rect 18799 16652 18865 16675
rect 18951 16652 19033 16675
rect 19119 16652 19185 16675
rect 18799 16612 18808 16652
rect 18848 16612 18865 16652
rect 18951 16612 18972 16652
rect 19012 16612 19033 16652
rect 19119 16612 19136 16652
rect 19176 16612 19185 16652
rect 18799 16589 18865 16612
rect 18951 16589 19033 16612
rect 19119 16589 19185 16612
rect 18799 16570 19185 16589
rect 931 16360 940 16400
rect 980 16360 17068 16400
rect 17108 16360 17117 16400
rect 9571 16276 9580 16316
rect 9620 16276 12844 16316
rect 12884 16276 12893 16316
rect 13027 16276 13036 16316
rect 13076 16276 15916 16316
rect 15956 16276 15965 16316
rect 4919 15919 5305 15938
rect 4919 15896 4985 15919
rect 5071 15896 5153 15919
rect 5239 15896 5305 15919
rect 20039 15919 20425 15938
rect 20039 15896 20105 15919
rect 20191 15896 20273 15919
rect 20359 15896 20425 15919
rect 4919 15856 4928 15896
rect 4968 15856 4985 15896
rect 5071 15856 5092 15896
rect 5132 15856 5153 15896
rect 5239 15856 5256 15896
rect 5296 15856 5305 15896
rect 13411 15856 13420 15896
rect 13460 15856 16972 15896
rect 17012 15856 17021 15896
rect 20039 15856 20048 15896
rect 20088 15856 20105 15896
rect 20191 15856 20212 15896
rect 20252 15856 20273 15896
rect 20359 15856 20376 15896
rect 20416 15856 20425 15896
rect 722 15835 846 15854
rect 722 15749 741 15835
rect 827 15812 846 15835
rect 4919 15833 4985 15856
rect 5071 15833 5153 15856
rect 5239 15833 5305 15856
rect 4919 15814 5305 15833
rect 20039 15833 20105 15856
rect 20191 15833 20273 15856
rect 20359 15833 20425 15856
rect 20039 15814 20425 15833
rect 827 15772 844 15812
rect 884 15772 893 15812
rect 7555 15772 7564 15812
rect 7604 15772 8620 15812
rect 8660 15772 8669 15812
rect 827 15749 846 15772
rect 722 15730 846 15749
rect 6307 15688 6316 15728
rect 6356 15688 7276 15728
rect 7316 15688 7325 15728
rect 13795 15688 13804 15728
rect 13844 15688 19372 15728
rect 19412 15688 19756 15728
rect 19796 15688 19805 15728
rect 8899 15604 8908 15644
rect 8948 15604 10828 15644
rect 10868 15604 10877 15644
rect 17138 15583 17262 15602
rect 17138 15497 17157 15583
rect 17243 15497 17262 15583
rect 17138 15478 17262 15497
rect 3619 15268 3628 15308
rect 3668 15268 16396 15308
rect 16436 15268 16445 15308
rect 7555 15184 7564 15224
rect 7604 15184 14668 15224
rect 14708 15184 14717 15224
rect 3679 15163 4065 15182
rect 3679 15140 3745 15163
rect 3831 15140 3913 15163
rect 3999 15140 4065 15163
rect 17180 15140 17220 15478
rect 3679 15100 3688 15140
rect 3728 15100 3745 15140
rect 3831 15100 3852 15140
rect 3892 15100 3913 15140
rect 3999 15100 4016 15140
rect 4056 15100 4065 15140
rect 16483 15100 16492 15140
rect 16532 15100 17220 15140
rect 18799 15163 19185 15182
rect 18799 15140 18865 15163
rect 18951 15140 19033 15163
rect 19119 15140 19185 15163
rect 18799 15100 18808 15140
rect 18848 15100 18865 15140
rect 18951 15100 18972 15140
rect 19012 15100 19033 15140
rect 19119 15100 19136 15140
rect 19176 15100 19185 15140
rect 3679 15077 3745 15100
rect 3831 15077 3913 15100
rect 3999 15077 4065 15100
rect 3679 15058 4065 15077
rect 18799 15077 18865 15100
rect 18951 15077 19033 15100
rect 19119 15077 19185 15100
rect 18799 15058 19185 15077
rect 1507 14848 1516 14888
rect 1556 14848 2540 14888
rect 17443 14848 17452 14888
rect 17492 14848 17588 14888
rect 2500 14720 2540 14848
rect 3715 14764 3724 14804
rect 3764 14764 9868 14804
rect 9908 14764 9917 14804
rect 2500 14680 17452 14720
rect 17492 14680 17501 14720
rect 4919 14407 5305 14426
rect 4919 14384 4985 14407
rect 5071 14384 5153 14407
rect 5239 14384 5305 14407
rect 16682 14407 16806 14426
rect 16682 14384 16701 14407
rect 4919 14344 4928 14384
rect 4968 14344 4985 14384
rect 5071 14344 5092 14384
rect 5132 14344 5153 14384
rect 5239 14344 5256 14384
rect 5296 14344 5305 14384
rect 16291 14344 16300 14384
rect 16340 14344 16701 14384
rect 4919 14321 4985 14344
rect 5071 14321 5153 14344
rect 5239 14321 5305 14344
rect 4919 14302 5305 14321
rect 16682 14321 16701 14344
rect 16787 14321 16806 14407
rect 16682 14302 16806 14321
rect 17548 14300 17588 14848
rect 20039 14407 20425 14426
rect 20039 14384 20105 14407
rect 20191 14384 20273 14407
rect 20359 14384 20425 14407
rect 20039 14344 20048 14384
rect 20088 14344 20105 14384
rect 20191 14344 20212 14384
rect 20252 14344 20273 14384
rect 20359 14344 20376 14384
rect 20416 14344 20425 14384
rect 20039 14321 20105 14344
rect 20191 14321 20273 14344
rect 20359 14321 20425 14344
rect 20039 14302 20425 14321
rect 17155 14260 17164 14300
rect 17204 14260 17588 14300
rect 10723 14008 10732 14048
rect 10772 14008 16108 14048
rect 16148 14008 16157 14048
rect 10147 13756 10156 13796
rect 10196 13756 10348 13796
rect 10388 13756 10397 13796
rect 3679 13651 4065 13670
rect 3679 13628 3745 13651
rect 3831 13628 3913 13651
rect 3999 13628 4065 13651
rect 3679 13588 3688 13628
rect 3728 13588 3745 13628
rect 3831 13588 3852 13628
rect 3892 13588 3913 13628
rect 3999 13588 4016 13628
rect 4056 13588 4065 13628
rect 3679 13565 3745 13588
rect 3831 13565 3913 13588
rect 3999 13565 4065 13588
rect 3679 13546 4065 13565
rect 18799 13651 19185 13670
rect 18799 13628 18865 13651
rect 18951 13628 19033 13651
rect 19119 13628 19185 13651
rect 18799 13588 18808 13628
rect 18848 13588 18865 13628
rect 18951 13588 18972 13628
rect 19012 13588 19033 13628
rect 19119 13588 19136 13628
rect 19176 13588 19185 13628
rect 18799 13565 18865 13588
rect 18951 13565 19033 13588
rect 19119 13565 19185 13588
rect 18799 13546 19185 13565
rect 2275 12916 2284 12956
rect 2324 12916 2540 12956
rect 2500 12872 2540 12916
rect 2467 12832 2476 12872
rect 2516 12832 2540 12872
rect 4919 12895 5305 12914
rect 4919 12872 4985 12895
rect 5071 12872 5153 12895
rect 5239 12872 5305 12895
rect 4919 12832 4928 12872
rect 4968 12832 4985 12872
rect 5071 12832 5092 12872
rect 5132 12832 5153 12872
rect 5239 12832 5256 12872
rect 5296 12832 5305 12872
rect 4919 12809 4985 12832
rect 5071 12809 5153 12832
rect 5239 12809 5305 12832
rect 4919 12790 5305 12809
rect 20039 12895 20425 12914
rect 20039 12872 20105 12895
rect 20191 12872 20273 12895
rect 20359 12872 20425 12895
rect 20039 12832 20048 12872
rect 20088 12832 20105 12872
rect 20191 12832 20212 12872
rect 20252 12832 20273 12872
rect 20359 12832 20376 12872
rect 20416 12832 20425 12872
rect 20039 12809 20105 12832
rect 20191 12809 20273 12832
rect 20359 12809 20425 12832
rect 20039 12790 20425 12809
rect 6403 12580 6412 12620
rect 6452 12580 7852 12620
rect 7892 12580 7901 12620
rect 16387 12580 16396 12620
rect 16436 12580 16588 12620
rect 16628 12580 16637 12620
rect 7363 12412 7372 12452
rect 7412 12412 12460 12452
rect 12500 12412 12509 12452
rect 3679 12139 4065 12158
rect 3679 12116 3745 12139
rect 3831 12116 3913 12139
rect 3999 12116 4065 12139
rect 3679 12076 3688 12116
rect 3728 12076 3745 12116
rect 3831 12076 3852 12116
rect 3892 12076 3913 12116
rect 3999 12076 4016 12116
rect 4056 12076 4065 12116
rect 3679 12053 3745 12076
rect 3831 12053 3913 12076
rect 3999 12053 4065 12076
rect 3679 12034 4065 12053
rect 18799 12139 19185 12158
rect 18799 12116 18865 12139
rect 18951 12116 19033 12139
rect 19119 12116 19185 12139
rect 18799 12076 18808 12116
rect 18848 12076 18865 12116
rect 18951 12076 18972 12116
rect 19012 12076 19033 12116
rect 19119 12076 19136 12116
rect 19176 12076 19185 12116
rect 18799 12053 18865 12076
rect 18951 12053 19033 12076
rect 19119 12053 19185 12076
rect 18799 12034 19185 12053
rect 7651 11992 7660 12032
rect 7700 11992 15916 12032
rect 15956 11992 15965 12032
rect 1123 11908 1132 11948
rect 1172 11908 9292 11948
rect 9332 11908 9341 11948
rect 17059 11824 17068 11864
rect 17108 11824 17356 11864
rect 17396 11824 17405 11864
rect 8035 11404 8044 11444
rect 8084 11404 13996 11444
rect 14036 11404 14045 11444
rect 4919 11383 5305 11402
rect 4919 11360 4985 11383
rect 5071 11360 5153 11383
rect 5239 11360 5305 11383
rect 4919 11320 4928 11360
rect 4968 11320 4985 11360
rect 5071 11320 5092 11360
rect 5132 11320 5153 11360
rect 5239 11320 5256 11360
rect 5296 11320 5305 11360
rect 4919 11297 4985 11320
rect 5071 11297 5153 11320
rect 5239 11297 5305 11320
rect 4919 11278 5305 11297
rect 20039 11383 20425 11402
rect 20039 11360 20105 11383
rect 20191 11360 20273 11383
rect 20359 11360 20425 11383
rect 20039 11320 20048 11360
rect 20088 11320 20105 11360
rect 20191 11320 20212 11360
rect 20252 11320 20273 11360
rect 20359 11320 20376 11360
rect 20416 11320 20425 11360
rect 20039 11297 20105 11320
rect 20191 11297 20273 11320
rect 20359 11297 20425 11320
rect 20039 11278 20425 11297
rect 12067 11152 12076 11192
rect 12116 11152 18124 11192
rect 18164 11152 18173 11192
rect 11779 10816 11788 10856
rect 11828 10816 12172 10856
rect 12212 10816 12221 10856
rect 5731 10732 5740 10772
rect 5780 10732 11980 10772
rect 12020 10732 12029 10772
rect 10051 10648 10060 10688
rect 10100 10648 11404 10688
rect 11444 10648 11453 10688
rect 3679 10627 4065 10646
rect 3679 10604 3745 10627
rect 3831 10604 3913 10627
rect 3999 10604 4065 10627
rect 3679 10564 3688 10604
rect 3728 10564 3745 10604
rect 3831 10564 3852 10604
rect 3892 10564 3913 10604
rect 3999 10564 4016 10604
rect 4056 10564 4065 10604
rect 3679 10541 3745 10564
rect 3831 10541 3913 10564
rect 3999 10541 4065 10564
rect 3679 10522 4065 10541
rect 18799 10627 19185 10646
rect 18799 10604 18865 10627
rect 18951 10604 19033 10627
rect 19119 10604 19185 10627
rect 18799 10564 18808 10604
rect 18848 10564 18865 10604
rect 18951 10564 18972 10604
rect 19012 10564 19033 10604
rect 19119 10564 19136 10604
rect 19176 10564 19185 10604
rect 18799 10541 18865 10564
rect 18951 10541 19033 10564
rect 19119 10541 19185 10564
rect 18799 10522 19185 10541
rect 11107 10480 11116 10520
rect 11156 10480 11308 10520
rect 11348 10480 11357 10520
rect 12547 10396 12556 10436
rect 12596 10396 12748 10436
rect 12788 10396 12797 10436
rect 3427 10312 3436 10352
rect 3476 10312 3820 10352
rect 3860 10312 3869 10352
rect 10531 10060 10540 10100
rect 10580 10060 11116 10100
rect 11156 10060 13900 10100
rect 13940 10060 13949 10100
rect 1219 9976 1228 10016
rect 1268 9976 13228 10016
rect 13268 9976 13277 10016
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 11107 9808 11116 9848
rect 11156 9808 13420 9848
rect 13460 9808 16108 9848
rect 16148 9808 16157 9848
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 1891 9724 1900 9764
rect 1940 9724 2284 9764
rect 2324 9724 2333 9764
rect 3139 9640 3148 9680
rect 3188 9640 7564 9680
rect 7604 9640 7613 9680
rect 1411 9472 1420 9512
rect 1460 9472 9580 9512
rect 9620 9472 14188 9512
rect 14228 9472 14237 9512
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 10531 8716 10540 8756
rect 10580 8716 12652 8756
rect 12692 8716 15436 8756
rect 15476 8716 15485 8756
rect 2179 8632 2188 8672
rect 2228 8632 15340 8672
rect 15380 8632 15389 8672
rect 1219 8548 1228 8588
rect 1268 8548 4780 8588
rect 4820 8548 4829 8588
rect 12355 8548 12364 8588
rect 12404 8548 17548 8588
rect 17588 8548 17597 8588
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 9955 8128 9964 8168
rect 10004 8128 19756 8168
rect 19796 8128 19805 8168
rect 10754 7855 10878 7874
rect 10754 7769 10773 7855
rect 10859 7832 10878 7855
rect 10859 7792 11884 7832
rect 11924 7792 11933 7832
rect 10859 7769 10878 7792
rect 10754 7750 10878 7769
rect 16682 7687 16806 7706
rect 16682 7664 16701 7687
rect 12259 7624 12268 7664
rect 12308 7624 16701 7664
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 16682 7601 16701 7624
rect 16787 7601 16806 7687
rect 16682 7582 16806 7601
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 12547 7540 12556 7580
rect 12596 7540 16492 7580
rect 16532 7540 16541 7580
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 4291 7120 4300 7160
rect 4340 7120 4780 7160
rect 4820 7120 14572 7160
rect 14612 7120 14621 7160
rect 3811 6952 3820 6992
rect 3860 6952 20524 6992
rect 20564 6952 20573 6992
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 4099 6448 4108 6488
rect 4148 6448 7564 6488
rect 7604 6448 13900 6488
rect 13940 6448 14092 6488
rect 14132 6448 15052 6488
rect 15092 6448 15101 6488
rect 7651 6280 7660 6320
rect 7700 6280 19468 6320
rect 19508 6280 19517 6320
rect 4675 6196 4684 6236
rect 4724 6196 10252 6236
rect 10292 6196 10301 6236
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 4919 5230 5305 5249
rect 11666 5251 11790 5270
rect 11666 5228 11685 5251
rect 7363 5188 7372 5228
rect 7412 5188 11685 5228
rect 11666 5165 11685 5188
rect 11771 5165 11790 5251
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 11666 5146 11790 5165
rect 9571 5020 9580 5060
rect 9620 5020 13804 5060
rect 13844 5020 13853 5060
rect 7171 4768 7180 4808
rect 7220 4768 13996 4808
rect 14036 4768 20044 4808
rect 20084 4768 20093 4808
rect 4963 4684 4972 4724
rect 5012 4684 7276 4724
rect 7316 4684 20812 4724
rect 20852 4684 20861 4724
rect 4579 4600 4588 4640
rect 4628 4600 9292 4640
rect 9332 4600 9341 4640
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 6691 4516 6700 4556
rect 6740 4516 7276 4556
rect 7316 4516 7325 4556
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 4195 4348 4204 4388
rect 4244 4348 17068 4388
rect 17108 4348 17117 4388
rect 8995 4264 9004 4304
rect 9044 4264 12076 4304
rect 12116 4264 12125 4304
rect 4771 4180 4780 4220
rect 4820 4180 7180 4220
rect 7220 4180 7229 4220
rect 11320 4180 11596 4220
rect 11636 4180 11645 4220
rect 11320 4136 11360 4180
rect 4099 4096 4108 4136
rect 4148 4096 4876 4136
rect 4916 4096 11360 4136
rect 11320 4012 16876 4052
rect 16916 4012 17548 4052
rect 17588 4012 17597 4052
rect 11320 3968 11360 4012
rect 4291 3928 4300 3968
rect 4340 3928 9676 3968
rect 9716 3928 11360 3968
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 1634 3655 1758 3674
rect 1634 3632 1653 3655
rect 1411 3592 1420 3632
rect 1460 3592 1653 3632
rect 1634 3569 1653 3592
rect 1739 3632 1758 3655
rect 1739 3592 6316 3632
rect 6356 3592 6365 3632
rect 1739 3569 1758 3592
rect 1634 3550 1758 3569
rect 11320 3508 19660 3548
rect 19700 3508 19709 3548
rect 11320 3464 11360 3508
rect 10147 3424 10156 3464
rect 10196 3424 11360 3464
rect 16483 3424 16492 3464
rect 16532 3424 17164 3464
rect 17204 3424 17213 3464
rect 9763 3340 9772 3380
rect 9812 3340 18316 3380
rect 18356 3340 20620 3380
rect 20660 3340 20669 3380
rect 14947 3256 14956 3296
rect 14996 3256 15628 3296
rect 15668 3256 15677 3296
rect 2179 3172 2188 3212
rect 2228 3172 12556 3212
rect 12596 3172 12605 3212
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 2659 2668 2668 2708
rect 2708 2668 7564 2708
rect 7604 2668 7613 2708
rect 5635 2584 5644 2624
rect 5684 2584 10060 2624
rect 10100 2584 10109 2624
rect 20131 2500 20140 2540
rect 20180 2500 20220 2540
rect 20140 2456 20180 2500
rect 9379 2416 9388 2456
rect 9428 2416 20180 2456
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 5539 1996 5548 2036
rect 5588 1996 13132 2036
rect 13172 1996 13181 2036
rect 6499 1912 6508 1952
rect 6548 1912 15820 1952
rect 15860 1912 20524 1952
rect 20564 1912 20573 1952
rect 6883 1828 6892 1868
rect 6932 1828 9924 1868
rect 10819 1828 10828 1868
rect 10868 1828 17740 1868
rect 17780 1828 17789 1868
rect 9884 1784 9924 1828
rect 9884 1744 14380 1784
rect 14420 1744 20716 1784
rect 20756 1744 20765 1784
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 3679 1450 4065 1469
rect 9842 1471 9966 1490
rect 9842 1448 9861 1471
rect 4291 1408 4300 1448
rect 4340 1408 9861 1448
rect 9842 1385 9861 1408
rect 9947 1385 9966 1471
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 9842 1366 9966 1385
rect 7106 1303 7230 1322
rect 722 1219 846 1238
rect 722 1133 741 1219
rect 827 1196 846 1219
rect 7106 1217 7125 1303
rect 7211 1280 7230 1303
rect 7220 1240 7230 1280
rect 14755 1240 14764 1280
rect 14804 1240 18700 1280
rect 18740 1240 18749 1280
rect 7211 1217 7230 1240
rect 7106 1198 7230 1217
rect 827 1156 1516 1196
rect 1556 1156 1565 1196
rect 5251 1156 5260 1196
rect 5300 1156 6732 1196
rect 827 1133 846 1156
rect 722 1114 846 1133
rect 6692 1112 6732 1156
rect 6692 1072 12364 1112
rect 12404 1072 12413 1112
rect 8018 883 8142 902
rect 8018 860 8037 883
rect 7939 820 7948 860
rect 7988 820 8037 860
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 8018 797 8037 820
rect 8123 797 8142 883
rect 8018 778 8142 797
rect 13034 883 13158 902
rect 13034 797 13053 883
rect 13139 860 13158 883
rect 13172 820 13181 860
rect 13139 797 13158 820
rect 13034 778 13158 797
rect 20039 799 20425 818
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 4919 694 5305 713
rect 13946 715 14070 734
rect 13946 692 13965 715
rect 13891 652 13900 692
rect 13940 652 13965 692
rect 13946 629 13965 652
rect 14051 629 14070 715
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 13946 610 14070 629
rect 11299 400 11308 440
rect 11348 400 18892 440
rect 18932 400 18941 440
rect 15770 295 15894 314
rect 15770 272 15789 295
rect 15619 232 15628 272
rect 15668 232 15789 272
rect 15770 209 15789 232
rect 15875 209 15894 295
rect 15770 190 15894 209
rect 5059 64 5068 104
rect 5108 64 11692 104
rect 11732 64 11741 104
rect 11875 64 11884 104
rect 11924 64 18124 104
rect 18164 64 18173 104
<< via5 >>
rect 4985 41600 5071 41623
rect 5153 41600 5239 41623
rect 20105 41600 20191 41623
rect 20273 41600 20359 41623
rect 4985 41560 5010 41600
rect 5010 41560 5050 41600
rect 5050 41560 5071 41600
rect 5153 41560 5174 41600
rect 5174 41560 5214 41600
rect 5214 41560 5239 41600
rect 20105 41560 20130 41600
rect 20130 41560 20170 41600
rect 20170 41560 20191 41600
rect 20273 41560 20294 41600
rect 20294 41560 20334 41600
rect 20334 41560 20359 41600
rect 4985 41537 5071 41560
rect 5153 41537 5239 41560
rect 20105 41537 20191 41560
rect 20273 41537 20359 41560
rect 3745 40844 3831 40867
rect 3913 40844 3999 40867
rect 3745 40804 3770 40844
rect 3770 40804 3810 40844
rect 3810 40804 3831 40844
rect 3913 40804 3934 40844
rect 3934 40804 3974 40844
rect 3974 40804 3999 40844
rect 3745 40781 3831 40804
rect 3913 40781 3999 40804
rect 18865 40844 18951 40867
rect 19033 40844 19119 40867
rect 18865 40804 18890 40844
rect 18890 40804 18930 40844
rect 18930 40804 18951 40844
rect 19033 40804 19054 40844
rect 19054 40804 19094 40844
rect 19094 40804 19119 40844
rect 18865 40781 18951 40804
rect 19033 40781 19119 40804
rect 2109 40277 2195 40363
rect 17157 40277 17243 40363
rect 4985 40088 5071 40111
rect 5153 40088 5239 40111
rect 4985 40048 5010 40088
rect 5010 40048 5050 40088
rect 5050 40048 5071 40088
rect 5153 40048 5174 40088
rect 5174 40048 5214 40088
rect 5214 40048 5239 40088
rect 4985 40025 5071 40048
rect 5153 40025 5239 40048
rect 20105 40088 20191 40111
rect 20273 40088 20359 40111
rect 20105 40048 20130 40088
rect 20130 40048 20170 40088
rect 20170 40048 20191 40088
rect 20273 40048 20294 40088
rect 20294 40048 20334 40088
rect 20334 40048 20359 40088
rect 20105 40025 20191 40048
rect 20273 40025 20359 40048
rect 3745 39332 3831 39355
rect 3913 39332 3999 39355
rect 3745 39292 3770 39332
rect 3770 39292 3810 39332
rect 3810 39292 3831 39332
rect 3913 39292 3934 39332
rect 3934 39292 3974 39332
rect 3974 39292 3999 39332
rect 3745 39269 3831 39292
rect 3913 39269 3999 39292
rect 13053 39269 13139 39355
rect 18865 39332 18951 39355
rect 19033 39332 19119 39355
rect 18865 39292 18890 39332
rect 18890 39292 18930 39332
rect 18930 39292 18951 39332
rect 19033 39292 19054 39332
rect 19054 39292 19094 39332
rect 19094 39292 19119 39332
rect 18865 39269 18951 39292
rect 19033 39269 19119 39292
rect 4985 38576 5071 38599
rect 5153 38576 5239 38599
rect 4985 38536 5010 38576
rect 5010 38536 5050 38576
rect 5050 38536 5071 38576
rect 5153 38536 5174 38576
rect 5174 38536 5214 38576
rect 5214 38536 5239 38576
rect 4985 38513 5071 38536
rect 5153 38513 5239 38536
rect 20105 38576 20191 38599
rect 20273 38576 20359 38599
rect 20105 38536 20130 38576
rect 20130 38536 20170 38576
rect 20170 38536 20191 38576
rect 20273 38536 20294 38576
rect 20294 38536 20334 38576
rect 20334 38536 20359 38576
rect 20105 38513 20191 38536
rect 20273 38513 20359 38536
rect 7125 38177 7211 38263
rect 3745 37820 3831 37843
rect 3913 37820 3999 37843
rect 3745 37780 3770 37820
rect 3770 37780 3810 37820
rect 3810 37780 3831 37820
rect 3913 37780 3934 37820
rect 3934 37780 3974 37820
rect 3974 37780 3999 37820
rect 3745 37757 3831 37780
rect 3913 37757 3999 37780
rect 18865 37820 18951 37843
rect 19033 37820 19119 37843
rect 18865 37780 18890 37820
rect 18890 37780 18930 37820
rect 18930 37780 18951 37820
rect 19033 37780 19054 37820
rect 19054 37780 19094 37820
rect 19094 37780 19119 37820
rect 18865 37757 18951 37780
rect 19033 37757 19119 37780
rect 8949 37421 9035 37507
rect 4985 37064 5071 37087
rect 5153 37064 5239 37087
rect 4985 37024 5010 37064
rect 5010 37024 5050 37064
rect 5050 37024 5071 37064
rect 5153 37024 5174 37064
rect 5174 37024 5214 37064
rect 5214 37024 5239 37064
rect 4985 37001 5071 37024
rect 5153 37001 5239 37024
rect 20105 37064 20191 37087
rect 20273 37064 20359 37087
rect 20105 37024 20130 37064
rect 20130 37024 20170 37064
rect 20170 37024 20191 37064
rect 20273 37024 20294 37064
rect 20294 37024 20334 37064
rect 20334 37024 20359 37064
rect 13965 36917 14051 37003
rect 20105 37001 20191 37024
rect 20273 37001 20359 37024
rect 3745 36308 3831 36331
rect 3913 36308 3999 36331
rect 3745 36268 3770 36308
rect 3770 36268 3810 36308
rect 3810 36268 3831 36308
rect 3913 36268 3934 36308
rect 3934 36268 3974 36308
rect 3974 36268 3999 36308
rect 3745 36245 3831 36268
rect 3913 36245 3999 36268
rect 18865 36308 18951 36331
rect 19033 36308 19119 36331
rect 18865 36268 18890 36308
rect 18890 36268 18930 36308
rect 18930 36268 18951 36308
rect 19033 36268 19054 36308
rect 19054 36268 19094 36308
rect 19094 36268 19119 36308
rect 18865 36245 18951 36268
rect 19033 36245 19119 36268
rect 4985 35552 5071 35575
rect 5153 35552 5239 35575
rect 4985 35512 5010 35552
rect 5010 35512 5050 35552
rect 5050 35512 5071 35552
rect 5153 35512 5174 35552
rect 5174 35512 5214 35552
rect 5214 35512 5239 35552
rect 4985 35489 5071 35512
rect 5153 35489 5239 35512
rect 20105 35552 20191 35575
rect 20273 35552 20359 35575
rect 20105 35512 20130 35552
rect 20130 35512 20170 35552
rect 20170 35512 20191 35552
rect 20273 35512 20294 35552
rect 20294 35512 20334 35552
rect 20334 35512 20359 35552
rect 20105 35489 20191 35512
rect 20273 35489 20359 35512
rect 3745 34796 3831 34819
rect 3913 34796 3999 34819
rect 3745 34756 3770 34796
rect 3770 34756 3810 34796
rect 3810 34756 3831 34796
rect 3913 34756 3934 34796
rect 3934 34756 3974 34796
rect 3974 34756 3999 34796
rect 3745 34733 3831 34756
rect 3913 34733 3999 34756
rect 18865 34796 18951 34819
rect 19033 34796 19119 34819
rect 18865 34756 18890 34796
rect 18890 34756 18930 34796
rect 18930 34756 18951 34796
rect 19033 34756 19054 34796
rect 19054 34756 19094 34796
rect 19094 34756 19119 34796
rect 18865 34733 18951 34756
rect 19033 34733 19119 34756
rect 4985 34040 5071 34063
rect 5153 34040 5239 34063
rect 20105 34040 20191 34063
rect 20273 34040 20359 34063
rect 4985 34000 5010 34040
rect 5010 34000 5050 34040
rect 5050 34000 5071 34040
rect 5153 34000 5174 34040
rect 5174 34000 5214 34040
rect 5214 34000 5239 34040
rect 20105 34000 20130 34040
rect 20130 34000 20170 34040
rect 20170 34000 20191 34040
rect 20273 34000 20294 34040
rect 20294 34000 20334 34040
rect 20334 34000 20359 34040
rect 4985 33977 5071 34000
rect 5153 33977 5239 34000
rect 20105 33977 20191 34000
rect 20273 33977 20359 34000
rect 3745 33284 3831 33307
rect 3913 33284 3999 33307
rect 3745 33244 3770 33284
rect 3770 33244 3810 33284
rect 3810 33244 3831 33284
rect 3913 33244 3934 33284
rect 3934 33244 3974 33284
rect 3974 33244 3999 33284
rect 3745 33221 3831 33244
rect 3913 33221 3999 33244
rect 18865 33284 18951 33307
rect 19033 33284 19119 33307
rect 18865 33244 18890 33284
rect 18890 33244 18930 33284
rect 18930 33244 18951 33284
rect 19033 33244 19054 33284
rect 19054 33244 19094 33284
rect 19094 33244 19119 33284
rect 18865 33221 18951 33244
rect 19033 33221 19119 33244
rect 15789 32801 15875 32887
rect 4985 32528 5071 32551
rect 5153 32528 5239 32551
rect 20105 32528 20191 32551
rect 20273 32528 20359 32551
rect 4985 32488 5010 32528
rect 5010 32488 5050 32528
rect 5050 32488 5071 32528
rect 5153 32488 5174 32528
rect 5174 32488 5214 32528
rect 5214 32488 5239 32528
rect 20105 32488 20130 32528
rect 20130 32488 20170 32528
rect 20170 32488 20191 32528
rect 20273 32488 20294 32528
rect 20294 32488 20334 32528
rect 20334 32488 20359 32528
rect 4985 32465 5071 32488
rect 5153 32465 5239 32488
rect 20105 32465 20191 32488
rect 20273 32465 20359 32488
rect 3745 31772 3831 31795
rect 3913 31772 3999 31795
rect 3745 31732 3770 31772
rect 3770 31732 3810 31772
rect 3810 31732 3831 31772
rect 3913 31732 3934 31772
rect 3934 31732 3974 31772
rect 3974 31732 3999 31772
rect 3745 31709 3831 31732
rect 3913 31709 3999 31732
rect 18865 31772 18951 31795
rect 19033 31772 19119 31795
rect 18865 31732 18890 31772
rect 18890 31732 18930 31772
rect 18930 31732 18951 31772
rect 19033 31732 19054 31772
rect 19054 31732 19094 31772
rect 19094 31732 19119 31772
rect 18865 31709 18951 31732
rect 19033 31709 19119 31732
rect 4985 31016 5071 31039
rect 5153 31016 5239 31039
rect 4985 30976 5010 31016
rect 5010 30976 5050 31016
rect 5050 30976 5071 31016
rect 5153 30976 5174 31016
rect 5174 30976 5214 31016
rect 5214 30976 5239 31016
rect 4985 30953 5071 30976
rect 5153 30953 5239 30976
rect 20105 31016 20191 31039
rect 20273 31016 20359 31039
rect 20105 30976 20130 31016
rect 20130 30976 20170 31016
rect 20170 30976 20191 31016
rect 20273 30976 20294 31016
rect 20294 30976 20334 31016
rect 20334 30976 20359 31016
rect 20105 30953 20191 30976
rect 20273 30953 20359 30976
rect 3745 30260 3831 30283
rect 3913 30260 3999 30283
rect 3745 30220 3770 30260
rect 3770 30220 3810 30260
rect 3810 30220 3831 30260
rect 3913 30220 3934 30260
rect 3934 30220 3974 30260
rect 3974 30220 3999 30260
rect 3745 30197 3831 30220
rect 3913 30197 3999 30220
rect 18865 30260 18951 30283
rect 19033 30260 19119 30283
rect 18865 30220 18890 30260
rect 18890 30220 18930 30260
rect 18930 30220 18951 30260
rect 19033 30220 19054 30260
rect 19054 30220 19094 30260
rect 19094 30220 19119 30260
rect 18865 30197 18951 30220
rect 19033 30197 19119 30220
rect 4985 29504 5071 29527
rect 5153 29504 5239 29527
rect 4985 29464 5010 29504
rect 5010 29464 5050 29504
rect 5050 29464 5071 29504
rect 5153 29464 5174 29504
rect 5174 29464 5214 29504
rect 5214 29464 5239 29504
rect 4985 29441 5071 29464
rect 5153 29441 5239 29464
rect 20105 29504 20191 29527
rect 20273 29504 20359 29527
rect 20105 29464 20130 29504
rect 20130 29464 20170 29504
rect 20170 29464 20191 29504
rect 20273 29464 20294 29504
rect 20294 29464 20334 29504
rect 20334 29464 20359 29504
rect 20105 29441 20191 29464
rect 20273 29441 20359 29464
rect 3745 28748 3831 28771
rect 3913 28748 3999 28771
rect 3745 28708 3770 28748
rect 3770 28708 3810 28748
rect 3810 28708 3831 28748
rect 3913 28708 3934 28748
rect 3934 28708 3974 28748
rect 3974 28708 3999 28748
rect 3745 28685 3831 28708
rect 3913 28685 3999 28708
rect 18865 28748 18951 28771
rect 19033 28748 19119 28771
rect 18865 28708 18890 28748
rect 18890 28708 18930 28748
rect 18930 28708 18951 28748
rect 19033 28708 19054 28748
rect 19054 28708 19094 28748
rect 19094 28708 19119 28748
rect 18865 28685 18951 28708
rect 19033 28685 19119 28708
rect 8037 28349 8123 28435
rect 11685 28181 11771 28267
rect 4985 27992 5071 28015
rect 5153 27992 5239 28015
rect 4985 27952 5010 27992
rect 5010 27952 5050 27992
rect 5050 27952 5071 27992
rect 5153 27952 5174 27992
rect 5174 27952 5214 27992
rect 5214 27952 5239 27992
rect 4985 27929 5071 27952
rect 5153 27929 5239 27952
rect 20105 27992 20191 28015
rect 20273 27992 20359 28015
rect 20105 27952 20130 27992
rect 20130 27952 20170 27992
rect 20170 27952 20191 27992
rect 20273 27952 20294 27992
rect 20294 27952 20334 27992
rect 20334 27952 20359 27992
rect 20105 27929 20191 27952
rect 20273 27929 20359 27952
rect 3745 27236 3831 27259
rect 3913 27236 3999 27259
rect 3745 27196 3770 27236
rect 3770 27196 3810 27236
rect 3810 27196 3831 27236
rect 3913 27196 3934 27236
rect 3934 27196 3974 27236
rect 3974 27196 3999 27236
rect 3745 27173 3831 27196
rect 3913 27173 3999 27196
rect 18865 27236 18951 27259
rect 19033 27236 19119 27259
rect 18865 27196 18890 27236
rect 18890 27196 18930 27236
rect 18930 27196 18951 27236
rect 19033 27196 19054 27236
rect 19054 27196 19094 27236
rect 19094 27196 19119 27236
rect 18865 27173 18951 27196
rect 19033 27173 19119 27196
rect 9861 26585 9947 26671
rect 4985 26480 5071 26503
rect 5153 26480 5239 26503
rect 4985 26440 5010 26480
rect 5010 26440 5050 26480
rect 5050 26440 5071 26480
rect 5153 26440 5174 26480
rect 5174 26440 5214 26480
rect 5214 26440 5239 26480
rect 4985 26417 5071 26440
rect 5153 26417 5239 26440
rect 8949 26480 9035 26503
rect 8949 26440 9004 26480
rect 9004 26440 9035 26480
rect 8949 26417 9035 26440
rect 20105 26480 20191 26503
rect 20273 26480 20359 26503
rect 20105 26440 20130 26480
rect 20130 26440 20170 26480
rect 20170 26440 20191 26480
rect 20273 26440 20294 26480
rect 20294 26440 20334 26480
rect 20334 26440 20359 26480
rect 20105 26417 20191 26440
rect 20273 26417 20359 26440
rect 3745 25724 3831 25747
rect 3913 25724 3999 25747
rect 3745 25684 3770 25724
rect 3770 25684 3810 25724
rect 3810 25684 3831 25724
rect 3913 25684 3934 25724
rect 3934 25684 3974 25724
rect 3974 25684 3999 25724
rect 3745 25661 3831 25684
rect 3913 25661 3999 25684
rect 18865 25724 18951 25747
rect 19033 25724 19119 25747
rect 18865 25684 18890 25724
rect 18890 25684 18930 25724
rect 18930 25684 18951 25724
rect 19033 25684 19054 25724
rect 19054 25684 19094 25724
rect 19094 25684 19119 25724
rect 18865 25661 18951 25684
rect 19033 25661 19119 25684
rect 4985 24968 5071 24991
rect 5153 24968 5239 24991
rect 4985 24928 5010 24968
rect 5010 24928 5050 24968
rect 5050 24928 5071 24968
rect 5153 24928 5174 24968
rect 5174 24928 5214 24968
rect 5214 24928 5239 24968
rect 4985 24905 5071 24928
rect 5153 24905 5239 24928
rect 20105 24968 20191 24991
rect 20273 24968 20359 24991
rect 20105 24928 20130 24968
rect 20130 24928 20170 24968
rect 20170 24928 20191 24968
rect 20273 24928 20294 24968
rect 20294 24928 20334 24968
rect 20334 24928 20359 24968
rect 20105 24905 20191 24928
rect 20273 24905 20359 24928
rect 7125 24653 7211 24739
rect 3745 24212 3831 24235
rect 3913 24212 3999 24235
rect 3745 24172 3770 24212
rect 3770 24172 3810 24212
rect 3810 24172 3831 24212
rect 3913 24172 3934 24212
rect 3934 24172 3974 24212
rect 3974 24172 3999 24212
rect 3745 24149 3831 24172
rect 3913 24149 3999 24172
rect 18865 24212 18951 24235
rect 19033 24212 19119 24235
rect 18865 24172 18890 24212
rect 18890 24172 18930 24212
rect 18930 24172 18951 24212
rect 19033 24172 19054 24212
rect 19054 24172 19094 24212
rect 19094 24172 19119 24212
rect 18865 24149 18951 24172
rect 19033 24149 19119 24172
rect 7125 23981 7211 24067
rect 1197 23645 1283 23731
rect 4985 23456 5071 23479
rect 5153 23456 5239 23479
rect 4985 23416 5010 23456
rect 5010 23416 5050 23456
rect 5050 23416 5071 23456
rect 5153 23416 5174 23456
rect 5174 23416 5214 23456
rect 5214 23416 5239 23456
rect 4985 23393 5071 23416
rect 5153 23393 5239 23416
rect 20105 23456 20191 23479
rect 20273 23456 20359 23479
rect 20105 23416 20130 23456
rect 20130 23416 20170 23456
rect 20170 23416 20191 23456
rect 20273 23416 20294 23456
rect 20294 23416 20334 23456
rect 20334 23416 20359 23456
rect 20105 23393 20191 23416
rect 20273 23393 20359 23416
rect 3745 22700 3831 22723
rect 3913 22700 3999 22723
rect 18865 22700 18951 22723
rect 19033 22700 19119 22723
rect 3745 22660 3770 22700
rect 3770 22660 3810 22700
rect 3810 22660 3831 22700
rect 3913 22660 3934 22700
rect 3934 22660 3974 22700
rect 3974 22660 3999 22700
rect 18865 22660 18890 22700
rect 18890 22660 18930 22700
rect 18930 22660 18951 22700
rect 19033 22660 19054 22700
rect 19054 22660 19094 22700
rect 19094 22660 19119 22700
rect 3745 22637 3831 22660
rect 3913 22637 3999 22660
rect 18865 22637 18951 22660
rect 19033 22637 19119 22660
rect 4985 21944 5071 21967
rect 5153 21944 5239 21967
rect 4985 21904 5010 21944
rect 5010 21904 5050 21944
rect 5050 21904 5071 21944
rect 5153 21904 5174 21944
rect 5174 21904 5214 21944
rect 5214 21904 5239 21944
rect 4985 21881 5071 21904
rect 5153 21881 5239 21904
rect 20105 21944 20191 21967
rect 20273 21944 20359 21967
rect 20105 21904 20130 21944
rect 20130 21904 20170 21944
rect 20170 21904 20191 21944
rect 20273 21904 20294 21944
rect 20294 21904 20334 21944
rect 20334 21904 20359 21944
rect 20105 21881 20191 21904
rect 20273 21881 20359 21904
rect 2109 21713 2195 21799
rect 3745 21188 3831 21211
rect 3913 21188 3999 21211
rect 3745 21148 3770 21188
rect 3770 21148 3810 21188
rect 3810 21148 3831 21188
rect 3913 21148 3934 21188
rect 3934 21148 3974 21188
rect 3974 21148 3999 21188
rect 3745 21125 3831 21148
rect 3913 21125 3999 21148
rect 18865 21188 18951 21211
rect 19033 21188 19119 21211
rect 18865 21148 18890 21188
rect 18890 21148 18930 21188
rect 18930 21148 18951 21188
rect 19033 21148 19054 21188
rect 19054 21148 19094 21188
rect 19094 21148 19119 21188
rect 18865 21125 18951 21148
rect 19033 21125 19119 21148
rect 4985 20432 5071 20455
rect 5153 20432 5239 20455
rect 4985 20392 5010 20432
rect 5010 20392 5050 20432
rect 5050 20392 5071 20432
rect 5153 20392 5174 20432
rect 5174 20392 5214 20432
rect 5214 20392 5239 20432
rect 4985 20369 5071 20392
rect 5153 20369 5239 20392
rect 20105 20432 20191 20455
rect 20273 20432 20359 20455
rect 20105 20392 20130 20432
rect 20130 20392 20170 20432
rect 20170 20392 20191 20432
rect 20273 20392 20294 20432
rect 20294 20392 20334 20432
rect 20334 20392 20359 20432
rect 20105 20369 20191 20392
rect 20273 20369 20359 20392
rect 3745 19676 3831 19699
rect 3913 19676 3999 19699
rect 3745 19636 3770 19676
rect 3770 19636 3810 19676
rect 3810 19636 3831 19676
rect 3913 19636 3934 19676
rect 3934 19636 3974 19676
rect 3974 19636 3999 19676
rect 3745 19613 3831 19636
rect 3913 19613 3999 19636
rect 18865 19676 18951 19699
rect 19033 19676 19119 19699
rect 18865 19636 18890 19676
rect 18890 19636 18930 19676
rect 18930 19636 18951 19676
rect 19033 19636 19054 19676
rect 19054 19636 19094 19676
rect 19094 19636 19119 19676
rect 18865 19613 18951 19636
rect 19033 19613 19119 19636
rect 10773 19025 10859 19111
rect 4985 18920 5071 18943
rect 5153 18920 5239 18943
rect 20105 18920 20191 18943
rect 20273 18920 20359 18943
rect 4985 18880 5010 18920
rect 5010 18880 5050 18920
rect 5050 18880 5071 18920
rect 5153 18880 5174 18920
rect 5174 18880 5214 18920
rect 5214 18880 5239 18920
rect 20105 18880 20130 18920
rect 20130 18880 20170 18920
rect 20170 18880 20191 18920
rect 20273 18880 20294 18920
rect 20294 18880 20334 18920
rect 20334 18880 20359 18920
rect 4985 18857 5071 18880
rect 5153 18857 5239 18880
rect 20105 18857 20191 18880
rect 20273 18857 20359 18880
rect 3745 18164 3831 18187
rect 3913 18164 3999 18187
rect 3745 18124 3770 18164
rect 3770 18124 3810 18164
rect 3810 18124 3831 18164
rect 3913 18124 3934 18164
rect 3934 18124 3974 18164
rect 3974 18124 3999 18164
rect 3745 18101 3831 18124
rect 3913 18101 3999 18124
rect 18865 18164 18951 18187
rect 19033 18164 19119 18187
rect 18865 18124 18890 18164
rect 18890 18124 18930 18164
rect 18930 18124 18951 18164
rect 19033 18124 19054 18164
rect 19054 18124 19094 18164
rect 19094 18124 19119 18164
rect 18865 18101 18951 18124
rect 19033 18101 19119 18124
rect 1197 17849 1283 17935
rect 2109 17681 2195 17767
rect 4985 17408 5071 17431
rect 5153 17408 5239 17431
rect 4985 17368 5010 17408
rect 5010 17368 5050 17408
rect 5050 17368 5071 17408
rect 5153 17368 5174 17408
rect 5174 17368 5214 17408
rect 5214 17368 5239 17408
rect 4985 17345 5071 17368
rect 5153 17345 5239 17368
rect 20105 17408 20191 17431
rect 20273 17408 20359 17431
rect 20105 17368 20130 17408
rect 20130 17368 20170 17408
rect 20170 17368 20191 17408
rect 20273 17368 20294 17408
rect 20294 17368 20334 17408
rect 20334 17368 20359 17408
rect 20105 17345 20191 17368
rect 20273 17345 20359 17368
rect 3745 16652 3831 16675
rect 3913 16652 3999 16675
rect 3745 16612 3770 16652
rect 3770 16612 3810 16652
rect 3810 16612 3831 16652
rect 3913 16612 3934 16652
rect 3934 16612 3974 16652
rect 3974 16612 3999 16652
rect 3745 16589 3831 16612
rect 3913 16589 3999 16612
rect 18865 16652 18951 16675
rect 19033 16652 19119 16675
rect 18865 16612 18890 16652
rect 18890 16612 18930 16652
rect 18930 16612 18951 16652
rect 19033 16612 19054 16652
rect 19054 16612 19094 16652
rect 19094 16612 19119 16652
rect 18865 16589 18951 16612
rect 19033 16589 19119 16612
rect 4985 15896 5071 15919
rect 5153 15896 5239 15919
rect 20105 15896 20191 15919
rect 20273 15896 20359 15919
rect 4985 15856 5010 15896
rect 5010 15856 5050 15896
rect 5050 15856 5071 15896
rect 5153 15856 5174 15896
rect 5174 15856 5214 15896
rect 5214 15856 5239 15896
rect 20105 15856 20130 15896
rect 20130 15856 20170 15896
rect 20170 15856 20191 15896
rect 20273 15856 20294 15896
rect 20294 15856 20334 15896
rect 20334 15856 20359 15896
rect 741 15749 827 15835
rect 4985 15833 5071 15856
rect 5153 15833 5239 15856
rect 20105 15833 20191 15856
rect 20273 15833 20359 15856
rect 17157 15497 17243 15583
rect 3745 15140 3831 15163
rect 3913 15140 3999 15163
rect 3745 15100 3770 15140
rect 3770 15100 3810 15140
rect 3810 15100 3831 15140
rect 3913 15100 3934 15140
rect 3934 15100 3974 15140
rect 3974 15100 3999 15140
rect 18865 15140 18951 15163
rect 19033 15140 19119 15163
rect 18865 15100 18890 15140
rect 18890 15100 18930 15140
rect 18930 15100 18951 15140
rect 19033 15100 19054 15140
rect 19054 15100 19094 15140
rect 19094 15100 19119 15140
rect 3745 15077 3831 15100
rect 3913 15077 3999 15100
rect 18865 15077 18951 15100
rect 19033 15077 19119 15100
rect 4985 14384 5071 14407
rect 5153 14384 5239 14407
rect 4985 14344 5010 14384
rect 5010 14344 5050 14384
rect 5050 14344 5071 14384
rect 5153 14344 5174 14384
rect 5174 14344 5214 14384
rect 5214 14344 5239 14384
rect 4985 14321 5071 14344
rect 5153 14321 5239 14344
rect 16701 14321 16787 14407
rect 20105 14384 20191 14407
rect 20273 14384 20359 14407
rect 20105 14344 20130 14384
rect 20130 14344 20170 14384
rect 20170 14344 20191 14384
rect 20273 14344 20294 14384
rect 20294 14344 20334 14384
rect 20334 14344 20359 14384
rect 20105 14321 20191 14344
rect 20273 14321 20359 14344
rect 3745 13628 3831 13651
rect 3913 13628 3999 13651
rect 3745 13588 3770 13628
rect 3770 13588 3810 13628
rect 3810 13588 3831 13628
rect 3913 13588 3934 13628
rect 3934 13588 3974 13628
rect 3974 13588 3999 13628
rect 3745 13565 3831 13588
rect 3913 13565 3999 13588
rect 18865 13628 18951 13651
rect 19033 13628 19119 13651
rect 18865 13588 18890 13628
rect 18890 13588 18930 13628
rect 18930 13588 18951 13628
rect 19033 13588 19054 13628
rect 19054 13588 19094 13628
rect 19094 13588 19119 13628
rect 18865 13565 18951 13588
rect 19033 13565 19119 13588
rect 4985 12872 5071 12895
rect 5153 12872 5239 12895
rect 4985 12832 5010 12872
rect 5010 12832 5050 12872
rect 5050 12832 5071 12872
rect 5153 12832 5174 12872
rect 5174 12832 5214 12872
rect 5214 12832 5239 12872
rect 4985 12809 5071 12832
rect 5153 12809 5239 12832
rect 20105 12872 20191 12895
rect 20273 12872 20359 12895
rect 20105 12832 20130 12872
rect 20130 12832 20170 12872
rect 20170 12832 20191 12872
rect 20273 12832 20294 12872
rect 20294 12832 20334 12872
rect 20334 12832 20359 12872
rect 20105 12809 20191 12832
rect 20273 12809 20359 12832
rect 3745 12116 3831 12139
rect 3913 12116 3999 12139
rect 3745 12076 3770 12116
rect 3770 12076 3810 12116
rect 3810 12076 3831 12116
rect 3913 12076 3934 12116
rect 3934 12076 3974 12116
rect 3974 12076 3999 12116
rect 3745 12053 3831 12076
rect 3913 12053 3999 12076
rect 18865 12116 18951 12139
rect 19033 12116 19119 12139
rect 18865 12076 18890 12116
rect 18890 12076 18930 12116
rect 18930 12076 18951 12116
rect 19033 12076 19054 12116
rect 19054 12076 19094 12116
rect 19094 12076 19119 12116
rect 18865 12053 18951 12076
rect 19033 12053 19119 12076
rect 4985 11360 5071 11383
rect 5153 11360 5239 11383
rect 4985 11320 5010 11360
rect 5010 11320 5050 11360
rect 5050 11320 5071 11360
rect 5153 11320 5174 11360
rect 5174 11320 5214 11360
rect 5214 11320 5239 11360
rect 4985 11297 5071 11320
rect 5153 11297 5239 11320
rect 20105 11360 20191 11383
rect 20273 11360 20359 11383
rect 20105 11320 20130 11360
rect 20130 11320 20170 11360
rect 20170 11320 20191 11360
rect 20273 11320 20294 11360
rect 20294 11320 20334 11360
rect 20334 11320 20359 11360
rect 20105 11297 20191 11320
rect 20273 11297 20359 11320
rect 3745 10604 3831 10627
rect 3913 10604 3999 10627
rect 3745 10564 3770 10604
rect 3770 10564 3810 10604
rect 3810 10564 3831 10604
rect 3913 10564 3934 10604
rect 3934 10564 3974 10604
rect 3974 10564 3999 10604
rect 3745 10541 3831 10564
rect 3913 10541 3999 10564
rect 18865 10604 18951 10627
rect 19033 10604 19119 10627
rect 18865 10564 18890 10604
rect 18890 10564 18930 10604
rect 18930 10564 18951 10604
rect 19033 10564 19054 10604
rect 19054 10564 19094 10604
rect 19094 10564 19119 10604
rect 18865 10541 18951 10564
rect 19033 10541 19119 10564
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 10773 7769 10859 7855
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 16701 7601 16787 7687
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 11685 5165 11771 5251
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 1653 3569 1739 3655
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 9861 1385 9947 1471
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 741 1133 827 1219
rect 7125 1280 7211 1303
rect 7125 1240 7180 1280
rect 7180 1240 7211 1280
rect 7125 1217 7211 1240
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 8037 797 8123 883
rect 13053 860 13139 883
rect 13053 820 13132 860
rect 13132 820 13139 860
rect 13053 797 13139 820
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 13965 629 14051 715
rect 20105 713 20191 736
rect 20273 713 20359 736
rect 15789 209 15875 295
<< metal6 >>
rect 3652 40867 4092 43008
rect 3652 40781 3745 40867
rect 3831 40781 3913 40867
rect 3999 40781 4092 40867
rect 1988 40363 2316 40484
rect 1988 40277 2109 40363
rect 2195 40277 2316 40363
rect 1076 23731 1404 23852
rect 1076 23645 1197 23731
rect 1283 23645 1404 23731
rect 1076 17935 1404 23645
rect 1988 21799 2316 40277
rect 1988 21713 2109 21799
rect 2195 21713 2316 21799
rect 1988 21592 2316 21713
rect 3652 39355 4092 40781
rect 3652 39269 3745 39355
rect 3831 39269 3913 39355
rect 3999 39269 4092 39355
rect 3652 37843 4092 39269
rect 3652 37757 3745 37843
rect 3831 37757 3913 37843
rect 3999 37757 4092 37843
rect 3652 36331 4092 37757
rect 3652 36245 3745 36331
rect 3831 36245 3913 36331
rect 3999 36245 4092 36331
rect 3652 34819 4092 36245
rect 3652 34733 3745 34819
rect 3831 34733 3913 34819
rect 3999 34733 4092 34819
rect 3652 33307 4092 34733
rect 3652 33221 3745 33307
rect 3831 33221 3913 33307
rect 3999 33221 4092 33307
rect 3652 31795 4092 33221
rect 3652 31709 3745 31795
rect 3831 31709 3913 31795
rect 3999 31709 4092 31795
rect 3652 30283 4092 31709
rect 3652 30197 3745 30283
rect 3831 30197 3913 30283
rect 3999 30197 4092 30283
rect 3652 28771 4092 30197
rect 3652 28685 3745 28771
rect 3831 28685 3913 28771
rect 3999 28685 4092 28771
rect 3652 27259 4092 28685
rect 3652 27173 3745 27259
rect 3831 27173 3913 27259
rect 3999 27173 4092 27259
rect 3652 25747 4092 27173
rect 3652 25661 3745 25747
rect 3831 25661 3913 25747
rect 3999 25661 4092 25747
rect 3652 24235 4092 25661
rect 3652 24149 3745 24235
rect 3831 24149 3913 24235
rect 3999 24149 4092 24235
rect 3652 22723 4092 24149
rect 3652 22637 3745 22723
rect 3831 22637 3913 22723
rect 3999 22637 4092 22723
rect 1076 17849 1197 17935
rect 1283 17849 1404 17935
rect 3652 21211 4092 22637
rect 3652 21125 3745 21211
rect 3831 21125 3913 21211
rect 3999 21125 4092 21211
rect 3652 19699 4092 21125
rect 3652 19613 3745 19699
rect 3831 19613 3913 19699
rect 3999 19613 4092 19699
rect 3652 18187 4092 19613
rect 3652 18101 3745 18187
rect 3831 18101 3913 18187
rect 3999 18101 4092 18187
rect 1076 17728 1404 17849
rect 1988 17767 2316 17888
rect 1988 17681 2109 17767
rect 2195 17681 2316 17767
rect 1988 17364 2316 17681
rect 1532 17036 2316 17364
rect 620 15835 948 15956
rect 620 15749 741 15835
rect 827 15749 948 15835
rect 620 1219 948 15749
rect 1532 3655 1860 17036
rect 1532 3569 1653 3655
rect 1739 3569 1860 3655
rect 1532 3448 1860 3569
rect 3652 16675 4092 18101
rect 3652 16589 3745 16675
rect 3831 16589 3913 16675
rect 3999 16589 4092 16675
rect 3652 15163 4092 16589
rect 3652 15077 3745 15163
rect 3831 15077 3913 15163
rect 3999 15077 4092 15163
rect 3652 13651 4092 15077
rect 3652 13565 3745 13651
rect 3831 13565 3913 13651
rect 3999 13565 4092 13651
rect 3652 12139 4092 13565
rect 3652 12053 3745 12139
rect 3831 12053 3913 12139
rect 3999 12053 4092 12139
rect 3652 10627 4092 12053
rect 3652 10541 3745 10627
rect 3831 10541 3913 10627
rect 3999 10541 4092 10627
rect 3652 9115 4092 10541
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 620 1133 741 1219
rect 827 1133 948 1219
rect 620 1012 948 1133
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 41623 5332 43008
rect 4892 41537 4985 41623
rect 5071 41537 5153 41623
rect 5239 41537 5332 41623
rect 4892 40111 5332 41537
rect 18772 40867 19212 43008
rect 18772 40781 18865 40867
rect 18951 40781 19033 40867
rect 19119 40781 19212 40867
rect 4892 40025 4985 40111
rect 5071 40025 5153 40111
rect 5239 40025 5332 40111
rect 4892 38599 5332 40025
rect 17036 40363 17364 40484
rect 17036 40277 17157 40363
rect 17243 40277 17364 40363
rect 4892 38513 4985 38599
rect 5071 38513 5153 38599
rect 5239 38513 5332 38599
rect 4892 37087 5332 38513
rect 12932 39355 13260 39476
rect 12932 39269 13053 39355
rect 13139 39269 13260 39355
rect 4892 37001 4985 37087
rect 5071 37001 5153 37087
rect 5239 37001 5332 37087
rect 4892 35575 5332 37001
rect 4892 35489 4985 35575
rect 5071 35489 5153 35575
rect 5239 35489 5332 35575
rect 4892 34063 5332 35489
rect 4892 33977 4985 34063
rect 5071 33977 5153 34063
rect 5239 33977 5332 34063
rect 4892 32551 5332 33977
rect 4892 32465 4985 32551
rect 5071 32465 5153 32551
rect 5239 32465 5332 32551
rect 4892 31039 5332 32465
rect 4892 30953 4985 31039
rect 5071 30953 5153 31039
rect 5239 30953 5332 31039
rect 4892 29527 5332 30953
rect 4892 29441 4985 29527
rect 5071 29441 5153 29527
rect 5239 29441 5332 29527
rect 4892 28015 5332 29441
rect 4892 27929 4985 28015
rect 5071 27929 5153 28015
rect 5239 27929 5332 28015
rect 4892 26503 5332 27929
rect 4892 26417 4985 26503
rect 5071 26417 5153 26503
rect 5239 26417 5332 26503
rect 4892 24991 5332 26417
rect 4892 24905 4985 24991
rect 5071 24905 5153 24991
rect 5239 24905 5332 24991
rect 4892 23479 5332 24905
rect 7004 38263 7332 38384
rect 7004 38177 7125 38263
rect 7211 38177 7332 38263
rect 7004 24739 7332 38177
rect 8828 37507 9156 37628
rect 8828 37421 8949 37507
rect 9035 37421 9156 37507
rect 7004 24653 7125 24739
rect 7211 24653 7332 24739
rect 7004 24532 7332 24653
rect 7916 28435 8244 28556
rect 7916 28349 8037 28435
rect 8123 28349 8244 28435
rect 4892 23393 4985 23479
rect 5071 23393 5153 23479
rect 5239 23393 5332 23479
rect 4892 21967 5332 23393
rect 4892 21881 4985 21967
rect 5071 21881 5153 21967
rect 5239 21881 5332 21967
rect 4892 20455 5332 21881
rect 4892 20369 4985 20455
rect 5071 20369 5153 20455
rect 5239 20369 5332 20455
rect 4892 18943 5332 20369
rect 4892 18857 4985 18943
rect 5071 18857 5153 18943
rect 5239 18857 5332 18943
rect 4892 17431 5332 18857
rect 4892 17345 4985 17431
rect 5071 17345 5153 17431
rect 5239 17345 5332 17431
rect 4892 15919 5332 17345
rect 4892 15833 4985 15919
rect 5071 15833 5153 15919
rect 5239 15833 5332 15919
rect 4892 14407 5332 15833
rect 4892 14321 4985 14407
rect 5071 14321 5153 14407
rect 5239 14321 5332 14407
rect 4892 12895 5332 14321
rect 4892 12809 4985 12895
rect 5071 12809 5153 12895
rect 5239 12809 5332 12895
rect 4892 11383 5332 12809
rect 4892 11297 4985 11383
rect 5071 11297 5153 11383
rect 5239 11297 5332 11383
rect 4892 9871 5332 11297
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 7004 24067 7332 24188
rect 7004 23981 7125 24067
rect 7211 23981 7332 24067
rect 7004 1303 7332 23981
rect 7004 1217 7125 1303
rect 7211 1217 7332 1303
rect 7004 1096 7332 1217
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 7916 883 8244 28349
rect 8828 26503 9156 37421
rect 11564 28267 11892 28388
rect 11564 28181 11685 28267
rect 11771 28181 11892 28267
rect 8828 26417 8949 26503
rect 9035 26417 9156 26503
rect 8828 26296 9156 26417
rect 9740 26671 10068 26792
rect 9740 26585 9861 26671
rect 9947 26585 10068 26671
rect 9740 1471 10068 26585
rect 10652 19111 10980 19232
rect 10652 19025 10773 19111
rect 10859 19025 10980 19111
rect 10652 7855 10980 19025
rect 10652 7769 10773 7855
rect 10859 7769 10980 7855
rect 10652 7648 10980 7769
rect 11564 5251 11892 28181
rect 11564 5165 11685 5251
rect 11771 5165 11892 5251
rect 11564 5044 11892 5165
rect 9740 1385 9861 1471
rect 9947 1385 10068 1471
rect 9740 1264 10068 1385
rect 7916 797 8037 883
rect 8123 797 8244 883
rect 7916 676 8244 797
rect 12932 883 13260 39269
rect 12932 797 13053 883
rect 13139 797 13260 883
rect 12932 676 13260 797
rect 13844 37003 14172 37124
rect 13844 36917 13965 37003
rect 14051 36917 14172 37003
rect 13844 715 14172 36917
rect 13844 629 13965 715
rect 14051 629 14172 715
rect 13844 508 14172 629
rect 15668 32887 15996 33008
rect 15668 32801 15789 32887
rect 15875 32801 15996 32887
rect 15668 295 15996 32801
rect 17036 15583 17364 40277
rect 17036 15497 17157 15583
rect 17243 15497 17364 15583
rect 17036 15376 17364 15497
rect 18772 39355 19212 40781
rect 18772 39269 18865 39355
rect 18951 39269 19033 39355
rect 19119 39269 19212 39355
rect 18772 37843 19212 39269
rect 18772 37757 18865 37843
rect 18951 37757 19033 37843
rect 19119 37757 19212 37843
rect 18772 36331 19212 37757
rect 18772 36245 18865 36331
rect 18951 36245 19033 36331
rect 19119 36245 19212 36331
rect 18772 34819 19212 36245
rect 18772 34733 18865 34819
rect 18951 34733 19033 34819
rect 19119 34733 19212 34819
rect 18772 33307 19212 34733
rect 18772 33221 18865 33307
rect 18951 33221 19033 33307
rect 19119 33221 19212 33307
rect 18772 31795 19212 33221
rect 18772 31709 18865 31795
rect 18951 31709 19033 31795
rect 19119 31709 19212 31795
rect 18772 30283 19212 31709
rect 18772 30197 18865 30283
rect 18951 30197 19033 30283
rect 19119 30197 19212 30283
rect 18772 28771 19212 30197
rect 18772 28685 18865 28771
rect 18951 28685 19033 28771
rect 19119 28685 19212 28771
rect 18772 27259 19212 28685
rect 18772 27173 18865 27259
rect 18951 27173 19033 27259
rect 19119 27173 19212 27259
rect 18772 25747 19212 27173
rect 18772 25661 18865 25747
rect 18951 25661 19033 25747
rect 19119 25661 19212 25747
rect 18772 24235 19212 25661
rect 18772 24149 18865 24235
rect 18951 24149 19033 24235
rect 19119 24149 19212 24235
rect 18772 22723 19212 24149
rect 18772 22637 18865 22723
rect 18951 22637 19033 22723
rect 19119 22637 19212 22723
rect 18772 21211 19212 22637
rect 18772 21125 18865 21211
rect 18951 21125 19033 21211
rect 19119 21125 19212 21211
rect 18772 19699 19212 21125
rect 18772 19613 18865 19699
rect 18951 19613 19033 19699
rect 19119 19613 19212 19699
rect 18772 18187 19212 19613
rect 18772 18101 18865 18187
rect 18951 18101 19033 18187
rect 19119 18101 19212 18187
rect 18772 16675 19212 18101
rect 18772 16589 18865 16675
rect 18951 16589 19033 16675
rect 19119 16589 19212 16675
rect 18772 15163 19212 16589
rect 18772 15077 18865 15163
rect 18951 15077 19033 15163
rect 19119 15077 19212 15163
rect 16580 14407 16908 14528
rect 16580 14321 16701 14407
rect 16787 14321 16908 14407
rect 16580 7687 16908 14321
rect 16580 7601 16701 7687
rect 16787 7601 16908 7687
rect 16580 7480 16908 7601
rect 18772 13651 19212 15077
rect 18772 13565 18865 13651
rect 18951 13565 19033 13651
rect 19119 13565 19212 13651
rect 18772 12139 19212 13565
rect 18772 12053 18865 12139
rect 18951 12053 19033 12139
rect 19119 12053 19212 12139
rect 18772 10627 19212 12053
rect 18772 10541 18865 10627
rect 18951 10541 19033 10627
rect 19119 10541 19212 10627
rect 18772 9115 19212 10541
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 15668 209 15789 295
rect 15875 209 15996 295
rect 15668 88 15996 209
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 41623 20452 43008
rect 20012 41537 20105 41623
rect 20191 41537 20273 41623
rect 20359 41537 20452 41623
rect 20012 40111 20452 41537
rect 20012 40025 20105 40111
rect 20191 40025 20273 40111
rect 20359 40025 20452 40111
rect 20012 38599 20452 40025
rect 20012 38513 20105 38599
rect 20191 38513 20273 38599
rect 20359 38513 20452 38599
rect 20012 37087 20452 38513
rect 20012 37001 20105 37087
rect 20191 37001 20273 37087
rect 20359 37001 20452 37087
rect 20012 35575 20452 37001
rect 20012 35489 20105 35575
rect 20191 35489 20273 35575
rect 20359 35489 20452 35575
rect 20012 34063 20452 35489
rect 20012 33977 20105 34063
rect 20191 33977 20273 34063
rect 20359 33977 20452 34063
rect 20012 32551 20452 33977
rect 20012 32465 20105 32551
rect 20191 32465 20273 32551
rect 20359 32465 20452 32551
rect 20012 31039 20452 32465
rect 20012 30953 20105 31039
rect 20191 30953 20273 31039
rect 20359 30953 20452 31039
rect 20012 29527 20452 30953
rect 20012 29441 20105 29527
rect 20191 29441 20273 29527
rect 20359 29441 20452 29527
rect 20012 28015 20452 29441
rect 20012 27929 20105 28015
rect 20191 27929 20273 28015
rect 20359 27929 20452 28015
rect 20012 26503 20452 27929
rect 20012 26417 20105 26503
rect 20191 26417 20273 26503
rect 20359 26417 20452 26503
rect 20012 24991 20452 26417
rect 20012 24905 20105 24991
rect 20191 24905 20273 24991
rect 20359 24905 20452 24991
rect 20012 23479 20452 24905
rect 20012 23393 20105 23479
rect 20191 23393 20273 23479
rect 20359 23393 20452 23479
rect 20012 21967 20452 23393
rect 20012 21881 20105 21967
rect 20191 21881 20273 21967
rect 20359 21881 20452 21967
rect 20012 20455 20452 21881
rect 20012 20369 20105 20455
rect 20191 20369 20273 20455
rect 20359 20369 20452 20455
rect 20012 18943 20452 20369
rect 20012 18857 20105 18943
rect 20191 18857 20273 18943
rect 20359 18857 20452 18943
rect 20012 17431 20452 18857
rect 20012 17345 20105 17431
rect 20191 17345 20273 17431
rect 20359 17345 20452 17431
rect 20012 15919 20452 17345
rect 20012 15833 20105 15919
rect 20191 15833 20273 15919
rect 20359 15833 20452 15919
rect 20012 14407 20452 15833
rect 20012 14321 20105 14407
rect 20191 14321 20273 14407
rect 20359 14321 20452 14407
rect 20012 12895 20452 14321
rect 20012 12809 20105 12895
rect 20191 12809 20273 12895
rect 20359 12809 20452 12895
rect 20012 11383 20452 12809
rect 20012 11297 20105 11383
rect 20191 11297 20273 11383
rect 20359 11297 20452 11383
rect 20012 9871 20452 11297
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_inv_1  _0381_
timestamp 1676382929
transform -1 0 8832 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _0382_
timestamp 1676382929
transform 1 0 15168 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0383_
timestamp 1676382929
transform -1 0 5664 0 -1 14364
box -48 -56 336 834
use sg13g2_inv_1  _0384_
timestamp 1676382929
transform 1 0 15744 0 -1 5292
box -48 -56 336 834
use sg13g2_inv_1  _0385_
timestamp 1676382929
transform -1 0 20352 0 1 40068
box -48 -56 336 834
use sg13g2_inv_1  _0386_
timestamp 1676382929
transform -1 0 1440 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0387_
timestamp 1676382929
transform 1 0 20064 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0388_
timestamp 1676382929
transform -1 0 1440 0 1 34020
box -48 -56 336 834
use sg13g2_inv_1  _0389_
timestamp 1676382929
transform 1 0 20064 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0390_
timestamp 1676382929
transform -1 0 8352 0 -1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0391_
timestamp 1676382929
transform -1 0 14976 0 -1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0392_
timestamp 1676382929
transform 1 0 20064 0 -1 2268
box -48 -56 336 834
use sg13g2_inv_1  _0393_
timestamp 1676382929
transform 1 0 20064 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _0394_
timestamp 1676382929
transform 1 0 12960 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0395_
timestamp 1676382929
transform -1 0 11328 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  _0396_
timestamp 1676382929
transform 1 0 19392 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0397_
timestamp 1676382929
transform -1 0 17376 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0398_
timestamp 1676382929
transform 1 0 17952 0 1 8316
box -48 -56 336 834
use sg13g2_inv_1  _0399_
timestamp 1676382929
transform -1 0 11904 0 1 6804
box -48 -56 336 834
use sg13g2_inv_1  _0400_
timestamp 1676382929
transform 1 0 17376 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0401_
timestamp 1676382929
transform 1 0 13152 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  _0402_
timestamp 1676382929
transform 1 0 12768 0 1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0403_
timestamp 1676382929
transform 1 0 2880 0 -1 12852
box -48 -56 336 834
use sg13g2_inv_1  _0404_
timestamp 1676382929
transform 1 0 9600 0 1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0405_
timestamp 1676382929
transform -1 0 12576 0 -1 24948
box -48 -56 336 834
use sg13g2_inv_1  _0406_
timestamp 1676382929
transform 1 0 4128 0 1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0407_
timestamp 1676382929
transform -1 0 9312 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0408_
timestamp 1676382929
transform -1 0 1440 0 1 11340
box -48 -56 336 834
use sg13g2_inv_1  _0409_
timestamp 1676382929
transform -1 0 9120 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _0410_
timestamp 1676382929
transform 1 0 6624 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _0411_
timestamp 1676382929
transform 1 0 11040 0 -1 15876
box -48 -56 336 834
use sg13g2_inv_1  _0412_
timestamp 1676382929
transform -1 0 7200 0 1 3780
box -48 -56 336 834
use sg13g2_inv_1  _0413_
timestamp 1676382929
transform 1 0 18720 0 1 38556
box -48 -56 336 834
use sg13g2_inv_1  _0414_
timestamp 1676382929
transform 1 0 20064 0 -1 9828
box -48 -56 336 834
use sg13g2_inv_1  _0415_
timestamp 1676382929
transform 1 0 14496 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0416_
timestamp 1676382929
transform -1 0 10368 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0417_
timestamp 1676382929
transform -1 0 4992 0 1 11340
box -48 -56 336 834
use sg13g2_mux4_1  _0418_
timestamp 1677257233
transform -1 0 5568 0 1 3780
box -48 -56 2064 834
use sg13g2_inv_1  _0419_
timestamp 1676382929
transform -1 0 2208 0 -1 18900
box -48 -56 336 834
use sg13g2_nor2_1  _0420_
timestamp 1676627187
transform 1 0 1152 0 -1 6804
box -48 -56 432 834
use sg13g2_mux4_1  _0421_
timestamp 1677257233
transform 1 0 4416 0 -1 3780
box -48 -56 2064 834
use sg13g2_a21oi_1  _0422_
timestamp 1683973020
transform -1 0 5856 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _0423_
timestamp 1685175443
transform -1 0 4032 0 -1 3780
box -48 -56 538 834
use sg13g2_o21ai_1  _0424_
timestamp 1685175443
transform 1 0 6432 0 1 3780
box -48 -56 538 834
use sg13g2_a22oi_1  _0425_
timestamp 1685173987
transform 1 0 5856 0 1 2268
box -48 -56 624 834
use sg13g2_nand3_1  _0426_
timestamp 1683988354
transform 1 0 7584 0 -1 5292
box -48 -56 528 834
use sg13g2_nand2b_1  _0427_
timestamp 1676567195
transform -1 0 4608 0 1 2268
box -48 -56 528 834
use sg13g2_a22oi_1  _0428_
timestamp 1685173987
transform -1 0 2688 0 1 5292
box -48 -56 624 834
use sg13g2_nand2b_1  _0429_
timestamp 1676567195
transform -1 0 9216 0 1 2268
box -48 -56 528 834
use sg13g2_a21oi_1  _0430_
timestamp 1683973020
transform -1 0 1632 0 1 5292
box -48 -56 528 834
use sg13g2_nand2_1  _0431_
timestamp 1676557249
transform 1 0 1152 0 -1 5292
box -48 -56 432 834
use sg13g2_o21ai_1  _0432_
timestamp 1685175443
transform 1 0 1440 0 1 3780
box -48 -56 538 834
use sg13g2_mux4_1  _0433_
timestamp 1677257233
transform 1 0 1632 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0434_
timestamp 1677257233
transform 1 0 4992 0 -1 20412
box -48 -56 2064 834
use sg13g2_inv_1  _0435_
timestamp 1676382929
transform 1 0 14976 0 1 8316
box -48 -56 336 834
use sg13g2_nand3_1  _0436_
timestamp 1683988354
transform 1 0 14880 0 1 6804
box -48 -56 528 834
use sg13g2_mux2_1  _0437_
timestamp 1677247768
transform 1 0 16032 0 1 5292
box -48 -56 1008 834
use sg13g2_nor2_1  _0438_
timestamp 1676627187
transform 1 0 16992 0 1 5292
box -48 -56 432 834
use sg13g2_a221oi_1  _0439_
timestamp 1685197497
transform 1 0 16224 0 -1 6804
box -48 -56 816 834
use sg13g2_mux2_1  _0440_
timestamp 1677247768
transform 1 0 16032 0 -1 5292
box -48 -56 1008 834
use sg13g2_a22oi_1  _0441_
timestamp 1685173987
transform -1 0 17568 0 -1 6804
box -48 -56 624 834
use sg13g2_a22oi_1  _0442_
timestamp 1685173987
transform 1 0 15360 0 1 6804
box -48 -56 624 834
use sg13g2_mux4_1  _0443_
timestamp 1677257233
transform -1 0 4704 0 1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0444_
timestamp 1677257233
transform 1 0 4704 0 -1 40068
box -48 -56 2064 834
use sg13g2_inv_1  _0445_
timestamp 1676382929
transform 1 0 20064 0 1 35532
box -48 -56 336 834
use sg13g2_nand3_1  _0446_
timestamp 1683988354
transform 1 0 17760 0 -1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _0447_
timestamp 1677247768
transform -1 0 19392 0 1 37044
box -48 -56 1008 834
use sg13g2_nor2_1  _0448_
timestamp 1676627187
transform 1 0 19008 0 -1 40068
box -48 -56 432 834
use sg13g2_a221oi_1  _0449_
timestamp 1685197497
transform 1 0 18144 0 -1 38556
box -48 -56 816 834
use sg13g2_mux2_1  _0450_
timestamp 1677247768
transform 1 0 17472 0 1 37044
box -48 -56 1008 834
use sg13g2_a22oi_1  _0451_
timestamp 1685173987
transform 1 0 18912 0 -1 38556
box -48 -56 624 834
use sg13g2_a22oi_1  _0452_
timestamp 1685173987
transform -1 0 18720 0 1 38556
box -48 -56 624 834
use sg13g2_mux4_1  _0453_
timestamp 1677257233
transform 1 0 5760 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0454_
timestamp 1677257233
transform -1 0 7008 0 -1 38556
box -48 -56 2064 834
use sg13g2_inv_1  _0455_
timestamp 1676382929
transform 1 0 17472 0 1 21924
box -48 -56 336 834
use sg13g2_nand3_1  _0456_
timestamp 1683988354
transform -1 0 20352 0 1 15876
box -48 -56 528 834
use sg13g2_mux2_1  _0457_
timestamp 1677247768
transform 1 0 19200 0 -1 15876
box -48 -56 1008 834
use sg13g2_nor2_1  _0458_
timestamp 1676627187
transform 1 0 16416 0 -1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  _0459_
timestamp 1685197497
transform 1 0 19104 0 1 15876
box -48 -56 816 834
use sg13g2_mux2_1  _0460_
timestamp 1677247768
transform 1 0 19008 0 1 14364
box -48 -56 1008 834
use sg13g2_a22oi_1  _0461_
timestamp 1685173987
transform -1 0 20064 0 -1 17388
box -48 -56 624 834
use sg13g2_a22oi_1  _0462_
timestamp 1685173987
transform 1 0 18912 0 -1 17388
box -48 -56 624 834
use sg13g2_mux4_1  _0463_
timestamp 1677257233
transform 1 0 5952 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _0464_
timestamp 1677257233
transform 1 0 3936 0 -1 23436
box -48 -56 2064 834
use sg13g2_inv_1  _0465_
timestamp 1676382929
transform -1 0 14016 0 1 5292
box -48 -56 336 834
use sg13g2_nand3_1  _0466_
timestamp 1683988354
transform 1 0 15456 0 1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _0467_
timestamp 1677247768
transform 1 0 16608 0 -1 11340
box -48 -56 1008 834
use sg13g2_nor2_1  _0468_
timestamp 1676627187
transform -1 0 17952 0 -1 11340
box -48 -56 432 834
use sg13g2_a221oi_1  _0469_
timestamp 1685197497
transform 1 0 16512 0 1 11340
box -48 -56 816 834
use sg13g2_mux2_1  _0470_
timestamp 1677247768
transform -1 0 17472 0 1 9828
box -48 -56 1008 834
use sg13g2_a22oi_1  _0471_
timestamp 1685173987
transform 1 0 15936 0 1 9828
box -48 -56 624 834
use sg13g2_a22oi_1  _0472_
timestamp 1685173987
transform 1 0 16224 0 -1 12852
box -48 -56 624 834
use sg13g2_mux4_1  _0473_
timestamp 1677257233
transform 1 0 6912 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0474_
timestamp 1677257233
transform 1 0 1824 0 1 756
box -48 -56 2064 834
use sg13g2_nand3_1  _0475_
timestamp 1683988354
transform 1 0 18336 0 -1 5292
box -48 -56 528 834
use sg13g2_mux2_1  _0476_
timestamp 1677247768
transform 1 0 19008 0 1 5292
box -48 -56 1008 834
use sg13g2_nor2_1  _0477_
timestamp 1676627187
transform 1 0 19968 0 1 5292
box -48 -56 432 834
use sg13g2_a221oi_1  _0478_
timestamp 1685197497
transform 1 0 19392 0 1 6804
box -48 -56 816 834
use sg13g2_mux2_1  _0479_
timestamp 1677247768
transform -1 0 20256 0 -1 6804
box -48 -56 1008 834
use sg13g2_a22oi_1  _0480_
timestamp 1685173987
transform 1 0 19392 0 -1 8316
box -48 -56 624 834
use sg13g2_a22oi_1  _0481_
timestamp 1685173987
transform 1 0 18816 0 -1 8316
box -48 -56 624 834
use sg13g2_mux4_1  _0482_
timestamp 1677257233
transform 1 0 8544 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0483_
timestamp 1677257233
transform 1 0 3840 0 -1 2268
box -48 -56 2064 834
use sg13g2_nand3_1  _0484_
timestamp 1683988354
transform 1 0 19776 0 -1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _0485_
timestamp 1677247768
transform 1 0 19296 0 1 18900
box -48 -56 1008 834
use sg13g2_nor2_1  _0486_
timestamp 1676627187
transform 1 0 19968 0 1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  _0487_
timestamp 1685197497
transform 1 0 19296 0 -1 18900
box -48 -56 816 834
use sg13g2_mux2_1  _0488_
timestamp 1677247768
transform -1 0 19776 0 -1 20412
box -48 -56 1008 834
use sg13g2_a22oi_1  _0489_
timestamp 1685173987
transform 1 0 19008 0 1 20412
box -48 -56 624 834
use sg13g2_a22oi_1  _0490_
timestamp 1685173987
transform 1 0 18240 0 -1 20412
box -48 -56 624 834
use sg13g2_mux4_1  _0491_
timestamp 1677257233
transform 1 0 7488 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0492_
timestamp 1677257233
transform -1 0 5472 0 1 34020
box -48 -56 2064 834
use sg13g2_nand3_1  _0493_
timestamp 1683988354
transform 1 0 11232 0 -1 18900
box -48 -56 528 834
use sg13g2_mux2_1  _0494_
timestamp 1677247768
transform -1 0 14208 0 1 17388
box -48 -56 1008 834
use sg13g2_nor2_1  _0495_
timestamp 1676627187
transform 1 0 14880 0 -1 20412
box -48 -56 432 834
use sg13g2_a221oi_1  _0496_
timestamp 1685197497
transform 1 0 12096 0 -1 20412
box -48 -56 816 834
use sg13g2_mux2_1  _0497_
timestamp 1677247768
transform 1 0 13248 0 -1 17388
box -48 -56 1008 834
use sg13g2_a22oi_1  _0498_
timestamp 1685173987
transform -1 0 16608 0 -1 17388
box -48 -56 624 834
use sg13g2_a22oi_1  _0499_
timestamp 1685173987
transform -1 0 14784 0 1 17388
box -48 -56 624 834
use sg13g2_mux4_1  _0500_
timestamp 1677257233
transform 1 0 6240 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0501_
timestamp 1677257233
transform 1 0 3648 0 -1 27972
box -48 -56 2064 834
use sg13g2_nand3_1  _0502_
timestamp 1683988354
transform -1 0 12480 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _0503_
timestamp 1677247768
transform 1 0 12288 0 1 8316
box -48 -56 1008 834
use sg13g2_nor2_1  _0504_
timestamp 1676627187
transform -1 0 14304 0 -1 8316
box -48 -56 432 834
use sg13g2_a221oi_1  _0505_
timestamp 1685197497
transform 1 0 12192 0 -1 9828
box -48 -56 816 834
use sg13g2_mux2_1  _0506_
timestamp 1677247768
transform -1 0 12288 0 1 8316
box -48 -56 1008 834
use sg13g2_a22oi_1  _0507_
timestamp 1685173987
transform 1 0 11712 0 1 9828
box -48 -56 624 834
use sg13g2_a22oi_1  _0508_
timestamp 1685173987
transform 1 0 11136 0 1 9828
box -48 -56 624 834
use sg13g2_nor2_1  _0509_
timestamp 1676627187
transform 1 0 19872 0 1 3780
box -48 -56 432 834
use sg13g2_mux4_1  _0510_
timestamp 1677257233
transform 1 0 6528 0 1 26460
box -48 -56 2064 834
use sg13g2_nand3b_1  _0511_
timestamp 1676573470
transform 1 0 16512 0 -1 3780
box -48 -56 720 834
use sg13g2_and2_1  _0512_
timestamp 1676901763
transform 1 0 17664 0 -1 5292
box -48 -56 528 834
use sg13g2_a21oi_1  _0513_
timestamp 1683973020
transform -1 0 20064 0 1 2268
box -48 -56 528 834
use sg13g2_nand2b_1  _0514_
timestamp 1676567195
transform 1 0 16992 0 -1 5292
box -48 -56 528 834
use sg13g2_mux4_1  _0515_
timestamp 1677257233
transform 1 0 15840 0 1 3780
box -48 -56 2064 834
use sg13g2_nor2_1  _0516_
timestamp 1676627187
transform -1 0 20256 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _0517_
timestamp 1683973020
transform -1 0 18336 0 1 3780
box -48 -56 528 834
use sg13g2_mux4_1  _0518_
timestamp 1677257233
transform 1 0 8448 0 1 38556
box -48 -56 2064 834
use sg13g2_nand3_1  _0519_
timestamp 1683988354
transform -1 0 16512 0 1 37044
box -48 -56 528 834
use sg13g2_mux2_1  _0520_
timestamp 1677247768
transform -1 0 17472 0 1 35532
box -48 -56 1008 834
use sg13g2_nor2_1  _0521_
timestamp 1676627187
transform 1 0 18240 0 -1 37044
box -48 -56 432 834
use sg13g2_a221oi_1  _0522_
timestamp 1685197497
transform 1 0 15840 0 -1 37044
box -48 -56 816 834
use sg13g2_mux2_1  _0523_
timestamp 1677247768
transform 1 0 15552 0 1 35532
box -48 -56 1008 834
use sg13g2_a22oi_1  _0524_
timestamp 1685173987
transform 1 0 16608 0 -1 37044
box -48 -56 624 834
use sg13g2_a22oi_1  _0525_
timestamp 1685173987
transform 1 0 15456 0 1 37044
box -48 -56 624 834
use sg13g2_mux4_1  _0526_
timestamp 1677257233
transform 1 0 7296 0 1 37044
box -48 -56 2064 834
use sg13g2_nand3_1  _0527_
timestamp 1683988354
transform 1 0 18432 0 1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _0528_
timestamp 1677247768
transform 1 0 19008 0 -1 12852
box -48 -56 1008 834
use sg13g2_nor2_1  _0529_
timestamp 1676627187
transform -1 0 18144 0 1 11340
box -48 -56 432 834
use sg13g2_a221oi_1  _0530_
timestamp 1685197497
transform 1 0 19584 0 1 12852
box -48 -56 816 834
use sg13g2_mux2_1  _0531_
timestamp 1677247768
transform 1 0 18624 0 1 12852
box -48 -56 1008 834
use sg13g2_a22oi_1  _0532_
timestamp 1685173987
transform 1 0 19392 0 -1 14364
box -48 -56 624 834
use sg13g2_a22oi_1  _0533_
timestamp 1685173987
transform 1 0 18816 0 -1 14364
box -48 -56 624 834
use sg13g2_mux4_1  _0534_
timestamp 1677257233
transform 1 0 5952 0 -1 21924
box -48 -56 2064 834
use sg13g2_nand3_1  _0535_
timestamp 1683988354
transform 1 0 16992 0 -1 8316
box -48 -56 528 834
use sg13g2_mux2_1  _0536_
timestamp 1677247768
transform 1 0 16992 0 1 8316
box -48 -56 1008 834
use sg13g2_nor2_1  _0537_
timestamp 1676627187
transform 1 0 17472 0 -1 8316
box -48 -56 432 834
use sg13g2_a221oi_1  _0538_
timestamp 1685197497
transform 1 0 17664 0 -1 9828
box -48 -56 816 834
use sg13g2_mux2_1  _0539_
timestamp 1677247768
transform -1 0 17664 0 -1 9828
box -48 -56 1008 834
use sg13g2_a22oi_1  _0540_
timestamp 1685173987
transform 1 0 15552 0 -1 9828
box -48 -56 624 834
use sg13g2_a22oi_1  _0541_
timestamp 1685173987
transform 1 0 16128 0 -1 9828
box -48 -56 624 834
use sg13g2_mux4_1  _0542_
timestamp 1677257233
transform 1 0 1632 0 -1 26460
box -48 -56 2064 834
use sg13g2_nand3_1  _0543_
timestamp 1683988354
transform -1 0 20064 0 -1 2268
box -48 -56 528 834
use sg13g2_mux2_1  _0544_
timestamp 1677247768
transform 1 0 18912 0 1 3780
box -48 -56 1008 834
use sg13g2_nor2_1  _0545_
timestamp 1676627187
transform 1 0 10656 0 1 3780
box -48 -56 432 834
use sg13g2_a221oi_1  _0546_
timestamp 1685197497
transform 1 0 19104 0 -1 3780
box -48 -56 816 834
use sg13g2_mux2_1  _0547_
timestamp 1677247768
transform -1 0 19776 0 -1 5292
box -48 -56 1008 834
use sg13g2_a22oi_1  _0548_
timestamp 1685173987
transform -1 0 18912 0 1 3780
box -48 -56 624 834
use sg13g2_a22oi_1  _0549_
timestamp 1685173987
transform 1 0 18528 0 -1 3780
box -48 -56 624 834
use sg13g2_mux4_1  _0550_
timestamp 1677257233
transform 1 0 3264 0 -1 37044
box -48 -56 2064 834
use sg13g2_nand3_1  _0551_
timestamp 1683988354
transform 1 0 15840 0 1 20412
box -48 -56 528 834
use sg13g2_mux2_1  _0552_
timestamp 1677247768
transform 1 0 16608 0 -1 18900
box -48 -56 1008 834
use sg13g2_nor2_1  _0553_
timestamp 1676627187
transform 1 0 15456 0 1 20412
box -48 -56 432 834
use sg13g2_a221oi_1  _0554_
timestamp 1685197497
transform 1 0 16512 0 1 18900
box -48 -56 816 834
use sg13g2_mux2_1  _0555_
timestamp 1677247768
transform -1 0 17376 0 1 17388
box -48 -56 1008 834
use sg13g2_a22oi_1  _0556_
timestamp 1685173987
transform 1 0 15360 0 -1 20412
box -48 -56 624 834
use sg13g2_a22oi_1  _0557_
timestamp 1685173987
transform 1 0 16608 0 -1 17388
box -48 -56 624 834
use sg13g2_mux4_1  _0558_
timestamp 1677257233
transform 1 0 7104 0 1 35532
box -48 -56 2064 834
use sg13g2_nand3_1  _0559_
timestamp 1683988354
transform 1 0 12480 0 -1 14364
box -48 -56 528 834
use sg13g2_mux2_1  _0560_
timestamp 1677247768
transform 1 0 13440 0 1 14364
box -48 -56 1008 834
use sg13g2_nor2_1  _0561_
timestamp 1676627187
transform -1 0 12480 0 -1 14364
box -48 -56 432 834
use sg13g2_a221oi_1  _0562_
timestamp 1685197497
transform -1 0 15264 0 -1 15876
box -48 -56 816 834
use sg13g2_mux2_1  _0563_
timestamp 1677247768
transform -1 0 14496 0 -1 15876
box -48 -56 1008 834
use sg13g2_a22oi_1  _0564_
timestamp 1685173987
transform 1 0 11328 0 -1 15876
box -48 -56 624 834
use sg13g2_a22oi_1  _0565_
timestamp 1685173987
transform 1 0 14400 0 1 14364
box -48 -56 624 834
use sg13g2_mux4_1  _0566_
timestamp 1677257233
transform 1 0 6528 0 1 21924
box -48 -56 2064 834
use sg13g2_nand3_1  _0567_
timestamp 1683988354
transform -1 0 12768 0 1 9828
box -48 -56 528 834
use sg13g2_mux2_1  _0568_
timestamp 1677247768
transform -1 0 11040 0 1 8316
box -48 -56 1008 834
use sg13g2_nor2_1  _0569_
timestamp 1676627187
transform 1 0 8352 0 -1 6804
box -48 -56 432 834
use sg13g2_a221oi_1  _0570_
timestamp 1685197497
transform 1 0 9696 0 -1 9828
box -48 -56 816 834
use sg13g2_mux2_1  _0571_
timestamp 1677247768
transform -1 0 10752 0 1 9828
box -48 -56 1008 834
use sg13g2_a22oi_1  _0572_
timestamp 1685173987
transform -1 0 9888 0 1 11340
box -48 -56 624 834
use sg13g2_a22oi_1  _0573_
timestamp 1685173987
transform 1 0 9600 0 -1 8316
box -48 -56 624 834
use sg13g2_o21ai_1  _0574_
timestamp 1685175443
transform 1 0 14592 0 -1 14364
box -48 -56 538 834
use sg13g2_a21oi_1  _0575_
timestamp 1683973020
transform 1 0 15072 0 -1 14364
box -48 -56 528 834
use sg13g2_nor2b_1  _0576_
timestamp 1685181386
transform 1 0 12480 0 1 12852
box -54 -56 528 834
use sg13g2_a21oi_1  _0577_
timestamp 1683973020
transform 1 0 13728 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _0578_
timestamp 1685175443
transform 1 0 15552 0 -1 14364
box -48 -56 538 834
use sg13g2_nor2_1  _0579_
timestamp 1676627187
transform 1 0 14976 0 1 12852
box -48 -56 432 834
use sg13g2_mux4_1  _0580_
timestamp 1677257233
transform 1 0 12960 0 1 12852
box -48 -56 2064 834
use sg13g2_nor2_1  _0581_
timestamp 1676627187
transform 1 0 15840 0 -1 12852
box -48 -56 432 834
use sg13g2_nor2_1  _0582_
timestamp 1676627187
transform 1 0 16032 0 -1 14364
box -48 -56 432 834
use sg13g2_o21ai_1  _0583_
timestamp 1685175443
transform 1 0 14976 0 -1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _0584_
timestamp 1683973020
transform 1 0 15456 0 -1 32508
box -48 -56 528 834
use sg13g2_nor2b_1  _0585_
timestamp 1685181386
transform 1 0 15264 0 -1 29484
box -54 -56 528 834
use sg13g2_a21oi_1  _0586_
timestamp 1683973020
transform 1 0 16320 0 1 29484
box -48 -56 528 834
use sg13g2_o21ai_1  _0587_
timestamp 1685175443
transform 1 0 16416 0 1 30996
box -48 -56 538 834
use sg13g2_nor2_1  _0588_
timestamp 1676627187
transform 1 0 16800 0 1 29484
box -48 -56 432 834
use sg13g2_mux4_1  _0589_
timestamp 1677257233
transform 1 0 14208 0 -1 30996
box -48 -56 2064 834
use sg13g2_nor2_1  _0590_
timestamp 1676627187
transform -1 0 18528 0 -1 32508
box -48 -56 432 834
use sg13g2_nor2_1  _0591_
timestamp 1676627187
transform 1 0 17760 0 -1 32508
box -48 -56 432 834
use sg13g2_o21ai_1  _0592_
timestamp 1685175443
transform -1 0 19872 0 -1 23436
box -48 -56 538 834
use sg13g2_a21oi_1  _0593_
timestamp 1683973020
transform -1 0 19488 0 1 23436
box -48 -56 528 834
use sg13g2_nor2b_1  _0594_
timestamp 1685181386
transform 1 0 18912 0 -1 23436
box -54 -56 528 834
use sg13g2_a21oi_1  _0595_
timestamp 1683973020
transform 1 0 19872 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _0596_
timestamp 1685175443
transform 1 0 19392 0 1 21924
box -48 -56 538 834
use sg13g2_nor2_1  _0597_
timestamp 1676627187
transform 1 0 19488 0 1 23436
box -48 -56 432 834
use sg13g2_mux4_1  _0598_
timestamp 1677257233
transform -1 0 19008 0 1 23436
box -48 -56 2064 834
use sg13g2_nor2_1  _0599_
timestamp 1676627187
transform -1 0 17280 0 -1 23436
box -48 -56 432 834
use sg13g2_nor2_1  _0600_
timestamp 1676627187
transform -1 0 20160 0 -1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  _0601_
timestamp 1685175443
transform -1 0 13344 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _0602_
timestamp 1683973020
transform 1 0 13632 0 -1 6804
box -48 -56 528 834
use sg13g2_nor2b_1  _0603_
timestamp 1685181386
transform 1 0 12960 0 -1 8316
box -54 -56 528 834
use sg13g2_a21oi_1  _0604_
timestamp 1683973020
transform 1 0 13920 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _0605_
timestamp 1685175443
transform 1 0 13440 0 -1 8316
box -48 -56 538 834
use sg13g2_nor2_1  _0606_
timestamp 1676627187
transform 1 0 13344 0 1 5292
box -48 -56 432 834
use sg13g2_mux4_1  _0607_
timestamp 1677257233
transform 1 0 11904 0 1 6804
box -48 -56 2064 834
use sg13g2_nor2_1  _0608_
timestamp 1676627187
transform 1 0 14208 0 -1 6804
box -48 -56 432 834
use sg13g2_nor2_1  _0609_
timestamp 1676627187
transform 1 0 14400 0 1 6804
box -48 -56 432 834
use sg13g2_o21ai_1  _0610_
timestamp 1685175443
transform 1 0 12288 0 1 5292
box -48 -56 538 834
use sg13g2_a21oi_1  _0611_
timestamp 1683973020
transform 1 0 13056 0 -1 5292
box -48 -56 528 834
use sg13g2_nor2b_1  _0612_
timestamp 1685181386
transform 1 0 10560 0 -1 5292
box -54 -56 528 834
use sg13g2_a21oi_1  _0613_
timestamp 1683973020
transform 1 0 11040 0 1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _0614_
timestamp 1685175443
transform 1 0 11424 0 -1 3780
box -48 -56 538 834
use sg13g2_nor2_1  _0615_
timestamp 1676627187
transform -1 0 12384 0 1 2268
box -48 -56 432 834
use sg13g2_mux4_1  _0616_
timestamp 1677257233
transform -1 0 13056 0 -1 5292
box -48 -56 2064 834
use sg13g2_nor2_1  _0617_
timestamp 1676627187
transform 1 0 10272 0 1 3780
box -48 -56 432 834
use sg13g2_nor2_1  _0618_
timestamp 1676627187
transform 1 0 15648 0 1 5292
box -48 -56 432 834
use sg13g2_o21ai_1  _0619_
timestamp 1685175443
transform 1 0 19200 0 -1 21924
box -48 -56 538 834
use sg13g2_a21oi_1  _0620_
timestamp 1683973020
transform 1 0 19680 0 -1 21924
box -48 -56 528 834
use sg13g2_nor2b_1  _0621_
timestamp 1685181386
transform 1 0 18720 0 -1 21924
box -54 -56 528 834
use sg13g2_a21oi_1  _0622_
timestamp 1683973020
transform -1 0 18240 0 -1 20412
box -48 -56 528 834
use sg13g2_o21ai_1  _0623_
timestamp 1685175443
transform -1 0 18816 0 1 20412
box -48 -56 538 834
use sg13g2_nor2_1  _0624_
timestamp 1676627187
transform 1 0 17280 0 1 18900
box -48 -56 432 834
use sg13g2_mux4_1  _0625_
timestamp 1677257233
transform 1 0 16320 0 1 20412
box -48 -56 2064 834
use sg13g2_nor2_1  _0626_
timestamp 1676627187
transform -1 0 20352 0 1 20412
box -48 -56 432 834
use sg13g2_nor2_1  _0627_
timestamp 1676627187
transform 1 0 19584 0 1 20412
box -48 -56 432 834
use sg13g2_o21ai_1  _0628_
timestamp 1685175443
transform 1 0 15552 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _0629_
timestamp 1683973020
transform 1 0 16032 0 1 32508
box -48 -56 528 834
use sg13g2_nor2b_1  _0630_
timestamp 1685181386
transform 1 0 13632 0 -1 32508
box -54 -56 528 834
use sg13g2_a21oi_1  _0631_
timestamp 1683973020
transform 1 0 14304 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _0632_
timestamp 1685175443
transform 1 0 14784 0 1 37044
box -48 -56 538 834
use sg13g2_nor2_1  _0633_
timestamp 1676627187
transform -1 0 15648 0 -1 35532
box -48 -56 432 834
use sg13g2_mux4_1  _0634_
timestamp 1677257233
transform 1 0 13536 0 1 32508
box -48 -56 2064 834
use sg13g2_nor2_1  _0635_
timestamp 1676627187
transform 1 0 17184 0 -1 37044
box -48 -56 432 834
use sg13g2_nor2_1  _0636_
timestamp 1676627187
transform 1 0 18816 0 1 32508
box -48 -56 432 834
use sg13g2_o21ai_1  _0637_
timestamp 1685175443
transform 1 0 11136 0 -1 12852
box -48 -56 538 834
use sg13g2_a21oi_1  _0638_
timestamp 1683973020
transform 1 0 11616 0 -1 12852
box -48 -56 528 834
use sg13g2_nor2b_1  _0639_
timestamp 1685181386
transform 1 0 8736 0 -1 11340
box -54 -56 528 834
use sg13g2_a21oi_1  _0640_
timestamp 1683973020
transform 1 0 11424 0 1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _0641_
timestamp 1685175443
transform 1 0 12000 0 1 12852
box -48 -56 538 834
use sg13g2_nor2_1  _0642_
timestamp 1676627187
transform -1 0 13344 0 -1 9828
box -48 -56 432 834
use sg13g2_mux4_1  _0643_
timestamp 1677257233
transform 1 0 10848 0 -1 11340
box -48 -56 2064 834
use sg13g2_nor2_1  _0644_
timestamp 1676627187
transform -1 0 12960 0 -1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _0645_
timestamp 1676627187
transform 1 0 10752 0 1 9828
box -48 -56 432 834
use sg13g2_nor3_1  _0646_
timestamp 1676639442
transform 1 0 6720 0 1 14364
box -48 -56 528 834
use sg13g2_nand2b_1  _0647_
timestamp 1676567195
transform 1 0 9120 0 1 14364
box -48 -56 528 834
use sg13g2_a221oi_1  _0648_
timestamp 1685197497
transform -1 0 6912 0 1 15876
box -48 -56 816 834
use sg13g2_mux4_1  _0649_
timestamp 1677257233
transform 1 0 9024 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0650_
timestamp 1677257233
transform 1 0 9024 0 1 15876
box -48 -56 2064 834
use sg13g2_mux2_1  _0651_
timestamp 1677247768
transform 1 0 8544 0 -1 17388
box -48 -56 1008 834
use sg13g2_nand2b_1  _0652_
timestamp 1676567195
transform -1 0 12960 0 1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _0653_
timestamp 1676557249
transform -1 0 17280 0 1 30996
box -48 -56 432 834
use sg13g2_a21oi_1  _0654_
timestamp 1683973020
transform 1 0 12096 0 -1 32508
box -48 -56 528 834
use sg13g2_nor3_1  _0655_
timestamp 1676639442
transform -1 0 1728 0 -1 34020
box -48 -56 528 834
use sg13g2_nand2b_1  _0656_
timestamp 1676567195
transform -1 0 4224 0 -1 34020
box -48 -56 528 834
use sg13g2_a221oi_1  _0657_
timestamp 1685197497
transform 1 0 1344 0 1 32508
box -48 -56 816 834
use sg13g2_inv_1  _0658_
timestamp 1676382929
transform 1 0 6144 0 -1 30996
box -48 -56 336 834
use sg13g2_o21ai_1  _0659_
timestamp 1685175443
transform -1 0 10272 0 1 34020
box -48 -56 538 834
use sg13g2_a21o_1  _0660_
timestamp 1677175127
transform -1 0 12480 0 1 32508
box -48 -56 720 834
use sg13g2_nor2b_1  _0661_
timestamp 1685181386
transform -1 0 13440 0 1 32508
box -54 -56 528 834
use sg13g2_a21oi_1  _0662_
timestamp 1683973020
transform 1 0 11616 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _0663_
timestamp 1685175443
transform 1 0 10272 0 1 34020
box -48 -56 538 834
use sg13g2_mux2_1  _0664_
timestamp 1677247768
transform 1 0 10656 0 -1 32508
box -48 -56 1008 834
use sg13g2_a21oi_1  _0665_
timestamp 1683973020
transform -1 0 13056 0 -1 32508
box -48 -56 528 834
use sg13g2_a22oi_1  _0666_
timestamp 1685173987
transform 1 0 11520 0 -1 30996
box -48 -56 624 834
use sg13g2_mux2_1  _0667_
timestamp 1677247768
transform 1 0 11904 0 -1 29484
box -48 -56 1008 834
use sg13g2_nand2b_1  _0668_
timestamp 1676567195
transform 1 0 12384 0 -1 27972
box -48 -56 528 834
use sg13g2_nand2b_1  _0669_
timestamp 1676567195
transform 1 0 1152 0 1 26460
box -48 -56 528 834
use sg13g2_nor3_1  _0670_
timestamp 1676639442
transform -1 0 1632 0 -1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  _0671_
timestamp 1685197497
transform 1 0 2784 0 1 27972
box -48 -56 816 834
use sg13g2_mux2_1  _0672_
timestamp 1677247768
transform -1 0 12672 0 1 29484
box -48 -56 1008 834
use sg13g2_a21oi_1  _0673_
timestamp 1683973020
transform -1 0 11424 0 1 27972
box -48 -56 528 834
use sg13g2_a21oi_1  _0674_
timestamp 1683973020
transform 1 0 11712 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _0675_
timestamp 1685175443
transform 1 0 11424 0 1 27972
box -48 -56 538 834
use sg13g2_mux2_1  _0676_
timestamp 1677247768
transform 1 0 11904 0 1 27972
box -48 -56 1008 834
use sg13g2_a21oi_1  _0677_
timestamp 1683973020
transform 1 0 12864 0 1 27972
box -48 -56 528 834
use sg13g2_a22oi_1  _0678_
timestamp 1685173987
transform -1 0 13440 0 -1 29484
box -48 -56 624 834
use sg13g2_mux2_1  _0679_
timestamp 1677247768
transform -1 0 6048 0 1 14364
box -48 -56 1008 834
use sg13g2_nand2b_1  _0680_
timestamp 1676567195
transform -1 0 3360 0 -1 11340
box -48 -56 528 834
use sg13g2_nand2b_1  _0681_
timestamp 1676567195
transform -1 0 2016 0 -1 6804
box -48 -56 528 834
use sg13g2_nor3_1  _0682_
timestamp 1676639442
transform 1 0 1632 0 1 5292
box -48 -56 528 834
use sg13g2_a221oi_1  _0683_
timestamp 1685197497
transform 1 0 4896 0 -1 8316
box -48 -56 816 834
use sg13g2_mux2_1  _0684_
timestamp 1677247768
transform -1 0 4128 0 -1 12852
box -48 -56 1008 834
use sg13g2_a21oi_1  _0685_
timestamp 1683973020
transform 1 0 1632 0 1 15876
box -48 -56 528 834
use sg13g2_a21oi_1  _0686_
timestamp 1683973020
transform 1 0 4320 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _0687_
timestamp 1685175443
transform -1 0 2208 0 -1 17388
box -48 -56 538 834
use sg13g2_mux2_1  _0688_
timestamp 1677247768
transform -1 0 3744 0 1 9828
box -48 -56 1008 834
use sg13g2_a21oi_1  _0689_
timestamp 1683973020
transform -1 0 1632 0 1 15876
box -48 -56 528 834
use sg13g2_a22oi_1  _0690_
timestamp 1685173987
transform -1 0 1824 0 1 14364
box -48 -56 624 834
use sg13g2_mux2_1  _0691_
timestamp 1677247768
transform -1 0 4320 0 -1 9828
box -48 -56 1008 834
use sg13g2_mux2_1  _0692_
timestamp 1677247768
transform -1 0 5376 0 -1 14364
box -48 -56 1008 834
use sg13g2_nand2b_1  _0693_
timestamp 1676567195
transform 1 0 2016 0 -1 6804
box -48 -56 528 834
use sg13g2_a21oi_1  _0694_
timestamp 1683973020
transform 1 0 1152 0 1 6804
box -48 -56 528 834
use sg13g2_a21oi_1  _0695_
timestamp 1683973020
transform 1 0 1248 0 -1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _0696_
timestamp 1685175443
transform 1 0 1632 0 1 6804
box -48 -56 538 834
use sg13g2_mux2_1  _0697_
timestamp 1677247768
transform -1 0 4128 0 1 8316
box -48 -56 1008 834
use sg13g2_a21oi_1  _0698_
timestamp 1683973020
transform 1 0 1248 0 -1 17388
box -48 -56 528 834
use sg13g2_a22oi_1  _0699_
timestamp 1685173987
transform -1 0 6624 0 1 14364
box -48 -56 624 834
use sg13g2_mux2_1  _0700_
timestamp 1677247768
transform 1 0 4800 0 -1 26460
box -48 -56 1008 834
use sg13g2_mux2_1  _0701_
timestamp 1677247768
transform 1 0 5184 0 -1 30996
box -48 -56 1008 834
use sg13g2_nand2b_1  _0702_
timestamp 1676567195
transform 1 0 5472 0 1 24948
box -48 -56 528 834
use sg13g2_a21oi_1  _0703_
timestamp 1683973020
transform -1 0 6912 0 -1 34020
box -48 -56 528 834
use sg13g2_a21oi_1  _0704_
timestamp 1683973020
transform -1 0 1728 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _0705_
timestamp 1685175443
transform 1 0 3936 0 1 26460
box -48 -56 538 834
use sg13g2_mux2_1  _0706_
timestamp 1677247768
transform -1 0 6624 0 -1 27972
box -48 -56 1008 834
use sg13g2_a21oi_1  _0707_
timestamp 1683973020
transform 1 0 4992 0 1 35532
box -48 -56 528 834
use sg13g2_a22oi_1  _0708_
timestamp 1685173987
transform -1 0 8736 0 1 30996
box -48 -56 624 834
use sg13g2_o21ai_1  _0709_
timestamp 1685175443
transform -1 0 7776 0 1 34020
box -48 -56 538 834
use sg13g2_a21o_1  _0710_
timestamp 1677175127
transform -1 0 9984 0 1 29484
box -48 -56 720 834
use sg13g2_nand2b_1  _0711_
timestamp 1676567195
transform -1 0 8928 0 1 32508
box -48 -56 528 834
use sg13g2_nand2_1  _0712_
timestamp 1676557249
transform 1 0 7776 0 -1 35532
box -48 -56 432 834
use sg13g2_a21oi_1  _0713_
timestamp 1683973020
transform -1 0 8544 0 -1 29484
box -48 -56 528 834
use sg13g2_nor2b_1  _0714_
timestamp 1685181386
transform -1 0 9120 0 1 26460
box -54 -56 528 834
use sg13g2_a21oi_1  _0715_
timestamp 1683973020
transform 1 0 9120 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _0716_
timestamp 1685175443
transform 1 0 9408 0 -1 27972
box -48 -56 538 834
use sg13g2_mux2_1  _0717_
timestamp 1677247768
transform 1 0 8352 0 1 29484
box -48 -56 1008 834
use sg13g2_a21oi_1  _0718_
timestamp 1683973020
transform 1 0 8928 0 -1 27972
box -48 -56 528 834
use sg13g2_a22oi_1  _0719_
timestamp 1685173987
transform -1 0 9888 0 -1 30996
box -48 -56 624 834
use sg13g2_nor2_1  _0720_
timestamp 1676627187
transform -1 0 9024 0 1 15876
box -48 -56 432 834
use sg13g2_nor2_1  _0721_
timestamp 1676627187
transform 1 0 11136 0 1 14364
box -48 -56 432 834
use sg13g2_nor3_1  _0722_
timestamp 1676639442
transform 1 0 10080 0 1 14364
box -48 -56 528 834
use sg13g2_o21ai_1  _0723_
timestamp 1685175443
transform -1 0 11040 0 -1 12852
box -48 -56 538 834
use sg13g2_a21o_1  _0724_
timestamp 1677175127
transform 1 0 10752 0 1 12852
box -48 -56 720 834
use sg13g2_nor2b_1  _0725_
timestamp 1685181386
transform -1 0 10752 0 1 12852
box -54 -56 528 834
use sg13g2_a21oi_1  _0726_
timestamp 1683973020
transform 1 0 9888 0 -1 12852
box -48 -56 528 834
use sg13g2_o21ai_1  _0727_
timestamp 1685175443
transform 1 0 9600 0 1 14364
box -48 -56 538 834
use sg13g2_mux2_1  _0728_
timestamp 1677247768
transform 1 0 10656 0 -1 14364
box -48 -56 1008 834
use sg13g2_a21oi_1  _0729_
timestamp 1683973020
transform 1 0 11616 0 -1 14364
box -48 -56 528 834
use sg13g2_a22oi_1  _0730_
timestamp 1685173987
transform -1 0 11136 0 1 14364
box -48 -56 624 834
use sg13g2_mux4_1  _0731_
timestamp 1677257233
transform 1 0 2112 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0732_
timestamp 1677257233
transform 1 0 2208 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux2_1  _0733_
timestamp 1677247768
transform 1 0 2784 0 -1 15876
box -48 -56 1008 834
use sg13g2_mux4_1  _0734_
timestamp 1677257233
transform 1 0 2496 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0735_
timestamp 1677257233
transform 1 0 2592 0 1 18900
box -48 -56 2064 834
use sg13g2_mux2_1  _0736_
timestamp 1677247768
transform 1 0 4512 0 -1 18900
box -48 -56 1008 834
use sg13g2_mux4_1  _0737_
timestamp 1677257233
transform 1 0 2208 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0738_
timestamp 1677257233
transform 1 0 2400 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux2_1  _0739_
timestamp 1677247768
transform 1 0 4416 0 -1 21924
box -48 -56 1008 834
use sg13g2_mux4_1  _0740_
timestamp 1677257233
transform 1 0 6048 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0741_
timestamp 1677257233
transform 1 0 6048 0 1 17388
box -48 -56 2064 834
use sg13g2_mux2_1  _0742_
timestamp 1677247768
transform 1 0 8064 0 1 17388
box -48 -56 1008 834
use sg13g2_o21ai_1  _0743_
timestamp 1685175443
transform 1 0 15168 0 -1 2268
box -48 -56 538 834
use sg13g2_a21oi_1  _0744_
timestamp 1683973020
transform 1 0 17664 0 -1 3780
box -48 -56 528 834
use sg13g2_or2_1  _0745_
timestamp 1684236171
transform -1 0 17760 0 1 2268
box -48 -56 528 834
use sg13g2_o21ai_1  _0746_
timestamp 1685175443
transform -1 0 14112 0 -1 5292
box -48 -56 538 834
use sg13g2_o21ai_1  _0747_
timestamp 1685175443
transform 1 0 13632 0 1 3780
box -48 -56 538 834
use sg13g2_nor2_1  _0748_
timestamp 1676627187
transform -1 0 18528 0 -1 3780
box -48 -56 432 834
use sg13g2_a21oi_1  _0749_
timestamp 1683973020
transform -1 0 17664 0 -1 3780
box -48 -56 528 834
use sg13g2_o21ai_1  _0750_
timestamp 1685175443
transform -1 0 13824 0 1 756
box -48 -56 538 834
use sg13g2_mux2_1  _0751_
timestamp 1677247768
transform 1 0 15264 0 -1 3780
box -48 -56 1008 834
use sg13g2_a21oi_1  _0752_
timestamp 1683973020
transform 1 0 17376 0 1 756
box -48 -56 528 834
use sg13g2_a21oi_1  _0753_
timestamp 1683973020
transform 1 0 12864 0 1 756
box -48 -56 528 834
use sg13g2_o21ai_1  _0754_
timestamp 1685175443
transform 1 0 14496 0 -1 38556
box -48 -56 538 834
use sg13g2_a21oi_1  _0755_
timestamp 1683973020
transform 1 0 15648 0 1 38556
box -48 -56 528 834
use sg13g2_or2_1  _0756_
timestamp 1684236171
transform 1 0 15168 0 1 38556
box -48 -56 528 834
use sg13g2_o21ai_1  _0757_
timestamp 1685175443
transform -1 0 17184 0 1 40068
box -48 -56 538 834
use sg13g2_o21ai_1  _0758_
timestamp 1685175443
transform -1 0 16992 0 1 37044
box -48 -56 538 834
use sg13g2_nor2_1  _0759_
timestamp 1676627187
transform 1 0 16128 0 1 38556
box -48 -56 432 834
use sg13g2_a21oi_1  _0760_
timestamp 1683973020
transform -1 0 14496 0 1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _0761_
timestamp 1685175443
transform -1 0 16224 0 1 40068
box -48 -56 538 834
use sg13g2_mux2_1  _0762_
timestamp 1677247768
transform 1 0 14976 0 -1 38556
box -48 -56 1008 834
use sg13g2_a21oi_1  _0763_
timestamp 1683973020
transform 1 0 17184 0 1 40068
box -48 -56 528 834
use sg13g2_a21oi_1  _0764_
timestamp 1683973020
transform -1 0 15936 0 -1 40068
box -48 -56 528 834
use sg13g2_mux4_1  _0765_
timestamp 1677257233
transform 1 0 15072 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0766_
timestamp 1677257233
transform 1 0 15552 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux2_1  _0767_
timestamp 1677247768
transform -1 0 17856 0 1 14364
box -48 -56 1008 834
use sg13g2_mux4_1  _0768_
timestamp 1677257233
transform 1 0 13056 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0769_
timestamp 1677257233
transform -1 0 15456 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux2_1  _0770_
timestamp 1677247768
transform 1 0 14400 0 -1 8316
box -48 -56 1008 834
use sg13g2_mux2_1  _0771_
timestamp 1677247768
transform 1 0 18624 0 -1 9828
box -48 -56 1008 834
use sg13g2_or2_1  _0772_
timestamp 1684236171
transform 1 0 17568 0 1 9828
box -48 -56 528 834
use sg13g2_o21ai_1  _0773_
timestamp 1685175443
transform -1 0 18816 0 -1 8316
box -48 -56 538 834
use sg13g2_o21ai_1  _0774_
timestamp 1685175443
transform 1 0 19680 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _0775_
timestamp 1683973020
transform -1 0 20064 0 -1 9828
box -48 -56 528 834
use sg13g2_mux4_1  _0776_
timestamp 1677257233
transform 1 0 18240 0 1 8316
box -48 -56 2064 834
use sg13g2_nor2_1  _0777_
timestamp 1676627187
transform 1 0 19968 0 -1 8316
box -48 -56 432 834
use sg13g2_nor2_1  _0778_
timestamp 1676627187
transform -1 0 18336 0 -1 11340
box -48 -56 432 834
use sg13g2_mux2_1  _0779_
timestamp 1677247768
transform 1 0 12192 0 -1 40068
box -48 -56 1008 834
use sg13g2_or2_1  _0780_
timestamp 1684236171
transform 1 0 13728 0 1 38556
box -48 -56 528 834
use sg13g2_o21ai_1  _0781_
timestamp 1685175443
transform 1 0 14208 0 1 38556
box -48 -56 538 834
use sg13g2_o21ai_1  _0782_
timestamp 1685175443
transform -1 0 16704 0 1 40068
box -48 -56 538 834
use sg13g2_a21oi_1  _0783_
timestamp 1683973020
transform -1 0 15360 0 -1 40068
box -48 -56 528 834
use sg13g2_a21oi_1  _0784_
timestamp 1683973020
transform -1 0 15168 0 1 38556
box -48 -56 528 834
use sg13g2_o21ai_1  _0785_
timestamp 1685175443
transform 1 0 15264 0 1 40068
box -48 -56 538 834
use sg13g2_mux2_1  _0786_
timestamp 1677247768
transform 1 0 12288 0 1 40068
box -48 -56 1008 834
use sg13g2_a21oi_1  _0787_
timestamp 1683973020
transform 1 0 16992 0 -1 41580
box -48 -56 528 834
use sg13g2_a21oi_1  _0788_
timestamp 1683973020
transform -1 0 5376 0 -1 41580
box -48 -56 528 834
use sg13g2_mux2_1  _0789_
timestamp 1677247768
transform 1 0 12672 0 -1 35532
box -48 -56 1008 834
use sg13g2_or2_1  _0790_
timestamp 1684236171
transform -1 0 13536 0 -1 32508
box -48 -56 528 834
use sg13g2_o21ai_1  _0791_
timestamp 1685175443
transform -1 0 10464 0 1 35532
box -48 -56 538 834
use sg13g2_o21ai_1  _0792_
timestamp 1685175443
transform -1 0 9984 0 1 35532
box -48 -56 538 834
use sg13g2_a21oi_1  _0793_
timestamp 1683973020
transform 1 0 14592 0 1 34020
box -48 -56 528 834
use sg13g2_mux4_1  _0794_
timestamp 1677257233
transform 1 0 10752 0 1 34020
box -48 -56 2064 834
use sg13g2_nor2_1  _0795_
timestamp 1676627187
transform -1 0 14016 0 1 37044
box -48 -56 432 834
use sg13g2_nor2_1  _0796_
timestamp 1676627187
transform 1 0 12480 0 -1 38556
box -48 -56 432 834
use sg13g2_mux2_1  _0797_
timestamp 1677247768
transform -1 0 9216 0 1 11340
box -48 -56 1008 834
use sg13g2_or2_1  _0798_
timestamp 1684236171
transform -1 0 8544 0 1 6804
box -48 -56 528 834
use sg13g2_o21ai_1  _0799_
timestamp 1685175443
transform 1 0 7584 0 1 6804
box -48 -56 538 834
use sg13g2_o21ai_1  _0800_
timestamp 1685175443
transform -1 0 8160 0 1 9828
box -48 -56 538 834
use sg13g2_a21oi_1  _0801_
timestamp 1683973020
transform 1 0 7776 0 -1 12852
box -48 -56 528 834
use sg13g2_mux4_1  _0802_
timestamp 1677257233
transform -1 0 8736 0 -1 11340
box -48 -56 2064 834
use sg13g2_nor2_1  _0803_
timestamp 1676627187
transform 1 0 3744 0 1 6804
box -48 -56 432 834
use sg13g2_nor2_1  _0804_
timestamp 1676627187
transform -1 0 7584 0 1 3780
box -48 -56 432 834
use sg13g2_o21ai_1  _0805_
timestamp 1685175443
transform -1 0 1728 0 1 23436
box -48 -56 538 834
use sg13g2_nand2b_1  _0806_
timestamp 1676567195
transform 1 0 3264 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _0807_
timestamp 1685175443
transform -1 0 2208 0 1 23436
box -48 -56 538 834
use sg13g2_mux4_1  _0808_
timestamp 1677257233
transform 1 0 12864 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0809_
timestamp 1677257233
transform 1 0 17280 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0810_
timestamp 1677257233
transform 1 0 16800 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0811_
timestamp 1677257233
transform 1 0 14880 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _0812_
timestamp 1677257233
transform 1 0 13632 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0813_
timestamp 1677257233
transform 1 0 17376 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0814_
timestamp 1677257233
transform 1 0 17376 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0815_
timestamp 1677257233
transform 1 0 13248 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0816_
timestamp 1677257233
transform 1 0 9024 0 -1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0817_
timestamp 1677257233
transform 1 0 11904 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0818_
timestamp 1677257233
transform 1 0 9888 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0819_
timestamp 1677257233
transform 1 0 9888 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0820_
timestamp 1677257233
transform 1 0 11040 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0821_
timestamp 1677257233
transform 1 0 15072 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0822_
timestamp 1677257233
transform 1 0 17088 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0823_
timestamp 1677257233
transform 1 0 12576 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0824_
timestamp 1677257233
transform 1 0 9792 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0825_
timestamp 1677257233
transform 1 0 17280 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0826_
timestamp 1677257233
transform 1 0 12480 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0827_
timestamp 1677257233
transform 1 0 10272 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0828_
timestamp 1677257233
transform 1 0 9504 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0829_
timestamp 1677257233
transform 1 0 17088 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0830_
timestamp 1677257233
transform 1 0 12672 0 -1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0831_
timestamp 1677257233
transform 1 0 9120 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _0832_
timestamp 1677257233
transform 1 0 9024 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0833_
timestamp 1677257233
transform 1 0 14784 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0834_
timestamp 1677257233
transform 1 0 17184 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0835_
timestamp 1677257233
transform 1 0 12864 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0836_
timestamp 1677257233
transform 1 0 8832 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0837_
timestamp 1677257233
transform 1 0 6240 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0838_
timestamp 1677257233
transform -1 0 10464 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0839_
timestamp 1677257233
transform -1 0 9696 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0840_
timestamp 1677257233
transform 1 0 6720 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0841_
timestamp 1677257233
transform -1 0 10272 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0842_
timestamp 1677257233
transform 1 0 7008 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0843_
timestamp 1677257233
transform 1 0 6432 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0844_
timestamp 1677257233
transform -1 0 8352 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0845_
timestamp 1677257233
transform 1 0 7776 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0846_
timestamp 1677257233
transform -1 0 8832 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0847_
timestamp 1677257233
transform 1 0 6432 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0848_
timestamp 1677257233
transform -1 0 7776 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0849_
timestamp 1677257233
transform -1 0 5184 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0850_
timestamp 1677257233
transform -1 0 5376 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0851_
timestamp 1677257233
transform -1 0 4512 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0852_
timestamp 1677257233
transform -1 0 5760 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0853_
timestamp 1677257233
transform -1 0 9024 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0854_
timestamp 1677257233
transform 1 0 2496 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0855_
timestamp 1677257233
transform 1 0 4128 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0856_
timestamp 1677257233
transform -1 0 4896 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0857_
timestamp 1677257233
transform -1 0 3552 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0858_
timestamp 1677257233
transform -1 0 8448 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0859_
timestamp 1677257233
transform -1 0 7776 0 -1 12852
box -48 -56 2064 834
use sg13g2_dlhq_1  _0860_
timestamp 1678805552
transform 1 0 4128 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0861_
timestamp 1678805552
transform -1 0 7296 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0862_
timestamp 1678805552
transform 1 0 4800 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0863_
timestamp 1678805552
transform 1 0 4800 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0864_
timestamp 1678805552
transform -1 0 13632 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _0865_
timestamp 1678805552
transform -1 0 12480 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _0866_
timestamp 1678805552
transform -1 0 9888 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0867_
timestamp 1678805552
transform -1 0 4320 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0868_
timestamp 1678805552
transform 1 0 2112 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0869_
timestamp 1678805552
transform 1 0 4128 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0870_
timestamp 1678805552
transform 1 0 1152 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _0871_
timestamp 1678805552
transform -1 0 16992 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _0872_
timestamp 1678805552
transform -1 0 8928 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0873_
timestamp 1678805552
transform 1 0 5472 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0874_
timestamp 1678805552
transform -1 0 5088 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0875_
timestamp 1678805552
transform 1 0 1728 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0876_
timestamp 1678805552
transform -1 0 15264 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0877_
timestamp 1678805552
transform -1 0 4416 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0878_
timestamp 1678805552
transform 1 0 1728 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _0879_
timestamp 1678805552
transform 1 0 1440 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0880_
timestamp 1678805552
transform 1 0 1440 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0881_
timestamp 1678805552
transform 1 0 1248 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _0882_
timestamp 1678805552
transform 1 0 4512 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0883_
timestamp 1678805552
transform -1 0 7392 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0884_
timestamp 1678805552
transform 1 0 5088 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0885_
timestamp 1678805552
transform -1 0 6624 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0886_
timestamp 1678805552
transform 1 0 5856 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0887_
timestamp 1678805552
transform 1 0 8832 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0888_
timestamp 1678805552
transform -1 0 11424 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _0889_
timestamp 1678805552
transform 1 0 10464 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0890_
timestamp 1678805552
transform 1 0 10560 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _0891_
timestamp 1678805552
transform 1 0 10656 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _0892_
timestamp 1678805552
transform 1 0 10464 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _0893_
timestamp 1678805552
transform 1 0 18048 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0894_
timestamp 1678805552
transform 1 0 18144 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0895_
timestamp 1678805552
transform 1 0 18336 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0896_
timestamp 1678805552
transform 1 0 4800 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0897_
timestamp 1678805552
transform 1 0 6624 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0898_
timestamp 1678805552
transform 1 0 5184 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0899_
timestamp 1678805552
transform -1 0 8640 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0900_
timestamp 1678805552
transform 1 0 5856 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _0901_
timestamp 1678805552
transform 1 0 8160 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _0902_
timestamp 1678805552
transform 1 0 4416 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0903_
timestamp 1678805552
transform 1 0 6048 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0904_
timestamp 1678805552
transform 1 0 4800 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0905_
timestamp 1678805552
transform 1 0 6432 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0906_
timestamp 1678805552
transform 1 0 5376 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0907_
timestamp 1678805552
transform 1 0 7392 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0908_
timestamp 1678805552
transform 1 0 7584 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0909_
timestamp 1678805552
transform 1 0 1920 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0910_
timestamp 1678805552
transform 1 0 3168 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0911_
timestamp 1678805552
transform 1 0 2112 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0912_
timestamp 1678805552
transform 1 0 6720 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0913_
timestamp 1678805552
transform 1 0 4800 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0914_
timestamp 1678805552
transform -1 0 11520 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0915_
timestamp 1678805552
transform 1 0 5952 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0916_
timestamp 1678805552
transform 1 0 1536 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0917_
timestamp 1678805552
transform -1 0 15744 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0918_
timestamp 1678805552
transform 1 0 8736 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0919_
timestamp 1678805552
transform 1 0 5664 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0920_
timestamp 1678805552
transform 1 0 12960 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0921_
timestamp 1678805552
transform 1 0 13344 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _0922_
timestamp 1678805552
transform -1 0 14784 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0923_
timestamp 1678805552
transform 1 0 13440 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0924_
timestamp 1678805552
transform 1 0 15264 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0925_
timestamp 1678805552
transform 1 0 14400 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0926_
timestamp 1678805552
transform 1 0 13248 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _0927_
timestamp 1678805552
transform 1 0 13632 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _0928_
timestamp 1678805552
transform 1 0 12864 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _0929_
timestamp 1678805552
transform 1 0 11232 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0930_
timestamp 1678805552
transform 1 0 13536 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0931_
timestamp 1678805552
transform -1 0 13536 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _0932_
timestamp 1678805552
transform 1 0 4416 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0933_
timestamp 1678805552
transform 1 0 4416 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0934_
timestamp 1678805552
transform 1 0 7008 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0935_
timestamp 1678805552
transform 1 0 1152 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _0936_
timestamp 1678805552
transform 1 0 1152 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _0937_
timestamp 1678805552
transform 1 0 1632 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _0938_
timestamp 1678805552
transform 1 0 1152 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _0939_
timestamp 1678805552
transform 1 0 1152 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0940_
timestamp 1678805552
transform 1 0 2784 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0941_
timestamp 1678805552
transform 1 0 1152 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0942_
timestamp 1678805552
transform 1 0 1824 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0943_
timestamp 1678805552
transform 1 0 1152 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0944_
timestamp 1678805552
transform 1 0 8256 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0945_
timestamp 1678805552
transform 1 0 8448 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0946_
timestamp 1678805552
transform 1 0 9024 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0947_
timestamp 1678805552
transform 1 0 6528 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0948_
timestamp 1678805552
transform 1 0 6432 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0949_
timestamp 1678805552
transform 1 0 6624 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0950_
timestamp 1678805552
transform 1 0 1824 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _0951_
timestamp 1678805552
transform 1 0 3072 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0952_
timestamp 1678805552
transform 1 0 1824 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0953_
timestamp 1678805552
transform 1 0 1152 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _0954_
timestamp 1678805552
transform -1 0 3072 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0955_
timestamp 1678805552
transform -1 0 2880 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0956_
timestamp 1678805552
transform 1 0 2784 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0957_
timestamp 1678805552
transform -1 0 5088 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0958_
timestamp 1678805552
transform 1 0 1152 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0959_
timestamp 1678805552
transform 1 0 9888 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0960_
timestamp 1678805552
transform 1 0 10080 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0961_
timestamp 1678805552
transform 1 0 10272 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0962_
timestamp 1678805552
transform 1 0 8928 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0963_
timestamp 1678805552
transform 1 0 9024 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _0964_
timestamp 1678805552
transform 1 0 9024 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0965_
timestamp 1678805552
transform 1 0 7488 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0966_
timestamp 1678805552
transform 1 0 9504 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0967_
timestamp 1678805552
transform -1 0 11136 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _0968_
timestamp 1678805552
transform -1 0 10848 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0969_
timestamp 1678805552
transform 1 0 9888 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0970_
timestamp 1678805552
transform 1 0 11520 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _0971_
timestamp 1678805552
transform 1 0 12288 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0972_
timestamp 1678805552
transform 1 0 12960 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0973_
timestamp 1678805552
transform 1 0 13920 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _0974_
timestamp 1678805552
transform 1 0 15456 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _0975_
timestamp 1678805552
transform 1 0 17088 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _0976_
timestamp 1678805552
transform 1 0 15936 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0977_
timestamp 1678805552
transform 1 0 7584 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0978_
timestamp 1678805552
transform 1 0 9600 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _0979_
timestamp 1678805552
transform -1 0 13632 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0980_
timestamp 1678805552
transform 1 0 12000 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _0981_
timestamp 1678805552
transform 1 0 10368 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _0982_
timestamp 1678805552
transform 1 0 12000 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _0983_
timestamp 1678805552
transform 1 0 17280 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _0984_
timestamp 1678805552
transform 1 0 15840 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _0985_
timestamp 1678805552
transform 1 0 17760 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _0986_
timestamp 1678805552
transform 1 0 13056 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0987_
timestamp 1678805552
transform 1 0 14688 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0988_
timestamp 1678805552
transform 1 0 14784 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0989_
timestamp 1678805552
transform 1 0 12096 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0990_
timestamp 1678805552
transform 1 0 12960 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _0991_
timestamp 1678805552
transform 1 0 14208 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _0992_
timestamp 1678805552
transform 1 0 13248 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _0993_
timestamp 1678805552
transform 1 0 11232 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _0994_
timestamp 1678805552
transform 1 0 17472 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _0995_
timestamp 1678805552
transform 1 0 16224 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _0996_
timestamp 1678805552
transform 1 0 15072 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _0997_
timestamp 1678805552
transform 1 0 13536 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _0998_
timestamp 1678805552
transform 1 0 9600 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _0999_
timestamp 1678805552
transform 1 0 7968 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1000_
timestamp 1678805552
transform 1 0 8640 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1001_
timestamp 1678805552
transform 1 0 7968 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1002_
timestamp 1678805552
transform -1 0 16320 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1003_
timestamp 1678805552
transform 1 0 11040 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1004_
timestamp 1678805552
transform 1 0 17760 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1005_
timestamp 1678805552
transform 1 0 16320 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1006_
timestamp 1678805552
transform 1 0 9600 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1007_
timestamp 1678805552
transform 1 0 7968 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1008_
timestamp 1678805552
transform 1 0 10656 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1009_
timestamp 1678805552
transform 1 0 7392 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1010_
timestamp 1678805552
transform 1 0 12480 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1011_
timestamp 1678805552
transform 1 0 10848 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1012_
timestamp 1678805552
transform 1 0 18048 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1013_
timestamp 1678805552
transform 1 0 15648 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1014_
timestamp 1678805552
transform 1 0 9600 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1015_
timestamp 1678805552
transform 1 0 7968 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1016_
timestamp 1678805552
transform 1 0 12672 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1017_
timestamp 1678805552
transform 1 0 11232 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1018_
timestamp 1678805552
transform 1 0 17760 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1019_
timestamp 1678805552
transform 1 0 15744 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1020_
timestamp 1678805552
transform 1 0 15264 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1021_
timestamp 1678805552
transform 1 0 13632 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1022_
timestamp 1678805552
transform 1 0 11328 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1023_
timestamp 1678805552
transform 1 0 9408 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1024_
timestamp 1678805552
transform 1 0 8544 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1025_
timestamp 1678805552
transform 1 0 10080 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1026_
timestamp 1678805552
transform 1 0 9216 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1027_
timestamp 1678805552
transform 1 0 10464 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1028_
timestamp 1678805552
transform 1 0 10368 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1029_
timestamp 1678805552
transform 1 0 12288 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1030_
timestamp 1678805552
transform 1 0 5760 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1031_
timestamp 1678805552
transform 1 0 9120 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1032_
timestamp 1678805552
transform 1 0 13440 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1033_
timestamp 1678805552
transform 1 0 11904 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1034_
timestamp 1678805552
transform 1 0 18144 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1035_
timestamp 1678805552
transform 1 0 16128 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1036_
timestamp 1678805552
transform 1 0 18624 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1037_
timestamp 1678805552
transform 1 0 15360 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1038_
timestamp 1678805552
transform 1 0 13824 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1039_
timestamp 1678805552
transform 1 0 12192 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1040_
timestamp 1678805552
transform 1 0 15168 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1041_
timestamp 1678805552
transform 1 0 13440 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1042_
timestamp 1678805552
transform 1 0 16992 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1043_
timestamp 1678805552
transform 1 0 15552 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1044_
timestamp 1678805552
transform 1 0 17664 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1045_
timestamp 1678805552
transform 1 0 15648 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1046_
timestamp 1678805552
transform 1 0 13344 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1047_
timestamp 1678805552
transform 1 0 11520 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1048_
timestamp 1678805552
transform 1 0 8160 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1049_
timestamp 1678805552
transform 1 0 8448 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1050_
timestamp 1678805552
transform 1 0 7968 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1051_
timestamp 1678805552
transform 1 0 11904 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1052_
timestamp 1678805552
transform 1 0 11520 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1053_
timestamp 1678805552
transform 1 0 11520 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1054_
timestamp 1678805552
transform 1 0 14784 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1055_
timestamp 1678805552
transform 1 0 14880 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1056_
timestamp 1678805552
transform 1 0 14976 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1057_
timestamp 1678805552
transform 1 0 17952 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1058_
timestamp 1678805552
transform 1 0 17952 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1059_
timestamp 1678805552
transform 1 0 17856 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1060_
timestamp 1678805552
transform 1 0 15264 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1061_
timestamp 1678805552
transform 1 0 15936 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1062_
timestamp 1678805552
transform 1 0 15360 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1063_
timestamp 1678805552
transform 1 0 17184 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1064_
timestamp 1678805552
transform 1 0 17184 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1065_
timestamp 1678805552
transform 1 0 16992 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1066_
timestamp 1678805552
transform 1 0 14016 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1067_
timestamp 1678805552
transform 1 0 13920 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1068_
timestamp 1678805552
transform 1 0 13632 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1069_
timestamp 1678805552
transform 1 0 14208 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1070_
timestamp 1678805552
transform 1 0 15840 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1071_
timestamp 1678805552
transform 1 0 15648 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1072_
timestamp 1678805552
transform 1 0 10560 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1073_
timestamp 1678805552
transform 1 0 10368 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1074_
timestamp 1678805552
transform 1 0 10368 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1075_
timestamp 1678805552
transform 1 0 11712 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1076_
timestamp 1678805552
transform 1 0 11328 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1077_
timestamp 1678805552
transform 1 0 11328 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1078_
timestamp 1678805552
transform 1 0 17664 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1079_
timestamp 1678805552
transform 1 0 17664 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1080_
timestamp 1678805552
transform 1 0 17664 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1081_
timestamp 1678805552
transform 1 0 17760 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1082_
timestamp 1678805552
transform 1 0 17664 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1083_
timestamp 1678805552
transform 1 0 17376 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1084_
timestamp 1678805552
transform 1 0 15360 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1085_
timestamp 1678805552
transform 1 0 14976 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1086_
timestamp 1678805552
transform -1 0 16416 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1087_
timestamp 1678805552
transform 1 0 17376 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1088_
timestamp 1678805552
transform 1 0 17568 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1089_
timestamp 1678805552
transform 1 0 17280 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1090_
timestamp 1678805552
transform 1 0 16320 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1091_
timestamp 1678805552
transform 1 0 16224 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1092_
timestamp 1678805552
transform 1 0 16512 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1093_
timestamp 1678805552
transform 1 0 14592 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1094_
timestamp 1678805552
transform 1 0 14112 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1095_
timestamp 1678805552
transform 1 0 14016 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1096_
timestamp 1678805552
transform 1 0 1152 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1097_
timestamp 1678805552
transform 1 0 1152 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1098_
timestamp 1678805552
transform -1 0 15648 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1099_
timestamp 1678805552
transform 1 0 1920 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1100_
timestamp 1678805552
transform 1 0 2112 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1101_
timestamp 1678805552
transform -1 0 9696 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1102_
timestamp 1678805552
transform 1 0 5280 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1103_
timestamp 1678805552
transform 1 0 7008 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1104_
timestamp 1678805552
transform 1 0 5280 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1105_
timestamp 1678805552
transform 1 0 5472 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1106_
timestamp 1678805552
transform -1 0 12096 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1107_
timestamp 1678805552
transform 1 0 2880 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1108_
timestamp 1678805552
transform 1 0 1152 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1109_
timestamp 1678805552
transform 1 0 1536 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1110_
timestamp 1678805552
transform 1 0 2304 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1111_
timestamp 1678805552
transform 1 0 4896 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1112_
timestamp 1678805552
transform 1 0 3072 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1113_
timestamp 1678805552
transform 1 0 6816 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1114_
timestamp 1678805552
transform 1 0 6816 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1115_
timestamp 1678805552
transform 1 0 8640 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1116_
timestamp 1678805552
transform 1 0 4800 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1117_
timestamp 1678805552
transform 1 0 6432 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1118_
timestamp 1678805552
transform 1 0 4608 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1119_
timestamp 1678805552
transform 1 0 6336 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1120_
timestamp 1678805552
transform 1 0 5184 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1121_
timestamp 1678805552
transform 1 0 7584 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1122_
timestamp 1678805552
transform 1 0 7008 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1123_
timestamp 1678805552
transform 1 0 8832 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1124_
timestamp 1678805552
transform 1 0 5184 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1125_
timestamp 1678805552
transform 1 0 7200 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1126_
timestamp 1678805552
transform 1 0 2976 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1127_
timestamp 1678805552
transform 1 0 4608 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1128_
timestamp 1678805552
transform 1 0 4128 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1129_
timestamp 1678805552
transform 1 0 5664 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1130_
timestamp 1678805552
transform -1 0 15360 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1131_
timestamp 1678805552
transform -1 0 13728 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1132_
timestamp 1678805552
transform 1 0 1152 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1133_
timestamp 1678805552
transform -1 0 4704 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1134_
timestamp 1678805552
transform -1 0 4800 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1135_
timestamp 1678805552
transform 1 0 3168 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1136_
timestamp 1678805552
transform -1 0 13728 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1137_
timestamp 1678805552
transform 1 0 1632 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1138_
timestamp 1678805552
transform -1 0 11136 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1139_
timestamp 1678805552
transform 1 0 3072 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1140_
timestamp 1678805552
transform -1 0 17376 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1141_
timestamp 1678805552
transform -1 0 14016 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1142_
timestamp 1678805552
transform 1 0 2208 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1143_
timestamp 1678805552
transform 1 0 4224 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1144_
timestamp 1678805552
transform 1 0 4800 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1145_
timestamp 1678805552
transform 1 0 3168 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1146_
timestamp 1678805552
transform -1 0 7008 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1147_
timestamp 1678805552
transform 1 0 1536 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1148_
timestamp 1678805552
transform 1 0 1440 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1149_
timestamp 1678805552
transform 1 0 3072 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1150_
timestamp 1678805552
transform 1 0 3744 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1151_
timestamp 1678805552
transform 1 0 4512 0 1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1152_
timestamp 1678805552
transform -1 0 3936 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1153_
timestamp 1678805552
transform -1 0 6336 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1154_
timestamp 1678805552
transform -1 0 6432 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1155_
timestamp 1678805552
transform 1 0 1632 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1156_
timestamp 1678805552
transform 1 0 1152 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1157_
timestamp 1678805552
transform 1 0 1152 0 1 8316
box -50 -56 1692 834
use sg13g2_buf_1  _1158_
timestamp 1676381911
transform -1 0 4320 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1159_
timestamp 1676381911
transform 1 0 16800 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1160_
timestamp 1676381911
transform 1 0 19296 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1161_
timestamp 1676381911
transform 1 0 18048 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1162_
timestamp 1676381911
transform 1 0 19968 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1163_
timestamp 1676381911
transform 1 0 19776 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1164_
timestamp 1676381911
transform 1 0 19392 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1165_
timestamp 1676381911
transform 1 0 19680 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1166_
timestamp 1676381911
transform 1 0 16800 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1167_
timestamp 1676381911
transform 1 0 19968 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1168_
timestamp 1676381911
transform 1 0 19680 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1169_
timestamp 1676381911
transform 1 0 18528 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1170_
timestamp 1676381911
transform 1 0 19968 0 -1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1171_
timestamp 1676381911
transform 1 0 17376 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1172_
timestamp 1676381911
transform 1 0 19680 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1173_
timestamp 1676381911
transform 1 0 19680 0 1 17388
box -48 -56 432 834
use sg13g2_buf_1  _1174_
timestamp 1676381911
transform 1 0 19776 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1175_
timestamp 1676381911
transform 1 0 17952 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1176_
timestamp 1676381911
transform 1 0 19872 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1177_
timestamp 1676381911
transform 1 0 19296 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1178_
timestamp 1676381911
transform 1 0 19872 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1179_
timestamp 1676381911
transform 1 0 17376 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1180_
timestamp 1676381911
transform 1 0 13728 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1181_
timestamp 1676381911
transform 1 0 10272 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1182_
timestamp 1676381911
transform 1 0 16992 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1183_
timestamp 1676381911
transform 1 0 19776 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1184_
timestamp 1676381911
transform 1 0 18912 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1185_
timestamp 1676381911
transform 1 0 19680 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1186_
timestamp 1676381911
transform 1 0 19680 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1187_
timestamp 1676381911
transform 1 0 19296 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1188_
timestamp 1676381911
transform 1 0 19296 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1189_
timestamp 1676381911
transform 1 0 3552 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1190_
timestamp 1676381911
transform 1 0 19776 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1191_
timestamp 1676381911
transform 1 0 19392 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1192_
timestamp 1676381911
transform 1 0 19776 0 1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1193_
timestamp 1676381911
transform 1 0 19680 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1194_
timestamp 1676381911
transform 1 0 19296 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1195_
timestamp 1676381911
transform 1 0 19680 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1196_
timestamp 1676381911
transform 1 0 19392 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1197_
timestamp 1676381911
transform 1 0 19680 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1198_
timestamp 1676381911
transform 1 0 15072 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _1199_
timestamp 1676381911
transform 1 0 19296 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1200_
timestamp 1676381911
transform 1 0 19680 0 -1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1201_
timestamp 1676381911
transform 1 0 19680 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1202_
timestamp 1676381911
transform 1 0 19776 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1203_
timestamp 1676381911
transform 1 0 19296 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1204_
timestamp 1676381911
transform 1 0 19680 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1205_
timestamp 1676381911
transform 1 0 19296 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1206_
timestamp 1676381911
transform 1 0 19296 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1207_
timestamp 1676381911
transform 1 0 19392 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1208_
timestamp 1676381911
transform 1 0 19488 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1209_
timestamp 1676381911
transform 1 0 19776 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1210_
timestamp 1676381911
transform 1 0 19872 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1211_
timestamp 1676381911
transform 1 0 19008 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1212_
timestamp 1676381911
transform 1 0 1248 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1213_
timestamp 1676381911
transform 1 0 19008 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1214_
timestamp 1676381911
transform 1 0 3264 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1215_
timestamp 1676381911
transform 1 0 13344 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1216_
timestamp 1676381911
transform 1 0 4224 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1217_
timestamp 1676381911
transform 1 0 13056 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1218_
timestamp 1676381911
transform 1 0 18624 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1219_
timestamp 1676381911
transform 1 0 5952 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1220_
timestamp 1676381911
transform 1 0 19392 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1221_
timestamp 1676381911
transform 1 0 1440 0 1 18900
box -48 -56 432 834
use sg13g2_buf_1  _1222_
timestamp 1676381911
transform 1 0 13248 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1223_
timestamp 1676381911
transform 1 0 14496 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1224_
timestamp 1676381911
transform 1 0 14112 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1225_
timestamp 1676381911
transform 1 0 12960 0 1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1226_
timestamp 1676381911
transform 1 0 12288 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1227_
timestamp 1676381911
transform 1 0 14688 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1228_
timestamp 1676381911
transform 1 0 15936 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1229_
timestamp 1676381911
transform 1 0 17856 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1230_
timestamp 1676381911
transform 1 0 13248 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1231_
timestamp 1676381911
transform 1 0 9120 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1232_
timestamp 1676381911
transform 1 0 12096 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1233_
timestamp 1676381911
transform 1 0 9696 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1234_
timestamp 1676381911
transform 1 0 17376 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1235_
timestamp 1676381911
transform 1 0 6912 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1236_
timestamp 1676381911
transform 1 0 16992 0 -1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1237_
timestamp 1676381911
transform 1 0 7200 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1238_
timestamp 1676381911
transform 1 0 12864 0 -1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1239_
timestamp 1676381911
transform -1 0 19776 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1240_
timestamp 1676381911
transform -1 0 20064 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1241_
timestamp 1676381911
transform -1 0 20160 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1242_
timestamp 1676381911
transform -1 0 20160 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1243_
timestamp 1676381911
transform -1 0 18816 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1244_
timestamp 1676381911
transform -1 0 17472 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1245_
timestamp 1676381911
transform -1 0 19776 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1246_
timestamp 1676381911
transform 1 0 7776 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1247_
timestamp 1676381911
transform 1 0 1728 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1248_
timestamp 1676381911
transform 1 0 1152 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1249_
timestamp 1676381911
transform -1 0 19776 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1250_
timestamp 1676381911
transform -1 0 20160 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1251_
timestamp 1676381911
transform 1 0 4224 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _1252_
timestamp 1676381911
transform 1 0 6432 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1253_
timestamp 1676381911
transform 1 0 7008 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1254_
timestamp 1676381911
transform 1 0 9504 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1255_
timestamp 1676381911
transform 1 0 9312 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1256_
timestamp 1676381911
transform 1 0 12672 0 1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1257_
timestamp 1676381911
transform 1 0 15264 0 1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1258_
timestamp 1676381911
transform 1 0 14400 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1259_
timestamp 1676381911
transform -1 0 2016 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1260_
timestamp 1676381911
transform 1 0 1248 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1261_
timestamp 1676381911
transform 1 0 1152 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1262_
timestamp 1676381911
transform -1 0 3168 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1263_
timestamp 1676381911
transform -1 0 5184 0 -1 30996
box -48 -56 432 834
use sg13g2_buf_1  _1264_
timestamp 1676381911
transform -1 0 3168 0 -1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1265_
timestamp 1676381911
transform 1 0 1440 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1266_
timestamp 1676381911
transform -1 0 4800 0 -1 26460
box -48 -56 432 834
use sg13g2_buf_1  _1267_
timestamp 1676381911
transform 1 0 1344 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1268_
timestamp 1676381911
transform 1 0 2304 0 1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1269_
timestamp 1676381911
transform -1 0 4704 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1270_
timestamp 1676381911
transform 1 0 1248 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1271_
timestamp 1676381911
transform 1 0 1248 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1272_
timestamp 1676381911
transform 1 0 3936 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1273_
timestamp 1676381911
transform 1 0 3072 0 1 34020
box -48 -56 432 834
use sg13g2_buf_1  _1274_
timestamp 1676381911
transform 1 0 1632 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1275_
timestamp 1676381911
transform 1 0 2112 0 1 32508
box -48 -56 432 834
use sg13g2_buf_1  _1276_
timestamp 1676381911
transform 1 0 1248 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1277_
timestamp 1676381911
transform 1 0 2016 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1278_
timestamp 1676381911
transform 1 0 4704 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1279_
timestamp 1676381911
transform -1 0 7776 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1280_
timestamp 1676381911
transform 1 0 1632 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1281_
timestamp 1676381911
transform 1 0 3936 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1282_
timestamp 1676381911
transform 1 0 3744 0 -1 35532
box -48 -56 432 834
use sg13g2_buf_1  _1283_
timestamp 1676381911
transform 1 0 1248 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1284_
timestamp 1676381911
transform 1 0 4224 0 1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1285_
timestamp 1676381911
transform 1 0 5952 0 1 24948
box -48 -56 432 834
use sg13g2_buf_1  _1286_
timestamp 1676381911
transform 1 0 5472 0 -1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1287_
timestamp 1676381911
transform 1 0 6816 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1288_
timestamp 1676381911
transform 1 0 1248 0 1 20412
box -48 -56 432 834
use sg13g2_buf_1  _1289_
timestamp 1676381911
transform 1 0 2784 0 -1 29484
box -48 -56 432 834
use sg13g2_buf_1  _1290_
timestamp 1676381911
transform -1 0 8544 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1291_
timestamp 1676381911
transform 1 0 3552 0 1 27972
box -48 -56 432 834
use sg13g2_buf_1  _1292_
timestamp 1676381911
transform -1 0 18240 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1293_
timestamp 1676381911
transform -1 0 10656 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1294_
timestamp 1676381911
transform 1 0 6336 0 -1 23436
box -48 -56 432 834
use sg13g2_buf_1  _1295_
timestamp 1676381911
transform 1 0 2784 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1296_
timestamp 1676381911
transform 1 0 1440 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1297_
timestamp 1676381911
transform -1 0 11232 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1298_
timestamp 1676381911
transform 1 0 1152 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1299_
timestamp 1676381911
transform -1 0 11616 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1300_
timestamp 1676381911
transform -1 0 17856 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1301_
timestamp 1676381911
transform 1 0 6912 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1302_
timestamp 1676381911
transform 1 0 9888 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1303_
timestamp 1676381911
transform 1 0 5856 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1304_
timestamp 1676381911
transform 1 0 9984 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1305_
timestamp 1676381911
transform 1 0 4800 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1306_
timestamp 1676381911
transform 1 0 4992 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1307_
timestamp 1676381911
transform 1 0 5568 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1308_
timestamp 1676381911
transform 1 0 9216 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1309_
timestamp 1676381911
transform 1 0 9504 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1310_
timestamp 1676381911
transform 1 0 10656 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1311_
timestamp 1676381911
transform -1 0 12000 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1312_
timestamp 1676381911
transform 1 0 11520 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1313_
timestamp 1676381911
transform 1 0 11136 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1314_
timestamp 1676381911
transform 1 0 11520 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1315_
timestamp 1676381911
transform -1 0 17856 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1316_
timestamp 1676381911
transform -1 0 18624 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1317_
timestamp 1676381911
transform -1 0 19008 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1318_
timestamp 1676381911
transform -1 0 19392 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1319_
timestamp 1676381911
transform -1 0 18432 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1320_
timestamp 1676381911
transform 1 0 4320 0 1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1321_
timestamp 1676381911
transform -1 0 18048 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1322_
timestamp 1676381911
transform 1 0 1152 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1323_
timestamp 1676381911
transform -1 0 19296 0 1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1324_
timestamp 1676381911
transform 1 0 4896 0 1 37044
box -48 -56 432 834
use sg13g2_buf_1  _1325_
timestamp 1676381911
transform -1 0 18624 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1326_
timestamp 1676381911
transform -1 0 19008 0 -1 40068
box -48 -56 432 834
use sg13g2_buf_1  _1327_
timestamp 1676381911
transform -1 0 19968 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1328_
timestamp 1676381911
transform 1 0 5184 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1329_
timestamp 1676381911
transform -1 0 20352 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1330_
timestamp 1676381911
transform 1 0 11040 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1331_
timestamp 1676381911
transform -1 0 19680 0 1 40068
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 20064 0 1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 20064 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 6240 0 1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform -1 0 1440 0 -1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 3360 0 -1 27972
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 4800 0 1 27972
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform -1 0 3936 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform -1 0 4800 0 1 27972
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform -1 0 4800 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform 1 0 1632 0 1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform -1 0 4992 0 1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 4224 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform 1 0 20064 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 6144 0 1 8316
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform 1 0 6144 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform -1 0 1440 0 1 18900
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 5856 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 1344 0 -1 18900
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform 1 0 9696 0 1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform -1 0 1440 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform 1 0 9216 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform -1 0 4224 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 7296 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform -1 0 4224 0 1 23436
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform 1 0 12000 0 1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 10272 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform -1 0 4992 0 -1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform 1 0 16224 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform -1 0 4800 0 1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform 1 0 15072 0 1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform -1 0 2304 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform 1 0 1536 0 -1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 1344 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform -1 0 1536 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform 1 0 1632 0 -1 18900
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform 1 0 19392 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform -1 0 1440 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform 1 0 4608 0 1 21924
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 1536 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform 1 0 15936 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform -1 0 14112 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform 1 0 8736 0 1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 9216 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform 1 0 4416 0 1 12852
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform -1 0 1440 0 -1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform 1 0 1632 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_47
timestamp 1679999689
transform -1 0 3072 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_48
timestamp 1679999689
transform 1 0 6432 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_49
timestamp 1679999689
transform 1 0 3648 0 1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_50
timestamp 1679999689
transform -1 0 4800 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_51
timestamp 1679999689
transform 1 0 6432 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_52
timestamp 1679999689
transform -1 0 3072 0 1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_53
timestamp 1679999689
transform 1 0 4704 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_54
timestamp 1679999689
transform 1 0 6432 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_55
timestamp 1679999689
transform 1 0 3648 0 -1 26460
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_56
timestamp 1679999689
transform 1 0 5568 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_57
timestamp 1679999689
transform 1 0 1824 0 -1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_58
timestamp 1679999689
transform -1 0 2304 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_59
timestamp 1679999689
transform 1 0 1824 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_60
timestamp 1679999689
transform 1 0 4608 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_61
timestamp 1679999689
transform 1 0 4992 0 1 18900
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_62
timestamp 1679999689
transform 1 0 4704 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_63
timestamp 1679999689
transform 1 0 4992 0 1 20412
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_64
timestamp 1679999689
transform -1 0 4800 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_65
timestamp 1679999689
transform 1 0 4128 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_66
timestamp 1679999689
transform -1 0 4128 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_67
timestamp 1679999689
transform -1 0 4416 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_68
timestamp 1679999689
transform -1 0 4128 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_69
timestamp 1679999689
transform -1 0 7008 0 -1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_70
timestamp 1679999689
transform 1 0 3456 0 -1 34020
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_71
timestamp 1679999689
transform -1 0 4224 0 1 37044
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_72
timestamp 1679999689
transform 1 0 3456 0 -1 35532
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_73
timestamp 1679999689
transform -1 0 4224 0 1 38556
box -48 -56 336 834
use sg13g2_buf_8  clkbuf_0_UserCLK
timestamp 1676451365
transform -1 0 11808 0 1 32508
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_UserCLK
timestamp 1676451365
transform -1 0 9312 0 -1 30996
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_UserCLK
timestamp 1676451365
transform 1 0 11424 0 -1 35532
box -48 -56 1296 834
use sg13g2_fill_1  FILLER_0_34
timestamp 1677579658
transform 1 0 4416 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_0_174
timestamp 1677579658
transform 1 0 17856 0 1 756
box -48 -56 144 834
use sg13g2_fill_1  FILLER_1_27
timestamp 1677579658
transform 1 0 3744 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_151
timestamp 1677580104
transform 1 0 15648 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_191
timestamp 1677579658
transform 1 0 19488 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_0
timestamp 1677579658
transform 1 0 1152 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_27
timestamp 1677579658
transform 1 0 3744 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_36
timestamp 1677579658
transform 1 0 4608 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_108
timestamp 1677579658
transform 1 0 11520 0 1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_173
timestamp 1677580104
transform 1 0 17760 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_3_0
timestamp 1677580104
transform 1 0 1152 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_30
timestamp 1677579658
transform 1 0 4032 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_75
timestamp 1677579658
transform 1 0 8352 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_97
timestamp 1677580104
transform 1 0 10464 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_112
timestamp 1677579658
transform 1 0 11904 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_199
timestamp 1677579658
transform 1 0 20256 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_112
timestamp 1677579658
transform 1 0 11904 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_135
timestamp 1677579658
transform 1 0 14112 0 1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_4_199
timestamp 1677579658
transform 1 0 20256 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_58
timestamp 1677580104
transform 1 0 6720 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_72
timestamp 1677580104
transform 1 0 8064 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_5_129
timestamp 1677579658
transform 1 0 13536 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_5_170
timestamp 1677580104
transform 1 0 17472 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_177
timestamp 1677580104
transform 1 0 18144 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_2  FILLER_5_198
timestamp 1677580104
transform 1 0 20160 0 -1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_33
timestamp 1677579658
transform 1 0 4320 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_121
timestamp 1677579658
transform 1 0 12768 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_52
timestamp 1677580104
transform 1 0 6144 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_135
timestamp 1677579658
transform 1 0 14112 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_171
timestamp 1677579658
transform 1 0 17568 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_199
timestamp 1677579658
transform 1 0 20256 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_65
timestamp 1677580104
transform 1 0 7392 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_142
timestamp 1677579658
transform 1 0 14784 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_171
timestamp 1677580104
transform 1 0 17568 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_8_198
timestamp 1677580104
transform 1 0 20160 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_17
timestamp 1677579658
transform 1 0 2784 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_47
timestamp 1677579658
transform 1 0 5664 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_9_69
timestamp 1677580104
transform 1 0 7776 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_94
timestamp 1677580104
transform 1 0 10176 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_9_118
timestamp 1677579658
transform 1 0 12480 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_137
timestamp 1677579658
transform 1 0 14304 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_9_174
timestamp 1677579658
transform 1 0 17856 0 -1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_126
timestamp 1677579658
transform 1 0 13248 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_164
timestamp 1677579658
transform 1 0 16896 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_10_199
timestamp 1677579658
transform 1 0 20256 0 1 8316
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_0
timestamp 1677579658
transform 1 0 1152 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_97
timestamp 1677579658
transform 1 0 10464 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_127
timestamp 1677579658
transform 1 0 13344 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_11_149
timestamp 1677579658
transform 1 0 15456 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_180
timestamp 1677580104
transform 1 0 18432 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_48
timestamp 1677579658
transform 1 0 5760 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_66
timestamp 1677580104
transform 1 0 7488 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_145
timestamp 1677579658
transform 1 0 15072 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_170
timestamp 1677579658
transform 1 0 17472 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_198
timestamp 1677580104
transform 1 0 20160 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_0
timestamp 1677579658
transform 1 0 1152 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_23
timestamp 1677579658
transform 1 0 3360 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_122
timestamp 1677579658
transform 1 0 12864 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_13_140
timestamp 1677579658
transform 1 0 14592 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_84
timestamp 1677579658
transform 1 0 9216 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_159
timestamp 1677579658
transform 1 0 16416 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_168
timestamp 1677579658
transform 1 0 17280 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_198
timestamp 1677580104
transform 1 0 20160 0 1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_17
timestamp 1677579658
transform 1 0 2784 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_96
timestamp 1677580104
transform 1 0 10368 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_103
timestamp 1677579658
transform 1 0 11040 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_184
timestamp 1677580104
transform 1 0 18816 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_37
timestamp 1677579658
transform 1 0 4704 0 1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_16_93
timestamp 1677580104
transform 1 0 10080 0 1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_16_112
timestamp 1677579658
transform 1 0 11904 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_17_64
timestamp 1677579658
transform 1 0 7296 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_0
timestamp 1677579658
transform 1 0 1152 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_57
timestamp 1677579658
transform 1 0 6624 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_63
timestamp 1677580104
transform 1 0 7200 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_65
timestamp 1677579658
transform 1 0 7392 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_144
timestamp 1677580104
transform 1 0 14976 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_146
timestamp 1677579658
transform 1 0 15168 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_174
timestamp 1677580104
transform 1 0 17856 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_185
timestamp 1677579658
transform 1 0 18912 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_147
timestamp 1677580104
transform 1 0 15264 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_19_149
timestamp 1677579658
transform 1 0 15456 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_198
timestamp 1677580104
transform 1 0 20160 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_34
timestamp 1677579658
transform 1 0 4416 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_60
timestamp 1677579658
transform 1 0 6912 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_103
timestamp 1679577901
transform 1 0 11040 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_107
timestamp 1677579658
transform 1 0 11424 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_125
timestamp 1677580104
transform 1 0 13152 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_127
timestamp 1677579658
transform 1 0 13344 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_20_186
timestamp 1677579658
transform 1 0 19008 0 1 15876
box -48 -56 144 834
use sg13g2_fill_1  FILLER_21_0
timestamp 1677579658
transform 1 0 1152 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_32
timestamp 1677580104
transform 1 0 4224 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_75
timestamp 1677580104
transform 1 0 8352 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_104
timestamp 1677580104
transform 1 0 11136 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_21_123
timestamp 1677580104
transform 1 0 12960 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_125
timestamp 1677579658
transform 1 0 13152 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_21_136
timestamp 1677580104
transform 1 0 14208 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_167
timestamp 1677579658
transform 1 0 17184 0 -1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_22_85
timestamp 1677580104
transform 1 0 9312 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_104
timestamp 1677580104
transform 1 0 11136 0 1 17388
box -48 -56 240 834
use sg13g2_fill_2  FILLER_22_197
timestamp 1677580104
transform 1 0 20064 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_199
timestamp 1677579658
transform 1 0 20256 0 1 17388
box -48 -56 144 834
use sg13g2_fill_2  FILLER_23_0
timestamp 1677580104
transform 1 0 1152 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_11
timestamp 1677580104
transform 1 0 2208 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_13
timestamp 1677579658
transform 1 0 2400 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_62
timestamp 1679581782
transform 1 0 7104 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_69
timestamp 1677580104
transform 1 0 7776 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_171
timestamp 1677579658
transform 1 0 17568 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_24_7
timestamp 1679581782
transform 1 0 1824 0 1 18900
box -48 -56 720 834
use sg13g2_fill_1  FILLER_24_14
timestamp 1677579658
transform 1 0 2496 0 1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_36
timestamp 1679577901
transform 1 0 4608 0 1 18900
box -48 -56 432 834
use sg13g2_decap_4  FILLER_24_43
timestamp 1679577901
transform 1 0 5280 0 1 18900
box -48 -56 432 834
use sg13g2_decap_4  FILLER_24_81
timestamp 1679577901
transform 1 0 8928 0 1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_24_85
timestamp 1677580104
transform 1 0 9312 0 1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_24_125
timestamp 1677579658
transform 1 0 13152 0 1 18900
box -48 -56 144 834
use sg13g2_fill_1  FILLER_24_199
timestamp 1677579658
transform 1 0 20256 0 1 18900
box -48 -56 144 834
use sg13g2_decap_8  FILLER_25_82
timestamp 1679581782
transform 1 0 9024 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_25_89
timestamp 1677579658
transform 1 0 9696 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_111
timestamp 1677580104
transform 1 0 11808 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_113
timestamp 1677579658
transform 1 0 12000 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_25_147
timestamp 1677579658
transform 1 0 15264 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_25_171
timestamp 1677580104
transform 1 0 17568 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_199
timestamp 1677579658
transform 1 0 20256 0 -1 20412
box -48 -56 144 834
use sg13g2_fill_1  FILLER_26_0
timestamp 1677579658
transform 1 0 1152 0 1 20412
box -48 -56 144 834
use sg13g2_fill_2  FILLER_26_8
timestamp 1677580104
transform 1 0 1920 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_10
timestamp 1677579658
transform 1 0 2112 0 1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_26_36
timestamp 1679577901
transform 1 0 4608 0 1 20412
box -48 -56 432 834
use sg13g2_decap_8  FILLER_26_60
timestamp 1679581782
transform 1 0 6912 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_67
timestamp 1679577901
transform 1 0 7584 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_143
timestamp 1677580104
transform 1 0 14880 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_184
timestamp 1677580104
transform 1 0 18816 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_0
timestamp 1677579658
transform 1 0 1152 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_44
timestamp 1679577901
transform 1 0 5376 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_2  FILLER_27_48
timestamp 1677580104
transform 1 0 5760 0 -1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_27_105
timestamp 1679581782
transform 1 0 11232 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_112
timestamp 1677580104
transform 1 0 11904 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_114
timestamp 1677579658
transform 1 0 12096 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_27_198
timestamp 1677580104
transform 1 0 20160 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_0
timestamp 1677579658
transform 1 0 1152 0 1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_28_77
timestamp 1679577901
transform 1 0 8544 0 1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_28_81
timestamp 1677579658
transform 1 0 8928 0 1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_124
timestamp 1677580104
transform 1 0 13056 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_151
timestamp 1677580104
transform 1 0 15648 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_199
timestamp 1677579658
transform 1 0 20256 0 1 21924
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_0
timestamp 1677579658
transform 1 0 1152 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_27
timestamp 1677580104
transform 1 0 3744 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_29_58
timestamp 1677580104
transform 1 0 6720 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_60
timestamp 1677579658
transform 1 0 6912 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_78
timestamp 1679581782
transform 1 0 8640 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_1  FILLER_29_85
timestamp 1677579658
transform 1 0 9312 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_29_103
timestamp 1677580104
transform 1 0 11040 0 -1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_29_105
timestamp 1677579658
transform 1 0 11232 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_123
timestamp 1677579658
transform 1 0 12960 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_145
timestamp 1677579658
transform 1 0 15072 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_163
timestamp 1677579658
transform 1 0 16800 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_0
timestamp 1677579658
transform 1 0 1152 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_28
timestamp 1677579658
transform 1 0 3840 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_49
timestamp 1677579658
transform 1 0 5856 0 1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_71
timestamp 1679581782
transform 1 0 7968 0 1 23436
box -48 -56 720 834
use sg13g2_decap_4  FILLER_30_78
timestamp 1679577901
transform 1 0 8640 0 1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_30_82
timestamp 1677579658
transform 1 0 9024 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_104
timestamp 1677579658
transform 1 0 11136 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_122
timestamp 1677579658
transform 1 0 12864 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_164
timestamp 1677579658
transform 1 0 16896 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_199
timestamp 1677579658
transform 1 0 20256 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_17
timestamp 1677580104
transform 1 0 2784 0 -1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_74
timestamp 1679577901
transform 1 0 8256 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_31_140
timestamp 1677579658
transform 1 0 14592 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_162
timestamp 1677580104
transform 1 0 16704 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_164
timestamp 1677579658
transform 1 0 16896 0 -1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_31_198
timestamp 1677580104
transform 1 0 20160 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_21
timestamp 1677580104
transform 1 0 3168 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_44
timestamp 1677579658
transform 1 0 5376 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_88
timestamp 1679581782
transform 1 0 9600 0 1 24948
box -48 -56 720 834
use sg13g2_fill_1  FILLER_32_137
timestamp 1677579658
transform 1 0 14304 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_163
timestamp 1677580104
transform 1 0 16800 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_165
timestamp 1677579658
transform 1 0 16992 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_32_187
timestamp 1677580104
transform 1 0 19104 0 1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_32_197
timestamp 1677580104
transform 1 0 20064 0 1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_32_199
timestamp 1677579658
transform 1 0 20256 0 1 24948
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_33
timestamp 1677579658
transform 1 0 4320 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_33_175
timestamp 1677579658
transform 1 0 17952 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_197
timestamp 1677580104
transform 1 0 20064 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_199
timestamp 1677579658
transform 1 0 20256 0 -1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_34
timestamp 1677580104
transform 1 0 4416 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_77
timestamp 1677579658
transform 1 0 8544 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_34_146
timestamp 1677579658
transform 1 0 15168 0 1 26460
box -48 -56 144 834
use sg13g2_fill_2  FILLER_34_197
timestamp 1677580104
transform 1 0 20064 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_199
timestamp 1677579658
transform 1 0 20256 0 1 26460
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_0
timestamp 1677579658
transform 1 0 1152 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_91
timestamp 1677580104
transform 1 0 9888 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_115
timestamp 1677580104
transform 1 0 12192 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_164
timestamp 1677579658
transform 1 0 16896 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_35_198
timestamp 1677580104
transform 1 0 20160 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_33
timestamp 1677580104
transform 1 0 4320 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_41
timestamp 1677579658
transform 1 0 5088 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_100
timestamp 1677580104
transform 1 0 10752 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_127
timestamp 1677579658
transform 1 0 13344 0 1 27972
box -48 -56 144 834
use sg13g2_fill_2  FILLER_36_187
timestamp 1677580104
transform 1 0 19104 0 1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_36_197
timestamp 1677580104
transform 1 0 20064 0 1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_36_199
timestamp 1677579658
transform 1 0 20256 0 1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_94
timestamp 1677579658
transform 1 0 10176 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_128
timestamp 1677580104
transform 1 0 13440 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_169
timestamp 1677579658
transform 1 0 17376 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_187
timestamp 1677580104
transform 1 0 19104 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_2  FILLER_37_197
timestamp 1677580104
transform 1 0 20064 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_199
timestamp 1677579658
transform 1 0 20256 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_37
timestamp 1677579658
transform 1 0 4704 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_55
timestamp 1677580104
transform 1 0 6432 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_74
timestamp 1677579658
transform 1 0 8256 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_92
timestamp 1677579658
transform 1 0 9984 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_188
timestamp 1677579658
transform 1 0 19200 0 1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_38_197
timestamp 1677580104
transform 1 0 20064 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_199
timestamp 1677579658
transform 1 0 20256 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_39_135
timestamp 1677579658
transform 1 0 14112 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_174
timestamp 1677580104
transform 1 0 17856 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_176
timestamp 1677579658
transform 1 0 18048 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_198
timestamp 1677580104
transform 1 0 20160 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_54
timestamp 1677580104
transform 1 0 6336 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_99
timestamp 1677580104
transform 1 0 10656 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_40_139
timestamp 1677580104
transform 1 0 14496 0 1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_40_141
timestamp 1677579658
transform 1 0 14688 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_168
timestamp 1677579658
transform 1 0 17280 0 1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_40_198
timestamp 1677580104
transform 1 0 20160 0 1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_80
timestamp 1677580104
transform 1 0 8832 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_129
timestamp 1677579658
transform 1 0 13536 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_41_135
timestamp 1677580104
transform 1 0 14112 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_142
timestamp 1677580104
transform 1 0 14784 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_154
timestamp 1677580104
transform 1 0 15936 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_197
timestamp 1677580104
transform 1 0 20064 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_199
timestamp 1677579658
transform 1 0 20256 0 -1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_0
timestamp 1677580104
transform 1 0 1152 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_128
timestamp 1677579658
transform 1 0 13440 0 1 32508
box -48 -56 144 834
use sg13g2_fill_2  FILLER_42_160
timestamp 1677580104
transform 1 0 16512 0 1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_42_162
timestamp 1677579658
transform 1 0 16704 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_42_188
timestamp 1677579658
transform 1 0 19200 0 1 32508
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_0
timestamp 1677579658
transform 1 0 1152 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_6
timestamp 1677579658
transform 1 0 1728 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_60
timestamp 1677579658
transform 1 0 6912 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_78
timestamp 1677580104
transform 1 0 8640 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_114
timestamp 1677580104
transform 1 0 12096 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_43_167
timestamp 1677580104
transform 1 0 17184 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_45
timestamp 1677580104
transform 1 0 5472 0 1 34020
box -48 -56 240 834
use sg13g2_fill_2  FILLER_44_121
timestamp 1677580104
transform 1 0 12768 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_199
timestamp 1677579658
transform 1 0 20256 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_45_189
timestamp 1677579658
transform 1 0 19296 0 -1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_45_198
timestamp 1677580104
transform 1 0 20160 0 -1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_0
timestamp 1677580104
transform 1 0 1152 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_10
timestamp 1677580104
transform 1 0 2112 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_114
timestamp 1677580104
transform 1 0 12096 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_170
timestamp 1677580104
transform 1 0 17472 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_0
timestamp 1677579658
transform 1 0 1152 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_43
timestamp 1677580104
transform 1 0 5280 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_133
timestamp 1677579658
transform 1 0 13920 0 -1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_151
timestamp 1677580104
transform 1 0 15648 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_171
timestamp 1677580104
transform 1 0 17568 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_198
timestamp 1677580104
transform 1 0 20160 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_48_147
timestamp 1677580104
transform 1 0 15264 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_165
timestamp 1677579658
transform 1 0 16992 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_0
timestamp 1677579658
transform 1 0 1152 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_61
timestamp 1677580104
transform 1 0 7008 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_2  FILLER_49_175
timestamp 1677580104
transform 1 0 17952 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_199
timestamp 1677579658
transform 1 0 20256 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_50_0
timestamp 1677579658
transform 1 0 1152 0 1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_50_32
timestamp 1677579658
transform 1 0 4224 0 1 38556
box -48 -56 144 834
use sg13g2_fill_1  FILLER_50_41
timestamp 1677579658
transform 1 0 5088 0 1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_198
timestamp 1677580104
transform 1 0 20160 0 1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_125
timestamp 1677579658
transform 1 0 13152 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_148
timestamp 1677579658
transform 1 0 15360 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_51_198
timestamp 1677580104
transform 1 0 20160 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_0
timestamp 1677579658
transform 1 0 1152 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_76
timestamp 1677580104
transform 1 0 8448 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_184
timestamp 1677579658
transform 1 0 18816 0 1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_53_38
timestamp 1677579658
transform 1 0 4800 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_78
timestamp 1677580104
transform 1 0 8640 0 -1 41580
box -48 -56 240 834
use sg13g2_fill_2  FILLER_53_198
timestamp 1677580104
transform 1 0 20160 0 -1 41580
box -48 -56 240 834
<< labels >>
flabel metal3 s 0 23396 80 23476 0 FreeSans 320 0 0 0 CLK_TT_PROJECT
port 0 nsew signal output
flabel metal3 s 21424 16172 21504 16252 0 FreeSans 320 0 0 0 E1BEG[0]
port 1 nsew signal output
flabel metal3 s 21424 16508 21504 16588 0 FreeSans 320 0 0 0 E1BEG[1]
port 2 nsew signal output
flabel metal3 s 21424 16844 21504 16924 0 FreeSans 320 0 0 0 E1BEG[2]
port 3 nsew signal output
flabel metal3 s 21424 17180 21504 17260 0 FreeSans 320 0 0 0 E1BEG[3]
port 4 nsew signal output
flabel metal3 s 21424 17516 21504 17596 0 FreeSans 320 0 0 0 E2BEG[0]
port 5 nsew signal output
flabel metal3 s 21424 17852 21504 17932 0 FreeSans 320 0 0 0 E2BEG[1]
port 6 nsew signal output
flabel metal3 s 21424 18188 21504 18268 0 FreeSans 320 0 0 0 E2BEG[2]
port 7 nsew signal output
flabel metal3 s 21424 18524 21504 18604 0 FreeSans 320 0 0 0 E2BEG[3]
port 8 nsew signal output
flabel metal3 s 21424 18860 21504 18940 0 FreeSans 320 0 0 0 E2BEG[4]
port 9 nsew signal output
flabel metal3 s 21424 19196 21504 19276 0 FreeSans 320 0 0 0 E2BEG[5]
port 10 nsew signal output
flabel metal3 s 21424 19532 21504 19612 0 FreeSans 320 0 0 0 E2BEG[6]
port 11 nsew signal output
flabel metal3 s 21424 19868 21504 19948 0 FreeSans 320 0 0 0 E2BEG[7]
port 12 nsew signal output
flabel metal3 s 21424 20204 21504 20284 0 FreeSans 320 0 0 0 E2BEGb[0]
port 13 nsew signal output
flabel metal3 s 21424 20540 21504 20620 0 FreeSans 320 0 0 0 E2BEGb[1]
port 14 nsew signal output
flabel metal3 s 21424 20876 21504 20956 0 FreeSans 320 0 0 0 E2BEGb[2]
port 15 nsew signal output
flabel metal3 s 21424 21212 21504 21292 0 FreeSans 320 0 0 0 E2BEGb[3]
port 16 nsew signal output
flabel metal3 s 21424 21548 21504 21628 0 FreeSans 320 0 0 0 E2BEGb[4]
port 17 nsew signal output
flabel metal3 s 21424 21884 21504 21964 0 FreeSans 320 0 0 0 E2BEGb[5]
port 18 nsew signal output
flabel metal3 s 21424 22220 21504 22300 0 FreeSans 320 0 0 0 E2BEGb[6]
port 19 nsew signal output
flabel metal3 s 21424 22556 21504 22636 0 FreeSans 320 0 0 0 E2BEGb[7]
port 20 nsew signal output
flabel metal3 s 21424 28268 21504 28348 0 FreeSans 320 0 0 0 E6BEG[0]
port 21 nsew signal output
flabel metal3 s 21424 31628 21504 31708 0 FreeSans 320 0 0 0 E6BEG[10]
port 22 nsew signal output
flabel metal3 s 21424 31964 21504 32044 0 FreeSans 320 0 0 0 E6BEG[11]
port 23 nsew signal output
flabel metal3 s 21424 28604 21504 28684 0 FreeSans 320 0 0 0 E6BEG[1]
port 24 nsew signal output
flabel metal3 s 21424 28940 21504 29020 0 FreeSans 320 0 0 0 E6BEG[2]
port 25 nsew signal output
flabel metal3 s 21424 29276 21504 29356 0 FreeSans 320 0 0 0 E6BEG[3]
port 26 nsew signal output
flabel metal3 s 21424 29612 21504 29692 0 FreeSans 320 0 0 0 E6BEG[4]
port 27 nsew signal output
flabel metal3 s 21424 29948 21504 30028 0 FreeSans 320 0 0 0 E6BEG[5]
port 28 nsew signal output
flabel metal3 s 21424 30284 21504 30364 0 FreeSans 320 0 0 0 E6BEG[6]
port 29 nsew signal output
flabel metal3 s 21424 30620 21504 30700 0 FreeSans 320 0 0 0 E6BEG[7]
port 30 nsew signal output
flabel metal3 s 21424 30956 21504 31036 0 FreeSans 320 0 0 0 E6BEG[8]
port 31 nsew signal output
flabel metal3 s 21424 31292 21504 31372 0 FreeSans 320 0 0 0 E6BEG[9]
port 32 nsew signal output
flabel metal3 s 21424 22892 21504 22972 0 FreeSans 320 0 0 0 EE4BEG[0]
port 33 nsew signal output
flabel metal3 s 21424 26252 21504 26332 0 FreeSans 320 0 0 0 EE4BEG[10]
port 34 nsew signal output
flabel metal3 s 21424 26588 21504 26668 0 FreeSans 320 0 0 0 EE4BEG[11]
port 35 nsew signal output
flabel metal3 s 21424 26924 21504 27004 0 FreeSans 320 0 0 0 EE4BEG[12]
port 36 nsew signal output
flabel metal3 s 21424 27260 21504 27340 0 FreeSans 320 0 0 0 EE4BEG[13]
port 37 nsew signal output
flabel metal3 s 21424 27596 21504 27676 0 FreeSans 320 0 0 0 EE4BEG[14]
port 38 nsew signal output
flabel metal3 s 21424 27932 21504 28012 0 FreeSans 320 0 0 0 EE4BEG[15]
port 39 nsew signal output
flabel metal3 s 21424 23228 21504 23308 0 FreeSans 320 0 0 0 EE4BEG[1]
port 40 nsew signal output
flabel metal3 s 21424 23564 21504 23644 0 FreeSans 320 0 0 0 EE4BEG[2]
port 41 nsew signal output
flabel metal3 s 21424 23900 21504 23980 0 FreeSans 320 0 0 0 EE4BEG[3]
port 42 nsew signal output
flabel metal3 s 21424 24236 21504 24316 0 FreeSans 320 0 0 0 EE4BEG[4]
port 43 nsew signal output
flabel metal3 s 21424 24572 21504 24652 0 FreeSans 320 0 0 0 EE4BEG[5]
port 44 nsew signal output
flabel metal3 s 21424 24908 21504 24988 0 FreeSans 320 0 0 0 EE4BEG[6]
port 45 nsew signal output
flabel metal3 s 21424 25244 21504 25324 0 FreeSans 320 0 0 0 EE4BEG[7]
port 46 nsew signal output
flabel metal3 s 21424 25580 21504 25660 0 FreeSans 320 0 0 0 EE4BEG[8]
port 47 nsew signal output
flabel metal3 s 21424 25916 21504 25996 0 FreeSans 320 0 0 0 EE4BEG[9]
port 48 nsew signal output
flabel metal3 s 0 22892 80 22972 0 FreeSans 320 0 0 0 ENA_TT_PROJECT
port 49 nsew signal output
flabel metal3 s 0 24404 80 24484 0 FreeSans 320 0 0 0 FrameData[0]
port 50 nsew signal input
flabel metal3 s 0 29444 80 29524 0 FreeSans 320 0 0 0 FrameData[10]
port 51 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 FrameData[11]
port 52 nsew signal input
flabel metal3 s 0 30452 80 30532 0 FreeSans 320 0 0 0 FrameData[12]
port 53 nsew signal input
flabel metal3 s 0 30956 80 31036 0 FreeSans 320 0 0 0 FrameData[13]
port 54 nsew signal input
flabel metal3 s 0 31460 80 31540 0 FreeSans 320 0 0 0 FrameData[14]
port 55 nsew signal input
flabel metal3 s 0 31964 80 32044 0 FreeSans 320 0 0 0 FrameData[15]
port 56 nsew signal input
flabel metal3 s 0 32468 80 32548 0 FreeSans 320 0 0 0 FrameData[16]
port 57 nsew signal input
flabel metal3 s 0 32972 80 33052 0 FreeSans 320 0 0 0 FrameData[17]
port 58 nsew signal input
flabel metal3 s 0 33476 80 33556 0 FreeSans 320 0 0 0 FrameData[18]
port 59 nsew signal input
flabel metal3 s 0 33980 80 34060 0 FreeSans 320 0 0 0 FrameData[19]
port 60 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 FrameData[1]
port 61 nsew signal input
flabel metal3 s 0 34484 80 34564 0 FreeSans 320 0 0 0 FrameData[20]
port 62 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 FrameData[21]
port 63 nsew signal input
flabel metal3 s 0 35492 80 35572 0 FreeSans 320 0 0 0 FrameData[22]
port 64 nsew signal input
flabel metal3 s 0 35996 80 36076 0 FreeSans 320 0 0 0 FrameData[23]
port 65 nsew signal input
flabel metal3 s 0 36500 80 36580 0 FreeSans 320 0 0 0 FrameData[24]
port 66 nsew signal input
flabel metal3 s 0 37004 80 37084 0 FreeSans 320 0 0 0 FrameData[25]
port 67 nsew signal input
flabel metal3 s 0 37508 80 37588 0 FreeSans 320 0 0 0 FrameData[26]
port 68 nsew signal input
flabel metal3 s 0 38012 80 38092 0 FreeSans 320 0 0 0 FrameData[27]
port 69 nsew signal input
flabel metal3 s 0 38516 80 38596 0 FreeSans 320 0 0 0 FrameData[28]
port 70 nsew signal input
flabel metal3 s 0 39020 80 39100 0 FreeSans 320 0 0 0 FrameData[29]
port 71 nsew signal input
flabel metal3 s 0 25412 80 25492 0 FreeSans 320 0 0 0 FrameData[2]
port 72 nsew signal input
flabel metal3 s 0 39524 80 39604 0 FreeSans 320 0 0 0 FrameData[30]
port 73 nsew signal input
flabel metal3 s 0 40028 80 40108 0 FreeSans 320 0 0 0 FrameData[31]
port 74 nsew signal input
flabel metal3 s 0 25916 80 25996 0 FreeSans 320 0 0 0 FrameData[3]
port 75 nsew signal input
flabel metal3 s 0 26420 80 26500 0 FreeSans 320 0 0 0 FrameData[4]
port 76 nsew signal input
flabel metal3 s 0 26924 80 27004 0 FreeSans 320 0 0 0 FrameData[5]
port 77 nsew signal input
flabel metal3 s 0 27428 80 27508 0 FreeSans 320 0 0 0 FrameData[6]
port 78 nsew signal input
flabel metal3 s 0 27932 80 28012 0 FreeSans 320 0 0 0 FrameData[7]
port 79 nsew signal input
flabel metal3 s 0 28436 80 28516 0 FreeSans 320 0 0 0 FrameData[8]
port 80 nsew signal input
flabel metal3 s 0 28940 80 29020 0 FreeSans 320 0 0 0 FrameData[9]
port 81 nsew signal input
flabel metal3 s 21424 32300 21504 32380 0 FreeSans 320 0 0 0 FrameData_O[0]
port 82 nsew signal output
flabel metal3 s 21424 35660 21504 35740 0 FreeSans 320 0 0 0 FrameData_O[10]
port 83 nsew signal output
flabel metal3 s 21424 35996 21504 36076 0 FreeSans 320 0 0 0 FrameData_O[11]
port 84 nsew signal output
flabel metal3 s 21424 36332 21504 36412 0 FreeSans 320 0 0 0 FrameData_O[12]
port 85 nsew signal output
flabel metal3 s 21424 36668 21504 36748 0 FreeSans 320 0 0 0 FrameData_O[13]
port 86 nsew signal output
flabel metal3 s 21424 37004 21504 37084 0 FreeSans 320 0 0 0 FrameData_O[14]
port 87 nsew signal output
flabel metal3 s 21424 37340 21504 37420 0 FreeSans 320 0 0 0 FrameData_O[15]
port 88 nsew signal output
flabel metal3 s 21424 37676 21504 37756 0 FreeSans 320 0 0 0 FrameData_O[16]
port 89 nsew signal output
flabel metal3 s 21424 38012 21504 38092 0 FreeSans 320 0 0 0 FrameData_O[17]
port 90 nsew signal output
flabel metal3 s 21424 38348 21504 38428 0 FreeSans 320 0 0 0 FrameData_O[18]
port 91 nsew signal output
flabel metal3 s 21424 38684 21504 38764 0 FreeSans 320 0 0 0 FrameData_O[19]
port 92 nsew signal output
flabel metal3 s 21424 32636 21504 32716 0 FreeSans 320 0 0 0 FrameData_O[1]
port 93 nsew signal output
flabel metal3 s 21424 39020 21504 39100 0 FreeSans 320 0 0 0 FrameData_O[20]
port 94 nsew signal output
flabel metal3 s 21424 39356 21504 39436 0 FreeSans 320 0 0 0 FrameData_O[21]
port 95 nsew signal output
flabel metal3 s 21424 39692 21504 39772 0 FreeSans 320 0 0 0 FrameData_O[22]
port 96 nsew signal output
flabel metal3 s 21424 40028 21504 40108 0 FreeSans 320 0 0 0 FrameData_O[23]
port 97 nsew signal output
flabel metal3 s 21424 40364 21504 40444 0 FreeSans 320 0 0 0 FrameData_O[24]
port 98 nsew signal output
flabel metal3 s 21424 40700 21504 40780 0 FreeSans 320 0 0 0 FrameData_O[25]
port 99 nsew signal output
flabel metal3 s 21424 41036 21504 41116 0 FreeSans 320 0 0 0 FrameData_O[26]
port 100 nsew signal output
flabel metal3 s 21424 41372 21504 41452 0 FreeSans 320 0 0 0 FrameData_O[27]
port 101 nsew signal output
flabel metal3 s 21424 41708 21504 41788 0 FreeSans 320 0 0 0 FrameData_O[28]
port 102 nsew signal output
flabel metal3 s 21424 42044 21504 42124 0 FreeSans 320 0 0 0 FrameData_O[29]
port 103 nsew signal output
flabel metal3 s 21424 32972 21504 33052 0 FreeSans 320 0 0 0 FrameData_O[2]
port 104 nsew signal output
flabel metal3 s 21424 42380 21504 42460 0 FreeSans 320 0 0 0 FrameData_O[30]
port 105 nsew signal output
flabel metal3 s 21424 42716 21504 42796 0 FreeSans 320 0 0 0 FrameData_O[31]
port 106 nsew signal output
flabel metal3 s 21424 33308 21504 33388 0 FreeSans 320 0 0 0 FrameData_O[3]
port 107 nsew signal output
flabel metal3 s 21424 33644 21504 33724 0 FreeSans 320 0 0 0 FrameData_O[4]
port 108 nsew signal output
flabel metal3 s 21424 33980 21504 34060 0 FreeSans 320 0 0 0 FrameData_O[5]
port 109 nsew signal output
flabel metal3 s 21424 34316 21504 34396 0 FreeSans 320 0 0 0 FrameData_O[6]
port 110 nsew signal output
flabel metal3 s 21424 34652 21504 34732 0 FreeSans 320 0 0 0 FrameData_O[7]
port 111 nsew signal output
flabel metal3 s 21424 34988 21504 35068 0 FreeSans 320 0 0 0 FrameData_O[8]
port 112 nsew signal output
flabel metal3 s 21424 35324 21504 35404 0 FreeSans 320 0 0 0 FrameData_O[9]
port 113 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 FrameStrobe[0]
port 114 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 FrameStrobe[10]
port 115 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 FrameStrobe[11]
port 116 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 FrameStrobe[12]
port 117 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 FrameStrobe[13]
port 118 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 FrameStrobe[14]
port 119 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 FrameStrobe[15]
port 120 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 FrameStrobe[16]
port 121 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 FrameStrobe[17]
port 122 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 FrameStrobe[18]
port 123 nsew signal input
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 FrameStrobe[19]
port 124 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 FrameStrobe[1]
port 125 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 FrameStrobe[2]
port 126 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 FrameStrobe[3]
port 127 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 FrameStrobe[4]
port 128 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 FrameStrobe[5]
port 129 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 FrameStrobe[6]
port 130 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 FrameStrobe[7]
port 131 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 FrameStrobe[8]
port 132 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 FrameStrobe[9]
port 133 nsew signal input
flabel metal2 s 15800 42928 15880 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[0]
port 134 nsew signal output
flabel metal2 s 17720 42928 17800 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[10]
port 135 nsew signal output
flabel metal2 s 17912 42928 17992 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[11]
port 136 nsew signal output
flabel metal2 s 18104 42928 18184 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[12]
port 137 nsew signal output
flabel metal2 s 18296 42928 18376 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[13]
port 138 nsew signal output
flabel metal2 s 18488 42928 18568 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[14]
port 139 nsew signal output
flabel metal2 s 18680 42928 18760 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[15]
port 140 nsew signal output
flabel metal2 s 18872 42928 18952 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[16]
port 141 nsew signal output
flabel metal2 s 19064 42928 19144 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[17]
port 142 nsew signal output
flabel metal2 s 19256 42928 19336 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[18]
port 143 nsew signal output
flabel metal2 s 19448 42928 19528 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[19]
port 144 nsew signal output
flabel metal2 s 15992 42928 16072 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[1]
port 145 nsew signal output
flabel metal2 s 16184 42928 16264 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[2]
port 146 nsew signal output
flabel metal2 s 16376 42928 16456 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[3]
port 147 nsew signal output
flabel metal2 s 16568 42928 16648 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[4]
port 148 nsew signal output
flabel metal2 s 16760 42928 16840 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[5]
port 149 nsew signal output
flabel metal2 s 16952 42928 17032 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[6]
port 150 nsew signal output
flabel metal2 s 17144 42928 17224 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[7]
port 151 nsew signal output
flabel metal2 s 17336 42928 17416 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[8]
port 152 nsew signal output
flabel metal2 s 17528 42928 17608 43008 0 FreeSans 320 0 0 0 FrameStrobe_O[9]
port 153 nsew signal output
flabel metal2 s 1784 42928 1864 43008 0 FreeSans 320 0 0 0 N1BEG[0]
port 154 nsew signal output
flabel metal2 s 1976 42928 2056 43008 0 FreeSans 320 0 0 0 N1BEG[1]
port 155 nsew signal output
flabel metal2 s 2168 42928 2248 43008 0 FreeSans 320 0 0 0 N1BEG[2]
port 156 nsew signal output
flabel metal2 s 2360 42928 2440 43008 0 FreeSans 320 0 0 0 N1BEG[3]
port 157 nsew signal output
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 N1END[0]
port 158 nsew signal input
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 N1END[1]
port 159 nsew signal input
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 N1END[2]
port 160 nsew signal input
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 N1END[3]
port 161 nsew signal input
flabel metal2 s 2552 42928 2632 43008 0 FreeSans 320 0 0 0 N2BEG[0]
port 162 nsew signal output
flabel metal2 s 2744 42928 2824 43008 0 FreeSans 320 0 0 0 N2BEG[1]
port 163 nsew signal output
flabel metal2 s 2936 42928 3016 43008 0 FreeSans 320 0 0 0 N2BEG[2]
port 164 nsew signal output
flabel metal2 s 3128 42928 3208 43008 0 FreeSans 320 0 0 0 N2BEG[3]
port 165 nsew signal output
flabel metal2 s 3320 42928 3400 43008 0 FreeSans 320 0 0 0 N2BEG[4]
port 166 nsew signal output
flabel metal2 s 3512 42928 3592 43008 0 FreeSans 320 0 0 0 N2BEG[5]
port 167 nsew signal output
flabel metal2 s 3704 42928 3784 43008 0 FreeSans 320 0 0 0 N2BEG[6]
port 168 nsew signal output
flabel metal2 s 3896 42928 3976 43008 0 FreeSans 320 0 0 0 N2BEG[7]
port 169 nsew signal output
flabel metal2 s 4088 42928 4168 43008 0 FreeSans 320 0 0 0 N2BEGb[0]
port 170 nsew signal output
flabel metal2 s 4280 42928 4360 43008 0 FreeSans 320 0 0 0 N2BEGb[1]
port 171 nsew signal output
flabel metal2 s 4472 42928 4552 43008 0 FreeSans 320 0 0 0 N2BEGb[2]
port 172 nsew signal output
flabel metal2 s 4664 42928 4744 43008 0 FreeSans 320 0 0 0 N2BEGb[3]
port 173 nsew signal output
flabel metal2 s 4856 42928 4936 43008 0 FreeSans 320 0 0 0 N2BEGb[4]
port 174 nsew signal output
flabel metal2 s 5048 42928 5128 43008 0 FreeSans 320 0 0 0 N2BEGb[5]
port 175 nsew signal output
flabel metal2 s 5240 42928 5320 43008 0 FreeSans 320 0 0 0 N2BEGb[6]
port 176 nsew signal output
flabel metal2 s 5432 42928 5512 43008 0 FreeSans 320 0 0 0 N2BEGb[7]
port 177 nsew signal output
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 N2END[0]
port 178 nsew signal input
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 N2END[1]
port 179 nsew signal input
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 N2END[2]
port 180 nsew signal input
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 N2END[3]
port 181 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 N2END[4]
port 182 nsew signal input
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 N2END[5]
port 183 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 N2END[6]
port 184 nsew signal input
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 N2END[7]
port 185 nsew signal input
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 N2MID[0]
port 186 nsew signal input
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 N2MID[1]
port 187 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 N2MID[2]
port 188 nsew signal input
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 N2MID[3]
port 189 nsew signal input
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 N2MID[4]
port 190 nsew signal input
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 N2MID[5]
port 191 nsew signal input
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 N2MID[6]
port 192 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 N2MID[7]
port 193 nsew signal input
flabel metal2 s 5624 42928 5704 43008 0 FreeSans 320 0 0 0 N4BEG[0]
port 194 nsew signal output
flabel metal2 s 7544 42928 7624 43008 0 FreeSans 320 0 0 0 N4BEG[10]
port 195 nsew signal output
flabel metal2 s 7736 42928 7816 43008 0 FreeSans 320 0 0 0 N4BEG[11]
port 196 nsew signal output
flabel metal2 s 7928 42928 8008 43008 0 FreeSans 320 0 0 0 N4BEG[12]
port 197 nsew signal output
flabel metal2 s 8120 42928 8200 43008 0 FreeSans 320 0 0 0 N4BEG[13]
port 198 nsew signal output
flabel metal2 s 8312 42928 8392 43008 0 FreeSans 320 0 0 0 N4BEG[14]
port 199 nsew signal output
flabel metal2 s 8504 42928 8584 43008 0 FreeSans 320 0 0 0 N4BEG[15]
port 200 nsew signal output
flabel metal2 s 5816 42928 5896 43008 0 FreeSans 320 0 0 0 N4BEG[1]
port 201 nsew signal output
flabel metal2 s 6008 42928 6088 43008 0 FreeSans 320 0 0 0 N4BEG[2]
port 202 nsew signal output
flabel metal2 s 6200 42928 6280 43008 0 FreeSans 320 0 0 0 N4BEG[3]
port 203 nsew signal output
flabel metal2 s 6392 42928 6472 43008 0 FreeSans 320 0 0 0 N4BEG[4]
port 204 nsew signal output
flabel metal2 s 6584 42928 6664 43008 0 FreeSans 320 0 0 0 N4BEG[5]
port 205 nsew signal output
flabel metal2 s 6776 42928 6856 43008 0 FreeSans 320 0 0 0 N4BEG[6]
port 206 nsew signal output
flabel metal2 s 6968 42928 7048 43008 0 FreeSans 320 0 0 0 N4BEG[7]
port 207 nsew signal output
flabel metal2 s 7160 42928 7240 43008 0 FreeSans 320 0 0 0 N4BEG[8]
port 208 nsew signal output
flabel metal2 s 7352 42928 7432 43008 0 FreeSans 320 0 0 0 N4BEG[9]
port 209 nsew signal output
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 N4END[0]
port 210 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 N4END[10]
port 211 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 N4END[11]
port 212 nsew signal input
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 N4END[12]
port 213 nsew signal input
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 N4END[13]
port 214 nsew signal input
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 N4END[14]
port 215 nsew signal input
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 N4END[15]
port 216 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 N4END[1]
port 217 nsew signal input
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 N4END[2]
port 218 nsew signal input
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 N4END[3]
port 219 nsew signal input
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 N4END[4]
port 220 nsew signal input
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 N4END[5]
port 221 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 N4END[6]
port 222 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 N4END[7]
port 223 nsew signal input
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 N4END[8]
port 224 nsew signal input
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 N4END[9]
port 225 nsew signal input
flabel metal3 s 0 23900 80 23980 0 FreeSans 320 0 0 0 RST_N_TT_PROJECT
port 226 nsew signal output
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 S1BEG[0]
port 227 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 S1BEG[1]
port 228 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 S1BEG[2]
port 229 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 S1BEG[3]
port 230 nsew signal output
flabel metal2 s 8696 42928 8776 43008 0 FreeSans 320 0 0 0 S1END[0]
port 231 nsew signal input
flabel metal2 s 8888 42928 8968 43008 0 FreeSans 320 0 0 0 S1END[1]
port 232 nsew signal input
flabel metal2 s 9080 42928 9160 43008 0 FreeSans 320 0 0 0 S1END[2]
port 233 nsew signal input
flabel metal2 s 9272 42928 9352 43008 0 FreeSans 320 0 0 0 S1END[3]
port 234 nsew signal input
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 S2BEG[0]
port 235 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 S2BEG[1]
port 236 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 S2BEG[2]
port 237 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 S2BEG[3]
port 238 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 S2BEG[4]
port 239 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 S2BEG[5]
port 240 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 S2BEG[6]
port 241 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 S2BEG[7]
port 242 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 S2BEGb[0]
port 243 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 S2BEGb[1]
port 244 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 S2BEGb[2]
port 245 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 S2BEGb[3]
port 246 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 S2BEGb[4]
port 247 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 S2BEGb[5]
port 248 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 S2BEGb[6]
port 249 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 S2BEGb[7]
port 250 nsew signal output
flabel metal2 s 11000 42928 11080 43008 0 FreeSans 320 0 0 0 S2END[0]
port 251 nsew signal input
flabel metal2 s 11192 42928 11272 43008 0 FreeSans 320 0 0 0 S2END[1]
port 252 nsew signal input
flabel metal2 s 11384 42928 11464 43008 0 FreeSans 320 0 0 0 S2END[2]
port 253 nsew signal input
flabel metal2 s 11576 42928 11656 43008 0 FreeSans 320 0 0 0 S2END[3]
port 254 nsew signal input
flabel metal2 s 11768 42928 11848 43008 0 FreeSans 320 0 0 0 S2END[4]
port 255 nsew signal input
flabel metal2 s 11960 42928 12040 43008 0 FreeSans 320 0 0 0 S2END[5]
port 256 nsew signal input
flabel metal2 s 12152 42928 12232 43008 0 FreeSans 320 0 0 0 S2END[6]
port 257 nsew signal input
flabel metal2 s 12344 42928 12424 43008 0 FreeSans 320 0 0 0 S2END[7]
port 258 nsew signal input
flabel metal2 s 9464 42928 9544 43008 0 FreeSans 320 0 0 0 S2MID[0]
port 259 nsew signal input
flabel metal2 s 9656 42928 9736 43008 0 FreeSans 320 0 0 0 S2MID[1]
port 260 nsew signal input
flabel metal2 s 9848 42928 9928 43008 0 FreeSans 320 0 0 0 S2MID[2]
port 261 nsew signal input
flabel metal2 s 10040 42928 10120 43008 0 FreeSans 320 0 0 0 S2MID[3]
port 262 nsew signal input
flabel metal2 s 10232 42928 10312 43008 0 FreeSans 320 0 0 0 S2MID[4]
port 263 nsew signal input
flabel metal2 s 10424 42928 10504 43008 0 FreeSans 320 0 0 0 S2MID[5]
port 264 nsew signal input
flabel metal2 s 10616 42928 10696 43008 0 FreeSans 320 0 0 0 S2MID[6]
port 265 nsew signal input
flabel metal2 s 10808 42928 10888 43008 0 FreeSans 320 0 0 0 S2MID[7]
port 266 nsew signal input
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 S4BEG[0]
port 267 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 S4BEG[10]
port 268 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 S4BEG[11]
port 269 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 S4BEG[12]
port 270 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 S4BEG[13]
port 271 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 S4BEG[14]
port 272 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 S4BEG[15]
port 273 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 S4BEG[1]
port 274 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 S4BEG[2]
port 275 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 S4BEG[3]
port 276 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 S4BEG[4]
port 277 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 S4BEG[5]
port 278 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 S4BEG[6]
port 279 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 S4BEG[7]
port 280 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 S4BEG[8]
port 281 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 S4BEG[9]
port 282 nsew signal output
flabel metal2 s 12536 42928 12616 43008 0 FreeSans 320 0 0 0 S4END[0]
port 283 nsew signal input
flabel metal2 s 14456 42928 14536 43008 0 FreeSans 320 0 0 0 S4END[10]
port 284 nsew signal input
flabel metal2 s 14648 42928 14728 43008 0 FreeSans 320 0 0 0 S4END[11]
port 285 nsew signal input
flabel metal2 s 14840 42928 14920 43008 0 FreeSans 320 0 0 0 S4END[12]
port 286 nsew signal input
flabel metal2 s 15032 42928 15112 43008 0 FreeSans 320 0 0 0 S4END[13]
port 287 nsew signal input
flabel metal2 s 15224 42928 15304 43008 0 FreeSans 320 0 0 0 S4END[14]
port 288 nsew signal input
flabel metal2 s 15416 42928 15496 43008 0 FreeSans 320 0 0 0 S4END[15]
port 289 nsew signal input
flabel metal2 s 12728 42928 12808 43008 0 FreeSans 320 0 0 0 S4END[1]
port 290 nsew signal input
flabel metal2 s 12920 42928 13000 43008 0 FreeSans 320 0 0 0 S4END[2]
port 291 nsew signal input
flabel metal2 s 13112 42928 13192 43008 0 FreeSans 320 0 0 0 S4END[3]
port 292 nsew signal input
flabel metal2 s 13304 42928 13384 43008 0 FreeSans 320 0 0 0 S4END[4]
port 293 nsew signal input
flabel metal2 s 13496 42928 13576 43008 0 FreeSans 320 0 0 0 S4END[5]
port 294 nsew signal input
flabel metal2 s 13688 42928 13768 43008 0 FreeSans 320 0 0 0 S4END[6]
port 295 nsew signal input
flabel metal2 s 13880 42928 13960 43008 0 FreeSans 320 0 0 0 S4END[7]
port 296 nsew signal input
flabel metal2 s 14072 42928 14152 43008 0 FreeSans 320 0 0 0 S4END[8]
port 297 nsew signal input
flabel metal2 s 14264 42928 14344 43008 0 FreeSans 320 0 0 0 S4END[9]
port 298 nsew signal input
flabel metal3 s 0 18860 80 18940 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT0
port 299 nsew signal output
flabel metal3 s 0 19364 80 19444 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT1
port 300 nsew signal output
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT2
port 301 nsew signal output
flabel metal3 s 0 20372 80 20452 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT3
port 302 nsew signal output
flabel metal3 s 0 20876 80 20956 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT4
port 303 nsew signal output
flabel metal3 s 0 21380 80 21460 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT5
port 304 nsew signal output
flabel metal3 s 0 21884 80 21964 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT6
port 305 nsew signal output
flabel metal3 s 0 22388 80 22468 0 FreeSans 320 0 0 0 UIO_IN_TT_PROJECT7
port 306 nsew signal output
flabel metal3 s 0 10796 80 10876 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT0
port 307 nsew signal input
flabel metal3 s 0 11300 80 11380 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT1
port 308 nsew signal input
flabel metal3 s 0 11804 80 11884 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT2
port 309 nsew signal input
flabel metal3 s 0 12308 80 12388 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT3
port 310 nsew signal input
flabel metal3 s 0 12812 80 12892 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT4
port 311 nsew signal input
flabel metal3 s 0 13316 80 13396 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT5
port 312 nsew signal input
flabel metal3 s 0 13820 80 13900 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT6
port 313 nsew signal input
flabel metal3 s 0 14324 80 14404 0 FreeSans 320 0 0 0 UIO_OE_TT_PROJECT7
port 314 nsew signal input
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT0
port 315 nsew signal input
flabel metal3 s 0 7268 80 7348 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT1
port 316 nsew signal input
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT2
port 317 nsew signal input
flabel metal3 s 0 8276 80 8356 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT3
port 318 nsew signal input
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT4
port 319 nsew signal input
flabel metal3 s 0 9284 80 9364 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT5
port 320 nsew signal input
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT6
port 321 nsew signal input
flabel metal3 s 0 10292 80 10372 0 FreeSans 320 0 0 0 UIO_OUT_TT_PROJECT7
port 322 nsew signal input
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT0
port 323 nsew signal output
flabel metal3 s 0 15332 80 15412 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT1
port 324 nsew signal output
flabel metal3 s 0 15836 80 15916 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT2
port 325 nsew signal output
flabel metal3 s 0 16340 80 16420 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT3
port 326 nsew signal output
flabel metal3 s 0 16844 80 16924 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT4
port 327 nsew signal output
flabel metal3 s 0 17348 80 17428 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT5
port 328 nsew signal output
flabel metal3 s 0 17852 80 17932 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT6
port 329 nsew signal output
flabel metal3 s 0 18356 80 18436 0 FreeSans 320 0 0 0 UI_IN_TT_PROJECT7
port 330 nsew signal output
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT0
port 331 nsew signal input
flabel metal3 s 0 3236 80 3316 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT1
port 332 nsew signal input
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT2
port 333 nsew signal input
flabel metal3 s 0 4244 80 4324 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT3
port 334 nsew signal input
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT4
port 335 nsew signal input
flabel metal3 s 0 5252 80 5332 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT5
port 336 nsew signal input
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT6
port 337 nsew signal input
flabel metal3 s 0 6260 80 6340 0 FreeSans 320 0 0 0 UO_OUT_TT_PROJECT7
port 338 nsew signal input
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 UserCLK
port 339 nsew signal input
flabel metal2 s 15608 42928 15688 43008 0 FreeSans 320 0 0 0 UserCLKo
port 340 nsew signal output
flabel metal6 s 4892 0 5332 43008 0 FreeSans 2624 90 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 4892 42680 5332 43008 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 0 20452 43008 0 FreeSans 2624 90 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 20012 42680 20452 43008 0 FreeSans 2624 0 0 0 VGND
port 341 nsew ground bidirectional
flabel metal6 s 3652 0 4092 43008 0 FreeSans 2624 90 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 3652 42680 4092 43008 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 0 19212 43008 0 FreeSans 2624 90 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal6 s 18772 42680 19212 43008 0 FreeSans 2624 0 0 0 VPWR
port 342 nsew power bidirectional
flabel metal3 s 21424 44 21504 124 0 FreeSans 320 0 0 0 W1END[0]
port 343 nsew signal input
flabel metal3 s 21424 380 21504 460 0 FreeSans 320 0 0 0 W1END[1]
port 344 nsew signal input
flabel metal3 s 21424 716 21504 796 0 FreeSans 320 0 0 0 W1END[2]
port 345 nsew signal input
flabel metal3 s 21424 1052 21504 1132 0 FreeSans 320 0 0 0 W1END[3]
port 346 nsew signal input
flabel metal3 s 21424 4076 21504 4156 0 FreeSans 320 0 0 0 W2END[0]
port 347 nsew signal input
flabel metal3 s 21424 4412 21504 4492 0 FreeSans 320 0 0 0 W2END[1]
port 348 nsew signal input
flabel metal3 s 21424 4748 21504 4828 0 FreeSans 320 0 0 0 W2END[2]
port 349 nsew signal input
flabel metal3 s 21424 5084 21504 5164 0 FreeSans 320 0 0 0 W2END[3]
port 350 nsew signal input
flabel metal3 s 21424 5420 21504 5500 0 FreeSans 320 0 0 0 W2END[4]
port 351 nsew signal input
flabel metal3 s 21424 5756 21504 5836 0 FreeSans 320 0 0 0 W2END[5]
port 352 nsew signal input
flabel metal3 s 21424 6092 21504 6172 0 FreeSans 320 0 0 0 W2END[6]
port 353 nsew signal input
flabel metal3 s 21424 6428 21504 6508 0 FreeSans 320 0 0 0 W2END[7]
port 354 nsew signal input
flabel metal3 s 21424 1388 21504 1468 0 FreeSans 320 0 0 0 W2MID[0]
port 355 nsew signal input
flabel metal3 s 21424 1724 21504 1804 0 FreeSans 320 0 0 0 W2MID[1]
port 356 nsew signal input
flabel metal3 s 21424 2060 21504 2140 0 FreeSans 320 0 0 0 W2MID[2]
port 357 nsew signal input
flabel metal3 s 21424 2396 21504 2476 0 FreeSans 320 0 0 0 W2MID[3]
port 358 nsew signal input
flabel metal3 s 21424 2732 21504 2812 0 FreeSans 320 0 0 0 W2MID[4]
port 359 nsew signal input
flabel metal3 s 21424 3068 21504 3148 0 FreeSans 320 0 0 0 W2MID[5]
port 360 nsew signal input
flabel metal3 s 21424 3404 21504 3484 0 FreeSans 320 0 0 0 W2MID[6]
port 361 nsew signal input
flabel metal3 s 21424 3740 21504 3820 0 FreeSans 320 0 0 0 W2MID[7]
port 362 nsew signal input
flabel metal3 s 21424 12140 21504 12220 0 FreeSans 320 0 0 0 W6END[0]
port 363 nsew signal input
flabel metal3 s 21424 15500 21504 15580 0 FreeSans 320 0 0 0 W6END[10]
port 364 nsew signal input
flabel metal3 s 21424 15836 21504 15916 0 FreeSans 320 0 0 0 W6END[11]
port 365 nsew signal input
flabel metal3 s 21424 12476 21504 12556 0 FreeSans 320 0 0 0 W6END[1]
port 366 nsew signal input
flabel metal3 s 21424 12812 21504 12892 0 FreeSans 320 0 0 0 W6END[2]
port 367 nsew signal input
flabel metal3 s 21424 13148 21504 13228 0 FreeSans 320 0 0 0 W6END[3]
port 368 nsew signal input
flabel metal3 s 21424 13484 21504 13564 0 FreeSans 320 0 0 0 W6END[4]
port 369 nsew signal input
flabel metal3 s 21424 13820 21504 13900 0 FreeSans 320 0 0 0 W6END[5]
port 370 nsew signal input
flabel metal3 s 21424 14156 21504 14236 0 FreeSans 320 0 0 0 W6END[6]
port 371 nsew signal input
flabel metal3 s 21424 14492 21504 14572 0 FreeSans 320 0 0 0 W6END[7]
port 372 nsew signal input
flabel metal3 s 21424 14828 21504 14908 0 FreeSans 320 0 0 0 W6END[8]
port 373 nsew signal input
flabel metal3 s 21424 15164 21504 15244 0 FreeSans 320 0 0 0 W6END[9]
port 374 nsew signal input
flabel metal3 s 21424 6764 21504 6844 0 FreeSans 320 0 0 0 WW4END[0]
port 375 nsew signal input
flabel metal3 s 21424 10124 21504 10204 0 FreeSans 320 0 0 0 WW4END[10]
port 376 nsew signal input
flabel metal3 s 21424 10460 21504 10540 0 FreeSans 320 0 0 0 WW4END[11]
port 377 nsew signal input
flabel metal3 s 21424 10796 21504 10876 0 FreeSans 320 0 0 0 WW4END[12]
port 378 nsew signal input
flabel metal3 s 21424 11132 21504 11212 0 FreeSans 320 0 0 0 WW4END[13]
port 379 nsew signal input
flabel metal3 s 21424 11468 21504 11548 0 FreeSans 320 0 0 0 WW4END[14]
port 380 nsew signal input
flabel metal3 s 21424 11804 21504 11884 0 FreeSans 320 0 0 0 WW4END[15]
port 381 nsew signal input
flabel metal3 s 21424 7100 21504 7180 0 FreeSans 320 0 0 0 WW4END[1]
port 382 nsew signal input
flabel metal3 s 21424 7436 21504 7516 0 FreeSans 320 0 0 0 WW4END[2]
port 383 nsew signal input
flabel metal3 s 21424 7772 21504 7852 0 FreeSans 320 0 0 0 WW4END[3]
port 384 nsew signal input
flabel metal3 s 21424 8108 21504 8188 0 FreeSans 320 0 0 0 WW4END[4]
port 385 nsew signal input
flabel metal3 s 21424 8444 21504 8524 0 FreeSans 320 0 0 0 WW4END[5]
port 386 nsew signal input
flabel metal3 s 21424 8780 21504 8860 0 FreeSans 320 0 0 0 WW4END[6]
port 387 nsew signal input
flabel metal3 s 21424 9116 21504 9196 0 FreeSans 320 0 0 0 WW4END[7]
port 388 nsew signal input
flabel metal3 s 21424 9452 21504 9532 0 FreeSans 320 0 0 0 WW4END[8]
port 389 nsew signal input
flabel metal3 s 21424 9788 21504 9868 0 FreeSans 320 0 0 0 WW4END[9]
port 390 nsew signal input
rlabel metal1 10802 41580 10802 41580 0 VGND
rlabel metal1 10752 40824 10752 40824 0 VPWR
rlabel metal2 4224 24654 4224 24654 0 CLK_TT_PROJECT
rlabel metal3 21138 16212 21138 16212 0 E1BEG[0]
rlabel metal2 19488 17052 19488 17052 0 E1BEG[1]
rlabel metal2 18336 15834 18336 15834 0 E1BEG[2]
rlabel metal2 20256 12390 20256 12390 0 E1BEG[3]
rlabel metal2 20016 11928 20016 11928 0 E2BEG[0]
rlabel metal3 19632 31164 19632 31164 0 E2BEG[1]
rlabel metal2 19968 31668 19968 31668 0 E2BEG[2]
rlabel metal3 21138 18564 21138 18564 0 E2BEG[3]
rlabel metal3 21186 18900 21186 18900 0 E2BEG[4]
rlabel metal3 20736 29148 20736 29148 0 E2BEG[5]
rlabel metal2 18720 31710 18720 31710 0 E2BEG[6]
rlabel metal2 20256 14154 20256 14154 0 E2BEG[7]
rlabel metal2 17664 12306 17664 12306 0 E2BEGb[0]
rlabel metal2 19968 35112 19968 35112 0 E2BEGb[1]
rlabel metal4 19968 19446 19968 19446 0 E2BEGb[2]
rlabel metal3 20832 4830 20832 4830 0 E2BEGb[3]
rlabel metal2 18288 13020 18288 13020 0 E2BEGb[4]
rlabel metal3 21378 21924 21378 21924 0 E2BEGb[5]
rlabel metal3 19632 31080 19632 31080 0 E2BEGb[6]
rlabel metal3 20994 22596 20994 22596 0 E2BEGb[7]
rlabel metal2 17664 27888 17664 27888 0 E6BEG[0]
rlabel metal3 20802 31668 20802 31668 0 E6BEG[10]
rlabel metal2 19872 32802 19872 32802 0 E6BEG[11]
rlabel metal2 14016 23982 14016 23982 0 E6BEG[1]
rlabel metal3 17136 30156 17136 30156 0 E6BEG[2]
rlabel metal3 17472 29274 17472 29274 0 E6BEG[3]
rlabel metal2 20064 30030 20064 30030 0 E6BEG[4]
rlabel metal3 20802 29988 20802 29988 0 E6BEG[5]
rlabel metal3 21234 30324 21234 30324 0 E6BEG[6]
rlabel metal2 19776 30996 19776 30996 0 E6BEG[7]
rlabel metal3 20544 31038 20544 31038 0 E6BEG[8]
rlabel metal3 21090 31332 21090 31332 0 E6BEG[9]
rlabel metal3 19680 23226 19680 23226 0 EE4BEG[0]
rlabel metal3 21186 26292 21186 26292 0 EE4BEG[10]
rlabel metal2 20064 27006 20064 27006 0 EE4BEG[11]
rlabel metal2 19584 27552 19584 27552 0 EE4BEG[12]
rlabel metal3 20064 28980 20064 28980 0 EE4BEG[13]
rlabel metal2 19728 29652 19728 29652 0 EE4BEG[14]
rlabel metal2 19680 28476 19680 28476 0 EE4BEG[15]
rlabel metal3 19920 29820 19920 29820 0 EE4BEG[1]
rlabel metal4 19872 24192 19872 24192 0 EE4BEG[2]
rlabel metal2 19584 24612 19584 24612 0 EE4BEG[3]
rlabel metal2 19968 24696 19968 24696 0 EE4BEG[4]
rlabel metal2 20064 25578 20064 25578 0 EE4BEG[5]
rlabel metal2 19968 26712 19968 26712 0 EE4BEG[6]
rlabel metal2 15312 21000 15312 21000 0 EE4BEG[7]
rlabel metal3 19584 26586 19584 26586 0 EE4BEG[8]
rlabel metal2 21216 33096 21216 33096 0 EE4BEG[9]
rlabel metal3 942 22932 942 22932 0 ENA_TT_PROJECT
rlabel metal5 2304 36624 2304 36624 0 FrameData[0]
rlabel metal2 1536 34482 1536 34482 0 FrameData[10]
rlabel metal2 1392 30660 1392 30660 0 FrameData[11]
rlabel metal2 11424 2016 11424 2016 0 FrameData[12]
rlabel metal3 19536 38976 19536 38976 0 FrameData[13]
rlabel metal2 1536 18984 1536 18984 0 FrameData[14]
rlabel metal2 1632 31332 1632 31332 0 FrameData[15]
rlabel via2 78 32508 78 32508 0 FrameData[16]
rlabel via2 78 33012 78 33012 0 FrameData[17]
rlabel metal2 1920 33642 1920 33642 0 FrameData[18]
rlabel metal2 1440 9702 1440 9702 0 FrameData[19]
rlabel metal3 15888 12516 15888 12516 0 FrameData[1]
rlabel metal3 14304 12096 14304 12096 0 FrameData[20]
rlabel metal3 750 35028 750 35028 0 FrameData[21]
rlabel metal2 1536 19908 1536 19908 0 FrameData[22]
rlabel metal3 654 36036 654 36036 0 FrameData[23]
rlabel metal2 1296 12516 1296 12516 0 FrameData[24]
rlabel metal2 14304 12264 14304 12264 0 FrameData[25]
rlabel metal2 17952 16842 17952 16842 0 FrameData[26]
rlabel metal2 11520 378 11520 378 0 FrameData[27]
rlabel metal2 13632 2016 13632 2016 0 FrameData[28]
rlabel metal2 1392 37380 1392 37380 0 FrameData[29]
rlabel metal2 1296 29148 1296 29148 0 FrameData[2]
rlabel metal2 2208 7896 2208 7896 0 FrameData[30]
rlabel metal2 12384 36036 12384 36036 0 FrameData[31]
rlabel metal2 17088 12936 17088 12936 0 FrameData[3]
rlabel metal2 1872 18648 1872 18648 0 FrameData[4]
rlabel metal4 2400 13272 2400 13272 0 FrameData[5]
rlabel metal2 1248 32214 1248 32214 0 FrameData[6]
rlabel metal4 2496 13398 2496 13398 0 FrameData[7]
rlabel metal5 2112 9744 2112 9744 0 FrameData[8]
rlabel metal2 2160 2352 2160 2352 0 FrameData[9]
rlabel metal2 19776 32550 19776 32550 0 FrameData_O[0]
rlabel metal3 21186 35700 21186 35700 0 FrameData_O[10]
rlabel metal3 20802 36036 20802 36036 0 FrameData_O[11]
rlabel metal3 19410 36372 19410 36372 0 FrameData_O[12]
rlabel metal3 19872 36750 19872 36750 0 FrameData_O[13]
rlabel metal3 21042 37044 21042 37044 0 FrameData_O[14]
rlabel metal3 20898 37380 20898 37380 0 FrameData_O[15]
rlabel metal3 20802 37716 20802 37716 0 FrameData_O[16]
rlabel metal3 14016 23940 14016 23940 0 FrameData_O[17]
rlabel metal3 14976 35448 14976 35448 0 FrameData_O[18]
rlabel metal4 12528 33348 12528 33348 0 FrameData_O[19]
rlabel metal3 21330 32676 21330 32676 0 FrameData_O[1]
rlabel metal5 15456 34020 15456 34020 0 FrameData_O[20]
rlabel metal2 16224 38094 16224 38094 0 FrameData_O[21]
rlabel metal2 18144 39648 18144 39648 0 FrameData_O[22]
rlabel metal2 13536 39900 13536 39900 0 FrameData_O[23]
rlabel metal3 15744 35574 15744 35574 0 FrameData_O[24]
rlabel metal3 14640 30828 14640 30828 0 FrameData_O[25]
rlabel metal4 12480 39480 12480 39480 0 FrameData_O[26]
rlabel metal2 21264 29400 21264 29400 0 FrameData_O[27]
rlabel metal4 16416 42000 16416 42000 0 FrameData_O[28]
rlabel metal4 17280 26040 17280 26040 0 FrameData_O[29]
rlabel metal3 20994 33012 20994 33012 0 FrameData_O[2]
rlabel metal2 7440 37968 7440 37968 0 FrameData_O[30]
rlabel metal2 13152 27552 13152 27552 0 FrameData_O[31]
rlabel metal3 21042 33348 21042 33348 0 FrameData_O[3]
rlabel metal3 21090 33684 21090 33684 0 FrameData_O[4]
rlabel metal3 21138 34020 21138 34020 0 FrameData_O[5]
rlabel metal3 20994 34356 20994 34356 0 FrameData_O[6]
rlabel metal3 20802 34692 20802 34692 0 FrameData_O[7]
rlabel metal3 20802 35028 20802 35028 0 FrameData_O[8]
rlabel metal4 17664 35910 17664 35910 0 FrameData_O[9]
rlabel metal2 2496 8694 2496 8694 0 FrameStrobe[0]
rlabel metal2 17760 492 17760 492 0 FrameStrobe[10]
rlabel metal2 17952 660 17952 660 0 FrameStrobe[11]
rlabel via2 18144 72 18144 72 0 FrameStrobe[12]
rlabel metal2 18336 366 18336 366 0 FrameStrobe[13]
rlabel metal2 18528 660 18528 660 0 FrameStrobe[14]
rlabel metal2 18720 660 18720 660 0 FrameStrobe[15]
rlabel metal2 18912 240 18912 240 0 FrameStrobe[16]
rlabel metal2 19104 492 19104 492 0 FrameStrobe[17]
rlabel metal2 19296 324 19296 324 0 FrameStrobe[18]
rlabel metal2 19488 408 19488 408 0 FrameStrobe[19]
rlabel metal2 16032 198 16032 198 0 FrameStrobe[1]
rlabel metal2 13056 18732 13056 18732 0 FrameStrobe[2]
rlabel metal2 19296 1260 19296 1260 0 FrameStrobe[3]
rlabel metal3 16512 10584 16512 10584 0 FrameStrobe[4]
rlabel metal2 14304 14406 14304 14406 0 FrameStrobe[5]
rlabel metal2 16992 660 16992 660 0 FrameStrobe[6]
rlabel metal2 14400 630 14400 630 0 FrameStrobe[7]
rlabel metal3 1872 35952 1872 35952 0 FrameStrobe[8]
rlabel metal2 17568 240 17568 240 0 FrameStrobe[9]
rlabel metal2 19488 39942 19488 39942 0 FrameStrobe_O[0]
rlabel metal3 18624 41412 18624 41412 0 FrameStrobe_O[10]
rlabel metal2 19872 41454 19872 41454 0 FrameStrobe_O[11]
rlabel metal2 18144 42768 18144 42768 0 FrameStrobe_O[12]
rlabel metal2 18336 42138 18336 42138 0 FrameStrobe_O[13]
rlabel metal2 18528 42600 18528 42600 0 FrameStrobe_O[14]
rlabel metal3 14688 36750 14688 36750 0 FrameStrobe_O[15]
rlabel metal2 18912 42810 18912 42810 0 FrameStrobe_O[16]
rlabel metal2 13008 30072 13008 30072 0 FrameStrobe_O[17]
rlabel via2 19296 42936 19296 42936 0 FrameStrobe_O[18]
rlabel metal3 14736 25536 14736 25536 0 FrameStrobe_O[19]
rlabel metal2 19776 40866 19776 40866 0 FrameStrobe_O[1]
rlabel metal2 19824 39060 19824 39060 0 FrameStrobe_O[2]
rlabel metal2 19872 40572 19872 40572 0 FrameStrobe_O[3]
rlabel metal3 17568 40656 17568 40656 0 FrameStrobe_O[4]
rlabel metal2 16800 41760 16800 41760 0 FrameStrobe_O[5]
rlabel metal3 18624 35028 18624 35028 0 FrameStrobe_O[6]
rlabel metal2 17184 42222 17184 42222 0 FrameStrobe_O[7]
rlabel metal3 2112 35700 2112 35700 0 FrameStrobe_O[8]
rlabel metal4 1440 40236 1440 40236 0 FrameStrobe_O[9]
rlabel metal2 6096 23772 6096 23772 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 7680 23863 7680 23863 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 12288 35700 12288 35700 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit10.Q
rlabel metal3 3456 37632 3456 37632 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 5568 2013 5568 2013 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit12.Q
rlabel metal4 2112 6720 2112 6720 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 15840 840 15840 840 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 2016 1554 2016 1554 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit15.Q
rlabel metal3 3936 23100 3936 23100 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit16.Q
rlabel via1 5712 23095 5712 23095 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 6816 38430 6816 38430 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 5280 38301 5280 38301 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit19.Q
rlabel metal3 5952 35154 5952 35154 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 4896 39774 4896 39774 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 6432 40401 6432 40401 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit21.Q
rlabel metal3 4080 20076 4080 20076 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 6720 19985 6720 19985 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 6672 16212 6672 16212 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit24.Q
rlabel metal2 6048 15372 6048 15372 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 1440 34230 1440 34230 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 1981 33019 1981 33019 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit27.Q
rlabel metal3 1680 26208 1680 26208 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 1248 26922 1248 26922 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 7200 34650 7200 34650 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 1920 5880 1920 5880 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 1925 6514 1925 6514 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 4512 35784 4512 35784 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 12288 39648 12288 39648 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 1872 27468 1872 27468 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit6.Q
rlabel metal3 3408 29400 3408 29400 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit7.Q
rlabel metal3 3600 29820 3600 29820 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 5376 28263 5376 28263 0 Inst_W_TT_IF_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 15552 5124 15552 5124 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit0.Q
rlabel metal3 15312 5880 15312 5880 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 7296 35952 7296 35952 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 8832 35828 8832 35828 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 3504 37128 3504 37128 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 4752 37380 4752 37380 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 1776 26124 1776 26124 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 3120 29484 3120 29484 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit15.Q
rlabel metal3 4992 21588 4992 21588 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 7680 21837 7680 21837 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit17.Q
rlabel metal3 6192 37632 6192 37632 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit18.Q
rlabel metal3 8688 37632 8688 37632 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 2880 24528 2880 24528 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 8592 38892 8592 38892 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 10176 39571 10176 39571 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 6720 27090 6720 27090 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 8256 27853 8256 27853 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 6384 24612 6384 24612 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit24.Q
rlabel metal2 7968 24861 7968 24861 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 7680 37254 7680 37254 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit26.Q
rlabel metal2 9216 36873 9216 36873 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 8688 39732 8688 39732 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 10272 40359 10272 40359 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 2112 24612 2112 24612 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 7104 27888 7104 27888 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit30.Q
rlabel via1 8688 27631 8688 27631 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 1728 4746 1728 4746 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 1152 5250 1152 5250 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 2304 5754 2304 5754 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 5760 2646 5760 2646 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 6816 21336 6816 21336 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 8304 22323 8304 22323 0 Inst_W_TT_IF_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 17184 8022 17184 8022 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit0.Q
rlabel metal3 19200 13188 19200 13188 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit1.Q
rlabel metal3 11808 9660 11808 9660 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit10.Q
rlabel metal3 13152 7980 13152 7980 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 12288 8022 12288 8022 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit12.Q
rlabel metal3 12720 18732 12720 18732 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 14016 18270 14016 18270 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit14.Q
rlabel metal3 12192 17640 12192 17640 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit15.Q
rlabel metal3 18912 18732 18912 18732 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 19200 19194 19200 19194 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 20160 18312 20160 18312 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 19296 7560 19296 7560 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit19.Q
rlabel metal3 18624 12516 18624 12516 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 19152 5628 19152 5628 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit20.Q
rlabel metal3 19337 1932 19337 1932 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 16608 12936 16608 12936 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 16512 10458 16512 10458 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit23.Q
rlabel metal3 15264 11004 15264 11004 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit24.Q
rlabel metal2 19200 16296 19200 16296 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit25.Q
rlabel metal3 17856 14700 17856 14700 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 20147 17099 20147 17099 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 18240 38262 18240 38262 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit28.Q
rlabel metal2 19104 39774 19104 39774 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 18624 14784 18624 14784 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 17952 36918 17952 36918 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 16128 6951 16128 6951 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 15936 36654 15936 36654 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 17280 36204 17280 36204 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit5.Q
rlabel metal3 15888 37380 15888 37380 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 16800 3780 16800 3780 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 17376 2142 17376 2142 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit8.Q
rlabel metal3 17664 2436 17664 2436 0 Inst_W_TT_IF_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 9216 26166 9216 26166 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 10752 27129 10752 27129 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 16704 23520 16704 23520 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 15024 23268 15024 23268 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 18528 33523 18528 33523 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit12.Q
rlabel metal2 16992 33138 16992 33138 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit13.Q
rlabel via1 19056 35191 19056 35191 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit14.Q
rlabel metal3 17472 35238 17472 35238 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 14880 18942 14880 18942 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 13056 19782 13056 19782 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 9744 9492 9744 9492 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 12384 10311 12384 10311 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 14976 27885 14976 27885 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 9360 7812 9360 7812 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 15168 15582 15168 15582 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit21.Q
rlabel metal3 13680 15540 13680 15540 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit22.Q
rlabel metal3 12864 14532 12864 14532 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit23.Q
rlabel metal3 16368 17976 16368 17976 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit24.Q
rlabel metal3 16560 18564 16560 18564 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit25.Q
rlabel metal3 16320 18396 16320 18396 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 19200 3528 19200 3528 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 19632 1932 19632 1932 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 19392 2184 19392 2184 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 13440 27332 13440 27332 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 16512 9450 16512 9450 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 17232 8652 17232 8652 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit31.Q
rlabel metal3 19440 30828 19440 30828 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit4.Q
rlabel metal2 17664 31962 17664 31962 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 19104 33933 19104 33933 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 17568 33936 17568 33936 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 15360 22010 15360 22010 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 13776 21756 13776 21756 0 Inst_W_TT_IF_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 11136 22008 11136 22008 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 9360 21756 9360 21756 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit1.Q
rlabel via1 12048 24586 12048 24586 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 10464 25242 10464 25242 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 14112 30828 14112 30828 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 12672 31290 12672 31290 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 19440 26292 19440 26292 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 17472 26880 17472 26880 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit15.Q
rlabel via2 11520 20073 11520 20073 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit16.Q
rlabel metal3 9792 20076 9792 20076 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 14304 24861 14304 24861 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 12768 24318 12768 24318 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 10848 24073 10848 24073 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit2.Q
rlabel metal3 19056 27720 19056 27720 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 17280 28602 17280 28602 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 16800 28058 16800 28058 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 15216 28308 15216 28308 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 12768 22351 12768 22351 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 11232 22554 11232 22554 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 10080 27846 10080 27846 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 11616 27097 11616 27097 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit27.Q
rlabel metal3 10416 37716 10416 37716 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit28.Q
rlabel metal3 11808 36120 11808 36120 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 9312 24444 9312 24444 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 12048 36708 12048 36708 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 13824 36372 13824 36372 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 14400 25991 14400 25991 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 12864 26166 12864 26166 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit5.Q
rlabel metal3 19056 24780 19056 24780 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 17280 25578 17280 25578 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 11184 18732 11184 18732 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 9504 18984 9504 18984 0 Inst_W_TT_IF_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 10752 16345 10752 16345 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 8736 17094 8736 17094 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 17472 20454 17472 20454 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 12864 4620 12864 4620 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 11520 3024 11520 3024 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 11712 3612 11712 3612 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 13248 4998 13248 4998 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 12096 7308 12096 7308 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 13536 6972 13536 6972 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit16.Q
rlabel via2 17280 23774 17280 23774 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 19488 22218 19488 22218 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit18.Q
rlabel metal3 18240 22512 18240 22512 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 11904 12474 11904 12474 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 15648 29484 15648 29484 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit20.Q
rlabel metal3 15888 31332 15888 31332 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 16704 31479 16704 31479 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit22.Q
rlabel metal2 14688 13986 14688 13986 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit23.Q
rlabel metal3 15264 14028 15264 14028 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 15792 12600 15792 12600 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 14832 19488 14832 19488 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit26.Q
rlabel metal3 13056 20706 13056 20706 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 19008 29568 19008 29568 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 17376 30114 17376 30114 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit29.Q
rlabel metal3 12000 11508 12000 11508 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 16608 25032 16608 25032 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 14976 25620 14976 25620 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 13056 12558 13056 12558 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 13728 33138 13728 33138 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 14496 35112 14496 35112 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 15072 36960 15072 36960 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit7.Q
rlabel metal3 16704 20748 16704 20748 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit8.Q
rlabel metal2 18624 21630 18624 21630 0 Inst_W_TT_IF_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 8544 16800 8544 16800 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 2400 21084 2400 21084 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 9792 14952 9792 14952 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 11904 14112 11904 14112 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 11616 13944 11616 13944 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 7680 34692 7680 34692 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 9216 27552 9216 27552 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 9024 27216 9024 27216 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 4992 26208 4992 26208 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit16.Q
rlabel metal3 5760 35868 5760 35868 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit17.Q
rlabel metal3 4944 35868 4944 35868 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 1632 10080 1632 10080 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 4128 21627 4128 21627 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 1536 12348 1536 12348 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit20.Q
rlabel metal3 1296 11676 1296 11676 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit21.Q
rlabel via2 4320 14700 4320 14700 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 3269 10957 3269 10957 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 1536 16128 1536 16128 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 12480 30114 12480 30114 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 11808 27678 11808 27678 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit26.Q
rlabel metal3 12048 29064 12048 29064 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 12864 32928 12864 32928 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 11712 32130 11712 32130 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 4416 21588 4416 21588 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 12960 32130 12960 32130 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 9216 15246 9216 15246 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit31.Q
rlabel metal2 2640 18564 2640 18564 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 4224 18305 4224 18305 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 4416 17976 4416 17976 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 2304 15036 2304 15036 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 3840 16088 3840 16088 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 2784 14196 2784 14196 0 Inst_W_TT_IF_ConfigMem.Inst_frame6_bit9.Q
rlabel metal3 7056 5880 7056 5880 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 7584 6090 7584 6090 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit1.Q
rlabel metal2 8256 4368 8256 4368 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 6336 5166 6336 5166 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit11.Q
rlabel metal3 10128 2100 10128 2100 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 7488 1218 7488 1218 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit13.Q
rlabel metal3 4752 3276 4752 3276 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 14208 756 14208 756 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 10272 6678 10272 6678 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit16.Q
rlabel metal3 8112 17724 8112 17724 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 14784 10213 14784 10213 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 14592 8148 14592 8148 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 6624 8946 6624 8946 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 13248 10836 13248 10836 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 15744 15792 15744 15792 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 17664 14658 17664 14658 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 15936 16380 15936 16380 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit23.Q
rlabel metal3 14592 37212 14592 37212 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit24.Q
rlabel metal3 17136 40404 17136 40404 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit25.Q
rlabel metal3 17376 38892 17376 38892 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit26.Q
rlabel metal3 13296 1764 13296 1764 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit27.Q
rlabel metal3 16272 1680 16272 1680 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 12000 2184 12000 2184 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 8160 8743 8160 8743 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 6240 17388 6240 17388 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit30.Q
rlabel metal2 7776 17684 7776 17684 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 7200 15582 7200 15582 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit4.Q
rlabel metal4 8928 14364 8928 14364 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 8640 3612 8640 3612 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 3456 4410 3456 4410 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 8448 2653 8448 2653 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit8.Q
rlabel metal3 5232 1764 5232 1764 0 Inst_W_TT_IF_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 2640 37380 2640 37380 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit0.Q
rlabel metal4 15456 38094 15456 38094 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit1.Q
rlabel metal2 3456 32883 3456 32883 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit10.Q
rlabel metal3 4608 32172 4608 32172 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit11.Q
rlabel metal3 6288 6636 6288 6636 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit12.Q
rlabel metal2 5856 7686 5856 7686 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit13.Q
rlabel metal2 8544 11046 8544 11046 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit14.Q
rlabel metal3 4176 7392 4176 7392 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit15.Q
rlabel metal3 5952 11676 5952 11676 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit16.Q
rlabel metal2 9936 35868 9936 35868 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit17.Q
rlabel metal3 13920 36078 13920 36078 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit18.Q
rlabel metal2 12048 33852 12048 33852 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit19.Q
rlabel metal2 7344 19488 7344 19488 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit2.Q
rlabel metal2 15072 39774 15072 39774 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit20.Q
rlabel metal3 16704 41244 16704 41244 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit21.Q
rlabel metal2 12000 38640 12000 38640 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit22.Q
rlabel metal2 19776 9072 19776 9072 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit23.Q
rlabel metal2 19680 11424 19680 11424 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 19872 10710 19872 10710 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 6624 13104 6624 13104 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit26.Q
rlabel metal2 8208 11844 8208 11844 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 8640 32214 8640 32214 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit28.Q
rlabel metal2 7104 32799 7104 32799 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit29.Q
rlabel metal3 7968 18732 7968 18732 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit3.Q
rlabel metal2 7968 34566 7968 34566 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit30.Q
rlabel metal2 9552 34419 9552 34419 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 4032 10255 4032 10255 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit4.Q
rlabel metal2 3264 9744 3264 9744 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit5.Q
rlabel metal2 13680 3192 13680 3192 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit6.Q
rlabel metal2 2736 10836 2736 10836 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit7.Q
rlabel metal3 3456 25284 3456 25284 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit8.Q
rlabel metal3 4176 26292 4176 26292 0 Inst_W_TT_IF_ConfigMem.Inst_frame8_bit9.Q
rlabel metal2 7584 12558 7584 12558 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit22.Q
rlabel via1 6000 12511 6000 12511 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit23.Q
rlabel metal2 8256 33138 8256 33138 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit24.Q
rlabel via1 6672 32874 6672 32874 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit25.Q
rlabel metal2 12096 37044 12096 37044 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit26.Q
rlabel metal2 1824 37681 1824 37681 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit27.Q
rlabel metal2 8304 2100 8304 2100 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit28.Q
rlabel metal2 2832 5880 2832 5880 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit29.Q
rlabel metal2 3600 7392 3600 7392 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit30.Q
rlabel metal4 5664 7812 5664 7812 0 Inst_W_TT_IF_ConfigMem.Inst_frame9_bit31.Q
rlabel metal3 10944 16716 10944 16716 0 Inst_W_TT_IF_switch_matrix.E1BEG0
rlabel metal3 18528 17808 18528 17808 0 Inst_W_TT_IF_switch_matrix.E1BEG1
rlabel metal2 18144 16422 18144 16422 0 Inst_W_TT_IF_switch_matrix.E1BEG2
rlabel metal4 16416 14028 16416 14028 0 Inst_W_TT_IF_switch_matrix.E1BEG3
rlabel metal3 15648 14322 15648 14322 0 Inst_W_TT_IF_switch_matrix.E2BEG0
rlabel metal3 18912 30366 18912 30366 0 Inst_W_TT_IF_switch_matrix.E2BEG1
rlabel metal2 19776 31878 19776 31878 0 Inst_W_TT_IF_switch_matrix.E2BEG2
rlabel metal2 16992 12894 16992 12894 0 Inst_W_TT_IF_switch_matrix.E2BEG3
rlabel metal4 17472 13062 17472 13062 0 Inst_W_TT_IF_switch_matrix.E2BEG4
rlabel metal3 16464 29652 16464 29652 0 Inst_W_TT_IF_switch_matrix.E2BEG5
rlabel metal2 18624 31962 18624 31962 0 Inst_W_TT_IF_switch_matrix.E2BEG6
rlabel metal4 17664 15246 17664 15246 0 Inst_W_TT_IF_switch_matrix.E2BEG7
rlabel metal3 14208 11760 14208 11760 0 Inst_W_TT_IF_switch_matrix.E2BEGb0
rlabel metal2 19248 33096 19248 33096 0 Inst_W_TT_IF_switch_matrix.E2BEGb1
rlabel metal4 19776 19194 19776 19194 0 Inst_W_TT_IF_switch_matrix.E2BEGb2
rlabel metal2 19872 5166 19872 5166 0 Inst_W_TT_IF_switch_matrix.E2BEGb3
rlabel metal2 14688 7476 14688 7476 0 Inst_W_TT_IF_switch_matrix.E2BEGb4
rlabel metal2 20016 22344 20016 22344 0 Inst_W_TT_IF_switch_matrix.E2BEGb5
rlabel metal2 19392 32046 19392 32046 0 Inst_W_TT_IF_switch_matrix.E2BEGb6
rlabel metal2 16128 14196 16128 14196 0 Inst_W_TT_IF_switch_matrix.E2BEGb7
rlabel metal2 17472 27468 17472 27468 0 Inst_W_TT_IF_switch_matrix.E6BEG0
rlabel metal3 12240 36792 12240 36792 0 Inst_W_TT_IF_switch_matrix.E6BEG1
rlabel metal3 19008 35280 19008 35280 0 Inst_W_TT_IF_switch_matrix.E6BEG10
rlabel metal3 18864 35112 18864 35112 0 Inst_W_TT_IF_switch_matrix.E6BEG11
rlabel metal2 13536 36078 13536 36078 0 Inst_W_TT_IF_switch_matrix.E6BEG2
rlabel metal2 17088 26922 17088 26922 0 Inst_W_TT_IF_switch_matrix.E6BEG3
rlabel metal2 19392 29652 19392 29652 0 Inst_W_TT_IF_switch_matrix.E6BEG4
rlabel metal2 19152 32088 19152 32088 0 Inst_W_TT_IF_switch_matrix.E6BEG5
rlabel metal2 19296 34986 19296 34986 0 Inst_W_TT_IF_switch_matrix.E6BEG6
rlabel metal3 17856 33180 17856 33180 0 Inst_W_TT_IF_switch_matrix.E6BEG7
rlabel metal2 19392 32844 19392 32844 0 Inst_W_TT_IF_switch_matrix.E6BEG8
rlabel metal3 19008 35952 19008 35952 0 Inst_W_TT_IF_switch_matrix.E6BEG9
rlabel metal2 19488 24486 19488 24486 0 Inst_W_TT_IF_switch_matrix.EE4BEG0
rlabel metal2 19872 31080 19872 31080 0 Inst_W_TT_IF_switch_matrix.EE4BEG1
rlabel metal2 19776 27804 19776 27804 0 Inst_W_TT_IF_switch_matrix.EE4BEG10
rlabel metal2 11712 20370 11712 20370 0 Inst_W_TT_IF_switch_matrix.EE4BEG11
rlabel metal2 14544 24780 14544 24780 0 Inst_W_TT_IF_switch_matrix.EE4BEG12
rlabel metal2 19632 29064 19632 29064 0 Inst_W_TT_IF_switch_matrix.EE4BEG13
rlabel metal3 18288 29904 18288 29904 0 Inst_W_TT_IF_switch_matrix.EE4BEG14
rlabel metal3 19392 27174 19392 27174 0 Inst_W_TT_IF_switch_matrix.EE4BEG15
rlabel metal3 18240 26040 18240 26040 0 Inst_W_TT_IF_switch_matrix.EE4BEG2
rlabel metal2 19392 25662 19392 25662 0 Inst_W_TT_IF_switch_matrix.EE4BEG3
rlabel metal2 19296 25746 19296 25746 0 Inst_W_TT_IF_switch_matrix.EE4BEG4
rlabel metal2 14592 26922 14592 26922 0 Inst_W_TT_IF_switch_matrix.EE4BEG5
rlabel metal2 19776 26544 19776 26544 0 Inst_W_TT_IF_switch_matrix.EE4BEG6
rlabel metal3 15312 19992 15312 19992 0 Inst_W_TT_IF_switch_matrix.EE4BEG7
rlabel metal2 19392 26670 19392 26670 0 Inst_W_TT_IF_switch_matrix.EE4BEG8
rlabel metal2 19728 33600 19728 33600 0 Inst_W_TT_IF_switch_matrix.EE4BEG9
rlabel metal3 1968 18984 1968 18984 0 Inst_W_TT_IF_switch_matrix.N1BEG0
rlabel metal3 6432 32508 6432 32508 0 Inst_W_TT_IF_switch_matrix.N1BEG1
rlabel metal3 1104 30576 1104 30576 0 Inst_W_TT_IF_switch_matrix.N1BEG2
rlabel metal2 3072 25074 3072 25074 0 Inst_W_TT_IF_switch_matrix.N1BEG3
rlabel metal3 864 8736 864 8736 0 Inst_W_TT_IF_switch_matrix.N2BEG0
rlabel metal2 3072 32382 3072 32382 0 Inst_W_TT_IF_switch_matrix.N2BEG1
rlabel metal3 1200 35112 1200 35112 0 Inst_W_TT_IF_switch_matrix.N2BEG2
rlabel metal3 6480 10836 6480 10836 0 Inst_W_TT_IF_switch_matrix.N2BEG3
rlabel metal3 912 35952 912 35952 0 Inst_W_TT_IF_switch_matrix.N2BEG4
rlabel metal3 1296 35364 1296 35364 0 Inst_W_TT_IF_switch_matrix.N2BEG5
rlabel metal3 3312 32340 3312 32340 0 Inst_W_TT_IF_switch_matrix.N2BEG6
rlabel metal2 1488 22344 1488 22344 0 Inst_W_TT_IF_switch_matrix.N2BEG7
rlabel metal6 11728 16716 11728 16716 0 Inst_W_TT_IF_switch_matrix.N4BEG0
rlabel via2 18143 38976 18143 38976 0 Inst_W_TT_IF_switch_matrix.N4BEG1
rlabel metal2 10560 40530 10560 40530 0 Inst_W_TT_IF_switch_matrix.N4BEG2
rlabel metal5 15120 11172 15120 11172 0 Inst_W_TT_IF_switch_matrix.N4BEG3
rlabel metal3 6480 13104 6480 13104 0 Inst_W_TT_IF_switch_matrix.S1BEG0
rlabel metal5 1160 1176 1160 1176 0 Inst_W_TT_IF_switch_matrix.S1BEG1
rlabel metal3 10512 13188 10512 13188 0 Inst_W_TT_IF_switch_matrix.S1BEG2
rlabel metal3 1104 3948 1104 3948 0 Inst_W_TT_IF_switch_matrix.S1BEG3
rlabel metal2 11520 7854 11520 7854 0 Inst_W_TT_IF_switch_matrix.S2BEG0
rlabel metal5 14304 1848 14304 1848 0 Inst_W_TT_IF_switch_matrix.S2BEG1
rlabel metal3 7680 4872 7680 4872 0 Inst_W_TT_IF_switch_matrix.S2BEG2
rlabel metal3 9312 2436 9312 2436 0 Inst_W_TT_IF_switch_matrix.S2BEG3
rlabel metal3 6816 2184 6816 2184 0 Inst_W_TT_IF_switch_matrix.S2BEG4
rlabel metal2 8496 3528 8496 3528 0 Inst_W_TT_IF_switch_matrix.S2BEG5
rlabel metal2 4896 1092 4896 1092 0 Inst_W_TT_IF_switch_matrix.S2BEG6
rlabel metal2 5088 2730 5088 2730 0 Inst_W_TT_IF_switch_matrix.S2BEG7
rlabel metal3 19248 1764 19248 1764 0 Inst_W_TT_IF_switch_matrix.S4BEG0
rlabel metal4 12384 1806 12384 1806 0 Inst_W_TT_IF_switch_matrix.S4BEG1
rlabel metal2 20448 1176 20448 1176 0 Inst_W_TT_IF_switch_matrix.S4BEG2
rlabel metal2 11088 1932 11088 1932 0 Inst_W_TT_IF_switch_matrix.S4BEG3
rlabel metal2 1728 22554 1728 22554 0 N1BEG[0]
rlabel metal3 1296 23268 1296 23268 0 N1BEG[1]
rlabel metal2 1440 31542 1440 31542 0 N1BEG[2]
rlabel metal3 1008 30156 1008 30156 0 N1BEG[3]
rlabel metal2 1872 3780 1872 3780 0 N1END[0]
rlabel metal2 2016 492 2016 492 0 N1END[1]
rlabel metal2 2208 828 2208 828 0 N1END[2]
rlabel metal2 2496 16548 2496 16548 0 N1END[3]
rlabel metal2 4800 30828 4800 30828 0 N2BEG[0]
rlabel metal2 2880 34566 2880 34566 0 N2BEG[1]
rlabel metal2 1728 35196 1728 35196 0 N2BEG[2]
rlabel metal2 4512 27006 4512 27006 0 N2BEG[3]
rlabel metal2 1776 36120 1776 36120 0 N2BEG[4]
rlabel metal2 2592 36288 2592 36288 0 N2BEG[5]
rlabel metal2 4416 38472 4416 38472 0 N2BEG[6]
rlabel metal3 1248 22512 1248 22512 0 N2BEG[7]
rlabel metal2 1536 36918 1536 36918 0 N2BEGb[0]
rlabel metal2 4272 38388 4272 38388 0 N2BEGb[1]
rlabel metal2 3360 34650 3360 34650 0 N2BEGb[2]
rlabel metal2 1920 40236 1920 40236 0 N2BEGb[3]
rlabel metal3 2352 33096 2352 33096 0 N2BEGb[4]
rlabel metal3 1344 21756 1344 21756 0 N2BEGb[5]
rlabel metal2 5280 42726 5280 42726 0 N2BEGb[6]
rlabel metal3 5280 39060 5280 39060 0 N2BEGb[7]
rlabel metal2 4128 576 4128 576 0 N2END[0]
rlabel metal2 4320 786 4320 786 0 N2END[1]
rlabel metal2 4608 1638 4608 1638 0 N2END[2]
rlabel metal2 4704 576 4704 576 0 N2END[3]
rlabel metal2 4896 324 4896 324 0 N2END[4]
rlabel metal4 11712 8946 11712 8946 0 N2END[5]
rlabel metal4 13152 20748 13152 20748 0 N2END[6]
rlabel metal2 5472 366 5472 366 0 N2END[7]
rlabel metal2 1392 19824 1392 19824 0 N2MID[0]
rlabel metal3 768 30408 768 30408 0 N2MID[1]
rlabel metal5 1968 18564 1968 18564 0 N2MID[2]
rlabel metal2 2112 1638 2112 1638 0 N2MID[3]
rlabel metal4 2208 27972 2208 27972 0 N2MID[4]
rlabel metal2 1344 21588 1344 21588 0 N2MID[5]
rlabel metal4 2112 30366 2112 30366 0 N2MID[6]
rlabel metal2 3936 408 3936 408 0 N2MID[7]
rlabel metal2 7488 40698 7488 40698 0 N4BEG[0]
rlabel metal3 4416 29064 4416 29064 0 N4BEG[10]
rlabel metal2 8256 40572 8256 40572 0 N4BEG[11]
rlabel metal3 5904 28476 5904 28476 0 N4BEG[12]
rlabel metal2 17904 41076 17904 41076 0 N4BEG[13]
rlabel metal2 10368 40740 10368 40740 0 N4BEG[14]
rlabel metal3 7248 23268 7248 23268 0 N4BEG[15]
rlabel metal5 2036 21756 2036 21756 0 N4BEG[1]
rlabel metal3 4992 28560 4992 28560 0 N4BEG[2]
rlabel metal3 5088 35364 5088 35364 0 N4BEG[3]
rlabel metal3 1968 38388 1968 38388 0 N4BEG[4]
rlabel metal3 5568 22512 5568 22512 0 N4BEG[5]
rlabel metal3 6336 25536 6336 25536 0 N4BEG[6]
rlabel metal2 5760 37296 5760 37296 0 N4BEG[7]
rlabel metal3 7152 32004 7152 32004 0 N4BEG[8]
rlabel metal4 1536 22554 1536 22554 0 N4BEG[9]
rlabel metal2 5664 534 5664 534 0 N4END[0]
rlabel metal2 7584 492 7584 492 0 N4END[10]
rlabel metal2 7776 660 7776 660 0 N4END[11]
rlabel metal2 7968 450 7968 450 0 N4END[12]
rlabel metal3 1392 20832 1392 20832 0 N4END[13]
rlabel metal2 8352 660 8352 660 0 N4END[14]
rlabel metal2 8544 660 8544 660 0 N4END[15]
rlabel metal2 5856 366 5856 366 0 N4END[1]
rlabel metal2 6048 492 6048 492 0 N4END[2]
rlabel metal2 6240 660 6240 660 0 N4END[3]
rlabel metal3 6192 33852 6192 33852 0 N4END[4]
rlabel metal2 1728 21042 1728 21042 0 N4END[5]
rlabel metal2 6816 660 6816 660 0 N4END[6]
rlabel metal2 7008 660 7008 660 0 N4END[7]
rlabel metal3 1440 38136 1440 38136 0 N4END[8]
rlabel metal2 7392 492 7392 492 0 N4END[9]
rlabel metal2 1824 4284 1824 4284 0 RST_N_TT_PROJECT
rlabel metal2 8736 1290 8736 1290 0 S1BEG[0]
rlabel metal2 1728 714 1728 714 0 S1BEG[1]
rlabel metal2 9120 576 9120 576 0 S1BEG[2]
rlabel metal2 1440 1554 1440 1554 0 S1BEG[3]
rlabel metal3 8256 17094 8256 17094 0 S1END[0]
rlabel metal2 1344 34524 1344 34524 0 S1END[1]
rlabel metal3 4320 36624 4320 36624 0 S1END[2]
rlabel metal2 2400 24822 2400 24822 0 S1END[3]
rlabel metal2 9504 408 9504 408 0 S2BEG[0]
rlabel metal2 17568 1512 17568 1512 0 S2BEG[1]
rlabel metal2 9888 114 9888 114 0 S2BEG[2]
rlabel metal2 10128 3948 10128 3948 0 S2BEG[3]
rlabel metal2 10272 870 10272 870 0 S2BEG[4]
rlabel metal2 10368 3612 10368 3612 0 S2BEG[5]
rlabel metal2 10656 156 10656 156 0 S2BEG[6]
rlabel metal3 5376 2436 5376 2436 0 S2BEG[7]
rlabel metal2 11040 282 11040 282 0 S2BEGb[0]
rlabel metal2 11232 492 11232 492 0 S2BEGb[1]
rlabel metal2 11424 114 11424 114 0 S2BEGb[2]
rlabel metal2 11616 828 11616 828 0 S2BEGb[3]
rlabel metal2 11712 1890 11712 1890 0 S2BEGb[4]
rlabel metal2 12000 660 12000 660 0 S2BEGb[5]
rlabel metal2 11472 2436 11472 2436 0 S2BEGb[6]
rlabel metal2 12384 786 12384 786 0 S2BEGb[7]
rlabel metal3 9984 27888 9984 27888 0 S2END[0]
rlabel metal3 11088 36120 11088 36120 0 S2END[1]
rlabel metal2 11424 42306 11424 42306 0 S2END[2]
rlabel metal2 1536 2100 1536 2100 0 S2END[3]
rlabel metal2 11808 42264 11808 42264 0 S2END[4]
rlabel metal2 12000 42726 12000 42726 0 S2END[5]
rlabel metal2 12192 42264 12192 42264 0 S2END[6]
rlabel metal2 12384 42264 12384 42264 0 S2END[7]
rlabel metal2 864 12516 864 12516 0 S2MID[0]
rlabel metal3 9360 1176 9360 1176 0 S2MID[1]
rlabel metal2 4512 2142 4512 2142 0 S2MID[2]
rlabel metal2 2496 1218 2496 1218 0 S2MID[3]
rlabel metal2 12192 4326 12192 4326 0 S2MID[4]
rlabel metal4 12576 35070 12576 35070 0 S2MID[5]
rlabel metal3 12336 1176 12336 1176 0 S2MID[6]
rlabel metal3 13968 2856 13968 2856 0 S2MID[7]
rlabel metal2 12576 492 12576 492 0 S4BEG[0]
rlabel metal2 14496 660 14496 660 0 S4BEG[10]
rlabel metal2 14688 660 14688 660 0 S4BEG[11]
rlabel metal2 14880 282 14880 282 0 S4BEG[12]
rlabel metal2 15072 240 15072 240 0 S4BEG[13]
rlabel metal2 15264 450 15264 450 0 S4BEG[14]
rlabel metal2 15456 744 15456 744 0 S4BEG[15]
rlabel metal2 12768 282 12768 282 0 S4BEG[1]
rlabel metal2 12960 492 12960 492 0 S4BEG[2]
rlabel metal2 13152 450 13152 450 0 S4BEG[3]
rlabel metal2 13344 660 13344 660 0 S4BEG[4]
rlabel metal2 13536 492 13536 492 0 S4BEG[5]
rlabel metal2 13728 492 13728 492 0 S4BEG[6]
rlabel metal2 13920 366 13920 366 0 S4BEG[7]
rlabel metal2 14112 744 14112 744 0 S4BEG[8]
rlabel metal2 14304 660 14304 660 0 S4BEG[9]
rlabel metal2 12576 42558 12576 42558 0 S4END[0]
rlabel metal2 14496 42306 14496 42306 0 S4END[10]
rlabel metal2 1248 42042 1248 42042 0 S4END[11]
rlabel metal2 14880 41886 14880 41886 0 S4END[12]
rlabel metal2 15072 42432 15072 42432 0 S4END[13]
rlabel metal2 18528 39858 18528 39858 0 S4END[14]
rlabel metal2 15456 42054 15456 42054 0 S4END[15]
rlabel metal2 8352 35700 8352 35700 0 S4END[1]
rlabel metal3 12480 36708 12480 36708 0 S4END[2]
rlabel metal2 13344 35364 13344 35364 0 S4END[3]
rlabel metal2 13344 42558 13344 42558 0 S4END[4]
rlabel metal2 13536 42516 13536 42516 0 S4END[5]
rlabel metal2 13728 42474 13728 42474 0 S4END[6]
rlabel metal2 13920 42600 13920 42600 0 S4END[7]
rlabel metal2 14112 41718 14112 41718 0 S4END[8]
rlabel metal2 14304 41676 14304 41676 0 S4END[9]
rlabel metal3 11664 10332 11664 10332 0 UIO_IN_TT_PROJECT0
rlabel metal3 702 19404 702 19404 0 UIO_IN_TT_PROJECT1
rlabel metal3 654 19908 654 19908 0 UIO_IN_TT_PROJECT2
rlabel metal3 174 20412 174 20412 0 UIO_IN_TT_PROJECT3
rlabel metal3 14448 13524 14448 13524 0 UIO_IN_TT_PROJECT4
rlabel metal2 12480 17808 12480 17808 0 UIO_IN_TT_PROJECT5
rlabel metal3 558 21924 558 21924 0 UIO_IN_TT_PROJECT6
rlabel metal3 11904 18900 11904 18900 0 UIO_IN_TT_PROJECT7
rlabel metal2 6336 17094 6336 17094 0 UIO_OE_TT_PROJECT0
rlabel metal4 1488 16296 1488 16296 0 UIO_OE_TT_PROJECT1
rlabel metal3 270 11844 270 11844 0 UIO_OE_TT_PROJECT2
rlabel metal3 3360 18480 3360 18480 0 UIO_OE_TT_PROJECT3
rlabel metal2 13632 19068 13632 19068 0 UIO_OE_TT_PROJECT4
rlabel metal3 894 13356 894 13356 0 UIO_OE_TT_PROJECT5
rlabel metal3 606 13860 606 13860 0 UIO_OE_TT_PROJECT6
rlabel metal3 606 14364 606 14364 0 UIO_OE_TT_PROJECT7
rlabel metal2 13632 13566 13632 13566 0 UIO_OUT_TT_PROJECT0
rlabel metal3 318 7308 318 7308 0 UIO_OUT_TT_PROJECT1
rlabel metal2 17568 34776 17568 34776 0 UIO_OUT_TT_PROJECT2
rlabel metal2 12384 18438 12384 18438 0 UIO_OUT_TT_PROJECT3
rlabel metal2 13488 18732 13488 18732 0 UIO_OUT_TT_PROJECT4
rlabel metal3 16416 12852 16416 12852 0 UIO_OUT_TT_PROJECT5
rlabel metal2 14784 33264 14784 33264 0 UIO_OUT_TT_PROJECT6
rlabel metal2 14160 18984 14160 18984 0 UIO_OUT_TT_PROJECT7
rlabel metal3 654 14868 654 14868 0 UI_IN_TT_PROJECT0
rlabel metal4 14688 15036 14688 15036 0 UI_IN_TT_PROJECT1
rlabel metal4 12576 16086 12576 16086 0 UI_IN_TT_PROJECT2
rlabel metal3 510 16380 510 16380 0 UI_IN_TT_PROJECT3
rlabel metal3 654 16884 654 16884 0 UI_IN_TT_PROJECT4
rlabel via2 78 17388 78 17388 0 UI_IN_TT_PROJECT5
rlabel metal3 318 17892 318 17892 0 UI_IN_TT_PROJECT6
rlabel metal3 654 18396 654 18396 0 UI_IN_TT_PROJECT7
rlabel metal3 1824 14406 1824 14406 0 UO_OUT_TT_PROJECT0
rlabel metal3 336 17304 336 17304 0 UO_OUT_TT_PROJECT1
rlabel metal3 720 17640 720 17640 0 UO_OUT_TT_PROJECT2
rlabel metal3 174 4284 174 4284 0 UO_OUT_TT_PROJECT3
rlabel metal2 2112 17010 2112 17010 0 UO_OUT_TT_PROJECT4
rlabel metal3 126 5292 126 5292 0 UO_OUT_TT_PROJECT5
rlabel metal3 270 5796 270 5796 0 UO_OUT_TT_PROJECT6
rlabel metal3 222 6300 222 6300 0 UO_OUT_TT_PROJECT7
rlabel metal2 15648 156 15648 156 0 UserCLK
rlabel metal2 19392 41118 19392 41118 0 UserCLKo
rlabel metal3 21330 84 21330 84 0 W1END[0]
rlabel metal3 20562 420 20562 420 0 W1END[1]
rlabel metal4 20544 1344 20544 1344 0 W1END[2]
rlabel metal3 20802 1092 20802 1092 0 W1END[3]
rlabel metal2 13248 11760 13248 11760 0 W2END[0]
rlabel metal2 14016 15498 14016 15498 0 W2END[1]
rlabel metal2 16896 17682 16896 17682 0 W2END[2]
rlabel metal2 12192 7056 12192 7056 0 W2END[3]
rlabel metal2 12768 3948 12768 3948 0 W2END[4]
rlabel metal3 14160 19572 14160 19572 0 W2END[5]
rlabel metal2 16032 36078 16032 36078 0 W2END[6]
rlabel metal2 16608 5964 16608 5964 0 W2END[7]
rlabel metal3 20802 1428 20802 1428 0 W2MID[0]
rlabel metal3 21090 1764 21090 1764 0 W2MID[1]
rlabel metal3 21042 2100 21042 2100 0 W2MID[2]
rlabel metal3 21138 2436 21138 2436 0 W2MID[3]
rlabel metal3 19296 3066 19296 3066 0 W2MID[4]
rlabel metal2 19488 12474 19488 12474 0 W2MID[5]
rlabel metal3 7248 15540 7248 15540 0 W2MID[6]
rlabel metal2 6720 8526 6720 8526 0 W2MID[7]
rlabel metal3 21138 12180 21138 12180 0 W6END[0]
rlabel metal3 14016 18900 14016 18900 0 W6END[10]
rlabel metal3 19536 7140 19536 7140 0 W6END[11]
rlabel metal3 19296 12474 19296 12474 0 W6END[1]
rlabel metal2 16704 19194 16704 19194 0 W6END[2]
rlabel metal3 20994 13188 20994 13188 0 W6END[3]
rlabel metal2 18480 12348 18480 12348 0 W6END[4]
rlabel metal2 15408 16212 15408 16212 0 W6END[5]
rlabel metal3 15696 36708 15696 36708 0 W6END[6]
rlabel metal2 17568 2562 17568 2562 0 W6END[7]
rlabel metal2 7296 12054 7296 12054 0 W6END[8]
rlabel metal3 13920 15414 13920 15414 0 W6END[9]
rlabel metal2 12864 8484 12864 8484 0 WW4END[0]
rlabel metal2 19296 19320 19296 19320 0 WW4END[10]
rlabel metal2 19680 5880 19680 5880 0 WW4END[11]
rlabel metal3 16704 10878 16704 10878 0 WW4END[12]
rlabel metal2 19296 13188 19296 13188 0 WW4END[13]
rlabel metal3 16752 14532 16752 14532 0 WW4END[14]
rlabel metal3 19074 11844 19074 11844 0 WW4END[15]
rlabel metal3 14544 14616 14544 14616 0 WW4END[1]
rlabel metal2 19872 19110 19872 19110 0 WW4END[2]
rlabel metal3 18912 8106 18912 8106 0 WW4END[3]
rlabel metal2 17568 8400 17568 8400 0 WW4END[4]
rlabel metal3 21042 8484 21042 8484 0 WW4END[5]
rlabel metal3 20256 33894 20256 33894 0 WW4END[6]
rlabel metal2 16608 5124 16608 5124 0 WW4END[7]
rlabel metal2 18528 8988 18528 8988 0 WW4END[8]
rlabel metal2 13920 15204 13920 15204 0 WW4END[9]
rlabel metal3 5568 5628 5568 5628 0 _0000_
rlabel metal2 17376 3696 17376 3696 0 _0001_
rlabel metal2 5424 13776 5424 13776 0 _0002_
rlabel metal3 16656 5628 16656 5628 0 _0003_
rlabel metal3 14928 38892 14928 38892 0 _0004_
rlabel metal2 1152 29358 1152 29358 0 _0005_
rlabel metal3 19680 37716 19680 37716 0 _0006_
rlabel metal3 1536 32844 1536 32844 0 _0007_
rlabel metal2 16800 14196 16800 14196 0 _0008_
rlabel metal3 7296 16212 7296 16212 0 _0009_
rlabel metal2 16320 10332 16320 10332 0 _0010_
rlabel metal2 20400 2100 20400 2100 0 _0011_
rlabel metal2 19776 18774 19776 18774 0 _0012_
rlabel metal3 13680 17556 13680 17556 0 _0013_
rlabel metal3 13344 8694 13344 8694 0 _0014_
rlabel metal3 19056 36708 19056 36708 0 _0015_
rlabel metal2 19776 14448 19776 14448 0 _0016_
rlabel metal2 18144 9534 18144 9534 0 _0017_
rlabel metal2 11712 4284 11712 4284 0 _0018_
rlabel metal2 16992 19278 16992 19278 0 _0019_
rlabel metal2 13344 15330 13344 15330 0 _0020_
rlabel metal2 8640 6552 8640 6552 0 _0021_
rlabel metal3 3312 11424 3312 11424 0 _0022_
rlabel metal2 12000 27720 12000 27720 0 _0023_
rlabel metal3 11136 28308 11136 28308 0 _0024_
rlabel metal3 3024 16212 3024 16212 0 _0025_
rlabel metal2 2016 9324 2016 9324 0 _0026_
rlabel metal2 1248 11424 1248 11424 0 _0027_
rlabel metal2 1440 27258 1440 27258 0 _0028_
rlabel metal2 6864 32424 6864 32424 0 _0029_
rlabel metal2 11232 14994 11232 14994 0 _0030_
rlabel metal3 13536 1596 13536 1596 0 _0031_
rlabel metal3 15600 37296 15600 37296 0 _0032_
rlabel metal2 18720 8022 18720 8022 0 _0033_
rlabel metal2 14304 39018 14304 39018 0 _0034_
rlabel metal2 12864 35532 12864 35532 0 _0035_
rlabel metal3 6192 11592 6192 11592 0 _0036_
rlabel metal3 1584 17304 1584 17304 0 _0037_
rlabel metal4 2304 15078 2304 15078 0 _0038_
rlabel metal2 2208 5922 2208 5922 0 _0039_
rlabel metal2 3840 3318 3840 3318 0 _0040_
rlabel metal2 5760 3150 5760 3150 0 _0041_
rlabel metal2 1728 3948 1728 3948 0 _0042_
rlabel metal2 6864 4116 6864 4116 0 _0043_
rlabel metal2 7680 4704 7680 4704 0 _0044_
rlabel metal2 1248 4872 1248 4872 0 _0045_
rlabel metal2 2496 4410 2496 4410 0 _0046_
rlabel metal3 1872 5628 1872 5628 0 _0047_
rlabel metal2 1248 5502 1248 5502 0 _0048_
rlabel metal2 1536 4788 1536 4788 0 _0049_
rlabel metal2 1632 4032 1632 4032 0 _0050_
rlabel metal2 13920 5082 13920 5082 0 _0051_
rlabel metal2 14976 7014 14976 7014 0 _0052_
rlabel metal2 15552 12684 15552 12684 0 _0053_
rlabel metal2 15456 7182 15456 7182 0 _0054_
rlabel via1 16852 6467 16852 6467 0 _0055_
rlabel metal2 17088 6300 17088 6300 0 _0056_
rlabel metal2 15840 6720 15840 6720 0 _0057_
rlabel metal2 16896 5124 16896 5124 0 _0058_
rlabel metal2 15552 7098 15552 7098 0 _0059_
rlabel metal2 16704 29946 16704 29946 0 _0060_
rlabel metal2 18480 35196 18480 35196 0 _0061_
rlabel metal3 16368 37548 16368 37548 0 _0062_
rlabel metal3 18288 36876 18288 36876 0 _0063_
rlabel metal2 18626 37884 18626 37884 0 _0064_
rlabel metal2 19392 39060 19392 39060 0 _0065_
rlabel metal2 18240 38682 18240 38682 0 _0066_
rlabel metal3 18528 37632 18528 37632 0 _0067_
rlabel metal3 18864 38976 18864 38976 0 _0068_
rlabel metal3 17904 17052 17904 17052 0 _0069_
rlabel metal3 15648 16212 15648 16212 0 _0070_
rlabel metal2 17664 21924 17664 21924 0 _0071_
rlabel metal2 19968 16632 19968 16632 0 _0072_
rlabel metal2 20064 15540 20064 15540 0 _0073_
rlabel metal2 19488 15834 19488 15834 0 _0074_
rlabel metal2 19392 16548 19392 16548 0 _0075_
rlabel metal2 19872 15960 19872 15960 0 _0076_
rlabel metal2 19104 16926 19104 16926 0 _0077_
rlabel metal3 7536 13272 7536 13272 0 _0078_
rlabel metal2 13920 5754 13920 5754 0 _0079_
rlabel metal2 13920 5460 13920 5460 0 _0080_
rlabel metal2 16080 11928 16080 11928 0 _0081_
rlabel metal2 17147 11508 17147 11508 0 _0082_
rlabel metal3 17040 10752 17040 10752 0 _0083_
rlabel metal2 16704 12222 16704 12222 0 _0084_
rlabel metal2 16128 10290 16128 10290 0 _0085_
rlabel metal2 16416 11886 16416 11886 0 _0086_
rlabel metal3 11664 4116 11664 4116 0 _0087_
rlabel metal2 19104 9366 19104 9366 0 _0088_
rlabel metal2 18576 4788 18576 4788 0 _0089_
rlabel via1 19970 7140 19970 7140 0 _0090_
rlabel metal2 19776 6930 19776 6930 0 _0091_
rlabel metal2 19344 7980 19344 7980 0 _0092_
rlabel metal2 19392 6846 19392 6846 0 _0093_
rlabel metal2 19008 7854 19008 7854 0 _0094_
rlabel metal2 18000 31416 18000 31416 0 _0095_
rlabel metal3 12528 37296 12528 37296 0 _0096_
rlabel metal2 18336 19929 18336 19929 0 _0097_
rlabel via1 19949 18564 19949 18564 0 _0098_
rlabel metal2 19680 18984 19680 18984 0 _0099_
rlabel metal2 18720 19488 18720 19488 0 _0100_
rlabel metal2 19008 19908 19008 19908 0 _0101_
rlabel metal2 18432 20013 18432 20013 0 _0102_
rlabel metal2 16512 17136 16512 17136 0 _0103_
rlabel metal2 12576 14154 12576 14154 0 _0104_
rlabel metal2 14688 17787 14688 17787 0 _0105_
rlabel metal2 12733 19900 12733 19900 0 _0106_
rlabel metal3 15600 19824 15600 19824 0 _0107_
rlabel metal2 14304 18165 14304 18165 0 _0108_
rlabel metal2 16416 16926 16416 16926 0 _0109_
rlabel metal3 16320 17766 16320 17766 0 _0110_
rlabel metal2 7488 10794 7488 10794 0 _0111_
rlabel metal2 14496 27426 14496 27426 0 _0112_
rlabel metal2 11424 9576 11424 9576 0 _0113_
rlabel metal2 13152 9030 13152 9030 0 _0114_
rlabel metal3 13344 8148 13344 8148 0 _0115_
rlabel metal3 12048 10164 12048 10164 0 _0116_
rlabel metal2 11520 8904 11520 8904 0 _0117_
rlabel metal2 11328 10374 11328 10374 0 _0118_
rlabel metal2 19968 2814 19968 2814 0 _0119_
rlabel metal2 13680 1764 13680 1764 0 _0120_
rlabel metal2 17088 3696 17088 3696 0 _0121_
rlabel metal2 18048 4410 18048 4410 0 _0122_
rlabel metal2 19872 2688 19872 2688 0 _0123_
rlabel metal3 17664 4116 17664 4116 0 _0124_
rlabel metal2 19968 3528 19968 3528 0 _0125_
rlabel metal3 20064 3612 20064 3612 0 _0126_
rlabel metal2 15456 40362 15456 40362 0 _0127_
rlabel metal2 15552 37506 15552 37506 0 _0128_
rlabel metal2 16477 36427 16477 36427 0 _0129_
rlabel metal2 17088 36666 17088 36666 0 _0130_
rlabel metal2 15936 37086 15936 37086 0 _0131_
rlabel metal2 16800 36498 16800 36498 0 _0132_
rlabel metal2 15648 37338 15648 37338 0 _0133_
rlabel metal2 16320 15372 16320 15372 0 _0134_
rlabel metal2 18864 14028 18864 14028 0 _0135_
rlabel metal2 19968 12894 19968 12894 0 _0136_
rlabel metal3 19968 13146 19968 13146 0 _0137_
rlabel metal2 19296 13650 19296 13650 0 _0138_
rlabel metal2 19584 13692 19584 13692 0 _0139_
rlabel metal2 19008 13902 19008 13902 0 _0140_
rlabel metal2 13536 19740 13536 19740 0 _0141_
rlabel metal2 16224 9450 16224 9450 0 _0142_
rlabel metal2 18245 9450 18245 9450 0 _0143_
rlabel metal2 18048 9618 18048 9618 0 _0144_
rlabel metal2 16608 9576 16608 9576 0 _0145_
rlabel metal2 15744 9324 15744 9324 0 _0146_
rlabel metal2 16320 9450 16320 9450 0 _0147_
rlabel metal2 15600 2268 15600 2268 0 _0148_
rlabel metal3 19152 2100 19152 2100 0 _0149_
rlabel via1 19732 3444 19732 3444 0 _0150_
rlabel metal2 18432 4368 18432 4368 0 _0151_
rlabel metal2 19008 3318 19008 3318 0 _0152_
rlabel metal2 18720 4452 18720 4452 0 _0153_
rlabel metal2 18720 3570 18720 3570 0 _0154_
rlabel metal3 15936 20076 15936 20076 0 _0155_
rlabel metal2 16560 18648 16560 18648 0 _0156_
rlabel metal2 17472 18606 17472 18606 0 _0157_
rlabel metal2 15840 19656 15840 19656 0 _0158_
rlabel metal2 17088 17556 17088 17556 0 _0159_
rlabel metal2 15552 19446 15552 19446 0 _0160_
rlabel metal2 16800 17220 16800 17220 0 _0161_
rlabel metal3 13632 16296 13632 16296 0 _0162_
rlabel metal2 12864 14238 12864 14238 0 _0163_
rlabel metal2 14626 15364 14626 15364 0 _0164_
rlabel metal2 11808 15414 11808 15414 0 _0165_
rlabel metal2 14928 14700 14928 14700 0 _0166_
rlabel metal2 11520 15414 11520 15414 0 _0167_
rlabel metal3 13104 14784 13104 14784 0 _0168_
rlabel metal3 13488 19992 13488 19992 0 _0169_
rlabel metal3 11856 8316 11856 8316 0 _0170_
rlabel via1 10274 9492 10274 9492 0 _0171_
rlabel metal3 10080 9450 10080 9450 0 _0172_
rlabel metal2 10080 8610 10080 8610 0 _0173_
rlabel metal2 9792 10416 9792 10416 0 _0174_
rlabel metal2 9552 9660 9552 9660 0 _0175_
rlabel metal2 15120 14028 15120 14028 0 _0176_
rlabel metal2 15120 13188 15120 13188 0 _0177_
rlabel metal3 13296 12516 13296 12516 0 _0178_
rlabel metal2 13920 13230 13920 13230 0 _0179_
rlabel metal2 15264 13398 15264 13398 0 _0180_
rlabel metal2 15264 13020 15264 13020 0 _0181_
rlabel metal2 16128 12768 16128 12768 0 _0182_
rlabel metal2 16176 12348 16176 12348 0 _0183_
rlabel metal2 15456 32172 15456 32172 0 _0184_
rlabel metal2 16896 29862 16896 29862 0 _0185_
rlabel metal2 16416 29568 16416 29568 0 _0186_
rlabel metal2 16416 30282 16416 30282 0 _0187_
rlabel metal2 17040 29820 17040 29820 0 _0188_
rlabel metal2 17184 30072 17184 30072 0 _0189_
rlabel metal2 16176 30828 16176 30828 0 _0190_
rlabel metal2 18096 32172 18096 32172 0 _0191_
rlabel metal2 19440 23268 19440 23268 0 _0192_
rlabel metal2 19584 23856 19584 23856 0 _0193_
rlabel metal2 19968 23052 19968 23052 0 _0194_
rlabel metal2 19584 22554 19584 22554 0 _0195_
rlabel metal2 19824 22260 19824 22260 0 _0196_
rlabel metal2 19776 24318 19776 24318 0 _0197_
rlabel metal2 16992 23352 16992 23352 0 _0198_
rlabel metal2 17136 23268 17136 23268 0 _0199_
rlabel metal2 12960 6132 12960 6132 0 _0200_
rlabel metal2 13440 5922 13440 5922 0 _0201_
rlabel metal3 13680 7140 13680 7140 0 _0202_
rlabel metal3 13824 7392 13824 7392 0 _0203_
rlabel metal2 13632 6216 13632 6216 0 _0204_
rlabel metal3 13872 5712 13872 5712 0 _0205_
rlabel metal3 14160 6468 14160 6468 0 _0206_
rlabel metal2 14544 6636 14544 6636 0 _0207_
rlabel metal2 13152 5082 13152 5082 0 _0208_
rlabel metal2 12336 2604 12336 2604 0 _0209_
rlabel metal2 11136 4452 11136 4452 0 _0210_
rlabel metal2 11616 3696 11616 3696 0 _0211_
rlabel metal2 12096 3030 12096 3030 0 _0212_
rlabel metal3 12336 2688 12336 2688 0 _0213_
rlabel metal2 10560 4578 10560 4578 0 _0214_
rlabel metal2 15936 5460 15936 5460 0 _0215_
rlabel metal2 19680 21588 19680 21588 0 _0216_
rlabel metal3 18576 21420 18576 21420 0 _0217_
rlabel metal3 18576 20076 18576 20076 0 _0218_
rlabel metal3 18336 20244 18336 20244 0 _0219_
rlabel metal2 18240 19698 18240 19698 0 _0220_
rlabel metal2 17568 19530 17568 19530 0 _0221_
rlabel metal2 20064 20706 20064 20706 0 _0222_
rlabel metal2 19872 20832 19872 20832 0 _0223_
rlabel metal2 16032 32844 16032 32844 0 _0224_
rlabel metal2 16128 33852 16128 33852 0 _0225_
rlabel metal2 14400 32214 14400 32214 0 _0226_
rlabel metal2 14496 33264 14496 33264 0 _0227_
rlabel metal2 15360 35406 15360 35406 0 _0228_
rlabel metal2 18912 32886 18912 32886 0 _0229_
rlabel metal2 17472 36036 17472 36036 0 _0230_
rlabel metal3 17952 32844 17952 32844 0 _0231_
rlabel metal2 11616 12516 11616 12516 0 _0232_
rlabel metal3 11760 10668 11760 10668 0 _0233_
rlabel metal2 11664 12684 11664 12684 0 _0234_
rlabel metal2 12192 13104 12192 13104 0 _0235_
rlabel metal3 12576 12852 12576 12852 0 _0236_
rlabel metal2 12960 9534 12960 9534 0 _0237_
rlabel metal3 12624 9072 12624 9072 0 _0238_
rlabel metal2 12768 8316 12768 8316 0 _0239_
rlabel metal2 6864 14868 6864 14868 0 _0240_
rlabel metal2 6528 15666 6528 15666 0 _0241_
rlabel metal2 6528 13020 6528 13020 0 _0242_
rlabel metal2 10992 15708 10992 15708 0 _0243_
rlabel metal3 9984 17052 9984 17052 0 _0244_
rlabel metal2 12384 32424 12384 32424 0 _0245_
rlabel metal2 17088 31668 17088 31668 0 _0246_
rlabel metal2 12288 32592 12288 32592 0 _0247_
rlabel metal2 1440 33180 1440 33180 0 _0248_
rlabel metal2 1728 33348 1728 33348 0 _0249_
rlabel metal2 1920 32550 1920 32550 0 _0250_
rlabel metal2 11424 31542 11424 31542 0 _0251_
rlabel metal3 12096 32886 12096 32886 0 _0252_
rlabel metal2 11616 31206 11616 31206 0 _0253_
rlabel metal2 12000 30786 12000 30786 0 _0254_
rlabel metal2 11664 31920 11664 31920 0 _0255_
rlabel metal2 11712 31038 11712 31038 0 _0256_
rlabel metal3 12096 32172 12096 32172 0 _0257_
rlabel metal3 12432 30576 12432 30576 0 _0258_
rlabel metal2 12624 27636 12624 27636 0 _0259_
rlabel metal2 13056 28056 13056 28056 0 _0260_
rlabel metal2 1536 27426 1536 27426 0 _0261_
rlabel metal3 2208 26292 2208 26292 0 _0262_
rlabel metal2 2352 32863 2352 32863 0 _0263_
rlabel metal2 11760 29988 11760 29988 0 _0264_
rlabel metal2 12960 28938 12960 28938 0 _0265_
rlabel metal2 11904 28056 11904 28056 0 _0266_
rlabel metal3 11904 28140 11904 28140 0 _0267_
rlabel metal2 13248 28224 13248 28224 0 _0268_
rlabel metal2 13008 28560 13008 28560 0 _0269_
rlabel metal3 5424 13188 5424 13188 0 _0270_
rlabel metal2 2976 11382 2976 11382 0 _0271_
rlabel metal2 1632 7056 1632 7056 0 _0272_
rlabel metal2 1776 5796 1776 5796 0 _0273_
rlabel metal2 5184 7980 5184 7980 0 _0274_
rlabel metal2 2016 15750 2016 15750 0 _0275_
rlabel metal2 1344 14658 1344 14658 0 _0276_
rlabel metal2 1920 16884 1920 16884 0 _0277_
rlabel metal2 1632 15582 1632 15582 0 _0278_
rlabel metal3 1104 15708 1104 15708 0 _0279_
rlabel metal2 1440 15414 1440 15414 0 _0280_
rlabel metal2 1536 7224 1536 7224 0 _0281_
rlabel metal2 2256 6468 2256 6468 0 _0282_
rlabel metal3 2208 6636 2208 6636 0 _0283_
rlabel metal2 2160 12348 2160 12348 0 _0284_
rlabel metal2 1920 7350 1920 7350 0 _0285_
rlabel metal2 2016 7266 2016 7266 0 _0286_
rlabel metal3 2112 12180 2112 12180 0 _0287_
rlabel metal2 6240 15288 6240 15288 0 _0288_
rlabel metal2 5616 28140 5616 28140 0 _0289_
rlabel metal2 6048 29694 6048 29694 0 _0290_
rlabel metal3 8160 31332 8160 31332 0 _0291_
rlabel metal2 8256 32004 8256 32004 0 _0292_
rlabel metal2 1632 27090 1632 27090 0 _0293_
rlabel metal2 4320 27048 4320 27048 0 _0294_
rlabel metal2 5472 32424 5472 32424 0 _0295_
rlabel metal2 5520 35364 5520 35364 0 _0296_
rlabel metal2 9600 29862 9600 29862 0 _0297_
rlabel metal2 9792 30366 9792 30366 0 _0298_
rlabel metal2 8256 29400 8256 29400 0 _0299_
rlabel metal2 8160 29190 8160 29190 0 _0300_
rlabel metal2 8592 26796 8592 26796 0 _0301_
rlabel metal2 9216 30240 9216 30240 0 _0302_
rlabel metal3 9456 27048 9456 27048 0 _0303_
rlabel metal2 9696 29778 9696 29778 0 _0304_
rlabel metal2 9264 29988 9264 29988 0 _0305_
rlabel metal2 9312 30156 9312 30156 0 _0306_
rlabel metal2 10368 14784 10368 14784 0 _0307_
rlabel metal2 10464 14658 10464 14658 0 _0308_
rlabel metal2 10320 13188 10320 13188 0 _0309_
rlabel metal2 10896 12684 10896 12684 0 _0310_
rlabel metal2 11040 14490 11040 14490 0 _0311_
rlabel metal2 10464 13314 10464 13314 0 _0312_
rlabel metal2 9936 12348 9936 12348 0 _0313_
rlabel metal2 9984 14742 9984 14742 0 _0314_
rlabel metal3 11760 14028 11760 14028 0 _0315_
rlabel metal2 10752 14448 10752 14448 0 _0316_
rlabel metal3 3696 15624 3696 15624 0 _0317_
rlabel metal3 3696 15540 3696 15540 0 _0318_
rlabel metal3 4752 18648 4752 18648 0 _0319_
rlabel metal2 4896 18564 4896 18564 0 _0320_
rlabel metal3 4560 20664 4560 20664 0 _0321_
rlabel metal2 4896 21630 4896 21630 0 _0322_
rlabel metal2 7968 17346 7968 17346 0 _0323_
rlabel metal3 8256 17640 8256 17640 0 _0324_
rlabel metal3 16656 2016 16656 2016 0 _0325_
rlabel metal2 18432 3360 18432 3360 0 _0326_
rlabel metal2 17280 2856 17280 2856 0 _0327_
rlabel metal2 13824 4326 13824 4326 0 _0328_
rlabel metal3 16128 3444 16128 3444 0 _0329_
rlabel metal3 15648 2184 15648 2184 0 _0330_
rlabel metal3 15552 3024 15552 3024 0 _0331_
rlabel metal3 13296 1092 13296 1092 0 _0332_
rlabel metal3 17040 1092 17040 1092 0 _0333_
rlabel metal2 13248 1050 13248 1050 0 _0334_
rlabel metal2 14880 38430 14880 38430 0 _0335_
rlabel metal2 16224 38976 16224 38976 0 _0336_
rlabel metal3 16224 39060 16224 39060 0 _0337_
rlabel metal2 16800 38808 16800 38808 0 _0338_
rlabel metal2 16560 37212 16560 37212 0 _0339_
rlabel metal2 16320 39102 16320 39102 0 _0340_
rlabel metal3 14880 37632 14880 37632 0 _0341_
rlabel metal2 15696 39732 15696 39732 0 _0342_
rlabel metal2 17568 40152 17568 40152 0 _0343_
rlabel metal2 15552 39984 15552 39984 0 _0344_
rlabel metal2 17280 14763 17280 14763 0 _0345_
rlabel metal2 17424 14700 17424 14700 0 _0346_
rlabel metal2 14976 9030 14976 9030 0 _0347_
rlabel metal2 14880 8064 14880 8064 0 _0348_
rlabel metal2 19680 9408 19680 9408 0 _0349_
rlabel metal3 18288 9996 18288 9996 0 _0350_
rlabel metal3 19296 10248 19296 10248 0 _0351_
rlabel metal2 19968 9744 19968 9744 0 _0352_
rlabel metal3 19632 9324 19632 9324 0 _0353_
rlabel metal2 20256 8064 20256 8064 0 _0354_
rlabel metal2 18240 9996 18240 9996 0 _0355_
rlabel metal3 14016 39732 14016 39732 0 _0356_
rlabel metal2 14496 38682 14496 38682 0 _0357_
rlabel metal2 14592 39144 14592 39144 0 _0358_
rlabel metal3 15744 39732 15744 39732 0 _0359_
rlabel metal3 14880 39480 14880 39480 0 _0360_
rlabel metal2 14976 38934 14976 38934 0 _0361_
rlabel metal2 5088 41328 5088 41328 0 _0362_
rlabel metal2 17376 40908 17376 40908 0 _0363_
rlabel metal4 7488 41076 7488 41076 0 _0364_
rlabel metal2 14976 34398 14976 34398 0 _0365_
rlabel metal2 13152 32382 13152 32382 0 _0366_
rlabel metal3 9936 35868 9936 35868 0 _0367_
rlabel metal2 14592 34818 14592 34818 0 _0368_
rlabel metal2 14688 35994 14688 35994 0 _0369_
rlabel metal3 13440 37380 13440 37380 0 _0370_
rlabel metal3 13296 37632 13296 37632 0 _0371_
rlabel metal2 8160 12432 8160 12432 0 _0372_
rlabel metal3 7968 7140 7968 7140 0 _0373_
rlabel metal2 7968 7854 7968 7854 0 _0374_
rlabel metal2 7824 12516 7824 12516 0 _0375_
rlabel metal2 8016 10332 8016 10332 0 _0376_
rlabel metal2 4032 7182 4032 7182 0 _0377_
rlabel metal2 7296 5544 7296 5544 0 _0378_
rlabel metal3 1536 23604 1536 23604 0 _0379_
rlabel metal2 2016 23520 2016 23520 0 _0380_
rlabel metal2 11424 33642 11424 33642 0 clknet_0_UserCLK
rlabel metal3 8352 30408 8352 30408 0 clknet_1_0__leaf_UserCLK
rlabel metal2 12480 36498 12480 36498 0 clknet_1_1__leaf_UserCLK
<< properties >>
string FIXED_BBOX 0 0 21504 43008
<< end >>
