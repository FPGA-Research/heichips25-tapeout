magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753465916
<< metal2 >>
rect 24536 366408 24616 366504
rect 25688 366408 25768 366504
rect 26840 366408 26920 366504
rect 27992 366408 28072 366504
rect 29144 366408 29224 366504
rect 30296 366408 30376 366504
rect 31448 366408 31528 366504
rect 32600 366408 32680 366504
rect 33752 366408 33832 366504
rect 34904 366408 34984 366504
rect 36056 366408 36136 366504
rect 37208 366408 37288 366504
rect 67544 366408 67624 366504
rect 68696 366408 68776 366504
rect 69848 366408 69928 366504
rect 71000 366408 71080 366504
rect 72152 366408 72232 366504
rect 73304 366408 73384 366504
rect 74456 366408 74536 366504
rect 75608 366408 75688 366504
rect 76760 366408 76840 366504
rect 77912 366408 77992 366504
rect 79064 366408 79144 366504
rect 80216 366408 80296 366504
rect 110552 366408 110632 366504
rect 111704 366408 111784 366504
rect 112856 366408 112936 366504
rect 114008 366408 114088 366504
rect 115160 366408 115240 366504
rect 116312 366408 116392 366504
rect 117464 366408 117544 366504
rect 118616 366408 118696 366504
rect 119768 366408 119848 366504
rect 120920 366408 121000 366504
rect 122072 366408 122152 366504
rect 123224 366408 123304 366504
rect 153560 366408 153640 366504
rect 154712 366408 154792 366504
rect 155864 366408 155944 366504
rect 157016 366408 157096 366504
rect 158168 366408 158248 366504
rect 159320 366408 159400 366504
rect 160472 366408 160552 366504
rect 161624 366408 161704 366504
rect 162776 366408 162856 366504
rect 163928 366408 164008 366504
rect 165080 366408 165160 366504
rect 166232 366408 166312 366504
rect 24556 366387 24596 366408
rect 25708 366387 25748 366408
rect 26860 366387 26900 366408
rect 28012 366387 28052 366408
rect 29164 366387 29204 366408
rect 30316 366387 30356 366408
rect 31468 366387 31508 366408
rect 32620 366387 32660 366408
rect 33772 366387 33812 366408
rect 34924 366387 34964 366408
rect 36076 366387 36116 366408
rect 37228 366387 37268 366408
rect 67564 366387 67604 366408
rect 68716 366387 68756 366408
rect 69868 366387 69908 366408
rect 71020 366387 71060 366408
rect 72172 366387 72212 366408
rect 73324 366387 73364 366408
rect 74476 366387 74516 366408
rect 75628 366387 75668 366408
rect 76780 366387 76820 366408
rect 77932 366387 77972 366408
rect 79084 366387 79124 366408
rect 80236 366387 80276 366408
rect 110572 366387 110612 366408
rect 111724 366387 111764 366408
rect 112876 366387 112916 366408
rect 114028 366387 114068 366408
rect 115180 366387 115220 366408
rect 116332 366387 116372 366408
rect 117484 366387 117524 366408
rect 118636 366387 118676 366408
rect 119788 366387 119828 366408
rect 120940 366387 120980 366408
rect 122092 366387 122132 366408
rect 123244 366387 123284 366408
rect 153580 366387 153620 366408
rect 154732 366387 154772 366408
rect 155884 366387 155924 366408
rect 157036 366387 157076 366408
rect 158188 366387 158228 366408
rect 159340 366387 159380 366408
rect 160492 366387 160532 366408
rect 161644 366387 161684 366408
rect 162796 366387 162836 366408
rect 163948 366387 163988 366408
rect 165100 366387 165140 366408
rect 166252 366387 166292 366408
rect 1132 197 1172 861
rect 1131 188 1173 197
rect 1131 148 1132 188
rect 1172 148 1173 188
rect 1131 139 1173 148
rect 1132 96 1172 139
rect 2092 96 2132 861
rect 3052 96 3092 861
rect 4012 96 4052 861
rect 4972 96 5012 861
rect 5932 96 5972 861
rect 6892 96 6932 861
rect 7852 96 7892 861
rect 8812 96 8852 861
rect 9772 96 9812 861
rect 10732 96 10772 861
rect 11692 96 11732 861
rect 12652 96 12692 861
rect 13612 96 13652 861
rect 14572 96 14612 861
rect 15532 96 15572 861
rect 16492 96 16532 861
rect 17452 96 17492 861
rect 18412 96 18452 861
rect 19372 96 19412 861
rect 20332 96 20372 861
rect 24556 96 24596 861
rect 25708 96 25748 861
rect 26860 96 26900 861
rect 28012 96 28052 861
rect 29164 96 29204 861
rect 30316 96 30356 861
rect 31468 96 31508 861
rect 32620 96 32660 861
rect 33772 96 33812 861
rect 34924 96 34964 861
rect 36076 96 36116 861
rect 37228 96 37268 861
rect 38399 785 38439 861
rect 38398 776 38440 785
rect 38380 736 38399 776
rect 38439 736 38440 776
rect 38380 727 38440 736
rect 38380 113 38420 727
rect 38379 104 38421 113
rect 1112 0 1192 96
rect 2072 0 2152 96
rect 3032 0 3112 96
rect 3992 0 4072 96
rect 4952 0 5032 96
rect 5912 0 5992 96
rect 6872 0 6952 96
rect 7832 0 7912 96
rect 8792 0 8872 96
rect 9752 0 9832 96
rect 10712 0 10792 96
rect 11672 0 11752 96
rect 12632 0 12712 96
rect 13592 0 13672 96
rect 14552 0 14632 96
rect 15512 0 15592 96
rect 16472 0 16552 96
rect 17432 0 17512 96
rect 18392 0 18472 96
rect 19352 0 19432 96
rect 20312 0 20392 96
rect 24536 0 24616 96
rect 25688 0 25768 96
rect 26840 0 26920 96
rect 27992 0 28072 96
rect 29144 0 29224 96
rect 30296 0 30376 96
rect 31448 0 31528 96
rect 32600 0 32680 96
rect 33752 0 33832 96
rect 34904 0 34984 96
rect 36056 0 36136 96
rect 37208 0 37288 96
rect 38379 64 38380 104
rect 38420 64 38421 104
rect 39532 96 39572 861
rect 40684 96 40724 861
rect 41836 96 41876 861
rect 42988 96 43028 861
rect 44140 96 44180 861
rect 45292 96 45332 861
rect 46444 96 46484 861
rect 47596 96 47636 861
rect 48748 96 48788 861
rect 49900 96 49940 861
rect 51052 96 51092 861
rect 52204 96 52244 861
rect 53356 96 53396 861
rect 54508 96 54548 861
rect 55660 96 55700 861
rect 56812 96 56852 861
rect 57964 96 58004 861
rect 59116 96 59156 861
rect 60268 96 60308 861
rect 61420 96 61460 861
rect 67564 96 67604 861
rect 68716 96 68756 861
rect 69868 96 69908 861
rect 71020 96 71060 861
rect 72172 96 72212 861
rect 73324 96 73364 861
rect 74476 96 74516 861
rect 75628 96 75668 861
rect 76780 96 76820 861
rect 77932 96 77972 861
rect 79084 96 79124 861
rect 80236 96 80276 861
rect 81407 785 81447 861
rect 81406 776 81448 785
rect 81406 736 81407 776
rect 81447 736 81448 776
rect 81406 727 81448 736
rect 82540 96 82580 861
rect 83692 96 83732 861
rect 84844 96 84884 861
rect 85996 96 86036 861
rect 87148 96 87188 861
rect 88300 96 88340 861
rect 89452 96 89492 861
rect 90604 96 90644 861
rect 91756 96 91796 861
rect 92908 96 92948 861
rect 94060 96 94100 861
rect 95212 96 95252 861
rect 96364 96 96404 861
rect 97516 96 97556 861
rect 98668 96 98708 861
rect 99820 96 99860 861
rect 100972 96 101012 861
rect 102124 96 102164 861
rect 103276 96 103316 861
rect 104428 96 104468 861
rect 110572 96 110612 861
rect 111724 96 111764 861
rect 112876 96 112916 861
rect 114028 96 114068 861
rect 115180 96 115220 861
rect 116332 96 116372 861
rect 117484 96 117524 861
rect 118636 96 118676 861
rect 119788 96 119828 861
rect 120940 96 120980 861
rect 122092 96 122132 861
rect 123244 96 123284 861
rect 124415 785 124455 861
rect 124414 776 124456 785
rect 124414 736 124415 776
rect 124455 736 124456 776
rect 124414 727 124456 736
rect 125548 96 125588 861
rect 126700 96 126740 861
rect 127852 96 127892 861
rect 129004 96 129044 861
rect 130156 96 130196 861
rect 131308 96 131348 861
rect 132460 96 132500 861
rect 133612 96 133652 861
rect 134764 96 134804 861
rect 135916 96 135956 861
rect 137068 96 137108 861
rect 138220 96 138260 861
rect 139372 96 139412 861
rect 140524 96 140564 861
rect 141676 96 141716 861
rect 142828 96 142868 861
rect 143980 96 144020 861
rect 145132 96 145172 861
rect 146284 96 146324 861
rect 147436 96 147476 861
rect 153580 96 153620 861
rect 154732 96 154772 861
rect 155884 96 155924 861
rect 157036 96 157076 861
rect 158188 96 158228 861
rect 159340 96 159380 861
rect 160492 96 160532 861
rect 161644 96 161684 861
rect 162796 96 162836 861
rect 163948 96 163988 861
rect 165100 96 165140 861
rect 166252 96 166292 861
rect 167385 785 167425 861
rect 167384 776 167426 785
rect 167384 736 167385 776
rect 167425 736 167426 776
rect 167384 727 167426 736
rect 168556 96 168596 861
rect 169708 96 169748 861
rect 170860 96 170900 861
rect 172012 96 172052 861
rect 173164 96 173204 861
rect 174316 96 174356 861
rect 175468 96 175508 861
rect 176620 96 176660 861
rect 177772 96 177812 861
rect 178924 96 178964 861
rect 180076 96 180116 861
rect 181228 96 181268 861
rect 182380 96 182420 861
rect 183532 96 183572 861
rect 184684 96 184724 861
rect 185836 96 185876 861
rect 186988 96 187028 861
rect 188140 96 188180 861
rect 189292 96 189332 861
rect 190444 96 190484 861
rect 194649 785 194689 861
rect 194648 776 194690 785
rect 194648 736 194649 776
rect 194689 736 194690 776
rect 194648 727 194690 736
rect 195628 96 195668 861
rect 196588 96 196628 861
rect 197548 96 197588 861
rect 198508 96 198548 861
rect 199468 96 199508 861
rect 200428 96 200468 861
rect 201388 96 201428 861
rect 202348 96 202388 861
rect 203308 96 203348 861
rect 204268 96 204308 861
rect 205228 96 205268 861
rect 206188 96 206228 861
rect 207148 96 207188 861
rect 208108 96 208148 861
rect 209068 96 209108 861
rect 210028 96 210068 861
rect 210988 96 211028 861
rect 211948 96 211988 861
rect 212908 96 212948 861
rect 213868 96 213908 861
rect 38379 55 38421 64
rect 39512 0 39592 96
rect 40664 0 40744 96
rect 41816 0 41896 96
rect 42968 0 43048 96
rect 44120 0 44200 96
rect 45272 0 45352 96
rect 46424 0 46504 96
rect 47576 0 47656 96
rect 48728 0 48808 96
rect 49880 0 49960 96
rect 51032 0 51112 96
rect 52184 0 52264 96
rect 53336 0 53416 96
rect 54488 0 54568 96
rect 55640 0 55720 96
rect 56792 0 56872 96
rect 57944 0 58024 96
rect 59096 0 59176 96
rect 60248 0 60328 96
rect 61400 0 61480 96
rect 67544 0 67624 96
rect 68696 0 68776 96
rect 69848 0 69928 96
rect 71000 0 71080 96
rect 72152 0 72232 96
rect 73304 0 73384 96
rect 74456 0 74536 96
rect 75608 0 75688 96
rect 76760 0 76840 96
rect 77912 0 77992 96
rect 79064 0 79144 96
rect 80216 0 80296 96
rect 82520 0 82600 96
rect 83672 0 83752 96
rect 84824 0 84904 96
rect 85976 0 86056 96
rect 87128 0 87208 96
rect 88280 0 88360 96
rect 89432 0 89512 96
rect 90584 0 90664 96
rect 91736 0 91816 96
rect 92888 0 92968 96
rect 94040 0 94120 96
rect 95192 0 95272 96
rect 96344 0 96424 96
rect 97496 0 97576 96
rect 98648 0 98728 96
rect 99800 0 99880 96
rect 100952 0 101032 96
rect 102104 0 102184 96
rect 103256 0 103336 96
rect 104408 0 104488 96
rect 110552 0 110632 96
rect 111704 0 111784 96
rect 112856 0 112936 96
rect 114008 0 114088 96
rect 115160 0 115240 96
rect 116312 0 116392 96
rect 117464 0 117544 96
rect 118616 0 118696 96
rect 119768 0 119848 96
rect 120920 0 121000 96
rect 122072 0 122152 96
rect 123224 0 123304 96
rect 125528 0 125608 96
rect 126680 0 126760 96
rect 127832 0 127912 96
rect 128984 0 129064 96
rect 130136 0 130216 96
rect 131288 0 131368 96
rect 132440 0 132520 96
rect 133592 0 133672 96
rect 134744 0 134824 96
rect 135896 0 135976 96
rect 137048 0 137128 96
rect 138200 0 138280 96
rect 139352 0 139432 96
rect 140504 0 140584 96
rect 141656 0 141736 96
rect 142808 0 142888 96
rect 143960 0 144040 96
rect 145112 0 145192 96
rect 146264 0 146344 96
rect 147416 0 147496 96
rect 153560 0 153640 96
rect 154712 0 154792 96
rect 155864 0 155944 96
rect 157016 0 157096 96
rect 158168 0 158248 96
rect 159320 0 159400 96
rect 160472 0 160552 96
rect 161624 0 161704 96
rect 162776 0 162856 96
rect 163928 0 164008 96
rect 165080 0 165160 96
rect 166232 0 166312 96
rect 168536 0 168616 96
rect 169688 0 169768 96
rect 170840 0 170920 96
rect 171992 0 172072 96
rect 173144 0 173224 96
rect 174296 0 174376 96
rect 175448 0 175528 96
rect 176600 0 176680 96
rect 177752 0 177832 96
rect 178904 0 178984 96
rect 180056 0 180136 96
rect 181208 0 181288 96
rect 182360 0 182440 96
rect 183512 0 183592 96
rect 184664 0 184744 96
rect 185816 0 185896 96
rect 186968 0 187048 96
rect 188120 0 188200 96
rect 189272 0 189352 96
rect 190424 0 190504 96
rect 195608 0 195688 96
rect 196568 0 196648 96
rect 197528 0 197608 96
rect 198488 0 198568 96
rect 199448 0 199528 96
rect 200408 0 200488 96
rect 201368 0 201448 96
rect 202328 0 202408 96
rect 203288 0 203368 96
rect 204248 0 204328 96
rect 205208 0 205288 96
rect 206168 0 206248 96
rect 207128 0 207208 96
rect 208088 0 208168 96
rect 209048 0 209128 96
rect 210008 0 210088 96
rect 210968 0 211048 96
rect 211928 0 212008 96
rect 212888 0 212968 96
rect 213848 0 213928 96
<< via2 >>
rect 1132 148 1172 188
rect 38399 736 38439 776
rect 38380 64 38420 104
rect 81407 736 81447 776
rect 124415 736 124455 776
rect 167385 736 167425 776
rect 194649 736 194689 776
<< metal3 >>
rect 0 366176 96 366196
rect 0 366136 117 366176
rect 0 366116 96 366136
rect 0 365840 96 365860
rect 0 365800 117 365840
rect 0 365780 96 365800
rect 0 365504 96 365524
rect 0 365464 117 365504
rect 0 365444 96 365464
rect 0 365168 96 365188
rect 0 365128 117 365168
rect 0 365108 96 365128
rect 0 364832 96 364852
rect 0 364792 117 364832
rect 0 364772 96 364792
rect 0 364496 96 364516
rect 0 364456 117 364496
rect 0 364436 96 364456
rect 0 364160 96 364180
rect 0 364120 117 364160
rect 0 364100 96 364120
rect 0 363824 96 363844
rect 0 363784 117 363824
rect 0 363764 96 363784
rect 0 363488 96 363508
rect 0 363448 117 363488
rect 0 363428 96 363448
rect 0 363152 96 363172
rect 0 363112 117 363152
rect 0 363092 96 363112
rect 0 362816 96 362836
rect 0 362776 117 362816
rect 0 362756 96 362776
rect 0 362480 96 362500
rect 0 362440 117 362480
rect 0 362420 96 362440
rect 0 362144 96 362164
rect 0 362104 117 362144
rect 0 362084 96 362104
rect 0 361808 96 361828
rect 0 361768 117 361808
rect 0 361748 96 361768
rect 0 361472 96 361492
rect 0 361432 117 361472
rect 0 361412 96 361432
rect 0 361136 96 361156
rect 0 361096 117 361136
rect 0 361076 96 361096
rect 0 360800 96 360820
rect 0 360760 117 360800
rect 0 360740 96 360760
rect 0 360464 96 360484
rect 0 360424 117 360464
rect 0 360404 96 360424
rect 0 360128 96 360148
rect 0 360088 117 360128
rect 0 360068 96 360088
rect 0 359792 96 359812
rect 0 359752 117 359792
rect 0 359732 96 359752
rect 0 359456 96 359476
rect 0 359416 117 359456
rect 0 359396 96 359416
rect 0 359120 96 359140
rect 0 359080 117 359120
rect 0 359060 96 359080
rect 0 358784 96 358804
rect 0 358744 117 358784
rect 0 358724 96 358744
rect 0 358448 96 358468
rect 0 358408 117 358448
rect 0 358388 96 358408
rect 0 358112 96 358132
rect 0 358072 117 358112
rect 0 358052 96 358072
rect 0 357776 96 357796
rect 0 357736 117 357776
rect 0 357716 96 357736
rect 0 357440 96 357460
rect 0 357400 117 357440
rect 0 357380 96 357400
rect 0 357104 96 357124
rect 0 357064 117 357104
rect 0 357044 96 357064
rect 0 356768 96 356788
rect 0 356728 117 356768
rect 0 356708 96 356728
rect 0 356432 96 356452
rect 0 356392 117 356432
rect 0 356372 96 356392
rect 0 356096 96 356116
rect 0 356056 117 356096
rect 0 356036 96 356056
rect 0 355760 96 355780
rect 0 355720 117 355760
rect 0 355700 96 355720
rect 0 352736 96 352756
rect 0 352696 117 352736
rect 0 352676 96 352696
rect 0 352232 96 352252
rect 0 352192 117 352232
rect 0 352172 96 352192
rect 0 351728 96 351748
rect 0 351688 117 351728
rect 0 351668 96 351688
rect 0 351224 96 351244
rect 0 351184 117 351224
rect 0 351164 96 351184
rect 0 350720 96 350740
rect 0 350680 117 350720
rect 0 350660 96 350680
rect 0 350216 96 350236
rect 0 350176 117 350216
rect 0 350156 96 350176
rect 0 349712 96 349732
rect 0 349672 117 349712
rect 0 349652 96 349672
rect 0 349208 96 349228
rect 0 349168 117 349208
rect 0 349148 96 349168
rect 0 348704 96 348724
rect 0 348664 117 348704
rect 0 348644 96 348664
rect 0 348200 96 348220
rect 0 348160 117 348200
rect 0 348140 96 348160
rect 0 347696 96 347716
rect 0 347656 117 347696
rect 0 347636 96 347656
rect 0 347192 96 347212
rect 0 347152 117 347192
rect 0 347132 96 347152
rect 0 346688 96 346708
rect 0 346648 117 346688
rect 0 346628 96 346648
rect 0 346184 96 346204
rect 0 346144 117 346184
rect 0 346124 96 346144
rect 0 345680 96 345700
rect 0 345640 117 345680
rect 0 345620 96 345640
rect 0 345176 96 345196
rect 0 345136 117 345176
rect 0 345116 96 345136
rect 0 344672 96 344692
rect 0 344632 117 344672
rect 0 344612 96 344632
rect 0 344168 96 344188
rect 0 344128 117 344168
rect 0 344108 96 344128
rect 0 343664 96 343684
rect 0 343624 117 343664
rect 0 343604 96 343624
rect 0 343160 96 343180
rect 0 343120 117 343160
rect 0 343100 96 343120
rect 0 342656 96 342676
rect 0 342616 117 342656
rect 0 342596 96 342616
rect 0 342152 96 342172
rect 0 342112 117 342152
rect 0 342092 96 342112
rect 0 341648 96 341668
rect 0 341608 117 341648
rect 0 341588 96 341608
rect 0 341144 96 341164
rect 0 341104 117 341144
rect 0 341084 96 341104
rect 0 340640 96 340660
rect 0 340600 117 340640
rect 0 340580 96 340600
rect 0 340136 96 340156
rect 0 340096 117 340136
rect 0 340076 96 340096
rect 0 339632 96 339652
rect 0 339592 117 339632
rect 0 339572 96 339592
rect 0 339128 96 339148
rect 0 339088 117 339128
rect 0 339068 96 339088
rect 0 338624 96 338644
rect 0 338584 117 338624
rect 0 338564 96 338584
rect 0 338120 96 338140
rect 0 338080 117 338120
rect 0 338060 96 338080
rect 0 337616 96 337636
rect 0 337576 117 337616
rect 0 337556 96 337576
rect 0 337112 96 337132
rect 0 337072 117 337112
rect 0 337052 96 337072
rect 0 336608 96 336628
rect 0 336568 117 336608
rect 0 336548 96 336568
rect 0 336104 96 336124
rect 0 336064 117 336104
rect 0 336044 96 336064
rect 0 335600 96 335620
rect 0 335560 117 335600
rect 0 335540 96 335560
rect 0 335096 96 335116
rect 0 335056 117 335096
rect 0 335036 96 335056
rect 0 334592 96 334612
rect 0 334552 117 334592
rect 0 334532 96 334552
rect 0 334088 96 334108
rect 0 334048 117 334088
rect 0 334028 96 334048
rect 0 333584 96 333604
rect 0 333544 117 333584
rect 0 333524 96 333544
rect 0 333080 96 333100
rect 0 333040 117 333080
rect 0 333020 96 333040
rect 0 332576 96 332596
rect 0 332536 117 332576
rect 0 332516 96 332536
rect 0 332072 96 332092
rect 0 332032 117 332072
rect 0 332012 96 332032
rect 0 331568 96 331588
rect 0 331528 117 331568
rect 0 331508 96 331528
rect 0 331064 96 331084
rect 0 331024 117 331064
rect 0 331004 96 331024
rect 0 330560 96 330580
rect 0 330520 117 330560
rect 0 330500 96 330520
rect 0 330056 96 330076
rect 0 330016 117 330056
rect 0 329996 96 330016
rect 0 329552 96 329572
rect 0 329512 117 329552
rect 0 329492 96 329512
rect 0 329048 96 329068
rect 0 329008 117 329048
rect 0 328988 96 329008
rect 0 328544 96 328564
rect 0 328504 117 328544
rect 0 328484 96 328504
rect 0 328040 96 328060
rect 0 328000 117 328040
rect 0 327980 96 328000
rect 0 327536 96 327556
rect 0 327496 117 327536
rect 0 327476 96 327496
rect 0 327032 96 327052
rect 0 326992 117 327032
rect 0 326972 96 326992
rect 0 326528 96 326548
rect 0 326488 117 326528
rect 0 326468 96 326488
rect 0 326024 96 326044
rect 0 325984 117 326024
rect 0 325964 96 325984
rect 0 325520 96 325540
rect 0 325480 117 325520
rect 0 325460 96 325480
rect 0 325016 96 325036
rect 0 324976 117 325016
rect 0 324956 96 324976
rect 0 324512 96 324532
rect 0 324472 117 324512
rect 0 324452 96 324472
rect 0 324008 96 324028
rect 0 323968 117 324008
rect 0 323948 96 323968
rect 0 323504 96 323524
rect 0 323464 117 323504
rect 0 323444 96 323464
rect 0 323000 96 323020
rect 0 322960 117 323000
rect 0 322940 96 322960
rect 0 322496 96 322516
rect 0 322456 117 322496
rect 0 322436 96 322456
rect 0 321992 96 322012
rect 0 321952 117 321992
rect 0 321932 96 321952
rect 0 321488 96 321508
rect 0 321448 117 321488
rect 0 321428 96 321448
rect 0 320984 96 321004
rect 0 320944 117 320984
rect 0 320924 96 320944
rect 215136 320648 215232 320668
rect 215115 320608 215232 320648
rect 215136 320588 215232 320608
rect 0 320480 96 320500
rect 0 320440 117 320480
rect 0 320420 96 320440
rect 215136 320312 215232 320332
rect 215115 320272 215232 320312
rect 215136 320252 215232 320272
rect 0 319976 96 319996
rect 215136 319976 215232 319996
rect 0 319936 117 319976
rect 215115 319936 215232 319976
rect 0 319916 96 319936
rect 215136 319916 215232 319936
rect 215136 319640 215232 319660
rect 215115 319600 215232 319640
rect 215136 319580 215232 319600
rect 0 319472 96 319492
rect 0 319432 117 319472
rect 0 319412 96 319432
rect 215136 319304 215232 319324
rect 215115 319264 215232 319304
rect 215136 319244 215232 319264
rect 0 318968 96 318988
rect 215136 318968 215232 318988
rect 0 318928 117 318968
rect 215115 318928 215232 318968
rect 0 318908 96 318928
rect 215136 318908 215232 318928
rect 215136 318632 215232 318652
rect 215115 318592 215232 318632
rect 215136 318572 215232 318592
rect 0 318464 96 318484
rect 0 318424 117 318464
rect 0 318404 96 318424
rect 215136 318296 215232 318316
rect 215115 318256 215232 318296
rect 215136 318236 215232 318256
rect 0 317960 96 317980
rect 215136 317960 215232 317980
rect 0 317920 117 317960
rect 215115 317920 215232 317960
rect 0 317900 96 317920
rect 215136 317900 215232 317920
rect 215136 317624 215232 317644
rect 215115 317584 215232 317624
rect 215136 317564 215232 317584
rect 0 317456 96 317476
rect 0 317416 117 317456
rect 0 317396 96 317416
rect 215136 317288 215232 317308
rect 215115 317248 215232 317288
rect 215136 317228 215232 317248
rect 0 316952 96 316972
rect 215136 316952 215232 316972
rect 0 316912 117 316952
rect 215115 316912 215232 316952
rect 0 316892 96 316912
rect 215136 316892 215232 316912
rect 215136 316616 215232 316636
rect 215115 316576 215232 316616
rect 215136 316556 215232 316576
rect 0 316448 96 316468
rect 0 316408 117 316448
rect 0 316388 96 316408
rect 215136 316280 215232 316300
rect 215115 316240 215232 316280
rect 215136 316220 215232 316240
rect 0 315944 96 315964
rect 215136 315944 215232 315964
rect 0 315904 117 315944
rect 215115 315904 215232 315944
rect 0 315884 96 315904
rect 215136 315884 215232 315904
rect 215136 315608 215232 315628
rect 215115 315568 215232 315608
rect 215136 315548 215232 315568
rect 0 315440 96 315460
rect 0 315400 117 315440
rect 0 315380 96 315400
rect 215136 315272 215232 315292
rect 215115 315232 215232 315272
rect 215136 315212 215232 315232
rect 215136 314936 215232 314956
rect 215115 314896 215232 314936
rect 215136 314876 215232 314896
rect 215136 314600 215232 314620
rect 215115 314560 215232 314600
rect 215136 314540 215232 314560
rect 215136 314264 215232 314284
rect 215115 314224 215232 314264
rect 215136 314204 215232 314224
rect 215136 313928 215232 313948
rect 215115 313888 215232 313928
rect 215136 313868 215232 313888
rect 215136 313592 215232 313612
rect 215115 313552 215232 313592
rect 215136 313532 215232 313552
rect 215136 313256 215232 313276
rect 215115 313216 215232 313256
rect 215136 313196 215232 313216
rect 215136 312920 215232 312940
rect 215115 312880 215232 312920
rect 215136 312860 215232 312880
rect 215136 312584 215232 312604
rect 215115 312544 215232 312584
rect 215136 312524 215232 312544
rect 215136 312248 215232 312268
rect 215115 312208 215232 312248
rect 215136 312188 215232 312208
rect 215136 311912 215232 311932
rect 215115 311872 215232 311912
rect 215136 311852 215232 311872
rect 215136 311576 215232 311596
rect 215115 311536 215232 311576
rect 215136 311516 215232 311536
rect 215136 311240 215232 311260
rect 215115 311200 215232 311240
rect 215136 311180 215232 311200
rect 215136 310904 215232 310924
rect 215115 310864 215232 310904
rect 215136 310844 215232 310864
rect 215136 310568 215232 310588
rect 215115 310528 215232 310568
rect 215136 310508 215232 310528
rect 215136 310232 215232 310252
rect 215115 310192 215232 310232
rect 215136 310172 215232 310192
rect 215136 309896 215232 309916
rect 215115 309856 215232 309896
rect 215136 309836 215232 309856
rect 0 309728 96 309748
rect 0 309688 117 309728
rect 0 309668 96 309688
rect 215136 309560 215232 309580
rect 215115 309520 215232 309560
rect 215136 309500 215232 309520
rect 0 309224 96 309244
rect 215136 309224 215232 309244
rect 0 309184 117 309224
rect 215115 309184 215232 309224
rect 0 309164 96 309184
rect 215136 309164 215232 309184
rect 215136 308888 215232 308908
rect 215115 308848 215232 308888
rect 215136 308828 215232 308848
rect 0 308720 96 308740
rect 0 308680 117 308720
rect 0 308660 96 308680
rect 215136 308552 215232 308572
rect 215115 308512 215232 308552
rect 215136 308492 215232 308512
rect 0 308216 96 308236
rect 215136 308216 215232 308236
rect 0 308176 117 308216
rect 215115 308176 215232 308216
rect 0 308156 96 308176
rect 215136 308156 215232 308176
rect 215136 307880 215232 307900
rect 215115 307840 215232 307880
rect 215136 307820 215232 307840
rect 0 307712 96 307732
rect 0 307672 117 307712
rect 0 307652 96 307672
rect 215136 307544 215232 307564
rect 215115 307504 215232 307544
rect 215136 307484 215232 307504
rect 0 307208 96 307228
rect 215136 307208 215232 307228
rect 0 307168 117 307208
rect 215115 307168 215232 307208
rect 0 307148 96 307168
rect 215136 307148 215232 307168
rect 215136 306872 215232 306892
rect 215115 306832 215232 306872
rect 215136 306812 215232 306832
rect 0 306704 96 306724
rect 0 306664 117 306704
rect 0 306644 96 306664
rect 215136 306536 215232 306556
rect 215115 306496 215232 306536
rect 215136 306476 215232 306496
rect 0 306200 96 306220
rect 215136 306200 215232 306220
rect 0 306160 117 306200
rect 215115 306160 215232 306200
rect 0 306140 96 306160
rect 215136 306140 215232 306160
rect 215136 305864 215232 305884
rect 215115 305824 215232 305864
rect 215136 305804 215232 305824
rect 0 305696 96 305716
rect 0 305656 117 305696
rect 0 305636 96 305656
rect 215136 305528 215232 305548
rect 215115 305488 215232 305528
rect 215136 305468 215232 305488
rect 0 305192 96 305212
rect 215136 305192 215232 305212
rect 0 305152 117 305192
rect 215115 305152 215232 305192
rect 0 305132 96 305152
rect 215136 305132 215232 305152
rect 215136 304856 215232 304876
rect 215115 304816 215232 304856
rect 215136 304796 215232 304816
rect 0 304688 96 304708
rect 0 304648 117 304688
rect 0 304628 96 304648
rect 215136 304520 215232 304540
rect 215115 304480 215232 304520
rect 215136 304460 215232 304480
rect 0 304184 96 304204
rect 215136 304184 215232 304204
rect 0 304144 117 304184
rect 215115 304144 215232 304184
rect 0 304124 96 304144
rect 215136 304124 215232 304144
rect 215136 303848 215232 303868
rect 215115 303808 215232 303848
rect 215136 303788 215232 303808
rect 0 303680 96 303700
rect 0 303640 117 303680
rect 0 303620 96 303640
rect 215136 303512 215232 303532
rect 215115 303472 215232 303512
rect 215136 303452 215232 303472
rect 0 303176 96 303196
rect 215136 303176 215232 303196
rect 0 303136 117 303176
rect 215115 303136 215232 303176
rect 0 303116 96 303136
rect 215136 303116 215232 303136
rect 215136 302840 215232 302860
rect 215115 302800 215232 302840
rect 215136 302780 215232 302800
rect 0 302672 96 302692
rect 0 302632 117 302672
rect 0 302612 96 302632
rect 215136 302504 215232 302524
rect 215115 302464 215232 302504
rect 215136 302444 215232 302464
rect 0 302168 96 302188
rect 215136 302168 215232 302188
rect 0 302128 117 302168
rect 215115 302128 215232 302168
rect 0 302108 96 302128
rect 215136 302108 215232 302128
rect 215136 301832 215232 301852
rect 215115 301792 215232 301832
rect 215136 301772 215232 301792
rect 0 301664 96 301684
rect 0 301624 117 301664
rect 0 301604 96 301624
rect 215136 301496 215232 301516
rect 215115 301456 215232 301496
rect 215136 301436 215232 301456
rect 0 301160 96 301180
rect 215136 301160 215232 301180
rect 0 301120 117 301160
rect 215115 301120 215232 301160
rect 0 301100 96 301120
rect 215136 301100 215232 301120
rect 215136 300824 215232 300844
rect 215115 300784 215232 300824
rect 215136 300764 215232 300784
rect 0 300656 96 300676
rect 0 300616 117 300656
rect 0 300596 96 300616
rect 215136 300488 215232 300508
rect 215115 300448 215232 300488
rect 215136 300428 215232 300448
rect 0 300152 96 300172
rect 215136 300152 215232 300172
rect 0 300112 117 300152
rect 215115 300112 215232 300152
rect 0 300092 96 300112
rect 215136 300092 215232 300112
rect 215136 299816 215232 299836
rect 215115 299776 215232 299816
rect 215136 299756 215232 299776
rect 0 299648 96 299668
rect 0 299608 117 299648
rect 0 299588 96 299608
rect 215136 299480 215232 299500
rect 215115 299440 215232 299480
rect 215136 299420 215232 299440
rect 0 299144 96 299164
rect 215136 299144 215232 299164
rect 0 299104 117 299144
rect 215115 299104 215232 299144
rect 0 299084 96 299104
rect 215136 299084 215232 299104
rect 215136 298808 215232 298828
rect 215115 298768 215232 298808
rect 215136 298748 215232 298768
rect 0 298640 96 298660
rect 0 298600 117 298640
rect 0 298580 96 298600
rect 215136 298472 215232 298492
rect 215115 298432 215232 298472
rect 215136 298412 215232 298432
rect 0 298136 96 298156
rect 215136 298136 215232 298156
rect 0 298096 117 298136
rect 215115 298096 215232 298136
rect 0 298076 96 298096
rect 215136 298076 215232 298096
rect 215136 297800 215232 297820
rect 215115 297760 215232 297800
rect 215136 297740 215232 297760
rect 0 297632 96 297652
rect 0 297592 117 297632
rect 0 297572 96 297592
rect 215136 297464 215232 297484
rect 215115 297424 215232 297464
rect 215136 297404 215232 297424
rect 0 297128 96 297148
rect 215136 297128 215232 297148
rect 0 297088 117 297128
rect 215115 297088 215232 297128
rect 0 297068 96 297088
rect 215136 297068 215232 297088
rect 215136 296792 215232 296812
rect 215115 296752 215232 296792
rect 215136 296732 215232 296752
rect 0 296624 96 296644
rect 0 296584 117 296624
rect 0 296564 96 296584
rect 215136 296456 215232 296476
rect 215115 296416 215232 296456
rect 215136 296396 215232 296416
rect 0 296120 96 296140
rect 215136 296120 215232 296140
rect 0 296080 117 296120
rect 215115 296080 215232 296120
rect 0 296060 96 296080
rect 215136 296060 215232 296080
rect 215136 295784 215232 295804
rect 215115 295744 215232 295784
rect 215136 295724 215232 295744
rect 0 295616 96 295636
rect 0 295576 117 295616
rect 0 295556 96 295576
rect 215136 295448 215232 295468
rect 215115 295408 215232 295448
rect 215136 295388 215232 295408
rect 0 295112 96 295132
rect 215136 295112 215232 295132
rect 0 295072 117 295112
rect 215115 295072 215232 295112
rect 0 295052 96 295072
rect 215136 295052 215232 295072
rect 215136 294776 215232 294796
rect 215115 294736 215232 294776
rect 215136 294716 215232 294736
rect 0 294608 96 294628
rect 0 294568 117 294608
rect 0 294548 96 294568
rect 215136 294440 215232 294460
rect 215115 294400 215232 294440
rect 215136 294380 215232 294400
rect 0 294104 96 294124
rect 215136 294104 215232 294124
rect 0 294064 117 294104
rect 215115 294064 215232 294104
rect 0 294044 96 294064
rect 215136 294044 215232 294064
rect 215136 293768 215232 293788
rect 215115 293728 215232 293768
rect 215136 293708 215232 293728
rect 0 293600 96 293620
rect 0 293560 117 293600
rect 0 293540 96 293560
rect 215136 293432 215232 293452
rect 215115 293392 215232 293432
rect 215136 293372 215232 293392
rect 0 293096 96 293116
rect 215136 293096 215232 293116
rect 0 293056 117 293096
rect 215115 293056 215232 293096
rect 0 293036 96 293056
rect 215136 293036 215232 293056
rect 215136 292760 215232 292780
rect 215115 292720 215232 292760
rect 215136 292700 215232 292720
rect 0 292592 96 292612
rect 0 292552 117 292592
rect 0 292532 96 292552
rect 215136 292424 215232 292444
rect 215115 292384 215232 292424
rect 215136 292364 215232 292384
rect 0 292088 96 292108
rect 215136 292088 215232 292108
rect 0 292048 117 292088
rect 215115 292048 215232 292088
rect 0 292028 96 292048
rect 215136 292028 215232 292048
rect 215136 291752 215232 291772
rect 215115 291712 215232 291752
rect 215136 291692 215232 291712
rect 0 291584 96 291604
rect 0 291544 117 291584
rect 0 291524 96 291544
rect 215136 291416 215232 291436
rect 215115 291376 215232 291416
rect 215136 291356 215232 291376
rect 0 291080 96 291100
rect 215136 291080 215232 291100
rect 0 291040 117 291080
rect 215115 291040 215232 291080
rect 0 291020 96 291040
rect 215136 291020 215232 291040
rect 215136 290744 215232 290764
rect 215115 290704 215232 290744
rect 215136 290684 215232 290704
rect 0 290576 96 290596
rect 0 290536 117 290576
rect 0 290516 96 290536
rect 215136 290408 215232 290428
rect 215115 290368 215232 290408
rect 215136 290348 215232 290368
rect 0 290072 96 290092
rect 215136 290072 215232 290092
rect 0 290032 117 290072
rect 215115 290032 215232 290072
rect 0 290012 96 290032
rect 215136 290012 215232 290032
rect 215136 289736 215232 289756
rect 215115 289696 215232 289736
rect 215136 289676 215232 289696
rect 0 289568 96 289588
rect 0 289528 117 289568
rect 0 289508 96 289528
rect 215136 289400 215232 289420
rect 215115 289360 215232 289400
rect 215136 289340 215232 289360
rect 0 289064 96 289084
rect 215136 289064 215232 289084
rect 0 289024 117 289064
rect 215115 289024 215232 289064
rect 0 289004 96 289024
rect 215136 289004 215232 289024
rect 215136 288728 215232 288748
rect 215115 288688 215232 288728
rect 215136 288668 215232 288688
rect 0 288560 96 288580
rect 0 288520 117 288560
rect 0 288500 96 288520
rect 215136 288392 215232 288412
rect 215115 288352 215232 288392
rect 215136 288332 215232 288352
rect 0 288056 96 288076
rect 215136 288056 215232 288076
rect 0 288016 117 288056
rect 215115 288016 215232 288056
rect 0 287996 96 288016
rect 215136 287996 215232 288016
rect 215136 287720 215232 287740
rect 215115 287680 215232 287720
rect 215136 287660 215232 287680
rect 0 287552 96 287572
rect 0 287512 117 287552
rect 0 287492 96 287512
rect 215136 287384 215232 287404
rect 215115 287344 215232 287384
rect 215136 287324 215232 287344
rect 0 287048 96 287068
rect 215136 287048 215232 287068
rect 0 287008 117 287048
rect 215115 287008 215232 287048
rect 0 286988 96 287008
rect 215136 286988 215232 287008
rect 215136 286712 215232 286732
rect 215115 286672 215232 286712
rect 215136 286652 215232 286672
rect 0 286544 96 286564
rect 0 286504 117 286544
rect 0 286484 96 286504
rect 215136 286376 215232 286396
rect 215115 286336 215232 286376
rect 215136 286316 215232 286336
rect 0 286040 96 286060
rect 215136 286040 215232 286060
rect 0 286000 117 286040
rect 215115 286000 215232 286040
rect 0 285980 96 286000
rect 215136 285980 215232 286000
rect 215136 285704 215232 285724
rect 215115 285664 215232 285704
rect 215136 285644 215232 285664
rect 0 285536 96 285556
rect 0 285496 117 285536
rect 0 285476 96 285496
rect 215136 285368 215232 285388
rect 215115 285328 215232 285368
rect 215136 285308 215232 285328
rect 0 285032 96 285052
rect 215136 285032 215232 285052
rect 0 284992 117 285032
rect 215115 284992 215232 285032
rect 0 284972 96 284992
rect 215136 284972 215232 284992
rect 215136 284696 215232 284716
rect 215115 284656 215232 284696
rect 215136 284636 215232 284656
rect 0 284528 96 284548
rect 0 284488 117 284528
rect 0 284468 96 284488
rect 215136 284360 215232 284380
rect 215115 284320 215232 284360
rect 215136 284300 215232 284320
rect 0 284024 96 284044
rect 215136 284024 215232 284044
rect 0 283984 117 284024
rect 215115 283984 215232 284024
rect 0 283964 96 283984
rect 215136 283964 215232 283984
rect 215136 283688 215232 283708
rect 215115 283648 215232 283688
rect 215136 283628 215232 283648
rect 0 283520 96 283540
rect 0 283480 117 283520
rect 0 283460 96 283480
rect 215136 283352 215232 283372
rect 215115 283312 215232 283352
rect 215136 283292 215232 283312
rect 0 283016 96 283036
rect 215136 283016 215232 283036
rect 0 282976 117 283016
rect 215115 282976 215232 283016
rect 0 282956 96 282976
rect 215136 282956 215232 282976
rect 0 282512 96 282532
rect 0 282472 117 282512
rect 0 282452 96 282472
rect 0 282008 96 282028
rect 0 281968 117 282008
rect 0 281948 96 281968
rect 0 281504 96 281524
rect 0 281464 117 281504
rect 0 281444 96 281464
rect 0 281000 96 281020
rect 0 280960 117 281000
rect 0 280940 96 280960
rect 0 280496 96 280516
rect 0 280456 117 280496
rect 0 280436 96 280456
rect 0 279992 96 280012
rect 0 279952 117 279992
rect 0 279932 96 279952
rect 0 279488 96 279508
rect 0 279448 117 279488
rect 0 279428 96 279448
rect 0 278984 96 279004
rect 0 278944 117 278984
rect 0 278924 96 278944
rect 0 278480 96 278500
rect 0 278440 117 278480
rect 0 278420 96 278440
rect 0 277976 96 277996
rect 0 277936 117 277976
rect 0 277916 96 277936
rect 0 277472 96 277492
rect 0 277432 117 277472
rect 0 277412 96 277432
rect 0 276968 96 276988
rect 0 276928 117 276968
rect 0 276908 96 276928
rect 0 276464 96 276484
rect 0 276424 117 276464
rect 0 276404 96 276424
rect 0 275960 96 275980
rect 0 275920 117 275960
rect 0 275900 96 275920
rect 0 275456 96 275476
rect 0 275416 117 275456
rect 0 275396 96 275416
rect 0 274952 96 274972
rect 0 274912 117 274952
rect 0 274892 96 274912
rect 0 274448 96 274468
rect 0 274408 117 274448
rect 0 274388 96 274408
rect 0 273944 96 273964
rect 0 273904 117 273944
rect 0 273884 96 273904
rect 0 273440 96 273460
rect 0 273400 117 273440
rect 0 273380 96 273400
rect 0 272936 96 272956
rect 0 272896 117 272936
rect 0 272876 96 272896
rect 0 272432 96 272452
rect 0 272392 117 272432
rect 0 272372 96 272392
rect 0 266720 96 266740
rect 0 266680 117 266720
rect 0 266660 96 266680
rect 0 266216 96 266236
rect 0 266176 117 266216
rect 0 266156 96 266176
rect 0 265712 96 265732
rect 0 265672 117 265712
rect 0 265652 96 265672
rect 0 265208 96 265228
rect 0 265168 117 265208
rect 0 265148 96 265168
rect 0 264704 96 264724
rect 0 264664 117 264704
rect 0 264644 96 264664
rect 0 264200 96 264220
rect 0 264160 117 264200
rect 0 264140 96 264160
rect 0 263696 96 263716
rect 0 263656 117 263696
rect 0 263636 96 263656
rect 0 263192 96 263212
rect 0 263152 117 263192
rect 0 263132 96 263152
rect 0 262688 96 262708
rect 0 262648 117 262688
rect 0 262628 96 262648
rect 0 262184 96 262204
rect 0 262144 117 262184
rect 0 262124 96 262144
rect 0 261680 96 261700
rect 0 261640 117 261680
rect 0 261620 96 261640
rect 0 261176 96 261196
rect 0 261136 117 261176
rect 0 261116 96 261136
rect 0 260672 96 260692
rect 0 260632 117 260672
rect 0 260612 96 260632
rect 0 260168 96 260188
rect 0 260128 117 260168
rect 0 260108 96 260128
rect 0 259664 96 259684
rect 0 259624 117 259664
rect 0 259604 96 259624
rect 0 259160 96 259180
rect 0 259120 117 259160
rect 0 259100 96 259120
rect 0 258656 96 258676
rect 0 258616 117 258656
rect 0 258596 96 258616
rect 0 258152 96 258172
rect 0 258112 117 258152
rect 0 258092 96 258112
rect 0 257648 96 257668
rect 0 257608 117 257648
rect 0 257588 96 257608
rect 0 257144 96 257164
rect 0 257104 117 257144
rect 0 257084 96 257104
rect 0 256640 96 256660
rect 0 256600 117 256640
rect 0 256580 96 256600
rect 0 256136 96 256156
rect 0 256096 117 256136
rect 0 256076 96 256096
rect 0 255632 96 255652
rect 0 255592 117 255632
rect 0 255572 96 255592
rect 0 255128 96 255148
rect 0 255088 117 255128
rect 0 255068 96 255088
rect 0 254624 96 254644
rect 0 254584 117 254624
rect 0 254564 96 254584
rect 0 254120 96 254140
rect 0 254080 117 254120
rect 0 254060 96 254080
rect 0 253616 96 253636
rect 0 253576 117 253616
rect 0 253556 96 253576
rect 0 253112 96 253132
rect 0 253072 117 253112
rect 0 253052 96 253072
rect 0 252608 96 252628
rect 0 252568 117 252608
rect 0 252548 96 252568
rect 0 252104 96 252124
rect 0 252064 117 252104
rect 0 252044 96 252064
rect 0 251600 96 251620
rect 0 251560 117 251600
rect 0 251540 96 251560
rect 0 251096 96 251116
rect 0 251056 117 251096
rect 0 251036 96 251056
rect 0 250592 96 250612
rect 215136 250592 215232 250612
rect 0 250552 117 250592
rect 215115 250552 215232 250592
rect 0 250532 96 250552
rect 215136 250532 215232 250552
rect 0 250088 96 250108
rect 215136 250088 215232 250108
rect 0 250048 117 250088
rect 215115 250048 215232 250088
rect 0 250028 96 250048
rect 215136 250028 215232 250048
rect 0 249584 96 249604
rect 215136 249584 215232 249604
rect 0 249544 117 249584
rect 215115 249544 215232 249584
rect 0 249524 96 249544
rect 215136 249524 215232 249544
rect 0 249080 96 249100
rect 215136 249080 215232 249100
rect 0 249040 117 249080
rect 215115 249040 215232 249080
rect 0 249020 96 249040
rect 215136 249020 215232 249040
rect 0 248576 96 248596
rect 215136 248576 215232 248596
rect 0 248536 117 248576
rect 215115 248536 215232 248576
rect 0 248516 96 248536
rect 215136 248516 215232 248536
rect 0 248072 96 248092
rect 215136 248072 215232 248092
rect 0 248032 117 248072
rect 215115 248032 215232 248072
rect 0 248012 96 248032
rect 215136 248012 215232 248032
rect 0 247568 96 247588
rect 215136 247568 215232 247588
rect 0 247528 117 247568
rect 215115 247528 215232 247568
rect 0 247508 96 247528
rect 215136 247508 215232 247528
rect 0 247064 96 247084
rect 215136 247064 215232 247084
rect 0 247024 117 247064
rect 215115 247024 215232 247064
rect 0 247004 96 247024
rect 215136 247004 215232 247024
rect 0 246560 96 246580
rect 215136 246560 215232 246580
rect 0 246520 117 246560
rect 215115 246520 215232 246560
rect 0 246500 96 246520
rect 215136 246500 215232 246520
rect 0 246056 96 246076
rect 215136 246056 215232 246076
rect 0 246016 117 246056
rect 215115 246016 215232 246056
rect 0 245996 96 246016
rect 215136 245996 215232 246016
rect 0 245552 96 245572
rect 215136 245552 215232 245572
rect 0 245512 117 245552
rect 215115 245512 215232 245552
rect 0 245492 96 245512
rect 215136 245492 215232 245512
rect 0 245048 96 245068
rect 215136 245048 215232 245068
rect 0 245008 117 245048
rect 215115 245008 215232 245048
rect 0 244988 96 245008
rect 215136 244988 215232 245008
rect 0 244544 96 244564
rect 215136 244544 215232 244564
rect 0 244504 117 244544
rect 215115 244504 215232 244544
rect 0 244484 96 244504
rect 215136 244484 215232 244504
rect 0 244040 96 244060
rect 215136 244040 215232 244060
rect 0 244000 117 244040
rect 215115 244000 215232 244040
rect 0 243980 96 244000
rect 215136 243980 215232 244000
rect 0 243536 96 243556
rect 215136 243536 215232 243556
rect 0 243496 117 243536
rect 215115 243496 215232 243536
rect 0 243476 96 243496
rect 215136 243476 215232 243496
rect 0 243032 96 243052
rect 215136 243032 215232 243052
rect 0 242992 117 243032
rect 215115 242992 215232 243032
rect 0 242972 96 242992
rect 215136 242972 215232 242992
rect 0 242528 96 242548
rect 215136 242528 215232 242548
rect 0 242488 117 242528
rect 215115 242488 215232 242528
rect 0 242468 96 242488
rect 215136 242468 215232 242488
rect 0 242024 96 242044
rect 215136 242024 215232 242044
rect 0 241984 117 242024
rect 215115 241984 215232 242024
rect 0 241964 96 241984
rect 215136 241964 215232 241984
rect 0 241520 96 241540
rect 215136 241520 215232 241540
rect 0 241480 117 241520
rect 215115 241480 215232 241520
rect 0 241460 96 241480
rect 215136 241460 215232 241480
rect 0 241016 96 241036
rect 215136 241016 215232 241036
rect 0 240976 117 241016
rect 215115 240976 215232 241016
rect 0 240956 96 240976
rect 215136 240956 215232 240976
rect 0 240512 96 240532
rect 215136 240512 215232 240532
rect 0 240472 117 240512
rect 215115 240472 215232 240512
rect 0 240452 96 240472
rect 215136 240452 215232 240472
rect 0 240008 96 240028
rect 215136 240008 215232 240028
rect 0 239968 117 240008
rect 215115 239968 215232 240008
rect 0 239948 96 239968
rect 215136 239948 215232 239968
rect 0 239504 96 239524
rect 215136 239504 215232 239524
rect 0 239464 117 239504
rect 215115 239464 215232 239504
rect 0 239444 96 239464
rect 215136 239444 215232 239464
rect 0 239000 96 239020
rect 215136 239000 215232 239020
rect 0 238960 117 239000
rect 215115 238960 215232 239000
rect 0 238940 96 238960
rect 215136 238940 215232 238960
rect 0 238496 96 238516
rect 215136 238496 215232 238516
rect 0 238456 117 238496
rect 215115 238456 215232 238496
rect 0 238436 96 238456
rect 215136 238436 215232 238456
rect 0 237992 96 238012
rect 215136 237992 215232 238012
rect 0 237952 117 237992
rect 215115 237952 215232 237992
rect 0 237932 96 237952
rect 215136 237932 215232 237952
rect 0 237488 96 237508
rect 215136 237488 215232 237508
rect 0 237448 117 237488
rect 215115 237448 215232 237488
rect 0 237428 96 237448
rect 215136 237428 215232 237448
rect 0 236984 96 237004
rect 215136 236984 215232 237004
rect 0 236944 117 236984
rect 215115 236944 215232 236984
rect 0 236924 96 236944
rect 215136 236924 215232 236944
rect 0 236480 96 236500
rect 215136 236480 215232 236500
rect 0 236440 117 236480
rect 215115 236440 215232 236480
rect 0 236420 96 236440
rect 215136 236420 215232 236440
rect 0 235976 96 235996
rect 215136 235976 215232 235996
rect 0 235936 117 235976
rect 215115 235936 215232 235976
rect 0 235916 96 235936
rect 215136 235916 215232 235936
rect 0 235472 96 235492
rect 215136 235472 215232 235492
rect 0 235432 117 235472
rect 215115 235432 215232 235472
rect 0 235412 96 235432
rect 215136 235412 215232 235432
rect 0 234968 96 234988
rect 215136 234968 215232 234988
rect 0 234928 117 234968
rect 215115 234928 215232 234968
rect 0 234908 96 234928
rect 215136 234908 215232 234928
rect 0 234464 96 234484
rect 215136 234464 215232 234484
rect 0 234424 117 234464
rect 215115 234424 215232 234464
rect 0 234404 96 234424
rect 215136 234404 215232 234424
rect 0 233960 96 233980
rect 215136 233960 215232 233980
rect 0 233920 117 233960
rect 215115 233920 215232 233960
rect 0 233900 96 233920
rect 215136 233900 215232 233920
rect 0 233456 96 233476
rect 215136 233456 215232 233476
rect 0 233416 117 233456
rect 215115 233416 215232 233456
rect 0 233396 96 233416
rect 215136 233396 215232 233416
rect 0 232952 96 232972
rect 215136 232952 215232 232972
rect 0 232912 117 232952
rect 215115 232912 215232 232952
rect 0 232892 96 232912
rect 215136 232892 215232 232912
rect 0 232448 96 232468
rect 215136 232448 215232 232468
rect 0 232408 117 232448
rect 215115 232408 215232 232448
rect 0 232388 96 232408
rect 215136 232388 215232 232408
rect 0 231944 96 231964
rect 215136 231944 215232 231964
rect 0 231904 117 231944
rect 215115 231904 215232 231944
rect 0 231884 96 231904
rect 215136 231884 215232 231904
rect 0 231440 96 231460
rect 215136 231440 215232 231460
rect 0 231400 117 231440
rect 215115 231400 215232 231440
rect 0 231380 96 231400
rect 215136 231380 215232 231400
rect 0 230936 96 230956
rect 215136 230936 215232 230956
rect 0 230896 117 230936
rect 215115 230896 215232 230936
rect 0 230876 96 230896
rect 215136 230876 215232 230896
rect 0 230432 96 230452
rect 215136 230432 215232 230452
rect 0 230392 117 230432
rect 215115 230392 215232 230432
rect 0 230372 96 230392
rect 215136 230372 215232 230392
rect 0 229928 96 229948
rect 215136 229928 215232 229948
rect 0 229888 117 229928
rect 215115 229888 215232 229928
rect 0 229868 96 229888
rect 215136 229868 215232 229888
rect 0 229424 96 229444
rect 215136 229424 215232 229444
rect 0 229384 117 229424
rect 215115 229384 215232 229424
rect 0 229364 96 229384
rect 215136 229364 215232 229384
rect 0 223712 96 223732
rect 0 223672 117 223712
rect 0 223652 96 223672
rect 0 223208 96 223228
rect 0 223168 117 223208
rect 0 223148 96 223168
rect 0 222704 96 222724
rect 0 222664 117 222704
rect 0 222644 96 222664
rect 0 222200 96 222220
rect 0 222160 117 222200
rect 0 222140 96 222160
rect 0 221696 96 221716
rect 0 221656 117 221696
rect 0 221636 96 221656
rect 0 221192 96 221212
rect 0 221152 117 221192
rect 0 221132 96 221152
rect 0 220688 96 220708
rect 0 220648 117 220688
rect 0 220628 96 220648
rect 0 220184 96 220204
rect 0 220144 117 220184
rect 0 220124 96 220144
rect 0 219680 96 219700
rect 0 219640 117 219680
rect 0 219620 96 219640
rect 0 219176 96 219196
rect 0 219136 117 219176
rect 0 219116 96 219136
rect 0 218672 96 218692
rect 0 218632 117 218672
rect 0 218612 96 218632
rect 0 218168 96 218188
rect 0 218128 117 218168
rect 0 218108 96 218128
rect 0 217664 96 217684
rect 0 217624 117 217664
rect 0 217604 96 217624
rect 0 217160 96 217180
rect 0 217120 117 217160
rect 0 217100 96 217120
rect 0 216656 96 216676
rect 0 216616 117 216656
rect 0 216596 96 216616
rect 0 216152 96 216172
rect 0 216112 117 216152
rect 0 216092 96 216112
rect 0 215648 96 215668
rect 0 215608 117 215648
rect 0 215588 96 215608
rect 0 215144 96 215164
rect 0 215104 117 215144
rect 0 215084 96 215104
rect 0 214640 96 214660
rect 0 214600 117 214640
rect 0 214580 96 214600
rect 0 214136 96 214156
rect 0 214096 117 214136
rect 0 214076 96 214096
rect 0 213632 96 213652
rect 0 213592 117 213632
rect 0 213572 96 213592
rect 0 213128 96 213148
rect 0 213088 117 213128
rect 0 213068 96 213088
rect 0 212624 96 212644
rect 0 212584 117 212624
rect 0 212564 96 212584
rect 0 212120 96 212140
rect 0 212080 117 212120
rect 0 212060 96 212080
rect 0 211616 96 211636
rect 0 211576 117 211616
rect 0 211556 96 211576
rect 0 211112 96 211132
rect 0 211072 117 211112
rect 0 211052 96 211072
rect 0 210608 96 210628
rect 0 210568 117 210608
rect 0 210548 96 210568
rect 0 210104 96 210124
rect 0 210064 117 210104
rect 0 210044 96 210064
rect 0 209600 96 209620
rect 0 209560 117 209600
rect 0 209540 96 209560
rect 0 209096 96 209116
rect 0 209056 117 209096
rect 0 209036 96 209056
rect 0 208592 96 208612
rect 0 208552 117 208592
rect 0 208532 96 208552
rect 0 208088 96 208108
rect 0 208048 117 208088
rect 0 208028 96 208048
rect 0 207584 96 207604
rect 215136 207584 215232 207604
rect 0 207544 117 207584
rect 215115 207544 215232 207584
rect 0 207524 96 207544
rect 215136 207524 215232 207544
rect 0 207080 96 207100
rect 215136 207080 215232 207100
rect 0 207040 117 207080
rect 215115 207040 215232 207080
rect 0 207020 96 207040
rect 215136 207020 215232 207040
rect 0 206576 96 206596
rect 215136 206576 215232 206596
rect 0 206536 117 206576
rect 215115 206536 215232 206576
rect 0 206516 96 206536
rect 215136 206516 215232 206536
rect 0 206072 96 206092
rect 215136 206072 215232 206092
rect 0 206032 117 206072
rect 215115 206032 215232 206072
rect 0 206012 96 206032
rect 215136 206012 215232 206032
rect 0 205568 96 205588
rect 215136 205568 215232 205588
rect 0 205528 117 205568
rect 215115 205528 215232 205568
rect 0 205508 96 205528
rect 215136 205508 215232 205528
rect 0 205064 96 205084
rect 215136 205064 215232 205084
rect 0 205024 117 205064
rect 215115 205024 215232 205064
rect 0 205004 96 205024
rect 215136 205004 215232 205024
rect 0 204560 96 204580
rect 215136 204560 215232 204580
rect 0 204520 117 204560
rect 215115 204520 215232 204560
rect 0 204500 96 204520
rect 215136 204500 215232 204520
rect 0 204056 96 204076
rect 215136 204056 215232 204076
rect 0 204016 117 204056
rect 215115 204016 215232 204056
rect 0 203996 96 204016
rect 215136 203996 215232 204016
rect 0 203552 96 203572
rect 215136 203552 215232 203572
rect 0 203512 117 203552
rect 215115 203512 215232 203552
rect 0 203492 96 203512
rect 215136 203492 215232 203512
rect 0 203048 96 203068
rect 215136 203048 215232 203068
rect 0 203008 117 203048
rect 215115 203008 215232 203048
rect 0 202988 96 203008
rect 215136 202988 215232 203008
rect 0 202544 96 202564
rect 215136 202544 215232 202564
rect 0 202504 117 202544
rect 215115 202504 215232 202544
rect 0 202484 96 202504
rect 215136 202484 215232 202504
rect 0 202040 96 202060
rect 215136 202040 215232 202060
rect 0 202000 117 202040
rect 215115 202000 215232 202040
rect 0 201980 96 202000
rect 215136 201980 215232 202000
rect 0 201536 96 201556
rect 215136 201536 215232 201556
rect 0 201496 117 201536
rect 215115 201496 215232 201536
rect 0 201476 96 201496
rect 215136 201476 215232 201496
rect 0 201032 96 201052
rect 215136 201032 215232 201052
rect 0 200992 117 201032
rect 215115 200992 215232 201032
rect 0 200972 96 200992
rect 215136 200972 215232 200992
rect 0 200528 96 200548
rect 215136 200528 215232 200548
rect 0 200488 117 200528
rect 215115 200488 215232 200528
rect 0 200468 96 200488
rect 215136 200468 215232 200488
rect 0 200024 96 200044
rect 215136 200024 215232 200044
rect 0 199984 117 200024
rect 215115 199984 215232 200024
rect 0 199964 96 199984
rect 215136 199964 215232 199984
rect 0 199520 96 199540
rect 215136 199520 215232 199540
rect 0 199480 117 199520
rect 215115 199480 215232 199520
rect 0 199460 96 199480
rect 215136 199460 215232 199480
rect 0 199016 96 199036
rect 215136 199016 215232 199036
rect 0 198976 117 199016
rect 215115 198976 215232 199016
rect 0 198956 96 198976
rect 215136 198956 215232 198976
rect 0 198512 96 198532
rect 215136 198512 215232 198532
rect 0 198472 117 198512
rect 215115 198472 215232 198512
rect 0 198452 96 198472
rect 215136 198452 215232 198472
rect 0 198008 96 198028
rect 215136 198008 215232 198028
rect 0 197968 117 198008
rect 215115 197968 215232 198008
rect 0 197948 96 197968
rect 215136 197948 215232 197968
rect 0 197504 96 197524
rect 215136 197504 215232 197524
rect 0 197464 117 197504
rect 215115 197464 215232 197504
rect 0 197444 96 197464
rect 215136 197444 215232 197464
rect 0 197000 96 197020
rect 215136 197000 215232 197020
rect 0 196960 117 197000
rect 215115 196960 215232 197000
rect 0 196940 96 196960
rect 215136 196940 215232 196960
rect 0 196496 96 196516
rect 215136 196496 215232 196516
rect 0 196456 117 196496
rect 215115 196456 215232 196496
rect 0 196436 96 196456
rect 215136 196436 215232 196456
rect 0 195992 96 196012
rect 215136 195992 215232 196012
rect 0 195952 117 195992
rect 215115 195952 215232 195992
rect 0 195932 96 195952
rect 215136 195932 215232 195952
rect 0 195488 96 195508
rect 215136 195488 215232 195508
rect 0 195448 117 195488
rect 215115 195448 215232 195488
rect 0 195428 96 195448
rect 215136 195428 215232 195448
rect 0 194984 96 195004
rect 215136 194984 215232 195004
rect 0 194944 117 194984
rect 215115 194944 215232 194984
rect 0 194924 96 194944
rect 215136 194924 215232 194944
rect 0 194480 96 194500
rect 215136 194480 215232 194500
rect 0 194440 117 194480
rect 215115 194440 215232 194480
rect 0 194420 96 194440
rect 215136 194420 215232 194440
rect 0 193976 96 193996
rect 215136 193976 215232 193996
rect 0 193936 117 193976
rect 215115 193936 215232 193976
rect 0 193916 96 193936
rect 215136 193916 215232 193936
rect 0 193472 96 193492
rect 215136 193472 215232 193492
rect 0 193432 117 193472
rect 215115 193432 215232 193472
rect 0 193412 96 193432
rect 215136 193412 215232 193432
rect 0 192968 96 192988
rect 215136 192968 215232 192988
rect 0 192928 117 192968
rect 215115 192928 215232 192968
rect 0 192908 96 192928
rect 215136 192908 215232 192928
rect 0 192464 96 192484
rect 215136 192464 215232 192484
rect 0 192424 117 192464
rect 215115 192424 215232 192464
rect 0 192404 96 192424
rect 215136 192404 215232 192424
rect 0 191960 96 191980
rect 215136 191960 215232 191980
rect 0 191920 117 191960
rect 215115 191920 215232 191960
rect 0 191900 96 191920
rect 215136 191900 215232 191920
rect 0 191456 96 191476
rect 215136 191456 215232 191476
rect 0 191416 117 191456
rect 215115 191416 215232 191456
rect 0 191396 96 191416
rect 215136 191396 215232 191416
rect 0 190952 96 190972
rect 215136 190952 215232 190972
rect 0 190912 117 190952
rect 215115 190912 215232 190952
rect 0 190892 96 190912
rect 215136 190892 215232 190912
rect 0 190448 96 190468
rect 215136 190448 215232 190468
rect 0 190408 117 190448
rect 215115 190408 215232 190448
rect 0 190388 96 190408
rect 215136 190388 215232 190408
rect 0 189944 96 189964
rect 215136 189944 215232 189964
rect 0 189904 117 189944
rect 215115 189904 215232 189944
rect 0 189884 96 189904
rect 215136 189884 215232 189904
rect 0 189440 96 189460
rect 215136 189440 215232 189460
rect 0 189400 117 189440
rect 215115 189400 215232 189440
rect 0 189380 96 189400
rect 215136 189380 215232 189400
rect 0 188936 96 188956
rect 215136 188936 215232 188956
rect 0 188896 117 188936
rect 215115 188896 215232 188936
rect 0 188876 96 188896
rect 215136 188876 215232 188896
rect 0 188432 96 188452
rect 215136 188432 215232 188452
rect 0 188392 117 188432
rect 215115 188392 215232 188432
rect 0 188372 96 188392
rect 215136 188372 215232 188392
rect 0 187928 96 187948
rect 215136 187928 215232 187948
rect 0 187888 117 187928
rect 215115 187888 215232 187928
rect 0 187868 96 187888
rect 215136 187868 215232 187888
rect 0 187424 96 187444
rect 215136 187424 215232 187444
rect 0 187384 117 187424
rect 215115 187384 215232 187424
rect 0 187364 96 187384
rect 215136 187364 215232 187384
rect 0 186920 96 186940
rect 215136 186920 215232 186940
rect 0 186880 117 186920
rect 215115 186880 215232 186920
rect 0 186860 96 186880
rect 215136 186860 215232 186880
rect 0 186416 96 186436
rect 215136 186416 215232 186436
rect 0 186376 117 186416
rect 215115 186376 215232 186416
rect 0 186356 96 186376
rect 215136 186356 215232 186376
rect 0 180704 96 180724
rect 0 180664 117 180704
rect 0 180644 96 180664
rect 0 180200 96 180220
rect 0 180160 117 180200
rect 0 180140 96 180160
rect 0 179696 96 179716
rect 0 179656 117 179696
rect 0 179636 96 179656
rect 0 179192 96 179212
rect 0 179152 117 179192
rect 0 179132 96 179152
rect 0 178688 96 178708
rect 0 178648 117 178688
rect 0 178628 96 178648
rect 0 178184 96 178204
rect 0 178144 117 178184
rect 0 178124 96 178144
rect 0 177680 96 177700
rect 0 177640 117 177680
rect 0 177620 96 177640
rect 0 177176 96 177196
rect 0 177136 117 177176
rect 0 177116 96 177136
rect 0 176672 96 176692
rect 0 176632 117 176672
rect 0 176612 96 176632
rect 0 176168 96 176188
rect 0 176128 117 176168
rect 0 176108 96 176128
rect 0 175664 96 175684
rect 0 175624 117 175664
rect 0 175604 96 175624
rect 0 175160 96 175180
rect 0 175120 117 175160
rect 0 175100 96 175120
rect 0 174656 96 174676
rect 0 174616 117 174656
rect 0 174596 96 174616
rect 0 174152 96 174172
rect 0 174112 117 174152
rect 0 174092 96 174112
rect 0 173648 96 173668
rect 0 173608 117 173648
rect 0 173588 96 173608
rect 0 173144 96 173164
rect 0 173104 117 173144
rect 0 173084 96 173104
rect 0 172640 96 172660
rect 0 172600 117 172640
rect 0 172580 96 172600
rect 0 172136 96 172156
rect 0 172096 117 172136
rect 0 172076 96 172096
rect 0 171632 96 171652
rect 0 171592 117 171632
rect 0 171572 96 171592
rect 0 171128 96 171148
rect 0 171088 117 171128
rect 0 171068 96 171088
rect 0 170624 96 170644
rect 0 170584 117 170624
rect 0 170564 96 170584
rect 0 170120 96 170140
rect 0 170080 117 170120
rect 0 170060 96 170080
rect 0 169616 96 169636
rect 0 169576 117 169616
rect 0 169556 96 169576
rect 0 169112 96 169132
rect 0 169072 117 169112
rect 0 169052 96 169072
rect 0 168608 96 168628
rect 0 168568 117 168608
rect 0 168548 96 168568
rect 0 168104 96 168124
rect 0 168064 117 168104
rect 0 168044 96 168064
rect 0 167600 96 167620
rect 0 167560 117 167600
rect 0 167540 96 167560
rect 0 167096 96 167116
rect 0 167056 117 167096
rect 0 167036 96 167056
rect 0 166592 96 166612
rect 0 166552 117 166592
rect 0 166532 96 166552
rect 0 166088 96 166108
rect 0 166048 117 166088
rect 0 166028 96 166048
rect 0 165584 96 165604
rect 0 165544 117 165584
rect 0 165524 96 165544
rect 0 165080 96 165100
rect 0 165040 117 165080
rect 0 165020 96 165040
rect 0 164576 96 164596
rect 215136 164576 215232 164596
rect 0 164536 117 164576
rect 215115 164536 215232 164576
rect 0 164516 96 164536
rect 215136 164516 215232 164536
rect 0 164072 96 164092
rect 215136 164072 215232 164092
rect 0 164032 117 164072
rect 215115 164032 215232 164072
rect 0 164012 96 164032
rect 215136 164012 215232 164032
rect 0 163568 96 163588
rect 215136 163568 215232 163588
rect 0 163528 117 163568
rect 215115 163528 215232 163568
rect 0 163508 96 163528
rect 215136 163508 215232 163528
rect 0 163064 96 163084
rect 215136 163064 215232 163084
rect 0 163024 117 163064
rect 215115 163024 215232 163064
rect 0 163004 96 163024
rect 215136 163004 215232 163024
rect 0 162560 96 162580
rect 215136 162560 215232 162580
rect 0 162520 117 162560
rect 215115 162520 215232 162560
rect 0 162500 96 162520
rect 215136 162500 215232 162520
rect 0 162056 96 162076
rect 215136 162056 215232 162076
rect 0 162016 117 162056
rect 215115 162016 215232 162056
rect 0 161996 96 162016
rect 215136 161996 215232 162016
rect 0 161552 96 161572
rect 215136 161552 215232 161572
rect 0 161512 117 161552
rect 215115 161512 215232 161552
rect 0 161492 96 161512
rect 215136 161492 215232 161512
rect 0 161048 96 161068
rect 215136 161048 215232 161068
rect 0 161008 117 161048
rect 215115 161008 215232 161048
rect 0 160988 96 161008
rect 215136 160988 215232 161008
rect 0 160544 96 160564
rect 215136 160544 215232 160564
rect 0 160504 117 160544
rect 215115 160504 215232 160544
rect 0 160484 96 160504
rect 215136 160484 215232 160504
rect 0 160040 96 160060
rect 215136 160040 215232 160060
rect 0 160000 117 160040
rect 215115 160000 215232 160040
rect 0 159980 96 160000
rect 215136 159980 215232 160000
rect 0 159536 96 159556
rect 215136 159536 215232 159556
rect 0 159496 117 159536
rect 215115 159496 215232 159536
rect 0 159476 96 159496
rect 215136 159476 215232 159496
rect 0 159032 96 159052
rect 215136 159032 215232 159052
rect 0 158992 117 159032
rect 215115 158992 215232 159032
rect 0 158972 96 158992
rect 215136 158972 215232 158992
rect 0 158528 96 158548
rect 215136 158528 215232 158548
rect 0 158488 117 158528
rect 215115 158488 215232 158528
rect 0 158468 96 158488
rect 215136 158468 215232 158488
rect 0 158024 96 158044
rect 215136 158024 215232 158044
rect 0 157984 117 158024
rect 215115 157984 215232 158024
rect 0 157964 96 157984
rect 215136 157964 215232 157984
rect 0 157520 96 157540
rect 215136 157520 215232 157540
rect 0 157480 117 157520
rect 215115 157480 215232 157520
rect 0 157460 96 157480
rect 215136 157460 215232 157480
rect 0 157016 96 157036
rect 215136 157016 215232 157036
rect 0 156976 117 157016
rect 215115 156976 215232 157016
rect 0 156956 96 156976
rect 215136 156956 215232 156976
rect 0 156512 96 156532
rect 215136 156512 215232 156532
rect 0 156472 117 156512
rect 215115 156472 215232 156512
rect 0 156452 96 156472
rect 215136 156452 215232 156472
rect 0 156008 96 156028
rect 215136 156008 215232 156028
rect 0 155968 117 156008
rect 215115 155968 215232 156008
rect 0 155948 96 155968
rect 215136 155948 215232 155968
rect 0 155504 96 155524
rect 215136 155504 215232 155524
rect 0 155464 117 155504
rect 215115 155464 215232 155504
rect 0 155444 96 155464
rect 215136 155444 215232 155464
rect 0 155000 96 155020
rect 215136 155000 215232 155020
rect 0 154960 117 155000
rect 215115 154960 215232 155000
rect 0 154940 96 154960
rect 215136 154940 215232 154960
rect 0 154496 96 154516
rect 215136 154496 215232 154516
rect 0 154456 117 154496
rect 215115 154456 215232 154496
rect 0 154436 96 154456
rect 215136 154436 215232 154456
rect 0 153992 96 154012
rect 215136 153992 215232 154012
rect 0 153952 117 153992
rect 215115 153952 215232 153992
rect 0 153932 96 153952
rect 215136 153932 215232 153952
rect 0 153488 96 153508
rect 215136 153488 215232 153508
rect 0 153448 117 153488
rect 215115 153448 215232 153488
rect 0 153428 96 153448
rect 215136 153428 215232 153448
rect 0 152984 96 153004
rect 215136 152984 215232 153004
rect 0 152944 117 152984
rect 215115 152944 215232 152984
rect 0 152924 96 152944
rect 215136 152924 215232 152944
rect 0 152480 96 152500
rect 215136 152480 215232 152500
rect 0 152440 117 152480
rect 215115 152440 215232 152480
rect 0 152420 96 152440
rect 215136 152420 215232 152440
rect 0 151976 96 151996
rect 215136 151976 215232 151996
rect 0 151936 117 151976
rect 215115 151936 215232 151976
rect 0 151916 96 151936
rect 215136 151916 215232 151936
rect 0 151472 96 151492
rect 215136 151472 215232 151492
rect 0 151432 117 151472
rect 215115 151432 215232 151472
rect 0 151412 96 151432
rect 215136 151412 215232 151432
rect 0 150968 96 150988
rect 215136 150968 215232 150988
rect 0 150928 117 150968
rect 215115 150928 215232 150968
rect 0 150908 96 150928
rect 215136 150908 215232 150928
rect 0 150464 96 150484
rect 215136 150464 215232 150484
rect 0 150424 117 150464
rect 215115 150424 215232 150464
rect 0 150404 96 150424
rect 215136 150404 215232 150424
rect 0 149960 96 149980
rect 215136 149960 215232 149980
rect 0 149920 117 149960
rect 215115 149920 215232 149960
rect 0 149900 96 149920
rect 215136 149900 215232 149920
rect 0 149456 96 149476
rect 215136 149456 215232 149476
rect 0 149416 117 149456
rect 215115 149416 215232 149456
rect 0 149396 96 149416
rect 215136 149396 215232 149416
rect 0 148952 96 148972
rect 215136 148952 215232 148972
rect 0 148912 117 148952
rect 215115 148912 215232 148952
rect 0 148892 96 148912
rect 215136 148892 215232 148912
rect 0 148448 96 148468
rect 215136 148448 215232 148468
rect 0 148408 117 148448
rect 215115 148408 215232 148448
rect 0 148388 96 148408
rect 215136 148388 215232 148408
rect 0 147944 96 147964
rect 215136 147944 215232 147964
rect 0 147904 117 147944
rect 215115 147904 215232 147944
rect 0 147884 96 147904
rect 215136 147884 215232 147904
rect 0 147440 96 147460
rect 215136 147440 215232 147460
rect 0 147400 117 147440
rect 215115 147400 215232 147440
rect 0 147380 96 147400
rect 215136 147380 215232 147400
rect 0 146936 96 146956
rect 215136 146936 215232 146956
rect 0 146896 117 146936
rect 215115 146896 215232 146936
rect 0 146876 96 146896
rect 215136 146876 215232 146896
rect 0 146432 96 146452
rect 215136 146432 215232 146452
rect 0 146392 117 146432
rect 215115 146392 215232 146432
rect 0 146372 96 146392
rect 215136 146372 215232 146392
rect 0 145928 96 145948
rect 215136 145928 215232 145948
rect 0 145888 117 145928
rect 215115 145888 215232 145928
rect 0 145868 96 145888
rect 215136 145868 215232 145888
rect 0 145424 96 145444
rect 215136 145424 215232 145444
rect 0 145384 117 145424
rect 215115 145384 215232 145424
rect 0 145364 96 145384
rect 215136 145364 215232 145384
rect 0 144920 96 144940
rect 215136 144920 215232 144940
rect 0 144880 117 144920
rect 215115 144880 215232 144920
rect 0 144860 96 144880
rect 215136 144860 215232 144880
rect 0 144416 96 144436
rect 215136 144416 215232 144436
rect 0 144376 117 144416
rect 215115 144376 215232 144416
rect 0 144356 96 144376
rect 215136 144356 215232 144376
rect 0 143912 96 143932
rect 215136 143912 215232 143932
rect 0 143872 117 143912
rect 215115 143872 215232 143912
rect 0 143852 96 143872
rect 215136 143852 215232 143872
rect 0 143408 96 143428
rect 215136 143408 215232 143428
rect 0 143368 117 143408
rect 215115 143368 215232 143408
rect 0 143348 96 143368
rect 215136 143348 215232 143368
rect 0 137696 96 137716
rect 0 137656 117 137696
rect 0 137636 96 137656
rect 0 137192 96 137212
rect 0 137152 117 137192
rect 0 137132 96 137152
rect 0 136688 96 136708
rect 0 136648 117 136688
rect 0 136628 96 136648
rect 0 136184 96 136204
rect 0 136144 117 136184
rect 0 136124 96 136144
rect 0 135680 96 135700
rect 0 135640 117 135680
rect 0 135620 96 135640
rect 0 135176 96 135196
rect 0 135136 117 135176
rect 0 135116 96 135136
rect 0 134672 96 134692
rect 0 134632 117 134672
rect 0 134612 96 134632
rect 0 134168 96 134188
rect 0 134128 117 134168
rect 0 134108 96 134128
rect 0 133664 96 133684
rect 0 133624 117 133664
rect 0 133604 96 133624
rect 0 133160 96 133180
rect 0 133120 117 133160
rect 0 133100 96 133120
rect 0 132656 96 132676
rect 0 132616 117 132656
rect 0 132596 96 132616
rect 0 132152 96 132172
rect 0 132112 117 132152
rect 0 132092 96 132112
rect 0 131648 96 131668
rect 0 131608 117 131648
rect 0 131588 96 131608
rect 0 131144 96 131164
rect 0 131104 117 131144
rect 0 131084 96 131104
rect 0 130640 96 130660
rect 0 130600 117 130640
rect 0 130580 96 130600
rect 0 130136 96 130156
rect 0 130096 117 130136
rect 0 130076 96 130096
rect 0 129632 96 129652
rect 0 129592 117 129632
rect 0 129572 96 129592
rect 0 129128 96 129148
rect 0 129088 117 129128
rect 0 129068 96 129088
rect 0 128624 96 128644
rect 0 128584 117 128624
rect 0 128564 96 128584
rect 0 128120 96 128140
rect 0 128080 117 128120
rect 0 128060 96 128080
rect 0 127616 96 127636
rect 0 127576 117 127616
rect 0 127556 96 127576
rect 0 127112 96 127132
rect 0 127072 117 127112
rect 0 127052 96 127072
rect 0 126608 96 126628
rect 0 126568 117 126608
rect 0 126548 96 126568
rect 0 126104 96 126124
rect 0 126064 117 126104
rect 0 126044 96 126064
rect 0 125600 96 125620
rect 0 125560 117 125600
rect 0 125540 96 125560
rect 0 125096 96 125116
rect 0 125056 117 125096
rect 0 125036 96 125056
rect 0 124592 96 124612
rect 0 124552 117 124592
rect 0 124532 96 124552
rect 0 124088 96 124108
rect 0 124048 117 124088
rect 0 124028 96 124048
rect 0 123584 96 123604
rect 0 123544 117 123584
rect 0 123524 96 123544
rect 0 123080 96 123100
rect 0 123040 117 123080
rect 0 123020 96 123040
rect 0 122576 96 122596
rect 0 122536 117 122576
rect 0 122516 96 122536
rect 0 122072 96 122092
rect 0 122032 117 122072
rect 0 122012 96 122032
rect 0 121568 96 121588
rect 215136 121568 215232 121588
rect 0 121528 117 121568
rect 215115 121528 215232 121568
rect 0 121508 96 121528
rect 215136 121508 215232 121528
rect 0 121064 96 121084
rect 215136 121064 215232 121084
rect 0 121024 117 121064
rect 215115 121024 215232 121064
rect 0 121004 96 121024
rect 215136 121004 215232 121024
rect 0 120560 96 120580
rect 215136 120560 215232 120580
rect 0 120520 117 120560
rect 215115 120520 215232 120560
rect 0 120500 96 120520
rect 215136 120500 215232 120520
rect 0 120056 96 120076
rect 215136 120056 215232 120076
rect 0 120016 117 120056
rect 215115 120016 215232 120056
rect 0 119996 96 120016
rect 215136 119996 215232 120016
rect 0 119552 96 119572
rect 215136 119552 215232 119572
rect 0 119512 117 119552
rect 215115 119512 215232 119552
rect 0 119492 96 119512
rect 215136 119492 215232 119512
rect 0 119048 96 119068
rect 215136 119048 215232 119068
rect 0 119008 117 119048
rect 215115 119008 215232 119048
rect 0 118988 96 119008
rect 215136 118988 215232 119008
rect 0 118544 96 118564
rect 215136 118544 215232 118564
rect 0 118504 117 118544
rect 215115 118504 215232 118544
rect 0 118484 96 118504
rect 215136 118484 215232 118504
rect 0 118040 96 118060
rect 215136 118040 215232 118060
rect 0 118000 117 118040
rect 215115 118000 215232 118040
rect 0 117980 96 118000
rect 215136 117980 215232 118000
rect 0 117536 96 117556
rect 215136 117536 215232 117556
rect 0 117496 117 117536
rect 215115 117496 215232 117536
rect 0 117476 96 117496
rect 215136 117476 215232 117496
rect 0 117032 96 117052
rect 215136 117032 215232 117052
rect 0 116992 117 117032
rect 215115 116992 215232 117032
rect 0 116972 96 116992
rect 215136 116972 215232 116992
rect 0 116528 96 116548
rect 215136 116528 215232 116548
rect 0 116488 117 116528
rect 215115 116488 215232 116528
rect 0 116468 96 116488
rect 215136 116468 215232 116488
rect 0 116024 96 116044
rect 215136 116024 215232 116044
rect 0 115984 117 116024
rect 215115 115984 215232 116024
rect 0 115964 96 115984
rect 215136 115964 215232 115984
rect 0 115520 96 115540
rect 215136 115520 215232 115540
rect 0 115480 117 115520
rect 215115 115480 215232 115520
rect 0 115460 96 115480
rect 215136 115460 215232 115480
rect 0 115016 96 115036
rect 215136 115016 215232 115036
rect 0 114976 117 115016
rect 215115 114976 215232 115016
rect 0 114956 96 114976
rect 215136 114956 215232 114976
rect 0 114512 96 114532
rect 215136 114512 215232 114532
rect 0 114472 117 114512
rect 215115 114472 215232 114512
rect 0 114452 96 114472
rect 215136 114452 215232 114472
rect 0 114008 96 114028
rect 215136 114008 215232 114028
rect 0 113968 117 114008
rect 215115 113968 215232 114008
rect 0 113948 96 113968
rect 215136 113948 215232 113968
rect 0 113504 96 113524
rect 215136 113504 215232 113524
rect 0 113464 117 113504
rect 215115 113464 215232 113504
rect 0 113444 96 113464
rect 215136 113444 215232 113464
rect 0 113000 96 113020
rect 215136 113000 215232 113020
rect 0 112960 117 113000
rect 215115 112960 215232 113000
rect 0 112940 96 112960
rect 215136 112940 215232 112960
rect 0 112496 96 112516
rect 215136 112496 215232 112516
rect 0 112456 117 112496
rect 215115 112456 215232 112496
rect 0 112436 96 112456
rect 215136 112436 215232 112456
rect 0 111992 96 112012
rect 215136 111992 215232 112012
rect 0 111952 117 111992
rect 215115 111952 215232 111992
rect 0 111932 96 111952
rect 215136 111932 215232 111952
rect 0 111488 96 111508
rect 215136 111488 215232 111508
rect 0 111448 117 111488
rect 215115 111448 215232 111488
rect 0 111428 96 111448
rect 215136 111428 215232 111448
rect 0 110984 96 111004
rect 215136 110984 215232 111004
rect 0 110944 117 110984
rect 215115 110944 215232 110984
rect 0 110924 96 110944
rect 215136 110924 215232 110944
rect 0 110480 96 110500
rect 215136 110480 215232 110500
rect 0 110440 117 110480
rect 215115 110440 215232 110480
rect 0 110420 96 110440
rect 215136 110420 215232 110440
rect 0 109976 96 109996
rect 215136 109976 215232 109996
rect 0 109936 117 109976
rect 215115 109936 215232 109976
rect 0 109916 96 109936
rect 215136 109916 215232 109936
rect 0 109472 96 109492
rect 215136 109472 215232 109492
rect 0 109432 117 109472
rect 215115 109432 215232 109472
rect 0 109412 96 109432
rect 215136 109412 215232 109432
rect 0 108968 96 108988
rect 215136 108968 215232 108988
rect 0 108928 117 108968
rect 215115 108928 215232 108968
rect 0 108908 96 108928
rect 215136 108908 215232 108928
rect 0 108464 96 108484
rect 215136 108464 215232 108484
rect 0 108424 117 108464
rect 215115 108424 215232 108464
rect 0 108404 96 108424
rect 215136 108404 215232 108424
rect 0 107960 96 107980
rect 215136 107960 215232 107980
rect 0 107920 117 107960
rect 215115 107920 215232 107960
rect 0 107900 96 107920
rect 215136 107900 215232 107920
rect 0 107456 96 107476
rect 215136 107456 215232 107476
rect 0 107416 117 107456
rect 215115 107416 215232 107456
rect 0 107396 96 107416
rect 215136 107396 215232 107416
rect 0 106952 96 106972
rect 215136 106952 215232 106972
rect 0 106912 117 106952
rect 215115 106912 215232 106952
rect 0 106892 96 106912
rect 215136 106892 215232 106912
rect 0 106448 96 106468
rect 215136 106448 215232 106468
rect 0 106408 117 106448
rect 215115 106408 215232 106448
rect 0 106388 96 106408
rect 215136 106388 215232 106408
rect 0 105944 96 105964
rect 215136 105944 215232 105964
rect 0 105904 117 105944
rect 215115 105904 215232 105944
rect 0 105884 96 105904
rect 215136 105884 215232 105904
rect 0 105440 96 105460
rect 215136 105440 215232 105460
rect 0 105400 117 105440
rect 215115 105400 215232 105440
rect 0 105380 96 105400
rect 215136 105380 215232 105400
rect 0 104936 96 104956
rect 215136 104936 215232 104956
rect 0 104896 117 104936
rect 215115 104896 215232 104936
rect 0 104876 96 104896
rect 215136 104876 215232 104896
rect 0 104432 96 104452
rect 215136 104432 215232 104452
rect 0 104392 117 104432
rect 215115 104392 215232 104432
rect 0 104372 96 104392
rect 215136 104372 215232 104392
rect 0 103928 96 103948
rect 215136 103928 215232 103948
rect 0 103888 117 103928
rect 215115 103888 215232 103928
rect 0 103868 96 103888
rect 215136 103868 215232 103888
rect 0 103424 96 103444
rect 215136 103424 215232 103444
rect 0 103384 117 103424
rect 215115 103384 215232 103424
rect 0 103364 96 103384
rect 215136 103364 215232 103384
rect 0 102920 96 102940
rect 215136 102920 215232 102940
rect 0 102880 117 102920
rect 215115 102880 215232 102920
rect 0 102860 96 102880
rect 215136 102860 215232 102880
rect 0 102416 96 102436
rect 215136 102416 215232 102436
rect 0 102376 117 102416
rect 215115 102376 215232 102416
rect 0 102356 96 102376
rect 215136 102356 215232 102376
rect 0 101912 96 101932
rect 215136 101912 215232 101932
rect 0 101872 117 101912
rect 215115 101872 215232 101912
rect 0 101852 96 101872
rect 215136 101852 215232 101872
rect 0 101408 96 101428
rect 215136 101408 215232 101428
rect 0 101368 117 101408
rect 215115 101368 215232 101408
rect 0 101348 96 101368
rect 215136 101348 215232 101368
rect 0 100904 96 100924
rect 215136 100904 215232 100924
rect 0 100864 117 100904
rect 215115 100864 215232 100904
rect 0 100844 96 100864
rect 215136 100844 215232 100864
rect 0 100400 96 100420
rect 215136 100400 215232 100420
rect 0 100360 117 100400
rect 215115 100360 215232 100400
rect 0 100340 96 100360
rect 215136 100340 215232 100360
rect 0 94688 96 94708
rect 0 94648 117 94688
rect 0 94628 96 94648
rect 0 94184 96 94204
rect 0 94144 117 94184
rect 0 94124 96 94144
rect 0 93680 96 93700
rect 0 93640 117 93680
rect 0 93620 96 93640
rect 0 93176 96 93196
rect 0 93136 117 93176
rect 0 93116 96 93136
rect 0 92672 96 92692
rect 0 92632 117 92672
rect 0 92612 96 92632
rect 0 92168 96 92188
rect 0 92128 117 92168
rect 0 92108 96 92128
rect 0 91664 96 91684
rect 0 91624 117 91664
rect 0 91604 96 91624
rect 0 91160 96 91180
rect 0 91120 117 91160
rect 0 91100 96 91120
rect 0 90656 96 90676
rect 0 90616 117 90656
rect 0 90596 96 90616
rect 0 90152 96 90172
rect 0 90112 117 90152
rect 0 90092 96 90112
rect 0 89648 96 89668
rect 0 89608 117 89648
rect 0 89588 96 89608
rect 0 89144 96 89164
rect 0 89104 117 89144
rect 0 89084 96 89104
rect 0 88640 96 88660
rect 0 88600 117 88640
rect 0 88580 96 88600
rect 0 88136 96 88156
rect 0 88096 117 88136
rect 0 88076 96 88096
rect 0 87632 96 87652
rect 0 87592 117 87632
rect 0 87572 96 87592
rect 0 87128 96 87148
rect 0 87088 117 87128
rect 0 87068 96 87088
rect 0 86624 96 86644
rect 0 86584 117 86624
rect 0 86564 96 86584
rect 0 86120 96 86140
rect 0 86080 117 86120
rect 0 86060 96 86080
rect 0 85616 96 85636
rect 0 85576 117 85616
rect 0 85556 96 85576
rect 0 85112 96 85132
rect 0 85072 117 85112
rect 0 85052 96 85072
rect 0 84608 96 84628
rect 0 84568 117 84608
rect 0 84548 96 84568
rect 0 84104 96 84124
rect 0 84064 117 84104
rect 0 84044 96 84064
rect 0 83600 96 83620
rect 0 83560 117 83600
rect 0 83540 96 83560
rect 0 83096 96 83116
rect 0 83056 117 83096
rect 0 83036 96 83056
rect 0 82592 96 82612
rect 0 82552 117 82592
rect 0 82532 96 82552
rect 0 82088 96 82108
rect 0 82048 117 82088
rect 0 82028 96 82048
rect 0 81584 96 81604
rect 0 81544 117 81584
rect 0 81524 96 81544
rect 0 81080 96 81100
rect 0 81040 117 81080
rect 0 81020 96 81040
rect 0 80576 96 80596
rect 0 80536 117 80576
rect 0 80516 96 80536
rect 0 80072 96 80092
rect 0 80032 117 80072
rect 0 80012 96 80032
rect 0 79568 96 79588
rect 0 79528 117 79568
rect 0 79508 96 79528
rect 0 79064 96 79084
rect 0 79024 117 79064
rect 0 79004 96 79024
rect 0 78560 96 78580
rect 215136 78560 215232 78580
rect 0 78520 117 78560
rect 215115 78520 215232 78560
rect 0 78500 96 78520
rect 215136 78500 215232 78520
rect 0 78056 96 78076
rect 215136 78056 215232 78076
rect 0 78016 117 78056
rect 215115 78016 215232 78056
rect 0 77996 96 78016
rect 215136 77996 215232 78016
rect 0 77552 96 77572
rect 215136 77552 215232 77572
rect 0 77512 117 77552
rect 215115 77512 215232 77552
rect 0 77492 96 77512
rect 215136 77492 215232 77512
rect 0 77048 96 77068
rect 215136 77048 215232 77068
rect 0 77008 117 77048
rect 215115 77008 215232 77048
rect 0 76988 96 77008
rect 215136 76988 215232 77008
rect 0 76544 96 76564
rect 215136 76544 215232 76564
rect 0 76504 117 76544
rect 215115 76504 215232 76544
rect 0 76484 96 76504
rect 215136 76484 215232 76504
rect 0 76040 96 76060
rect 215136 76040 215232 76060
rect 0 76000 117 76040
rect 215115 76000 215232 76040
rect 0 75980 96 76000
rect 215136 75980 215232 76000
rect 0 75536 96 75556
rect 215136 75536 215232 75556
rect 0 75496 117 75536
rect 215115 75496 215232 75536
rect 0 75476 96 75496
rect 215136 75476 215232 75496
rect 0 75032 96 75052
rect 215136 75032 215232 75052
rect 0 74992 117 75032
rect 215115 74992 215232 75032
rect 0 74972 96 74992
rect 215136 74972 215232 74992
rect 0 74528 96 74548
rect 215136 74528 215232 74548
rect 0 74488 117 74528
rect 215115 74488 215232 74528
rect 0 74468 96 74488
rect 215136 74468 215232 74488
rect 0 74024 96 74044
rect 215136 74024 215232 74044
rect 0 73984 117 74024
rect 215115 73984 215232 74024
rect 0 73964 96 73984
rect 215136 73964 215232 73984
rect 0 73520 96 73540
rect 215136 73520 215232 73540
rect 0 73480 117 73520
rect 215115 73480 215232 73520
rect 0 73460 96 73480
rect 215136 73460 215232 73480
rect 0 73016 96 73036
rect 215136 73016 215232 73036
rect 0 72976 117 73016
rect 215115 72976 215232 73016
rect 0 72956 96 72976
rect 215136 72956 215232 72976
rect 0 72512 96 72532
rect 215136 72512 215232 72532
rect 0 72472 117 72512
rect 215115 72472 215232 72512
rect 0 72452 96 72472
rect 215136 72452 215232 72472
rect 0 72008 96 72028
rect 215136 72008 215232 72028
rect 0 71968 117 72008
rect 215115 71968 215232 72008
rect 0 71948 96 71968
rect 215136 71948 215232 71968
rect 0 71504 96 71524
rect 215136 71504 215232 71524
rect 0 71464 117 71504
rect 215115 71464 215232 71504
rect 0 71444 96 71464
rect 215136 71444 215232 71464
rect 0 71000 96 71020
rect 215136 71000 215232 71020
rect 0 70960 117 71000
rect 215115 70960 215232 71000
rect 0 70940 96 70960
rect 215136 70940 215232 70960
rect 0 70496 96 70516
rect 215136 70496 215232 70516
rect 0 70456 117 70496
rect 215115 70456 215232 70496
rect 0 70436 96 70456
rect 215136 70436 215232 70456
rect 0 69992 96 70012
rect 215136 69992 215232 70012
rect 0 69952 117 69992
rect 215115 69952 215232 69992
rect 0 69932 96 69952
rect 215136 69932 215232 69952
rect 0 69488 96 69508
rect 215136 69488 215232 69508
rect 0 69448 117 69488
rect 215115 69448 215232 69488
rect 0 69428 96 69448
rect 215136 69428 215232 69448
rect 0 68984 96 69004
rect 215136 68984 215232 69004
rect 0 68944 117 68984
rect 215115 68944 215232 68984
rect 0 68924 96 68944
rect 215136 68924 215232 68944
rect 0 68480 96 68500
rect 215136 68480 215232 68500
rect 0 68440 117 68480
rect 215115 68440 215232 68480
rect 0 68420 96 68440
rect 215136 68420 215232 68440
rect 0 67976 96 67996
rect 215136 67976 215232 67996
rect 0 67936 117 67976
rect 215115 67936 215232 67976
rect 0 67916 96 67936
rect 215136 67916 215232 67936
rect 0 67472 96 67492
rect 215136 67472 215232 67492
rect 0 67432 117 67472
rect 215115 67432 215232 67472
rect 0 67412 96 67432
rect 215136 67412 215232 67432
rect 0 66968 96 66988
rect 215136 66968 215232 66988
rect 0 66928 117 66968
rect 215115 66928 215232 66968
rect 0 66908 96 66928
rect 215136 66908 215232 66928
rect 0 66464 96 66484
rect 215136 66464 215232 66484
rect 0 66424 117 66464
rect 215115 66424 215232 66464
rect 0 66404 96 66424
rect 215136 66404 215232 66424
rect 0 65960 96 65980
rect 215136 65960 215232 65980
rect 0 65920 117 65960
rect 215115 65920 215232 65960
rect 0 65900 96 65920
rect 215136 65900 215232 65920
rect 0 65456 96 65476
rect 215136 65456 215232 65476
rect 0 65416 117 65456
rect 215115 65416 215232 65456
rect 0 65396 96 65416
rect 215136 65396 215232 65416
rect 0 64952 96 64972
rect 215136 64952 215232 64972
rect 0 64912 117 64952
rect 215115 64912 215232 64952
rect 0 64892 96 64912
rect 215136 64892 215232 64912
rect 0 64448 96 64468
rect 215136 64448 215232 64468
rect 0 64408 117 64448
rect 215115 64408 215232 64448
rect 0 64388 96 64408
rect 215136 64388 215232 64408
rect 0 63944 96 63964
rect 215136 63944 215232 63964
rect 0 63904 117 63944
rect 215115 63904 215232 63944
rect 0 63884 96 63904
rect 215136 63884 215232 63904
rect 0 63440 96 63460
rect 215136 63440 215232 63460
rect 0 63400 117 63440
rect 215115 63400 215232 63440
rect 0 63380 96 63400
rect 215136 63380 215232 63400
rect 0 62936 96 62956
rect 215136 62936 215232 62956
rect 0 62896 117 62936
rect 215115 62896 215232 62936
rect 0 62876 96 62896
rect 215136 62876 215232 62896
rect 0 62432 96 62452
rect 215136 62432 215232 62452
rect 0 62392 117 62432
rect 215115 62392 215232 62432
rect 0 62372 96 62392
rect 215136 62372 215232 62392
rect 0 61928 96 61948
rect 215136 61928 215232 61948
rect 0 61888 117 61928
rect 215115 61888 215232 61928
rect 0 61868 96 61888
rect 215136 61868 215232 61888
rect 0 61424 96 61444
rect 215136 61424 215232 61444
rect 0 61384 117 61424
rect 215115 61384 215232 61424
rect 0 61364 96 61384
rect 215136 61364 215232 61384
rect 0 60920 96 60940
rect 215136 60920 215232 60940
rect 0 60880 117 60920
rect 215115 60880 215232 60920
rect 0 60860 96 60880
rect 215136 60860 215232 60880
rect 0 60416 96 60436
rect 215136 60416 215232 60436
rect 0 60376 117 60416
rect 215115 60376 215232 60416
rect 0 60356 96 60376
rect 215136 60356 215232 60376
rect 0 59912 96 59932
rect 215136 59912 215232 59932
rect 0 59872 117 59912
rect 215115 59872 215232 59912
rect 0 59852 96 59872
rect 215136 59852 215232 59872
rect 0 59408 96 59428
rect 215136 59408 215232 59428
rect 0 59368 117 59408
rect 215115 59368 215232 59408
rect 0 59348 96 59368
rect 215136 59348 215232 59368
rect 0 58904 96 58924
rect 215136 58904 215232 58924
rect 0 58864 117 58904
rect 215115 58864 215232 58904
rect 0 58844 96 58864
rect 215136 58844 215232 58864
rect 0 58400 96 58420
rect 215136 58400 215232 58420
rect 0 58360 117 58400
rect 215115 58360 215232 58400
rect 0 58340 96 58360
rect 215136 58340 215232 58360
rect 0 57896 96 57916
rect 215136 57896 215232 57916
rect 0 57856 117 57896
rect 215115 57856 215232 57896
rect 0 57836 96 57856
rect 215136 57836 215232 57856
rect 0 57392 96 57412
rect 215136 57392 215232 57412
rect 0 57352 117 57392
rect 215115 57352 215232 57392
rect 0 57332 96 57352
rect 215136 57332 215232 57352
rect 0 51680 96 51700
rect 0 51640 117 51680
rect 0 51620 96 51640
rect 0 51176 96 51196
rect 0 51136 117 51176
rect 0 51116 96 51136
rect 0 50672 96 50692
rect 0 50632 117 50672
rect 0 50612 96 50632
rect 0 50168 96 50188
rect 0 50128 117 50168
rect 0 50108 96 50128
rect 0 49664 96 49684
rect 0 49624 117 49664
rect 0 49604 96 49624
rect 0 49160 96 49180
rect 0 49120 117 49160
rect 0 49100 96 49120
rect 0 48656 96 48676
rect 0 48616 117 48656
rect 0 48596 96 48616
rect 0 48152 96 48172
rect 0 48112 117 48152
rect 0 48092 96 48112
rect 0 47648 96 47668
rect 0 47608 117 47648
rect 0 47588 96 47608
rect 0 47144 96 47164
rect 0 47104 117 47144
rect 0 47084 96 47104
rect 0 46640 96 46660
rect 0 46600 117 46640
rect 0 46580 96 46600
rect 0 46136 96 46156
rect 0 46096 117 46136
rect 0 46076 96 46096
rect 0 45632 96 45652
rect 0 45592 117 45632
rect 0 45572 96 45592
rect 0 45128 96 45148
rect 0 45088 117 45128
rect 0 45068 96 45088
rect 0 44624 96 44644
rect 0 44584 117 44624
rect 0 44564 96 44584
rect 0 44120 96 44140
rect 0 44080 117 44120
rect 0 44060 96 44080
rect 0 43616 96 43636
rect 0 43576 117 43616
rect 0 43556 96 43576
rect 0 43112 96 43132
rect 0 43072 117 43112
rect 0 43052 96 43072
rect 0 42608 96 42628
rect 0 42568 117 42608
rect 0 42548 96 42568
rect 0 42104 96 42124
rect 0 42064 117 42104
rect 0 42044 96 42064
rect 0 41600 96 41620
rect 0 41560 117 41600
rect 0 41540 96 41560
rect 0 41096 96 41116
rect 0 41056 117 41096
rect 0 41036 96 41056
rect 0 40592 96 40612
rect 0 40552 117 40592
rect 0 40532 96 40552
rect 0 40088 96 40108
rect 0 40048 117 40088
rect 0 40028 96 40048
rect 0 39584 96 39604
rect 0 39544 117 39584
rect 0 39524 96 39544
rect 0 39080 96 39100
rect 0 39040 117 39080
rect 0 39020 96 39040
rect 0 38576 96 38596
rect 0 38536 117 38576
rect 0 38516 96 38536
rect 0 38072 96 38092
rect 0 38032 117 38072
rect 0 38012 96 38032
rect 0 37568 96 37588
rect 0 37528 117 37568
rect 0 37508 96 37528
rect 0 37064 96 37084
rect 0 37024 117 37064
rect 0 37004 96 37024
rect 0 36560 96 36580
rect 0 36520 117 36560
rect 0 36500 96 36520
rect 0 36056 96 36076
rect 0 36016 117 36056
rect 0 35996 96 36016
rect 0 35552 96 35572
rect 215136 35552 215232 35572
rect 0 35512 117 35552
rect 215115 35512 215232 35552
rect 0 35492 96 35512
rect 215136 35492 215232 35512
rect 0 35048 96 35068
rect 215136 35048 215232 35068
rect 0 35008 117 35048
rect 215115 35008 215232 35048
rect 0 34988 96 35008
rect 215136 34988 215232 35008
rect 0 34544 96 34564
rect 215136 34544 215232 34564
rect 0 34504 117 34544
rect 215115 34504 215232 34544
rect 0 34484 96 34504
rect 215136 34484 215232 34504
rect 0 34040 96 34060
rect 215136 34040 215232 34060
rect 0 34000 117 34040
rect 215115 34000 215232 34040
rect 0 33980 96 34000
rect 215136 33980 215232 34000
rect 0 33536 96 33556
rect 215136 33536 215232 33556
rect 0 33496 117 33536
rect 215115 33496 215232 33536
rect 0 33476 96 33496
rect 215136 33476 215232 33496
rect 0 33032 96 33052
rect 215136 33032 215232 33052
rect 0 32992 117 33032
rect 215115 32992 215232 33032
rect 0 32972 96 32992
rect 215136 32972 215232 32992
rect 0 32528 96 32548
rect 215136 32528 215232 32548
rect 0 32488 117 32528
rect 215115 32488 215232 32528
rect 0 32468 96 32488
rect 215136 32468 215232 32488
rect 0 32024 96 32044
rect 215136 32024 215232 32044
rect 0 31984 117 32024
rect 215115 31984 215232 32024
rect 0 31964 96 31984
rect 215136 31964 215232 31984
rect 0 31520 96 31540
rect 215136 31520 215232 31540
rect 0 31480 117 31520
rect 215115 31480 215232 31520
rect 0 31460 96 31480
rect 215136 31460 215232 31480
rect 0 31016 96 31036
rect 215136 31016 215232 31036
rect 0 30976 117 31016
rect 215115 30976 215232 31016
rect 0 30956 96 30976
rect 215136 30956 215232 30976
rect 0 30512 96 30532
rect 215136 30512 215232 30532
rect 0 30472 117 30512
rect 215115 30472 215232 30512
rect 0 30452 96 30472
rect 215136 30452 215232 30472
rect 0 30008 96 30028
rect 215136 30008 215232 30028
rect 0 29968 117 30008
rect 215115 29968 215232 30008
rect 0 29948 96 29968
rect 215136 29948 215232 29968
rect 0 29504 96 29524
rect 215136 29504 215232 29524
rect 0 29464 117 29504
rect 215115 29464 215232 29504
rect 0 29444 96 29464
rect 215136 29444 215232 29464
rect 0 29000 96 29020
rect 215136 29000 215232 29020
rect 0 28960 117 29000
rect 215115 28960 215232 29000
rect 0 28940 96 28960
rect 215136 28940 215232 28960
rect 0 28496 96 28516
rect 215136 28496 215232 28516
rect 0 28456 117 28496
rect 215115 28456 215232 28496
rect 0 28436 96 28456
rect 215136 28436 215232 28456
rect 0 27992 96 28012
rect 215136 27992 215232 28012
rect 0 27952 117 27992
rect 215115 27952 215232 27992
rect 0 27932 96 27952
rect 215136 27932 215232 27952
rect 0 27488 96 27508
rect 215136 27488 215232 27508
rect 0 27448 117 27488
rect 215115 27448 215232 27488
rect 0 27428 96 27448
rect 215136 27428 215232 27448
rect 0 26984 96 27004
rect 215136 26984 215232 27004
rect 0 26944 117 26984
rect 215115 26944 215232 26984
rect 0 26924 96 26944
rect 215136 26924 215232 26944
rect 0 26480 96 26500
rect 215136 26480 215232 26500
rect 0 26440 117 26480
rect 215115 26440 215232 26480
rect 0 26420 96 26440
rect 215136 26420 215232 26440
rect 0 25976 96 25996
rect 215136 25976 215232 25996
rect 0 25936 117 25976
rect 215115 25936 215232 25976
rect 0 25916 96 25936
rect 215136 25916 215232 25936
rect 0 25472 96 25492
rect 215136 25472 215232 25492
rect 0 25432 117 25472
rect 215115 25432 215232 25472
rect 0 25412 96 25432
rect 215136 25412 215232 25432
rect 0 24968 96 24988
rect 215136 24968 215232 24988
rect 0 24928 117 24968
rect 215115 24928 215232 24968
rect 0 24908 96 24928
rect 215136 24908 215232 24928
rect 0 24464 96 24484
rect 215136 24464 215232 24484
rect 0 24424 117 24464
rect 215115 24424 215232 24464
rect 0 24404 96 24424
rect 215136 24404 215232 24424
rect 0 23960 96 23980
rect 215136 23960 215232 23980
rect 0 23920 117 23960
rect 215115 23920 215232 23960
rect 0 23900 96 23920
rect 215136 23900 215232 23920
rect 0 23456 96 23476
rect 215136 23456 215232 23476
rect 0 23416 117 23456
rect 215115 23416 215232 23456
rect 0 23396 96 23416
rect 215136 23396 215232 23416
rect 0 22952 96 22972
rect 215136 22952 215232 22972
rect 0 22912 117 22952
rect 215115 22912 215232 22952
rect 0 22892 96 22912
rect 215136 22892 215232 22912
rect 0 22448 96 22468
rect 215136 22448 215232 22468
rect 0 22408 117 22448
rect 215115 22408 215232 22448
rect 0 22388 96 22408
rect 215136 22388 215232 22408
rect 0 21944 96 21964
rect 215136 21944 215232 21964
rect 0 21904 117 21944
rect 215115 21904 215232 21944
rect 0 21884 96 21904
rect 215136 21884 215232 21904
rect 0 21440 96 21460
rect 215136 21440 215232 21460
rect 0 21400 117 21440
rect 215115 21400 215232 21440
rect 0 21380 96 21400
rect 215136 21380 215232 21400
rect 0 20936 96 20956
rect 215136 20936 215232 20956
rect 0 20896 117 20936
rect 215115 20896 215232 20936
rect 0 20876 96 20896
rect 215136 20876 215232 20896
rect 0 20432 96 20452
rect 215136 20432 215232 20452
rect 0 20392 117 20432
rect 215115 20392 215232 20432
rect 0 20372 96 20392
rect 215136 20372 215232 20392
rect 0 19928 96 19948
rect 215136 19928 215232 19948
rect 0 19888 117 19928
rect 215115 19888 215232 19928
rect 0 19868 96 19888
rect 215136 19868 215232 19888
rect 0 19424 96 19444
rect 215136 19424 215232 19444
rect 0 19384 117 19424
rect 215115 19384 215232 19424
rect 0 19364 96 19384
rect 215136 19364 215232 19384
rect 0 18920 96 18940
rect 215136 18920 215232 18940
rect 0 18880 117 18920
rect 215115 18880 215232 18920
rect 0 18860 96 18880
rect 215136 18860 215232 18880
rect 0 18416 96 18436
rect 215136 18416 215232 18436
rect 0 18376 117 18416
rect 215115 18376 215232 18416
rect 0 18356 96 18376
rect 215136 18356 215232 18376
rect 0 17912 96 17932
rect 215136 17912 215232 17932
rect 0 17872 117 17912
rect 215115 17872 215232 17912
rect 0 17852 96 17872
rect 215136 17852 215232 17872
rect 0 17408 96 17428
rect 215136 17408 215232 17428
rect 0 17368 117 17408
rect 215115 17368 215232 17408
rect 0 17348 96 17368
rect 215136 17348 215232 17368
rect 0 16904 96 16924
rect 215136 16904 215232 16924
rect 0 16864 117 16904
rect 215115 16864 215232 16904
rect 0 16844 96 16864
rect 215136 16844 215232 16864
rect 0 16400 96 16420
rect 215136 16400 215232 16420
rect 0 16360 117 16400
rect 215115 16360 215232 16400
rect 0 16340 96 16360
rect 215136 16340 215232 16360
rect 0 15896 96 15916
rect 215136 15896 215232 15916
rect 0 15856 117 15896
rect 215115 15856 215232 15896
rect 0 15836 96 15856
rect 215136 15836 215232 15856
rect 0 15392 96 15412
rect 215136 15392 215232 15412
rect 0 15352 117 15392
rect 215115 15352 215232 15392
rect 0 15332 96 15352
rect 215136 15332 215232 15352
rect 0 14888 96 14908
rect 215136 14888 215232 14908
rect 0 14848 117 14888
rect 215115 14848 215232 14888
rect 0 14828 96 14848
rect 215136 14828 215232 14848
rect 0 14384 96 14404
rect 215136 14384 215232 14404
rect 0 14344 117 14384
rect 215115 14344 215232 14384
rect 0 14324 96 14344
rect 215136 14324 215232 14344
rect 0 11360 96 11380
rect 0 11320 117 11360
rect 0 11300 96 11320
rect 0 11024 96 11044
rect 0 10984 117 11024
rect 0 10964 96 10984
rect 0 10688 96 10708
rect 0 10648 117 10688
rect 0 10628 96 10648
rect 0 10352 96 10372
rect 0 10312 117 10352
rect 0 10292 96 10312
rect 0 10016 96 10036
rect 0 9976 117 10016
rect 0 9956 96 9976
rect 0 9680 96 9700
rect 0 9640 117 9680
rect 0 9620 96 9640
rect 0 9344 96 9364
rect 0 9304 117 9344
rect 0 9284 96 9304
rect 0 9008 96 9028
rect 0 8968 117 9008
rect 0 8948 96 8968
rect 0 8672 96 8692
rect 0 8632 117 8672
rect 0 8612 96 8632
rect 0 8336 96 8356
rect 0 8296 117 8336
rect 0 8276 96 8296
rect 0 8000 96 8020
rect 0 7960 117 8000
rect 0 7940 96 7960
rect 0 7664 96 7684
rect 0 7624 117 7664
rect 0 7604 96 7624
rect 0 7328 96 7348
rect 0 7288 117 7328
rect 0 7268 96 7288
rect 0 6992 96 7012
rect 0 6952 117 6992
rect 0 6932 96 6952
rect 0 6656 96 6676
rect 0 6616 117 6656
rect 0 6596 96 6616
rect 0 6320 96 6340
rect 0 6280 117 6320
rect 0 6260 96 6280
rect 0 5984 96 6004
rect 0 5944 117 5984
rect 0 5924 96 5944
rect 0 5648 96 5668
rect 0 5608 117 5648
rect 0 5588 96 5608
rect 0 5312 96 5332
rect 0 5272 117 5312
rect 0 5252 96 5272
rect 0 4976 96 4996
rect 0 4936 117 4976
rect 0 4916 96 4936
rect 0 4640 96 4660
rect 0 4600 117 4640
rect 0 4580 96 4600
rect 0 4304 96 4324
rect 0 4264 117 4304
rect 0 4244 96 4264
rect 0 3968 96 3988
rect 0 3928 117 3968
rect 0 3908 96 3928
rect 0 3632 96 3652
rect 0 3592 117 3632
rect 0 3572 96 3592
rect 0 3296 96 3316
rect 0 3256 117 3296
rect 0 3236 96 3256
rect 0 2960 96 2980
rect 0 2920 117 2960
rect 0 2900 96 2920
rect 0 2624 96 2644
rect 0 2584 117 2624
rect 0 2564 96 2584
rect 0 2288 96 2308
rect 0 2248 117 2288
rect 0 2228 96 2248
rect 0 1952 96 1972
rect 0 1912 117 1952
rect 0 1892 96 1912
rect 0 1616 96 1636
rect 0 1576 117 1616
rect 0 1556 96 1576
rect 0 1280 96 1300
rect 0 1240 117 1280
rect 0 1220 96 1240
rect 0 944 96 964
rect 0 904 117 944
rect 0 884 96 904
rect 38390 736 38399 776
rect 38439 736 81407 776
rect 81447 736 124415 776
rect 124455 736 167385 776
rect 167425 736 194649 776
rect 194689 736 194698 776
rect 1123 148 1132 188
rect 1172 148 1181 188
rect 1132 104 1172 148
rect 1132 64 38380 104
rect 38420 64 38429 104
<< metal6 >>
rect 3748 840 4188 366408
rect 4988 840 5428 366408
rect 18868 840 19308 366408
rect 25252 840 25692 366408
rect 26492 840 26932 366408
rect 40372 840 40812 366408
rect 41612 840 42052 366408
rect 55492 840 55932 366408
rect 56732 840 57172 366408
rect 68260 840 68700 366408
rect 69500 840 69940 366408
rect 83380 840 83820 366408
rect 84620 840 85060 366408
rect 98500 840 98940 366408
rect 99740 840 100180 366408
rect 111268 840 111708 366408
rect 112508 840 112948 366408
rect 126388 840 126828 366408
rect 127628 840 128068 366408
rect 141508 840 141948 366408
rect 142748 840 143188 366408
rect 154276 840 154716 366408
rect 155516 840 155956 366408
rect 169396 840 169836 366408
rect 170636 840 171076 366408
rect 184516 840 184956 366408
rect 185756 840 186196 366408
rect 197284 840 197724 366408
rect 198524 840 198964 366408
rect 212404 840 212844 366408
use NW_term  Tile_X0Y0_NW_term
timestamp 0
transform 1 0 96 0 1 355656
box 0 0 1 1
use W_TT_IF  Tile_X0Y1_W_TT_IF
timestamp 0
transform 1 0 96 0 1 312648
box 0 0 1 1
use W_TT_IF  Tile_X0Y2_W_TT_IF
timestamp 0
transform 1 0 96 0 1 269640
box 0 0 1 1
use W_TT_IF  Tile_X0Y3_W_TT_IF
timestamp 0
transform 1 0 96 0 1 226632
box 0 0 1 1
use W_TT_IF  Tile_X0Y4_W_TT_IF
timestamp 0
transform 1 0 96 0 1 183624
box 0 0 1 1
use W_TT_IF  Tile_X0Y5_W_TT_IF
timestamp 0
transform 1 0 96 0 1 140616
box 0 0 1 1
use W_TT_IF  Tile_X0Y6_W_TT_IF
timestamp 0
transform 1 0 96 0 1 97608
box 0 0 1 1
use W_TT_IF  Tile_X0Y7_W_TT_IF
timestamp 0
transform 1 0 96 0 1 54600
box 0 0 1 1
use W_TT_IF  Tile_X0Y8_W_TT_IF
timestamp 0
transform 1 0 96 0 1 11592
box 0 0 1 1
use SW_term  Tile_X0Y9_SW_term
timestamp 0
transform 1 0 96 0 1 840
box 0 0 1 1
use N_IO4  Tile_X1Y0_N_IO4
timestamp 0
transform 1 0 21600 0 1 355656
box 0 0 1 1
use LUT4AB  Tile_X1Y1_LUT4AB
timestamp 0
transform 1 0 21600 0 1 312648
box 0 0 1 1
use LUT4AB  Tile_X1Y2_LUT4AB
timestamp 0
transform 1 0 21600 0 1 269640
box 0 0 1 1
use LUT4AB  Tile_X1Y3_LUT4AB
timestamp 0
transform 1 0 21600 0 1 226632
box 0 0 1 1
use LUT4AB  Tile_X1Y4_LUT4AB
timestamp 0
transform 1 0 21600 0 1 183624
box 0 0 1 1
use LUT4AB  Tile_X1Y5_LUT4AB
timestamp 0
transform 1 0 21600 0 1 140616
box 0 0 1 1
use LUT4AB  Tile_X1Y6_LUT4AB
timestamp 0
transform 1 0 21600 0 1 97608
box 0 0 1 1
use LUT4AB  Tile_X1Y7_LUT4AB
timestamp 0
transform 1 0 21600 0 1 54600
box 0 0 1 1
use LUT4AB  Tile_X1Y8_LUT4AB
timestamp 0
transform 1 0 21600 0 1 11592
box 0 0 1 1
use S_IO4  Tile_X1Y9_S_IO4
timestamp 0
transform 1 0 21600 0 1 840
box 0 0 1 1
use N_IO4  Tile_X2Y0_N_IO4
timestamp 0
transform 1 0 64608 0 1 355656
box 0 0 1 1
use LUT4AB  Tile_X2Y1_LUT4AB
timestamp 0
transform 1 0 64608 0 1 312648
box 0 0 1 1
use LUT4AB  Tile_X2Y2_LUT4AB
timestamp 0
transform 1 0 64608 0 1 269640
box 0 0 1 1
use LUT4AB  Tile_X2Y3_LUT4AB
timestamp 0
transform 1 0 64608 0 1 226632
box 0 0 1 1
use LUT4AB  Tile_X2Y4_LUT4AB
timestamp 0
transform 1 0 64608 0 1 183624
box 0 0 1 1
use LUT4AB  Tile_X2Y5_LUT4AB
timestamp 0
transform 1 0 64608 0 1 140616
box 0 0 1 1
use LUT4AB  Tile_X2Y6_LUT4AB
timestamp 0
transform 1 0 64608 0 1 97608
box 0 0 1 1
use LUT4AB  Tile_X2Y7_LUT4AB
timestamp 0
transform 1 0 64608 0 1 54600
box 0 0 1 1
use LUT4AB  Tile_X2Y8_LUT4AB
timestamp 0
transform 1 0 64608 0 1 11592
box 0 0 1 1
use S_IO4  Tile_X2Y9_S_IO4
timestamp 0
transform 1 0 64608 0 1 840
box 0 0 1 1
use N_IO4  Tile_X3Y0_N_IO4
timestamp 0
transform 1 0 107616 0 1 355656
box 0 0 1 1
use LUT4AB  Tile_X3Y1_LUT4AB
timestamp 0
transform 1 0 107616 0 1 312648
box 0 0 1 1
use LUT4AB  Tile_X3Y2_LUT4AB
timestamp 0
transform 1 0 107616 0 1 269640
box 0 0 1 1
use LUT4AB  Tile_X3Y3_LUT4AB
timestamp 0
transform 1 0 107616 0 1 226632
box 0 0 1 1
use LUT4AB  Tile_X3Y4_LUT4AB
timestamp 0
transform 1 0 107616 0 1 183624
box 0 0 1 1
use LUT4AB  Tile_X3Y5_LUT4AB
timestamp 0
transform 1 0 107616 0 1 140616
box 0 0 1 1
use LUT4AB  Tile_X3Y6_LUT4AB
timestamp 0
transform 1 0 107616 0 1 97608
box 0 0 1 1
use LUT4AB  Tile_X3Y7_LUT4AB
timestamp 0
transform 1 0 107616 0 1 54600
box 0 0 1 1
use LUT4AB  Tile_X3Y8_LUT4AB
timestamp 0
transform 1 0 107616 0 1 11592
box 0 0 1 1
use S_IO4  Tile_X3Y9_S_IO4
timestamp 0
transform 1 0 107616 0 1 840
box 0 0 1 1
use N_IO4  Tile_X4Y0_N_IO4
timestamp 0
transform 1 0 150624 0 1 355656
box 0 0 1 1
use LUT4AB  Tile_X4Y1_LUT4AB
timestamp 0
transform 1 0 150624 0 1 312648
box 0 0 1 1
use LUT4AB  Tile_X4Y2_LUT4AB
timestamp 0
transform 1 0 150624 0 1 269640
box 0 0 1 1
use LUT4AB  Tile_X4Y3_LUT4AB
timestamp 0
transform 1 0 150624 0 1 226632
box 0 0 1 1
use LUT4AB  Tile_X4Y4_LUT4AB
timestamp 0
transform 1 0 150624 0 1 183624
box 0 0 1 1
use LUT4AB  Tile_X4Y5_LUT4AB
timestamp 0
transform 1 0 150624 0 1 140616
box 0 0 1 1
use LUT4AB  Tile_X4Y6_LUT4AB
timestamp 0
transform 1 0 150624 0 1 97608
box 0 0 1 1
use LUT4AB  Tile_X4Y7_LUT4AB
timestamp 0
transform 1 0 150624 0 1 54600
box 0 0 1 1
use LUT4AB  Tile_X4Y8_LUT4AB
timestamp 0
transform 1 0 150624 0 1 11592
box 0 0 1 1
use S_IO4  Tile_X4Y9_S_IO4
timestamp 0
transform 1 0 150624 0 1 840
box 0 0 1 1
use NE_term  Tile_X5Y0_NE_term
timestamp 0
transform 1 0 193632 0 1 355656
box 0 0 1 1
use IHP_SRAM  Tile_X5Y1_IHP_SRAM
timestamp 0
transform 1 0 193632 0 1 269640
box 0 0 1 1
use E_TT_IF  Tile_X5Y3_E_TT_IF
timestamp 0
transform 1 0 193632 0 1 226632
box 0 0 1 1
use E_TT_IF  Tile_X5Y4_E_TT_IF
timestamp 0
transform 1 0 193632 0 1 183624
box 0 0 1 1
use E_TT_IF  Tile_X5Y5_E_TT_IF
timestamp 0
transform 1 0 193632 0 1 140616
box 0 0 1 1
use E_TT_IF  Tile_X5Y6_E_TT_IF
timestamp 0
transform 1 0 193632 0 1 97608
box 0 0 1 1
use E_TT_IF  Tile_X5Y7_E_TT_IF
timestamp 0
transform 1 0 193632 0 1 54600
box 0 0 1 1
use E_TT_IF  Tile_X5Y8_E_TT_IF
timestamp 0
transform 1 0 193632 0 1 11592
box 0 0 1 1
use SE_term  Tile_X5Y9_SE_term
timestamp 0
transform 1 0 193632 0 1 840
box 0 0 1 1
<< labels >>
flabel metal3 s 0 355700 96 355780 0 FreeSans 320 0 0 0 FrameData[0]
port 0 nsew signal input
flabel metal3 s 0 253052 96 253132 0 FreeSans 320 0 0 0 FrameData[100]
port 1 nsew signal input
flabel metal3 s 0 253556 96 253636 0 FreeSans 320 0 0 0 FrameData[101]
port 2 nsew signal input
flabel metal3 s 0 254060 96 254140 0 FreeSans 320 0 0 0 FrameData[102]
port 3 nsew signal input
flabel metal3 s 0 254564 96 254644 0 FreeSans 320 0 0 0 FrameData[103]
port 4 nsew signal input
flabel metal3 s 0 255068 96 255148 0 FreeSans 320 0 0 0 FrameData[104]
port 5 nsew signal input
flabel metal3 s 0 255572 96 255652 0 FreeSans 320 0 0 0 FrameData[105]
port 6 nsew signal input
flabel metal3 s 0 256076 96 256156 0 FreeSans 320 0 0 0 FrameData[106]
port 7 nsew signal input
flabel metal3 s 0 256580 96 256660 0 FreeSans 320 0 0 0 FrameData[107]
port 8 nsew signal input
flabel metal3 s 0 257084 96 257164 0 FreeSans 320 0 0 0 FrameData[108]
port 9 nsew signal input
flabel metal3 s 0 257588 96 257668 0 FreeSans 320 0 0 0 FrameData[109]
port 10 nsew signal input
flabel metal3 s 0 359060 96 359140 0 FreeSans 320 0 0 0 FrameData[10]
port 11 nsew signal input
flabel metal3 s 0 258092 96 258172 0 FreeSans 320 0 0 0 FrameData[110]
port 12 nsew signal input
flabel metal3 s 0 258596 96 258676 0 FreeSans 320 0 0 0 FrameData[111]
port 13 nsew signal input
flabel metal3 s 0 259100 96 259180 0 FreeSans 320 0 0 0 FrameData[112]
port 14 nsew signal input
flabel metal3 s 0 259604 96 259684 0 FreeSans 320 0 0 0 FrameData[113]
port 15 nsew signal input
flabel metal3 s 0 260108 96 260188 0 FreeSans 320 0 0 0 FrameData[114]
port 16 nsew signal input
flabel metal3 s 0 260612 96 260692 0 FreeSans 320 0 0 0 FrameData[115]
port 17 nsew signal input
flabel metal3 s 0 261116 96 261196 0 FreeSans 320 0 0 0 FrameData[116]
port 18 nsew signal input
flabel metal3 s 0 261620 96 261700 0 FreeSans 320 0 0 0 FrameData[117]
port 19 nsew signal input
flabel metal3 s 0 262124 96 262204 0 FreeSans 320 0 0 0 FrameData[118]
port 20 nsew signal input
flabel metal3 s 0 262628 96 262708 0 FreeSans 320 0 0 0 FrameData[119]
port 21 nsew signal input
flabel metal3 s 0 359396 96 359476 0 FreeSans 320 0 0 0 FrameData[11]
port 22 nsew signal input
flabel metal3 s 0 263132 96 263212 0 FreeSans 320 0 0 0 FrameData[120]
port 23 nsew signal input
flabel metal3 s 0 263636 96 263716 0 FreeSans 320 0 0 0 FrameData[121]
port 24 nsew signal input
flabel metal3 s 0 264140 96 264220 0 FreeSans 320 0 0 0 FrameData[122]
port 25 nsew signal input
flabel metal3 s 0 264644 96 264724 0 FreeSans 320 0 0 0 FrameData[123]
port 26 nsew signal input
flabel metal3 s 0 265148 96 265228 0 FreeSans 320 0 0 0 FrameData[124]
port 27 nsew signal input
flabel metal3 s 0 265652 96 265732 0 FreeSans 320 0 0 0 FrameData[125]
port 28 nsew signal input
flabel metal3 s 0 266156 96 266236 0 FreeSans 320 0 0 0 FrameData[126]
port 29 nsew signal input
flabel metal3 s 0 266660 96 266740 0 FreeSans 320 0 0 0 FrameData[127]
port 30 nsew signal input
flabel metal3 s 0 208028 96 208108 0 FreeSans 320 0 0 0 FrameData[128]
port 31 nsew signal input
flabel metal3 s 0 208532 96 208612 0 FreeSans 320 0 0 0 FrameData[129]
port 32 nsew signal input
flabel metal3 s 0 359732 96 359812 0 FreeSans 320 0 0 0 FrameData[12]
port 33 nsew signal input
flabel metal3 s 0 209036 96 209116 0 FreeSans 320 0 0 0 FrameData[130]
port 34 nsew signal input
flabel metal3 s 0 209540 96 209620 0 FreeSans 320 0 0 0 FrameData[131]
port 35 nsew signal input
flabel metal3 s 0 210044 96 210124 0 FreeSans 320 0 0 0 FrameData[132]
port 36 nsew signal input
flabel metal3 s 0 210548 96 210628 0 FreeSans 320 0 0 0 FrameData[133]
port 37 nsew signal input
flabel metal3 s 0 211052 96 211132 0 FreeSans 320 0 0 0 FrameData[134]
port 38 nsew signal input
flabel metal3 s 0 211556 96 211636 0 FreeSans 320 0 0 0 FrameData[135]
port 39 nsew signal input
flabel metal3 s 0 212060 96 212140 0 FreeSans 320 0 0 0 FrameData[136]
port 40 nsew signal input
flabel metal3 s 0 212564 96 212644 0 FreeSans 320 0 0 0 FrameData[137]
port 41 nsew signal input
flabel metal3 s 0 213068 96 213148 0 FreeSans 320 0 0 0 FrameData[138]
port 42 nsew signal input
flabel metal3 s 0 213572 96 213652 0 FreeSans 320 0 0 0 FrameData[139]
port 43 nsew signal input
flabel metal3 s 0 360068 96 360148 0 FreeSans 320 0 0 0 FrameData[13]
port 44 nsew signal input
flabel metal3 s 0 214076 96 214156 0 FreeSans 320 0 0 0 FrameData[140]
port 45 nsew signal input
flabel metal3 s 0 214580 96 214660 0 FreeSans 320 0 0 0 FrameData[141]
port 46 nsew signal input
flabel metal3 s 0 215084 96 215164 0 FreeSans 320 0 0 0 FrameData[142]
port 47 nsew signal input
flabel metal3 s 0 215588 96 215668 0 FreeSans 320 0 0 0 FrameData[143]
port 48 nsew signal input
flabel metal3 s 0 216092 96 216172 0 FreeSans 320 0 0 0 FrameData[144]
port 49 nsew signal input
flabel metal3 s 0 216596 96 216676 0 FreeSans 320 0 0 0 FrameData[145]
port 50 nsew signal input
flabel metal3 s 0 217100 96 217180 0 FreeSans 320 0 0 0 FrameData[146]
port 51 nsew signal input
flabel metal3 s 0 217604 96 217684 0 FreeSans 320 0 0 0 FrameData[147]
port 52 nsew signal input
flabel metal3 s 0 218108 96 218188 0 FreeSans 320 0 0 0 FrameData[148]
port 53 nsew signal input
flabel metal3 s 0 218612 96 218692 0 FreeSans 320 0 0 0 FrameData[149]
port 54 nsew signal input
flabel metal3 s 0 360404 96 360484 0 FreeSans 320 0 0 0 FrameData[14]
port 55 nsew signal input
flabel metal3 s 0 219116 96 219196 0 FreeSans 320 0 0 0 FrameData[150]
port 56 nsew signal input
flabel metal3 s 0 219620 96 219700 0 FreeSans 320 0 0 0 FrameData[151]
port 57 nsew signal input
flabel metal3 s 0 220124 96 220204 0 FreeSans 320 0 0 0 FrameData[152]
port 58 nsew signal input
flabel metal3 s 0 220628 96 220708 0 FreeSans 320 0 0 0 FrameData[153]
port 59 nsew signal input
flabel metal3 s 0 221132 96 221212 0 FreeSans 320 0 0 0 FrameData[154]
port 60 nsew signal input
flabel metal3 s 0 221636 96 221716 0 FreeSans 320 0 0 0 FrameData[155]
port 61 nsew signal input
flabel metal3 s 0 222140 96 222220 0 FreeSans 320 0 0 0 FrameData[156]
port 62 nsew signal input
flabel metal3 s 0 222644 96 222724 0 FreeSans 320 0 0 0 FrameData[157]
port 63 nsew signal input
flabel metal3 s 0 223148 96 223228 0 FreeSans 320 0 0 0 FrameData[158]
port 64 nsew signal input
flabel metal3 s 0 223652 96 223732 0 FreeSans 320 0 0 0 FrameData[159]
port 65 nsew signal input
flabel metal3 s 0 360740 96 360820 0 FreeSans 320 0 0 0 FrameData[15]
port 66 nsew signal input
flabel metal3 s 0 165020 96 165100 0 FreeSans 320 0 0 0 FrameData[160]
port 67 nsew signal input
flabel metal3 s 0 165524 96 165604 0 FreeSans 320 0 0 0 FrameData[161]
port 68 nsew signal input
flabel metal3 s 0 166028 96 166108 0 FreeSans 320 0 0 0 FrameData[162]
port 69 nsew signal input
flabel metal3 s 0 166532 96 166612 0 FreeSans 320 0 0 0 FrameData[163]
port 70 nsew signal input
flabel metal3 s 0 167036 96 167116 0 FreeSans 320 0 0 0 FrameData[164]
port 71 nsew signal input
flabel metal3 s 0 167540 96 167620 0 FreeSans 320 0 0 0 FrameData[165]
port 72 nsew signal input
flabel metal3 s 0 168044 96 168124 0 FreeSans 320 0 0 0 FrameData[166]
port 73 nsew signal input
flabel metal3 s 0 168548 96 168628 0 FreeSans 320 0 0 0 FrameData[167]
port 74 nsew signal input
flabel metal3 s 0 169052 96 169132 0 FreeSans 320 0 0 0 FrameData[168]
port 75 nsew signal input
flabel metal3 s 0 169556 96 169636 0 FreeSans 320 0 0 0 FrameData[169]
port 76 nsew signal input
flabel metal3 s 0 361076 96 361156 0 FreeSans 320 0 0 0 FrameData[16]
port 77 nsew signal input
flabel metal3 s 0 170060 96 170140 0 FreeSans 320 0 0 0 FrameData[170]
port 78 nsew signal input
flabel metal3 s 0 170564 96 170644 0 FreeSans 320 0 0 0 FrameData[171]
port 79 nsew signal input
flabel metal3 s 0 171068 96 171148 0 FreeSans 320 0 0 0 FrameData[172]
port 80 nsew signal input
flabel metal3 s 0 171572 96 171652 0 FreeSans 320 0 0 0 FrameData[173]
port 81 nsew signal input
flabel metal3 s 0 172076 96 172156 0 FreeSans 320 0 0 0 FrameData[174]
port 82 nsew signal input
flabel metal3 s 0 172580 96 172660 0 FreeSans 320 0 0 0 FrameData[175]
port 83 nsew signal input
flabel metal3 s 0 173084 96 173164 0 FreeSans 320 0 0 0 FrameData[176]
port 84 nsew signal input
flabel metal3 s 0 173588 96 173668 0 FreeSans 320 0 0 0 FrameData[177]
port 85 nsew signal input
flabel metal3 s 0 174092 96 174172 0 FreeSans 320 0 0 0 FrameData[178]
port 86 nsew signal input
flabel metal3 s 0 174596 96 174676 0 FreeSans 320 0 0 0 FrameData[179]
port 87 nsew signal input
flabel metal3 s 0 361412 96 361492 0 FreeSans 320 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s 0 175100 96 175180 0 FreeSans 320 0 0 0 FrameData[180]
port 89 nsew signal input
flabel metal3 s 0 175604 96 175684 0 FreeSans 320 0 0 0 FrameData[181]
port 90 nsew signal input
flabel metal3 s 0 176108 96 176188 0 FreeSans 320 0 0 0 FrameData[182]
port 91 nsew signal input
flabel metal3 s 0 176612 96 176692 0 FreeSans 320 0 0 0 FrameData[183]
port 92 nsew signal input
flabel metal3 s 0 177116 96 177196 0 FreeSans 320 0 0 0 FrameData[184]
port 93 nsew signal input
flabel metal3 s 0 177620 96 177700 0 FreeSans 320 0 0 0 FrameData[185]
port 94 nsew signal input
flabel metal3 s 0 178124 96 178204 0 FreeSans 320 0 0 0 FrameData[186]
port 95 nsew signal input
flabel metal3 s 0 178628 96 178708 0 FreeSans 320 0 0 0 FrameData[187]
port 96 nsew signal input
flabel metal3 s 0 179132 96 179212 0 FreeSans 320 0 0 0 FrameData[188]
port 97 nsew signal input
flabel metal3 s 0 179636 96 179716 0 FreeSans 320 0 0 0 FrameData[189]
port 98 nsew signal input
flabel metal3 s 0 361748 96 361828 0 FreeSans 320 0 0 0 FrameData[18]
port 99 nsew signal input
flabel metal3 s 0 180140 96 180220 0 FreeSans 320 0 0 0 FrameData[190]
port 100 nsew signal input
flabel metal3 s 0 180644 96 180724 0 FreeSans 320 0 0 0 FrameData[191]
port 101 nsew signal input
flabel metal3 s 0 122012 96 122092 0 FreeSans 320 0 0 0 FrameData[192]
port 102 nsew signal input
flabel metal3 s 0 122516 96 122596 0 FreeSans 320 0 0 0 FrameData[193]
port 103 nsew signal input
flabel metal3 s 0 123020 96 123100 0 FreeSans 320 0 0 0 FrameData[194]
port 104 nsew signal input
flabel metal3 s 0 123524 96 123604 0 FreeSans 320 0 0 0 FrameData[195]
port 105 nsew signal input
flabel metal3 s 0 124028 96 124108 0 FreeSans 320 0 0 0 FrameData[196]
port 106 nsew signal input
flabel metal3 s 0 124532 96 124612 0 FreeSans 320 0 0 0 FrameData[197]
port 107 nsew signal input
flabel metal3 s 0 125036 96 125116 0 FreeSans 320 0 0 0 FrameData[198]
port 108 nsew signal input
flabel metal3 s 0 125540 96 125620 0 FreeSans 320 0 0 0 FrameData[199]
port 109 nsew signal input
flabel metal3 s 0 362084 96 362164 0 FreeSans 320 0 0 0 FrameData[19]
port 110 nsew signal input
flabel metal3 s 0 356036 96 356116 0 FreeSans 320 0 0 0 FrameData[1]
port 111 nsew signal input
flabel metal3 s 0 126044 96 126124 0 FreeSans 320 0 0 0 FrameData[200]
port 112 nsew signal input
flabel metal3 s 0 126548 96 126628 0 FreeSans 320 0 0 0 FrameData[201]
port 113 nsew signal input
flabel metal3 s 0 127052 96 127132 0 FreeSans 320 0 0 0 FrameData[202]
port 114 nsew signal input
flabel metal3 s 0 127556 96 127636 0 FreeSans 320 0 0 0 FrameData[203]
port 115 nsew signal input
flabel metal3 s 0 128060 96 128140 0 FreeSans 320 0 0 0 FrameData[204]
port 116 nsew signal input
flabel metal3 s 0 128564 96 128644 0 FreeSans 320 0 0 0 FrameData[205]
port 117 nsew signal input
flabel metal3 s 0 129068 96 129148 0 FreeSans 320 0 0 0 FrameData[206]
port 118 nsew signal input
flabel metal3 s 0 129572 96 129652 0 FreeSans 320 0 0 0 FrameData[207]
port 119 nsew signal input
flabel metal3 s 0 130076 96 130156 0 FreeSans 320 0 0 0 FrameData[208]
port 120 nsew signal input
flabel metal3 s 0 130580 96 130660 0 FreeSans 320 0 0 0 FrameData[209]
port 121 nsew signal input
flabel metal3 s 0 362420 96 362500 0 FreeSans 320 0 0 0 FrameData[20]
port 122 nsew signal input
flabel metal3 s 0 131084 96 131164 0 FreeSans 320 0 0 0 FrameData[210]
port 123 nsew signal input
flabel metal3 s 0 131588 96 131668 0 FreeSans 320 0 0 0 FrameData[211]
port 124 nsew signal input
flabel metal3 s 0 132092 96 132172 0 FreeSans 320 0 0 0 FrameData[212]
port 125 nsew signal input
flabel metal3 s 0 132596 96 132676 0 FreeSans 320 0 0 0 FrameData[213]
port 126 nsew signal input
flabel metal3 s 0 133100 96 133180 0 FreeSans 320 0 0 0 FrameData[214]
port 127 nsew signal input
flabel metal3 s 0 133604 96 133684 0 FreeSans 320 0 0 0 FrameData[215]
port 128 nsew signal input
flabel metal3 s 0 134108 96 134188 0 FreeSans 320 0 0 0 FrameData[216]
port 129 nsew signal input
flabel metal3 s 0 134612 96 134692 0 FreeSans 320 0 0 0 FrameData[217]
port 130 nsew signal input
flabel metal3 s 0 135116 96 135196 0 FreeSans 320 0 0 0 FrameData[218]
port 131 nsew signal input
flabel metal3 s 0 135620 96 135700 0 FreeSans 320 0 0 0 FrameData[219]
port 132 nsew signal input
flabel metal3 s 0 362756 96 362836 0 FreeSans 320 0 0 0 FrameData[21]
port 133 nsew signal input
flabel metal3 s 0 136124 96 136204 0 FreeSans 320 0 0 0 FrameData[220]
port 134 nsew signal input
flabel metal3 s 0 136628 96 136708 0 FreeSans 320 0 0 0 FrameData[221]
port 135 nsew signal input
flabel metal3 s 0 137132 96 137212 0 FreeSans 320 0 0 0 FrameData[222]
port 136 nsew signal input
flabel metal3 s 0 137636 96 137716 0 FreeSans 320 0 0 0 FrameData[223]
port 137 nsew signal input
flabel metal3 s 0 79004 96 79084 0 FreeSans 320 0 0 0 FrameData[224]
port 138 nsew signal input
flabel metal3 s 0 79508 96 79588 0 FreeSans 320 0 0 0 FrameData[225]
port 139 nsew signal input
flabel metal3 s 0 80012 96 80092 0 FreeSans 320 0 0 0 FrameData[226]
port 140 nsew signal input
flabel metal3 s 0 80516 96 80596 0 FreeSans 320 0 0 0 FrameData[227]
port 141 nsew signal input
flabel metal3 s 0 81020 96 81100 0 FreeSans 320 0 0 0 FrameData[228]
port 142 nsew signal input
flabel metal3 s 0 81524 96 81604 0 FreeSans 320 0 0 0 FrameData[229]
port 143 nsew signal input
flabel metal3 s 0 363092 96 363172 0 FreeSans 320 0 0 0 FrameData[22]
port 144 nsew signal input
flabel metal3 s 0 82028 96 82108 0 FreeSans 320 0 0 0 FrameData[230]
port 145 nsew signal input
flabel metal3 s 0 82532 96 82612 0 FreeSans 320 0 0 0 FrameData[231]
port 146 nsew signal input
flabel metal3 s 0 83036 96 83116 0 FreeSans 320 0 0 0 FrameData[232]
port 147 nsew signal input
flabel metal3 s 0 83540 96 83620 0 FreeSans 320 0 0 0 FrameData[233]
port 148 nsew signal input
flabel metal3 s 0 84044 96 84124 0 FreeSans 320 0 0 0 FrameData[234]
port 149 nsew signal input
flabel metal3 s 0 84548 96 84628 0 FreeSans 320 0 0 0 FrameData[235]
port 150 nsew signal input
flabel metal3 s 0 85052 96 85132 0 FreeSans 320 0 0 0 FrameData[236]
port 151 nsew signal input
flabel metal3 s 0 85556 96 85636 0 FreeSans 320 0 0 0 FrameData[237]
port 152 nsew signal input
flabel metal3 s 0 86060 96 86140 0 FreeSans 320 0 0 0 FrameData[238]
port 153 nsew signal input
flabel metal3 s 0 86564 96 86644 0 FreeSans 320 0 0 0 FrameData[239]
port 154 nsew signal input
flabel metal3 s 0 363428 96 363508 0 FreeSans 320 0 0 0 FrameData[23]
port 155 nsew signal input
flabel metal3 s 0 87068 96 87148 0 FreeSans 320 0 0 0 FrameData[240]
port 156 nsew signal input
flabel metal3 s 0 87572 96 87652 0 FreeSans 320 0 0 0 FrameData[241]
port 157 nsew signal input
flabel metal3 s 0 88076 96 88156 0 FreeSans 320 0 0 0 FrameData[242]
port 158 nsew signal input
flabel metal3 s 0 88580 96 88660 0 FreeSans 320 0 0 0 FrameData[243]
port 159 nsew signal input
flabel metal3 s 0 89084 96 89164 0 FreeSans 320 0 0 0 FrameData[244]
port 160 nsew signal input
flabel metal3 s 0 89588 96 89668 0 FreeSans 320 0 0 0 FrameData[245]
port 161 nsew signal input
flabel metal3 s 0 90092 96 90172 0 FreeSans 320 0 0 0 FrameData[246]
port 162 nsew signal input
flabel metal3 s 0 90596 96 90676 0 FreeSans 320 0 0 0 FrameData[247]
port 163 nsew signal input
flabel metal3 s 0 91100 96 91180 0 FreeSans 320 0 0 0 FrameData[248]
port 164 nsew signal input
flabel metal3 s 0 91604 96 91684 0 FreeSans 320 0 0 0 FrameData[249]
port 165 nsew signal input
flabel metal3 s 0 363764 96 363844 0 FreeSans 320 0 0 0 FrameData[24]
port 166 nsew signal input
flabel metal3 s 0 92108 96 92188 0 FreeSans 320 0 0 0 FrameData[250]
port 167 nsew signal input
flabel metal3 s 0 92612 96 92692 0 FreeSans 320 0 0 0 FrameData[251]
port 168 nsew signal input
flabel metal3 s 0 93116 96 93196 0 FreeSans 320 0 0 0 FrameData[252]
port 169 nsew signal input
flabel metal3 s 0 93620 96 93700 0 FreeSans 320 0 0 0 FrameData[253]
port 170 nsew signal input
flabel metal3 s 0 94124 96 94204 0 FreeSans 320 0 0 0 FrameData[254]
port 171 nsew signal input
flabel metal3 s 0 94628 96 94708 0 FreeSans 320 0 0 0 FrameData[255]
port 172 nsew signal input
flabel metal3 s 0 35996 96 36076 0 FreeSans 320 0 0 0 FrameData[256]
port 173 nsew signal input
flabel metal3 s 0 36500 96 36580 0 FreeSans 320 0 0 0 FrameData[257]
port 174 nsew signal input
flabel metal3 s 0 37004 96 37084 0 FreeSans 320 0 0 0 FrameData[258]
port 175 nsew signal input
flabel metal3 s 0 37508 96 37588 0 FreeSans 320 0 0 0 FrameData[259]
port 176 nsew signal input
flabel metal3 s 0 364100 96 364180 0 FreeSans 320 0 0 0 FrameData[25]
port 177 nsew signal input
flabel metal3 s 0 38012 96 38092 0 FreeSans 320 0 0 0 FrameData[260]
port 178 nsew signal input
flabel metal3 s 0 38516 96 38596 0 FreeSans 320 0 0 0 FrameData[261]
port 179 nsew signal input
flabel metal3 s 0 39020 96 39100 0 FreeSans 320 0 0 0 FrameData[262]
port 180 nsew signal input
flabel metal3 s 0 39524 96 39604 0 FreeSans 320 0 0 0 FrameData[263]
port 181 nsew signal input
flabel metal3 s 0 40028 96 40108 0 FreeSans 320 0 0 0 FrameData[264]
port 182 nsew signal input
flabel metal3 s 0 40532 96 40612 0 FreeSans 320 0 0 0 FrameData[265]
port 183 nsew signal input
flabel metal3 s 0 41036 96 41116 0 FreeSans 320 0 0 0 FrameData[266]
port 184 nsew signal input
flabel metal3 s 0 41540 96 41620 0 FreeSans 320 0 0 0 FrameData[267]
port 185 nsew signal input
flabel metal3 s 0 42044 96 42124 0 FreeSans 320 0 0 0 FrameData[268]
port 186 nsew signal input
flabel metal3 s 0 42548 96 42628 0 FreeSans 320 0 0 0 FrameData[269]
port 187 nsew signal input
flabel metal3 s 0 364436 96 364516 0 FreeSans 320 0 0 0 FrameData[26]
port 188 nsew signal input
flabel metal3 s 0 43052 96 43132 0 FreeSans 320 0 0 0 FrameData[270]
port 189 nsew signal input
flabel metal3 s 0 43556 96 43636 0 FreeSans 320 0 0 0 FrameData[271]
port 190 nsew signal input
flabel metal3 s 0 44060 96 44140 0 FreeSans 320 0 0 0 FrameData[272]
port 191 nsew signal input
flabel metal3 s 0 44564 96 44644 0 FreeSans 320 0 0 0 FrameData[273]
port 192 nsew signal input
flabel metal3 s 0 45068 96 45148 0 FreeSans 320 0 0 0 FrameData[274]
port 193 nsew signal input
flabel metal3 s 0 45572 96 45652 0 FreeSans 320 0 0 0 FrameData[275]
port 194 nsew signal input
flabel metal3 s 0 46076 96 46156 0 FreeSans 320 0 0 0 FrameData[276]
port 195 nsew signal input
flabel metal3 s 0 46580 96 46660 0 FreeSans 320 0 0 0 FrameData[277]
port 196 nsew signal input
flabel metal3 s 0 47084 96 47164 0 FreeSans 320 0 0 0 FrameData[278]
port 197 nsew signal input
flabel metal3 s 0 47588 96 47668 0 FreeSans 320 0 0 0 FrameData[279]
port 198 nsew signal input
flabel metal3 s 0 364772 96 364852 0 FreeSans 320 0 0 0 FrameData[27]
port 199 nsew signal input
flabel metal3 s 0 48092 96 48172 0 FreeSans 320 0 0 0 FrameData[280]
port 200 nsew signal input
flabel metal3 s 0 48596 96 48676 0 FreeSans 320 0 0 0 FrameData[281]
port 201 nsew signal input
flabel metal3 s 0 49100 96 49180 0 FreeSans 320 0 0 0 FrameData[282]
port 202 nsew signal input
flabel metal3 s 0 49604 96 49684 0 FreeSans 320 0 0 0 FrameData[283]
port 203 nsew signal input
flabel metal3 s 0 50108 96 50188 0 FreeSans 320 0 0 0 FrameData[284]
port 204 nsew signal input
flabel metal3 s 0 50612 96 50692 0 FreeSans 320 0 0 0 FrameData[285]
port 205 nsew signal input
flabel metal3 s 0 51116 96 51196 0 FreeSans 320 0 0 0 FrameData[286]
port 206 nsew signal input
flabel metal3 s 0 51620 96 51700 0 FreeSans 320 0 0 0 FrameData[287]
port 207 nsew signal input
flabel metal3 s 0 884 96 964 0 FreeSans 320 0 0 0 FrameData[288]
port 208 nsew signal input
flabel metal3 s 0 1220 96 1300 0 FreeSans 320 0 0 0 FrameData[289]
port 209 nsew signal input
flabel metal3 s 0 365108 96 365188 0 FreeSans 320 0 0 0 FrameData[28]
port 210 nsew signal input
flabel metal3 s 0 1556 96 1636 0 FreeSans 320 0 0 0 FrameData[290]
port 211 nsew signal input
flabel metal3 s 0 1892 96 1972 0 FreeSans 320 0 0 0 FrameData[291]
port 212 nsew signal input
flabel metal3 s 0 2228 96 2308 0 FreeSans 320 0 0 0 FrameData[292]
port 213 nsew signal input
flabel metal3 s 0 2564 96 2644 0 FreeSans 320 0 0 0 FrameData[293]
port 214 nsew signal input
flabel metal3 s 0 2900 96 2980 0 FreeSans 320 0 0 0 FrameData[294]
port 215 nsew signal input
flabel metal3 s 0 3236 96 3316 0 FreeSans 320 0 0 0 FrameData[295]
port 216 nsew signal input
flabel metal3 s 0 3572 96 3652 0 FreeSans 320 0 0 0 FrameData[296]
port 217 nsew signal input
flabel metal3 s 0 3908 96 3988 0 FreeSans 320 0 0 0 FrameData[297]
port 218 nsew signal input
flabel metal3 s 0 4244 96 4324 0 FreeSans 320 0 0 0 FrameData[298]
port 219 nsew signal input
flabel metal3 s 0 4580 96 4660 0 FreeSans 320 0 0 0 FrameData[299]
port 220 nsew signal input
flabel metal3 s 0 365444 96 365524 0 FreeSans 320 0 0 0 FrameData[29]
port 221 nsew signal input
flabel metal3 s 0 356372 96 356452 0 FreeSans 320 0 0 0 FrameData[2]
port 222 nsew signal input
flabel metal3 s 0 4916 96 4996 0 FreeSans 320 0 0 0 FrameData[300]
port 223 nsew signal input
flabel metal3 s 0 5252 96 5332 0 FreeSans 320 0 0 0 FrameData[301]
port 224 nsew signal input
flabel metal3 s 0 5588 96 5668 0 FreeSans 320 0 0 0 FrameData[302]
port 225 nsew signal input
flabel metal3 s 0 5924 96 6004 0 FreeSans 320 0 0 0 FrameData[303]
port 226 nsew signal input
flabel metal3 s 0 6260 96 6340 0 FreeSans 320 0 0 0 FrameData[304]
port 227 nsew signal input
flabel metal3 s 0 6596 96 6676 0 FreeSans 320 0 0 0 FrameData[305]
port 228 nsew signal input
flabel metal3 s 0 6932 96 7012 0 FreeSans 320 0 0 0 FrameData[306]
port 229 nsew signal input
flabel metal3 s 0 7268 96 7348 0 FreeSans 320 0 0 0 FrameData[307]
port 230 nsew signal input
flabel metal3 s 0 7604 96 7684 0 FreeSans 320 0 0 0 FrameData[308]
port 231 nsew signal input
flabel metal3 s 0 7940 96 8020 0 FreeSans 320 0 0 0 FrameData[309]
port 232 nsew signal input
flabel metal3 s 0 365780 96 365860 0 FreeSans 320 0 0 0 FrameData[30]
port 233 nsew signal input
flabel metal3 s 0 8276 96 8356 0 FreeSans 320 0 0 0 FrameData[310]
port 234 nsew signal input
flabel metal3 s 0 8612 96 8692 0 FreeSans 320 0 0 0 FrameData[311]
port 235 nsew signal input
flabel metal3 s 0 8948 96 9028 0 FreeSans 320 0 0 0 FrameData[312]
port 236 nsew signal input
flabel metal3 s 0 9284 96 9364 0 FreeSans 320 0 0 0 FrameData[313]
port 237 nsew signal input
flabel metal3 s 0 9620 96 9700 0 FreeSans 320 0 0 0 FrameData[314]
port 238 nsew signal input
flabel metal3 s 0 9956 96 10036 0 FreeSans 320 0 0 0 FrameData[315]
port 239 nsew signal input
flabel metal3 s 0 10292 96 10372 0 FreeSans 320 0 0 0 FrameData[316]
port 240 nsew signal input
flabel metal3 s 0 10628 96 10708 0 FreeSans 320 0 0 0 FrameData[317]
port 241 nsew signal input
flabel metal3 s 0 10964 96 11044 0 FreeSans 320 0 0 0 FrameData[318]
port 242 nsew signal input
flabel metal3 s 0 11300 96 11380 0 FreeSans 320 0 0 0 FrameData[319]
port 243 nsew signal input
flabel metal3 s 0 366116 96 366196 0 FreeSans 320 0 0 0 FrameData[31]
port 244 nsew signal input
flabel metal3 s 0 337052 96 337132 0 FreeSans 320 0 0 0 FrameData[32]
port 245 nsew signal input
flabel metal3 s 0 337556 96 337636 0 FreeSans 320 0 0 0 FrameData[33]
port 246 nsew signal input
flabel metal3 s 0 338060 96 338140 0 FreeSans 320 0 0 0 FrameData[34]
port 247 nsew signal input
flabel metal3 s 0 338564 96 338644 0 FreeSans 320 0 0 0 FrameData[35]
port 248 nsew signal input
flabel metal3 s 0 339068 96 339148 0 FreeSans 320 0 0 0 FrameData[36]
port 249 nsew signal input
flabel metal3 s 0 339572 96 339652 0 FreeSans 320 0 0 0 FrameData[37]
port 250 nsew signal input
flabel metal3 s 0 340076 96 340156 0 FreeSans 320 0 0 0 FrameData[38]
port 251 nsew signal input
flabel metal3 s 0 340580 96 340660 0 FreeSans 320 0 0 0 FrameData[39]
port 252 nsew signal input
flabel metal3 s 0 356708 96 356788 0 FreeSans 320 0 0 0 FrameData[3]
port 253 nsew signal input
flabel metal3 s 0 341084 96 341164 0 FreeSans 320 0 0 0 FrameData[40]
port 254 nsew signal input
flabel metal3 s 0 341588 96 341668 0 FreeSans 320 0 0 0 FrameData[41]
port 255 nsew signal input
flabel metal3 s 0 342092 96 342172 0 FreeSans 320 0 0 0 FrameData[42]
port 256 nsew signal input
flabel metal3 s 0 342596 96 342676 0 FreeSans 320 0 0 0 FrameData[43]
port 257 nsew signal input
flabel metal3 s 0 343100 96 343180 0 FreeSans 320 0 0 0 FrameData[44]
port 258 nsew signal input
flabel metal3 s 0 343604 96 343684 0 FreeSans 320 0 0 0 FrameData[45]
port 259 nsew signal input
flabel metal3 s 0 344108 96 344188 0 FreeSans 320 0 0 0 FrameData[46]
port 260 nsew signal input
flabel metal3 s 0 344612 96 344692 0 FreeSans 320 0 0 0 FrameData[47]
port 261 nsew signal input
flabel metal3 s 0 345116 96 345196 0 FreeSans 320 0 0 0 FrameData[48]
port 262 nsew signal input
flabel metal3 s 0 345620 96 345700 0 FreeSans 320 0 0 0 FrameData[49]
port 263 nsew signal input
flabel metal3 s 0 357044 96 357124 0 FreeSans 320 0 0 0 FrameData[4]
port 264 nsew signal input
flabel metal3 s 0 346124 96 346204 0 FreeSans 320 0 0 0 FrameData[50]
port 265 nsew signal input
flabel metal3 s 0 346628 96 346708 0 FreeSans 320 0 0 0 FrameData[51]
port 266 nsew signal input
flabel metal3 s 0 347132 96 347212 0 FreeSans 320 0 0 0 FrameData[52]
port 267 nsew signal input
flabel metal3 s 0 347636 96 347716 0 FreeSans 320 0 0 0 FrameData[53]
port 268 nsew signal input
flabel metal3 s 0 348140 96 348220 0 FreeSans 320 0 0 0 FrameData[54]
port 269 nsew signal input
flabel metal3 s 0 348644 96 348724 0 FreeSans 320 0 0 0 FrameData[55]
port 270 nsew signal input
flabel metal3 s 0 349148 96 349228 0 FreeSans 320 0 0 0 FrameData[56]
port 271 nsew signal input
flabel metal3 s 0 349652 96 349732 0 FreeSans 320 0 0 0 FrameData[57]
port 272 nsew signal input
flabel metal3 s 0 350156 96 350236 0 FreeSans 320 0 0 0 FrameData[58]
port 273 nsew signal input
flabel metal3 s 0 350660 96 350740 0 FreeSans 320 0 0 0 FrameData[59]
port 274 nsew signal input
flabel metal3 s 0 357380 96 357460 0 FreeSans 320 0 0 0 FrameData[5]
port 275 nsew signal input
flabel metal3 s 0 351164 96 351244 0 FreeSans 320 0 0 0 FrameData[60]
port 276 nsew signal input
flabel metal3 s 0 351668 96 351748 0 FreeSans 320 0 0 0 FrameData[61]
port 277 nsew signal input
flabel metal3 s 0 352172 96 352252 0 FreeSans 320 0 0 0 FrameData[62]
port 278 nsew signal input
flabel metal3 s 0 352676 96 352756 0 FreeSans 320 0 0 0 FrameData[63]
port 279 nsew signal input
flabel metal3 s 0 294044 96 294124 0 FreeSans 320 0 0 0 FrameData[64]
port 280 nsew signal input
flabel metal3 s 0 294548 96 294628 0 FreeSans 320 0 0 0 FrameData[65]
port 281 nsew signal input
flabel metal3 s 0 295052 96 295132 0 FreeSans 320 0 0 0 FrameData[66]
port 282 nsew signal input
flabel metal3 s 0 295556 96 295636 0 FreeSans 320 0 0 0 FrameData[67]
port 283 nsew signal input
flabel metal3 s 0 296060 96 296140 0 FreeSans 320 0 0 0 FrameData[68]
port 284 nsew signal input
flabel metal3 s 0 296564 96 296644 0 FreeSans 320 0 0 0 FrameData[69]
port 285 nsew signal input
flabel metal3 s 0 357716 96 357796 0 FreeSans 320 0 0 0 FrameData[6]
port 286 nsew signal input
flabel metal3 s 0 297068 96 297148 0 FreeSans 320 0 0 0 FrameData[70]
port 287 nsew signal input
flabel metal3 s 0 297572 96 297652 0 FreeSans 320 0 0 0 FrameData[71]
port 288 nsew signal input
flabel metal3 s 0 298076 96 298156 0 FreeSans 320 0 0 0 FrameData[72]
port 289 nsew signal input
flabel metal3 s 0 298580 96 298660 0 FreeSans 320 0 0 0 FrameData[73]
port 290 nsew signal input
flabel metal3 s 0 299084 96 299164 0 FreeSans 320 0 0 0 FrameData[74]
port 291 nsew signal input
flabel metal3 s 0 299588 96 299668 0 FreeSans 320 0 0 0 FrameData[75]
port 292 nsew signal input
flabel metal3 s 0 300092 96 300172 0 FreeSans 320 0 0 0 FrameData[76]
port 293 nsew signal input
flabel metal3 s 0 300596 96 300676 0 FreeSans 320 0 0 0 FrameData[77]
port 294 nsew signal input
flabel metal3 s 0 301100 96 301180 0 FreeSans 320 0 0 0 FrameData[78]
port 295 nsew signal input
flabel metal3 s 0 301604 96 301684 0 FreeSans 320 0 0 0 FrameData[79]
port 296 nsew signal input
flabel metal3 s 0 358052 96 358132 0 FreeSans 320 0 0 0 FrameData[7]
port 297 nsew signal input
flabel metal3 s 0 302108 96 302188 0 FreeSans 320 0 0 0 FrameData[80]
port 298 nsew signal input
flabel metal3 s 0 302612 96 302692 0 FreeSans 320 0 0 0 FrameData[81]
port 299 nsew signal input
flabel metal3 s 0 303116 96 303196 0 FreeSans 320 0 0 0 FrameData[82]
port 300 nsew signal input
flabel metal3 s 0 303620 96 303700 0 FreeSans 320 0 0 0 FrameData[83]
port 301 nsew signal input
flabel metal3 s 0 304124 96 304204 0 FreeSans 320 0 0 0 FrameData[84]
port 302 nsew signal input
flabel metal3 s 0 304628 96 304708 0 FreeSans 320 0 0 0 FrameData[85]
port 303 nsew signal input
flabel metal3 s 0 305132 96 305212 0 FreeSans 320 0 0 0 FrameData[86]
port 304 nsew signal input
flabel metal3 s 0 305636 96 305716 0 FreeSans 320 0 0 0 FrameData[87]
port 305 nsew signal input
flabel metal3 s 0 306140 96 306220 0 FreeSans 320 0 0 0 FrameData[88]
port 306 nsew signal input
flabel metal3 s 0 306644 96 306724 0 FreeSans 320 0 0 0 FrameData[89]
port 307 nsew signal input
flabel metal3 s 0 358388 96 358468 0 FreeSans 320 0 0 0 FrameData[8]
port 308 nsew signal input
flabel metal3 s 0 307148 96 307228 0 FreeSans 320 0 0 0 FrameData[90]
port 309 nsew signal input
flabel metal3 s 0 307652 96 307732 0 FreeSans 320 0 0 0 FrameData[91]
port 310 nsew signal input
flabel metal3 s 0 308156 96 308236 0 FreeSans 320 0 0 0 FrameData[92]
port 311 nsew signal input
flabel metal3 s 0 308660 96 308740 0 FreeSans 320 0 0 0 FrameData[93]
port 312 nsew signal input
flabel metal3 s 0 309164 96 309244 0 FreeSans 320 0 0 0 FrameData[94]
port 313 nsew signal input
flabel metal3 s 0 309668 96 309748 0 FreeSans 320 0 0 0 FrameData[95]
port 314 nsew signal input
flabel metal3 s 0 251036 96 251116 0 FreeSans 320 0 0 0 FrameData[96]
port 315 nsew signal input
flabel metal3 s 0 251540 96 251620 0 FreeSans 320 0 0 0 FrameData[97]
port 316 nsew signal input
flabel metal3 s 0 252044 96 252124 0 FreeSans 320 0 0 0 FrameData[98]
port 317 nsew signal input
flabel metal3 s 0 252548 96 252628 0 FreeSans 320 0 0 0 FrameData[99]
port 318 nsew signal input
flabel metal3 s 0 358724 96 358804 0 FreeSans 320 0 0 0 FrameData[9]
port 319 nsew signal input
flabel metal2 s 2072 0 2152 96 0 FreeSans 640 0 0 0 FrameStrobe[0]
port 320 nsew signal input
flabel metal2 s 195608 0 195688 96 0 FreeSans 640 0 0 0 FrameStrobe[100]
port 321 nsew signal input
flabel metal2 s 196568 0 196648 96 0 FreeSans 640 0 0 0 FrameStrobe[101]
port 322 nsew signal input
flabel metal2 s 197528 0 197608 96 0 FreeSans 640 0 0 0 FrameStrobe[102]
port 323 nsew signal input
flabel metal2 s 198488 0 198568 96 0 FreeSans 640 0 0 0 FrameStrobe[103]
port 324 nsew signal input
flabel metal2 s 199448 0 199528 96 0 FreeSans 640 0 0 0 FrameStrobe[104]
port 325 nsew signal input
flabel metal2 s 200408 0 200488 96 0 FreeSans 640 0 0 0 FrameStrobe[105]
port 326 nsew signal input
flabel metal2 s 201368 0 201448 96 0 FreeSans 640 0 0 0 FrameStrobe[106]
port 327 nsew signal input
flabel metal2 s 202328 0 202408 96 0 FreeSans 640 0 0 0 FrameStrobe[107]
port 328 nsew signal input
flabel metal2 s 203288 0 203368 96 0 FreeSans 640 0 0 0 FrameStrobe[108]
port 329 nsew signal input
flabel metal2 s 204248 0 204328 96 0 FreeSans 640 0 0 0 FrameStrobe[109]
port 330 nsew signal input
flabel metal2 s 11672 0 11752 96 0 FreeSans 640 0 0 0 FrameStrobe[10]
port 331 nsew signal input
flabel metal2 s 205208 0 205288 96 0 FreeSans 640 0 0 0 FrameStrobe[110]
port 332 nsew signal input
flabel metal2 s 206168 0 206248 96 0 FreeSans 640 0 0 0 FrameStrobe[111]
port 333 nsew signal input
flabel metal2 s 207128 0 207208 96 0 FreeSans 640 0 0 0 FrameStrobe[112]
port 334 nsew signal input
flabel metal2 s 208088 0 208168 96 0 FreeSans 640 0 0 0 FrameStrobe[113]
port 335 nsew signal input
flabel metal2 s 209048 0 209128 96 0 FreeSans 640 0 0 0 FrameStrobe[114]
port 336 nsew signal input
flabel metal2 s 210008 0 210088 96 0 FreeSans 640 0 0 0 FrameStrobe[115]
port 337 nsew signal input
flabel metal2 s 210968 0 211048 96 0 FreeSans 640 0 0 0 FrameStrobe[116]
port 338 nsew signal input
flabel metal2 s 211928 0 212008 96 0 FreeSans 640 0 0 0 FrameStrobe[117]
port 339 nsew signal input
flabel metal2 s 212888 0 212968 96 0 FreeSans 640 0 0 0 FrameStrobe[118]
port 340 nsew signal input
flabel metal2 s 213848 0 213928 96 0 FreeSans 640 0 0 0 FrameStrobe[119]
port 341 nsew signal input
flabel metal2 s 12632 0 12712 96 0 FreeSans 640 0 0 0 FrameStrobe[11]
port 342 nsew signal input
flabel metal2 s 13592 0 13672 96 0 FreeSans 640 0 0 0 FrameStrobe[12]
port 343 nsew signal input
flabel metal2 s 14552 0 14632 96 0 FreeSans 640 0 0 0 FrameStrobe[13]
port 344 nsew signal input
flabel metal2 s 15512 0 15592 96 0 FreeSans 640 0 0 0 FrameStrobe[14]
port 345 nsew signal input
flabel metal2 s 16472 0 16552 96 0 FreeSans 640 0 0 0 FrameStrobe[15]
port 346 nsew signal input
flabel metal2 s 17432 0 17512 96 0 FreeSans 640 0 0 0 FrameStrobe[16]
port 347 nsew signal input
flabel metal2 s 18392 0 18472 96 0 FreeSans 640 0 0 0 FrameStrobe[17]
port 348 nsew signal input
flabel metal2 s 19352 0 19432 96 0 FreeSans 640 0 0 0 FrameStrobe[18]
port 349 nsew signal input
flabel metal2 s 20312 0 20392 96 0 FreeSans 640 0 0 0 FrameStrobe[19]
port 350 nsew signal input
flabel metal2 s 3032 0 3112 96 0 FreeSans 640 0 0 0 FrameStrobe[1]
port 351 nsew signal input
flabel metal2 s 39512 0 39592 96 0 FreeSans 640 0 0 0 FrameStrobe[20]
port 352 nsew signal input
flabel metal2 s 40664 0 40744 96 0 FreeSans 640 0 0 0 FrameStrobe[21]
port 353 nsew signal input
flabel metal2 s 41816 0 41896 96 0 FreeSans 640 0 0 0 FrameStrobe[22]
port 354 nsew signal input
flabel metal2 s 42968 0 43048 96 0 FreeSans 640 0 0 0 FrameStrobe[23]
port 355 nsew signal input
flabel metal2 s 44120 0 44200 96 0 FreeSans 640 0 0 0 FrameStrobe[24]
port 356 nsew signal input
flabel metal2 s 45272 0 45352 96 0 FreeSans 640 0 0 0 FrameStrobe[25]
port 357 nsew signal input
flabel metal2 s 46424 0 46504 96 0 FreeSans 640 0 0 0 FrameStrobe[26]
port 358 nsew signal input
flabel metal2 s 47576 0 47656 96 0 FreeSans 640 0 0 0 FrameStrobe[27]
port 359 nsew signal input
flabel metal2 s 48728 0 48808 96 0 FreeSans 640 0 0 0 FrameStrobe[28]
port 360 nsew signal input
flabel metal2 s 49880 0 49960 96 0 FreeSans 640 0 0 0 FrameStrobe[29]
port 361 nsew signal input
flabel metal2 s 3992 0 4072 96 0 FreeSans 640 0 0 0 FrameStrobe[2]
port 362 nsew signal input
flabel metal2 s 51032 0 51112 96 0 FreeSans 640 0 0 0 FrameStrobe[30]
port 363 nsew signal input
flabel metal2 s 52184 0 52264 96 0 FreeSans 640 0 0 0 FrameStrobe[31]
port 364 nsew signal input
flabel metal2 s 53336 0 53416 96 0 FreeSans 640 0 0 0 FrameStrobe[32]
port 365 nsew signal input
flabel metal2 s 54488 0 54568 96 0 FreeSans 640 0 0 0 FrameStrobe[33]
port 366 nsew signal input
flabel metal2 s 55640 0 55720 96 0 FreeSans 640 0 0 0 FrameStrobe[34]
port 367 nsew signal input
flabel metal2 s 56792 0 56872 96 0 FreeSans 640 0 0 0 FrameStrobe[35]
port 368 nsew signal input
flabel metal2 s 57944 0 58024 96 0 FreeSans 640 0 0 0 FrameStrobe[36]
port 369 nsew signal input
flabel metal2 s 59096 0 59176 96 0 FreeSans 640 0 0 0 FrameStrobe[37]
port 370 nsew signal input
flabel metal2 s 60248 0 60328 96 0 FreeSans 640 0 0 0 FrameStrobe[38]
port 371 nsew signal input
flabel metal2 s 61400 0 61480 96 0 FreeSans 640 0 0 0 FrameStrobe[39]
port 372 nsew signal input
flabel metal2 s 4952 0 5032 96 0 FreeSans 640 0 0 0 FrameStrobe[3]
port 373 nsew signal input
flabel metal2 s 82520 0 82600 96 0 FreeSans 640 0 0 0 FrameStrobe[40]
port 374 nsew signal input
flabel metal2 s 83672 0 83752 96 0 FreeSans 640 0 0 0 FrameStrobe[41]
port 375 nsew signal input
flabel metal2 s 84824 0 84904 96 0 FreeSans 640 0 0 0 FrameStrobe[42]
port 376 nsew signal input
flabel metal2 s 85976 0 86056 96 0 FreeSans 640 0 0 0 FrameStrobe[43]
port 377 nsew signal input
flabel metal2 s 87128 0 87208 96 0 FreeSans 640 0 0 0 FrameStrobe[44]
port 378 nsew signal input
flabel metal2 s 88280 0 88360 96 0 FreeSans 640 0 0 0 FrameStrobe[45]
port 379 nsew signal input
flabel metal2 s 89432 0 89512 96 0 FreeSans 640 0 0 0 FrameStrobe[46]
port 380 nsew signal input
flabel metal2 s 90584 0 90664 96 0 FreeSans 640 0 0 0 FrameStrobe[47]
port 381 nsew signal input
flabel metal2 s 91736 0 91816 96 0 FreeSans 640 0 0 0 FrameStrobe[48]
port 382 nsew signal input
flabel metal2 s 92888 0 92968 96 0 FreeSans 640 0 0 0 FrameStrobe[49]
port 383 nsew signal input
flabel metal2 s 5912 0 5992 96 0 FreeSans 640 0 0 0 FrameStrobe[4]
port 384 nsew signal input
flabel metal2 s 94040 0 94120 96 0 FreeSans 640 0 0 0 FrameStrobe[50]
port 385 nsew signal input
flabel metal2 s 95192 0 95272 96 0 FreeSans 640 0 0 0 FrameStrobe[51]
port 386 nsew signal input
flabel metal2 s 96344 0 96424 96 0 FreeSans 640 0 0 0 FrameStrobe[52]
port 387 nsew signal input
flabel metal2 s 97496 0 97576 96 0 FreeSans 640 0 0 0 FrameStrobe[53]
port 388 nsew signal input
flabel metal2 s 98648 0 98728 96 0 FreeSans 640 0 0 0 FrameStrobe[54]
port 389 nsew signal input
flabel metal2 s 99800 0 99880 96 0 FreeSans 640 0 0 0 FrameStrobe[55]
port 390 nsew signal input
flabel metal2 s 100952 0 101032 96 0 FreeSans 640 0 0 0 FrameStrobe[56]
port 391 nsew signal input
flabel metal2 s 102104 0 102184 96 0 FreeSans 640 0 0 0 FrameStrobe[57]
port 392 nsew signal input
flabel metal2 s 103256 0 103336 96 0 FreeSans 640 0 0 0 FrameStrobe[58]
port 393 nsew signal input
flabel metal2 s 104408 0 104488 96 0 FreeSans 640 0 0 0 FrameStrobe[59]
port 394 nsew signal input
flabel metal2 s 6872 0 6952 96 0 FreeSans 640 0 0 0 FrameStrobe[5]
port 395 nsew signal input
flabel metal2 s 125528 0 125608 96 0 FreeSans 640 0 0 0 FrameStrobe[60]
port 396 nsew signal input
flabel metal2 s 126680 0 126760 96 0 FreeSans 640 0 0 0 FrameStrobe[61]
port 397 nsew signal input
flabel metal2 s 127832 0 127912 96 0 FreeSans 640 0 0 0 FrameStrobe[62]
port 398 nsew signal input
flabel metal2 s 128984 0 129064 96 0 FreeSans 640 0 0 0 FrameStrobe[63]
port 399 nsew signal input
flabel metal2 s 130136 0 130216 96 0 FreeSans 640 0 0 0 FrameStrobe[64]
port 400 nsew signal input
flabel metal2 s 131288 0 131368 96 0 FreeSans 640 0 0 0 FrameStrobe[65]
port 401 nsew signal input
flabel metal2 s 132440 0 132520 96 0 FreeSans 640 0 0 0 FrameStrobe[66]
port 402 nsew signal input
flabel metal2 s 133592 0 133672 96 0 FreeSans 640 0 0 0 FrameStrobe[67]
port 403 nsew signal input
flabel metal2 s 134744 0 134824 96 0 FreeSans 640 0 0 0 FrameStrobe[68]
port 404 nsew signal input
flabel metal2 s 135896 0 135976 96 0 FreeSans 640 0 0 0 FrameStrobe[69]
port 405 nsew signal input
flabel metal2 s 7832 0 7912 96 0 FreeSans 640 0 0 0 FrameStrobe[6]
port 406 nsew signal input
flabel metal2 s 137048 0 137128 96 0 FreeSans 640 0 0 0 FrameStrobe[70]
port 407 nsew signal input
flabel metal2 s 138200 0 138280 96 0 FreeSans 640 0 0 0 FrameStrobe[71]
port 408 nsew signal input
flabel metal2 s 139352 0 139432 96 0 FreeSans 640 0 0 0 FrameStrobe[72]
port 409 nsew signal input
flabel metal2 s 140504 0 140584 96 0 FreeSans 640 0 0 0 FrameStrobe[73]
port 410 nsew signal input
flabel metal2 s 141656 0 141736 96 0 FreeSans 640 0 0 0 FrameStrobe[74]
port 411 nsew signal input
flabel metal2 s 142808 0 142888 96 0 FreeSans 640 0 0 0 FrameStrobe[75]
port 412 nsew signal input
flabel metal2 s 143960 0 144040 96 0 FreeSans 640 0 0 0 FrameStrobe[76]
port 413 nsew signal input
flabel metal2 s 145112 0 145192 96 0 FreeSans 640 0 0 0 FrameStrobe[77]
port 414 nsew signal input
flabel metal2 s 146264 0 146344 96 0 FreeSans 640 0 0 0 FrameStrobe[78]
port 415 nsew signal input
flabel metal2 s 147416 0 147496 96 0 FreeSans 640 0 0 0 FrameStrobe[79]
port 416 nsew signal input
flabel metal2 s 8792 0 8872 96 0 FreeSans 640 0 0 0 FrameStrobe[7]
port 417 nsew signal input
flabel metal2 s 168536 0 168616 96 0 FreeSans 640 0 0 0 FrameStrobe[80]
port 418 nsew signal input
flabel metal2 s 169688 0 169768 96 0 FreeSans 640 0 0 0 FrameStrobe[81]
port 419 nsew signal input
flabel metal2 s 170840 0 170920 96 0 FreeSans 640 0 0 0 FrameStrobe[82]
port 420 nsew signal input
flabel metal2 s 171992 0 172072 96 0 FreeSans 640 0 0 0 FrameStrobe[83]
port 421 nsew signal input
flabel metal2 s 173144 0 173224 96 0 FreeSans 640 0 0 0 FrameStrobe[84]
port 422 nsew signal input
flabel metal2 s 174296 0 174376 96 0 FreeSans 640 0 0 0 FrameStrobe[85]
port 423 nsew signal input
flabel metal2 s 175448 0 175528 96 0 FreeSans 640 0 0 0 FrameStrobe[86]
port 424 nsew signal input
flabel metal2 s 176600 0 176680 96 0 FreeSans 640 0 0 0 FrameStrobe[87]
port 425 nsew signal input
flabel metal2 s 177752 0 177832 96 0 FreeSans 640 0 0 0 FrameStrobe[88]
port 426 nsew signal input
flabel metal2 s 178904 0 178984 96 0 FreeSans 640 0 0 0 FrameStrobe[89]
port 427 nsew signal input
flabel metal2 s 9752 0 9832 96 0 FreeSans 640 0 0 0 FrameStrobe[8]
port 428 nsew signal input
flabel metal2 s 180056 0 180136 96 0 FreeSans 640 0 0 0 FrameStrobe[90]
port 429 nsew signal input
flabel metal2 s 181208 0 181288 96 0 FreeSans 640 0 0 0 FrameStrobe[91]
port 430 nsew signal input
flabel metal2 s 182360 0 182440 96 0 FreeSans 640 0 0 0 FrameStrobe[92]
port 431 nsew signal input
flabel metal2 s 183512 0 183592 96 0 FreeSans 640 0 0 0 FrameStrobe[93]
port 432 nsew signal input
flabel metal2 s 184664 0 184744 96 0 FreeSans 640 0 0 0 FrameStrobe[94]
port 433 nsew signal input
flabel metal2 s 185816 0 185896 96 0 FreeSans 640 0 0 0 FrameStrobe[95]
port 434 nsew signal input
flabel metal2 s 186968 0 187048 96 0 FreeSans 640 0 0 0 FrameStrobe[96]
port 435 nsew signal input
flabel metal2 s 188120 0 188200 96 0 FreeSans 640 0 0 0 FrameStrobe[97]
port 436 nsew signal input
flabel metal2 s 189272 0 189352 96 0 FreeSans 640 0 0 0 FrameStrobe[98]
port 437 nsew signal input
flabel metal2 s 190424 0 190504 96 0 FreeSans 640 0 0 0 FrameStrobe[99]
port 438 nsew signal input
flabel metal2 s 10712 0 10792 96 0 FreeSans 640 0 0 0 FrameStrobe[9]
port 439 nsew signal input
flabel metal3 s 0 336044 96 336124 0 FreeSans 320 0 0 0 Tile_X0Y1_CLK_TT_PROJECT
port 440 nsew signal output
flabel metal3 s 0 335540 96 335620 0 FreeSans 320 0 0 0 Tile_X0Y1_ENA_TT_PROJECT
port 441 nsew signal output
flabel metal3 s 0 336548 96 336628 0 FreeSans 320 0 0 0 Tile_X0Y1_RST_N_TT_PROJECT
port 442 nsew signal output
flabel metal3 s 0 331508 96 331588 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_IN_TT_PROJECT0
port 443 nsew signal output
flabel metal3 s 0 332012 96 332092 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_IN_TT_PROJECT1
port 444 nsew signal output
flabel metal3 s 0 332516 96 332596 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_IN_TT_PROJECT2
port 445 nsew signal output
flabel metal3 s 0 333020 96 333100 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_IN_TT_PROJECT3
port 446 nsew signal output
flabel metal3 s 0 333524 96 333604 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_IN_TT_PROJECT4
port 447 nsew signal output
flabel metal3 s 0 334028 96 334108 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_IN_TT_PROJECT5
port 448 nsew signal output
flabel metal3 s 0 334532 96 334612 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_IN_TT_PROJECT6
port 449 nsew signal output
flabel metal3 s 0 335036 96 335116 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_IN_TT_PROJECT7
port 450 nsew signal output
flabel metal3 s 0 323444 96 323524 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OE_TT_PROJECT0
port 451 nsew signal input
flabel metal3 s 0 323948 96 324028 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OE_TT_PROJECT1
port 452 nsew signal input
flabel metal3 s 0 324452 96 324532 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OE_TT_PROJECT2
port 453 nsew signal input
flabel metal3 s 0 324956 96 325036 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OE_TT_PROJECT3
port 454 nsew signal input
flabel metal3 s 0 325460 96 325540 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OE_TT_PROJECT4
port 455 nsew signal input
flabel metal3 s 0 325964 96 326044 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OE_TT_PROJECT5
port 456 nsew signal input
flabel metal3 s 0 326468 96 326548 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OE_TT_PROJECT6
port 457 nsew signal input
flabel metal3 s 0 326972 96 327052 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OE_TT_PROJECT7
port 458 nsew signal input
flabel metal3 s 0 319412 96 319492 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OUT_TT_PROJECT0
port 459 nsew signal input
flabel metal3 s 0 319916 96 319996 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OUT_TT_PROJECT1
port 460 nsew signal input
flabel metal3 s 0 320420 96 320500 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OUT_TT_PROJECT2
port 461 nsew signal input
flabel metal3 s 0 320924 96 321004 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OUT_TT_PROJECT3
port 462 nsew signal input
flabel metal3 s 0 321428 96 321508 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OUT_TT_PROJECT4
port 463 nsew signal input
flabel metal3 s 0 321932 96 322012 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OUT_TT_PROJECT5
port 464 nsew signal input
flabel metal3 s 0 322436 96 322516 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OUT_TT_PROJECT6
port 465 nsew signal input
flabel metal3 s 0 322940 96 323020 0 FreeSans 320 0 0 0 Tile_X0Y1_UIO_OUT_TT_PROJECT7
port 466 nsew signal input
flabel metal3 s 0 327476 96 327556 0 FreeSans 320 0 0 0 Tile_X0Y1_UI_IN_TT_PROJECT0
port 467 nsew signal output
flabel metal3 s 0 327980 96 328060 0 FreeSans 320 0 0 0 Tile_X0Y1_UI_IN_TT_PROJECT1
port 468 nsew signal output
flabel metal3 s 0 328484 96 328564 0 FreeSans 320 0 0 0 Tile_X0Y1_UI_IN_TT_PROJECT2
port 469 nsew signal output
flabel metal3 s 0 328988 96 329068 0 FreeSans 320 0 0 0 Tile_X0Y1_UI_IN_TT_PROJECT3
port 470 nsew signal output
flabel metal3 s 0 329492 96 329572 0 FreeSans 320 0 0 0 Tile_X0Y1_UI_IN_TT_PROJECT4
port 471 nsew signal output
flabel metal3 s 0 329996 96 330076 0 FreeSans 320 0 0 0 Tile_X0Y1_UI_IN_TT_PROJECT5
port 472 nsew signal output
flabel metal3 s 0 330500 96 330580 0 FreeSans 320 0 0 0 Tile_X0Y1_UI_IN_TT_PROJECT6
port 473 nsew signal output
flabel metal3 s 0 331004 96 331084 0 FreeSans 320 0 0 0 Tile_X0Y1_UI_IN_TT_PROJECT7
port 474 nsew signal output
flabel metal3 s 0 315380 96 315460 0 FreeSans 320 0 0 0 Tile_X0Y1_UO_OUT_TT_PROJECT0
port 475 nsew signal input
flabel metal3 s 0 315884 96 315964 0 FreeSans 320 0 0 0 Tile_X0Y1_UO_OUT_TT_PROJECT1
port 476 nsew signal input
flabel metal3 s 0 316388 96 316468 0 FreeSans 320 0 0 0 Tile_X0Y1_UO_OUT_TT_PROJECT2
port 477 nsew signal input
flabel metal3 s 0 316892 96 316972 0 FreeSans 320 0 0 0 Tile_X0Y1_UO_OUT_TT_PROJECT3
port 478 nsew signal input
flabel metal3 s 0 317396 96 317476 0 FreeSans 320 0 0 0 Tile_X0Y1_UO_OUT_TT_PROJECT4
port 479 nsew signal input
flabel metal3 s 0 317900 96 317980 0 FreeSans 320 0 0 0 Tile_X0Y1_UO_OUT_TT_PROJECT5
port 480 nsew signal input
flabel metal3 s 0 318404 96 318484 0 FreeSans 320 0 0 0 Tile_X0Y1_UO_OUT_TT_PROJECT6
port 481 nsew signal input
flabel metal3 s 0 318908 96 318988 0 FreeSans 320 0 0 0 Tile_X0Y1_UO_OUT_TT_PROJECT7
port 482 nsew signal input
flabel metal3 s 0 293036 96 293116 0 FreeSans 320 0 0 0 Tile_X0Y2_CLK_TT_PROJECT
port 483 nsew signal output
flabel metal3 s 0 292532 96 292612 0 FreeSans 320 0 0 0 Tile_X0Y2_ENA_TT_PROJECT
port 484 nsew signal output
flabel metal3 s 0 293540 96 293620 0 FreeSans 320 0 0 0 Tile_X0Y2_RST_N_TT_PROJECT
port 485 nsew signal output
flabel metal3 s 0 288500 96 288580 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_IN_TT_PROJECT0
port 486 nsew signal output
flabel metal3 s 0 289004 96 289084 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_IN_TT_PROJECT1
port 487 nsew signal output
flabel metal3 s 0 289508 96 289588 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_IN_TT_PROJECT2
port 488 nsew signal output
flabel metal3 s 0 290012 96 290092 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_IN_TT_PROJECT3
port 489 nsew signal output
flabel metal3 s 0 290516 96 290596 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_IN_TT_PROJECT4
port 490 nsew signal output
flabel metal3 s 0 291020 96 291100 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_IN_TT_PROJECT5
port 491 nsew signal output
flabel metal3 s 0 291524 96 291604 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_IN_TT_PROJECT6
port 492 nsew signal output
flabel metal3 s 0 292028 96 292108 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_IN_TT_PROJECT7
port 493 nsew signal output
flabel metal3 s 0 280436 96 280516 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OE_TT_PROJECT0
port 494 nsew signal input
flabel metal3 s 0 280940 96 281020 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OE_TT_PROJECT1
port 495 nsew signal input
flabel metal3 s 0 281444 96 281524 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OE_TT_PROJECT2
port 496 nsew signal input
flabel metal3 s 0 281948 96 282028 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OE_TT_PROJECT3
port 497 nsew signal input
flabel metal3 s 0 282452 96 282532 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OE_TT_PROJECT4
port 498 nsew signal input
flabel metal3 s 0 282956 96 283036 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OE_TT_PROJECT5
port 499 nsew signal input
flabel metal3 s 0 283460 96 283540 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OE_TT_PROJECT6
port 500 nsew signal input
flabel metal3 s 0 283964 96 284044 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OE_TT_PROJECT7
port 501 nsew signal input
flabel metal3 s 0 276404 96 276484 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OUT_TT_PROJECT0
port 502 nsew signal input
flabel metal3 s 0 276908 96 276988 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OUT_TT_PROJECT1
port 503 nsew signal input
flabel metal3 s 0 277412 96 277492 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OUT_TT_PROJECT2
port 504 nsew signal input
flabel metal3 s 0 277916 96 277996 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OUT_TT_PROJECT3
port 505 nsew signal input
flabel metal3 s 0 278420 96 278500 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OUT_TT_PROJECT4
port 506 nsew signal input
flabel metal3 s 0 278924 96 279004 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OUT_TT_PROJECT5
port 507 nsew signal input
flabel metal3 s 0 279428 96 279508 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OUT_TT_PROJECT6
port 508 nsew signal input
flabel metal3 s 0 279932 96 280012 0 FreeSans 320 0 0 0 Tile_X0Y2_UIO_OUT_TT_PROJECT7
port 509 nsew signal input
flabel metal3 s 0 284468 96 284548 0 FreeSans 320 0 0 0 Tile_X0Y2_UI_IN_TT_PROJECT0
port 510 nsew signal output
flabel metal3 s 0 284972 96 285052 0 FreeSans 320 0 0 0 Tile_X0Y2_UI_IN_TT_PROJECT1
port 511 nsew signal output
flabel metal3 s 0 285476 96 285556 0 FreeSans 320 0 0 0 Tile_X0Y2_UI_IN_TT_PROJECT2
port 512 nsew signal output
flabel metal3 s 0 285980 96 286060 0 FreeSans 320 0 0 0 Tile_X0Y2_UI_IN_TT_PROJECT3
port 513 nsew signal output
flabel metal3 s 0 286484 96 286564 0 FreeSans 320 0 0 0 Tile_X0Y2_UI_IN_TT_PROJECT4
port 514 nsew signal output
flabel metal3 s 0 286988 96 287068 0 FreeSans 320 0 0 0 Tile_X0Y2_UI_IN_TT_PROJECT5
port 515 nsew signal output
flabel metal3 s 0 287492 96 287572 0 FreeSans 320 0 0 0 Tile_X0Y2_UI_IN_TT_PROJECT6
port 516 nsew signal output
flabel metal3 s 0 287996 96 288076 0 FreeSans 320 0 0 0 Tile_X0Y2_UI_IN_TT_PROJECT7
port 517 nsew signal output
flabel metal3 s 0 272372 96 272452 0 FreeSans 320 0 0 0 Tile_X0Y2_UO_OUT_TT_PROJECT0
port 518 nsew signal input
flabel metal3 s 0 272876 96 272956 0 FreeSans 320 0 0 0 Tile_X0Y2_UO_OUT_TT_PROJECT1
port 519 nsew signal input
flabel metal3 s 0 273380 96 273460 0 FreeSans 320 0 0 0 Tile_X0Y2_UO_OUT_TT_PROJECT2
port 520 nsew signal input
flabel metal3 s 0 273884 96 273964 0 FreeSans 320 0 0 0 Tile_X0Y2_UO_OUT_TT_PROJECT3
port 521 nsew signal input
flabel metal3 s 0 274388 96 274468 0 FreeSans 320 0 0 0 Tile_X0Y2_UO_OUT_TT_PROJECT4
port 522 nsew signal input
flabel metal3 s 0 274892 96 274972 0 FreeSans 320 0 0 0 Tile_X0Y2_UO_OUT_TT_PROJECT5
port 523 nsew signal input
flabel metal3 s 0 275396 96 275476 0 FreeSans 320 0 0 0 Tile_X0Y2_UO_OUT_TT_PROJECT6
port 524 nsew signal input
flabel metal3 s 0 275900 96 275980 0 FreeSans 320 0 0 0 Tile_X0Y2_UO_OUT_TT_PROJECT7
port 525 nsew signal input
flabel metal3 s 0 250028 96 250108 0 FreeSans 320 0 0 0 Tile_X0Y3_CLK_TT_PROJECT
port 526 nsew signal output
flabel metal3 s 0 249524 96 249604 0 FreeSans 320 0 0 0 Tile_X0Y3_ENA_TT_PROJECT
port 527 nsew signal output
flabel metal3 s 0 250532 96 250612 0 FreeSans 320 0 0 0 Tile_X0Y3_RST_N_TT_PROJECT
port 528 nsew signal output
flabel metal3 s 0 245492 96 245572 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_IN_TT_PROJECT0
port 529 nsew signal output
flabel metal3 s 0 245996 96 246076 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_IN_TT_PROJECT1
port 530 nsew signal output
flabel metal3 s 0 246500 96 246580 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_IN_TT_PROJECT2
port 531 nsew signal output
flabel metal3 s 0 247004 96 247084 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_IN_TT_PROJECT3
port 532 nsew signal output
flabel metal3 s 0 247508 96 247588 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_IN_TT_PROJECT4
port 533 nsew signal output
flabel metal3 s 0 248012 96 248092 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_IN_TT_PROJECT5
port 534 nsew signal output
flabel metal3 s 0 248516 96 248596 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_IN_TT_PROJECT6
port 535 nsew signal output
flabel metal3 s 0 249020 96 249100 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_IN_TT_PROJECT7
port 536 nsew signal output
flabel metal3 s 0 237428 96 237508 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OE_TT_PROJECT0
port 537 nsew signal input
flabel metal3 s 0 237932 96 238012 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OE_TT_PROJECT1
port 538 nsew signal input
flabel metal3 s 0 238436 96 238516 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OE_TT_PROJECT2
port 539 nsew signal input
flabel metal3 s 0 238940 96 239020 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OE_TT_PROJECT3
port 540 nsew signal input
flabel metal3 s 0 239444 96 239524 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OE_TT_PROJECT4
port 541 nsew signal input
flabel metal3 s 0 239948 96 240028 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OE_TT_PROJECT5
port 542 nsew signal input
flabel metal3 s 0 240452 96 240532 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OE_TT_PROJECT6
port 543 nsew signal input
flabel metal3 s 0 240956 96 241036 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OE_TT_PROJECT7
port 544 nsew signal input
flabel metal3 s 0 233396 96 233476 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OUT_TT_PROJECT0
port 545 nsew signal input
flabel metal3 s 0 233900 96 233980 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OUT_TT_PROJECT1
port 546 nsew signal input
flabel metal3 s 0 234404 96 234484 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OUT_TT_PROJECT2
port 547 nsew signal input
flabel metal3 s 0 234908 96 234988 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OUT_TT_PROJECT3
port 548 nsew signal input
flabel metal3 s 0 235412 96 235492 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OUT_TT_PROJECT4
port 549 nsew signal input
flabel metal3 s 0 235916 96 235996 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OUT_TT_PROJECT5
port 550 nsew signal input
flabel metal3 s 0 236420 96 236500 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OUT_TT_PROJECT6
port 551 nsew signal input
flabel metal3 s 0 236924 96 237004 0 FreeSans 320 0 0 0 Tile_X0Y3_UIO_OUT_TT_PROJECT7
port 552 nsew signal input
flabel metal3 s 0 241460 96 241540 0 FreeSans 320 0 0 0 Tile_X0Y3_UI_IN_TT_PROJECT0
port 553 nsew signal output
flabel metal3 s 0 241964 96 242044 0 FreeSans 320 0 0 0 Tile_X0Y3_UI_IN_TT_PROJECT1
port 554 nsew signal output
flabel metal3 s 0 242468 96 242548 0 FreeSans 320 0 0 0 Tile_X0Y3_UI_IN_TT_PROJECT2
port 555 nsew signal output
flabel metal3 s 0 242972 96 243052 0 FreeSans 320 0 0 0 Tile_X0Y3_UI_IN_TT_PROJECT3
port 556 nsew signal output
flabel metal3 s 0 243476 96 243556 0 FreeSans 320 0 0 0 Tile_X0Y3_UI_IN_TT_PROJECT4
port 557 nsew signal output
flabel metal3 s 0 243980 96 244060 0 FreeSans 320 0 0 0 Tile_X0Y3_UI_IN_TT_PROJECT5
port 558 nsew signal output
flabel metal3 s 0 244484 96 244564 0 FreeSans 320 0 0 0 Tile_X0Y3_UI_IN_TT_PROJECT6
port 559 nsew signal output
flabel metal3 s 0 244988 96 245068 0 FreeSans 320 0 0 0 Tile_X0Y3_UI_IN_TT_PROJECT7
port 560 nsew signal output
flabel metal3 s 0 229364 96 229444 0 FreeSans 320 0 0 0 Tile_X0Y3_UO_OUT_TT_PROJECT0
port 561 nsew signal input
flabel metal3 s 0 229868 96 229948 0 FreeSans 320 0 0 0 Tile_X0Y3_UO_OUT_TT_PROJECT1
port 562 nsew signal input
flabel metal3 s 0 230372 96 230452 0 FreeSans 320 0 0 0 Tile_X0Y3_UO_OUT_TT_PROJECT2
port 563 nsew signal input
flabel metal3 s 0 230876 96 230956 0 FreeSans 320 0 0 0 Tile_X0Y3_UO_OUT_TT_PROJECT3
port 564 nsew signal input
flabel metal3 s 0 231380 96 231460 0 FreeSans 320 0 0 0 Tile_X0Y3_UO_OUT_TT_PROJECT4
port 565 nsew signal input
flabel metal3 s 0 231884 96 231964 0 FreeSans 320 0 0 0 Tile_X0Y3_UO_OUT_TT_PROJECT5
port 566 nsew signal input
flabel metal3 s 0 232388 96 232468 0 FreeSans 320 0 0 0 Tile_X0Y3_UO_OUT_TT_PROJECT6
port 567 nsew signal input
flabel metal3 s 0 232892 96 232972 0 FreeSans 320 0 0 0 Tile_X0Y3_UO_OUT_TT_PROJECT7
port 568 nsew signal input
flabel metal3 s 0 207020 96 207100 0 FreeSans 320 0 0 0 Tile_X0Y4_CLK_TT_PROJECT
port 569 nsew signal output
flabel metal3 s 0 206516 96 206596 0 FreeSans 320 0 0 0 Tile_X0Y4_ENA_TT_PROJECT
port 570 nsew signal output
flabel metal3 s 0 207524 96 207604 0 FreeSans 320 0 0 0 Tile_X0Y4_RST_N_TT_PROJECT
port 571 nsew signal output
flabel metal3 s 0 202484 96 202564 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_IN_TT_PROJECT0
port 572 nsew signal output
flabel metal3 s 0 202988 96 203068 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_IN_TT_PROJECT1
port 573 nsew signal output
flabel metal3 s 0 203492 96 203572 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_IN_TT_PROJECT2
port 574 nsew signal output
flabel metal3 s 0 203996 96 204076 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_IN_TT_PROJECT3
port 575 nsew signal output
flabel metal3 s 0 204500 96 204580 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_IN_TT_PROJECT4
port 576 nsew signal output
flabel metal3 s 0 205004 96 205084 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_IN_TT_PROJECT5
port 577 nsew signal output
flabel metal3 s 0 205508 96 205588 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_IN_TT_PROJECT6
port 578 nsew signal output
flabel metal3 s 0 206012 96 206092 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_IN_TT_PROJECT7
port 579 nsew signal output
flabel metal3 s 0 194420 96 194500 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OE_TT_PROJECT0
port 580 nsew signal input
flabel metal3 s 0 194924 96 195004 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OE_TT_PROJECT1
port 581 nsew signal input
flabel metal3 s 0 195428 96 195508 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OE_TT_PROJECT2
port 582 nsew signal input
flabel metal3 s 0 195932 96 196012 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OE_TT_PROJECT3
port 583 nsew signal input
flabel metal3 s 0 196436 96 196516 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OE_TT_PROJECT4
port 584 nsew signal input
flabel metal3 s 0 196940 96 197020 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OE_TT_PROJECT5
port 585 nsew signal input
flabel metal3 s 0 197444 96 197524 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OE_TT_PROJECT6
port 586 nsew signal input
flabel metal3 s 0 197948 96 198028 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OE_TT_PROJECT7
port 587 nsew signal input
flabel metal3 s 0 190388 96 190468 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OUT_TT_PROJECT0
port 588 nsew signal input
flabel metal3 s 0 190892 96 190972 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OUT_TT_PROJECT1
port 589 nsew signal input
flabel metal3 s 0 191396 96 191476 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OUT_TT_PROJECT2
port 590 nsew signal input
flabel metal3 s 0 191900 96 191980 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OUT_TT_PROJECT3
port 591 nsew signal input
flabel metal3 s 0 192404 96 192484 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OUT_TT_PROJECT4
port 592 nsew signal input
flabel metal3 s 0 192908 96 192988 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OUT_TT_PROJECT5
port 593 nsew signal input
flabel metal3 s 0 193412 96 193492 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OUT_TT_PROJECT6
port 594 nsew signal input
flabel metal3 s 0 193916 96 193996 0 FreeSans 320 0 0 0 Tile_X0Y4_UIO_OUT_TT_PROJECT7
port 595 nsew signal input
flabel metal3 s 0 198452 96 198532 0 FreeSans 320 0 0 0 Tile_X0Y4_UI_IN_TT_PROJECT0
port 596 nsew signal output
flabel metal3 s 0 198956 96 199036 0 FreeSans 320 0 0 0 Tile_X0Y4_UI_IN_TT_PROJECT1
port 597 nsew signal output
flabel metal3 s 0 199460 96 199540 0 FreeSans 320 0 0 0 Tile_X0Y4_UI_IN_TT_PROJECT2
port 598 nsew signal output
flabel metal3 s 0 199964 96 200044 0 FreeSans 320 0 0 0 Tile_X0Y4_UI_IN_TT_PROJECT3
port 599 nsew signal output
flabel metal3 s 0 200468 96 200548 0 FreeSans 320 0 0 0 Tile_X0Y4_UI_IN_TT_PROJECT4
port 600 nsew signal output
flabel metal3 s 0 200972 96 201052 0 FreeSans 320 0 0 0 Tile_X0Y4_UI_IN_TT_PROJECT5
port 601 nsew signal output
flabel metal3 s 0 201476 96 201556 0 FreeSans 320 0 0 0 Tile_X0Y4_UI_IN_TT_PROJECT6
port 602 nsew signal output
flabel metal3 s 0 201980 96 202060 0 FreeSans 320 0 0 0 Tile_X0Y4_UI_IN_TT_PROJECT7
port 603 nsew signal output
flabel metal3 s 0 186356 96 186436 0 FreeSans 320 0 0 0 Tile_X0Y4_UO_OUT_TT_PROJECT0
port 604 nsew signal input
flabel metal3 s 0 186860 96 186940 0 FreeSans 320 0 0 0 Tile_X0Y4_UO_OUT_TT_PROJECT1
port 605 nsew signal input
flabel metal3 s 0 187364 96 187444 0 FreeSans 320 0 0 0 Tile_X0Y4_UO_OUT_TT_PROJECT2
port 606 nsew signal input
flabel metal3 s 0 187868 96 187948 0 FreeSans 320 0 0 0 Tile_X0Y4_UO_OUT_TT_PROJECT3
port 607 nsew signal input
flabel metal3 s 0 188372 96 188452 0 FreeSans 320 0 0 0 Tile_X0Y4_UO_OUT_TT_PROJECT4
port 608 nsew signal input
flabel metal3 s 0 188876 96 188956 0 FreeSans 320 0 0 0 Tile_X0Y4_UO_OUT_TT_PROJECT5
port 609 nsew signal input
flabel metal3 s 0 189380 96 189460 0 FreeSans 320 0 0 0 Tile_X0Y4_UO_OUT_TT_PROJECT6
port 610 nsew signal input
flabel metal3 s 0 189884 96 189964 0 FreeSans 320 0 0 0 Tile_X0Y4_UO_OUT_TT_PROJECT7
port 611 nsew signal input
flabel metal3 s 0 164012 96 164092 0 FreeSans 320 0 0 0 Tile_X0Y5_CLK_TT_PROJECT
port 612 nsew signal output
flabel metal3 s 0 163508 96 163588 0 FreeSans 320 0 0 0 Tile_X0Y5_ENA_TT_PROJECT
port 613 nsew signal output
flabel metal3 s 0 164516 96 164596 0 FreeSans 320 0 0 0 Tile_X0Y5_RST_N_TT_PROJECT
port 614 nsew signal output
flabel metal3 s 0 159476 96 159556 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_IN_TT_PROJECT0
port 615 nsew signal output
flabel metal3 s 0 159980 96 160060 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_IN_TT_PROJECT1
port 616 nsew signal output
flabel metal3 s 0 160484 96 160564 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_IN_TT_PROJECT2
port 617 nsew signal output
flabel metal3 s 0 160988 96 161068 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_IN_TT_PROJECT3
port 618 nsew signal output
flabel metal3 s 0 161492 96 161572 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_IN_TT_PROJECT4
port 619 nsew signal output
flabel metal3 s 0 161996 96 162076 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_IN_TT_PROJECT5
port 620 nsew signal output
flabel metal3 s 0 162500 96 162580 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_IN_TT_PROJECT6
port 621 nsew signal output
flabel metal3 s 0 163004 96 163084 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_IN_TT_PROJECT7
port 622 nsew signal output
flabel metal3 s 0 151412 96 151492 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OE_TT_PROJECT0
port 623 nsew signal input
flabel metal3 s 0 151916 96 151996 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OE_TT_PROJECT1
port 624 nsew signal input
flabel metal3 s 0 152420 96 152500 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OE_TT_PROJECT2
port 625 nsew signal input
flabel metal3 s 0 152924 96 153004 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OE_TT_PROJECT3
port 626 nsew signal input
flabel metal3 s 0 153428 96 153508 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OE_TT_PROJECT4
port 627 nsew signal input
flabel metal3 s 0 153932 96 154012 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OE_TT_PROJECT5
port 628 nsew signal input
flabel metal3 s 0 154436 96 154516 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OE_TT_PROJECT6
port 629 nsew signal input
flabel metal3 s 0 154940 96 155020 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OE_TT_PROJECT7
port 630 nsew signal input
flabel metal3 s 0 147380 96 147460 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OUT_TT_PROJECT0
port 631 nsew signal input
flabel metal3 s 0 147884 96 147964 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OUT_TT_PROJECT1
port 632 nsew signal input
flabel metal3 s 0 148388 96 148468 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OUT_TT_PROJECT2
port 633 nsew signal input
flabel metal3 s 0 148892 96 148972 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OUT_TT_PROJECT3
port 634 nsew signal input
flabel metal3 s 0 149396 96 149476 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OUT_TT_PROJECT4
port 635 nsew signal input
flabel metal3 s 0 149900 96 149980 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OUT_TT_PROJECT5
port 636 nsew signal input
flabel metal3 s 0 150404 96 150484 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OUT_TT_PROJECT6
port 637 nsew signal input
flabel metal3 s 0 150908 96 150988 0 FreeSans 320 0 0 0 Tile_X0Y5_UIO_OUT_TT_PROJECT7
port 638 nsew signal input
flabel metal3 s 0 155444 96 155524 0 FreeSans 320 0 0 0 Tile_X0Y5_UI_IN_TT_PROJECT0
port 639 nsew signal output
flabel metal3 s 0 155948 96 156028 0 FreeSans 320 0 0 0 Tile_X0Y5_UI_IN_TT_PROJECT1
port 640 nsew signal output
flabel metal3 s 0 156452 96 156532 0 FreeSans 320 0 0 0 Tile_X0Y5_UI_IN_TT_PROJECT2
port 641 nsew signal output
flabel metal3 s 0 156956 96 157036 0 FreeSans 320 0 0 0 Tile_X0Y5_UI_IN_TT_PROJECT3
port 642 nsew signal output
flabel metal3 s 0 157460 96 157540 0 FreeSans 320 0 0 0 Tile_X0Y5_UI_IN_TT_PROJECT4
port 643 nsew signal output
flabel metal3 s 0 157964 96 158044 0 FreeSans 320 0 0 0 Tile_X0Y5_UI_IN_TT_PROJECT5
port 644 nsew signal output
flabel metal3 s 0 158468 96 158548 0 FreeSans 320 0 0 0 Tile_X0Y5_UI_IN_TT_PROJECT6
port 645 nsew signal output
flabel metal3 s 0 158972 96 159052 0 FreeSans 320 0 0 0 Tile_X0Y5_UI_IN_TT_PROJECT7
port 646 nsew signal output
flabel metal3 s 0 143348 96 143428 0 FreeSans 320 0 0 0 Tile_X0Y5_UO_OUT_TT_PROJECT0
port 647 nsew signal input
flabel metal3 s 0 143852 96 143932 0 FreeSans 320 0 0 0 Tile_X0Y5_UO_OUT_TT_PROJECT1
port 648 nsew signal input
flabel metal3 s 0 144356 96 144436 0 FreeSans 320 0 0 0 Tile_X0Y5_UO_OUT_TT_PROJECT2
port 649 nsew signal input
flabel metal3 s 0 144860 96 144940 0 FreeSans 320 0 0 0 Tile_X0Y5_UO_OUT_TT_PROJECT3
port 650 nsew signal input
flabel metal3 s 0 145364 96 145444 0 FreeSans 320 0 0 0 Tile_X0Y5_UO_OUT_TT_PROJECT4
port 651 nsew signal input
flabel metal3 s 0 145868 96 145948 0 FreeSans 320 0 0 0 Tile_X0Y5_UO_OUT_TT_PROJECT5
port 652 nsew signal input
flabel metal3 s 0 146372 96 146452 0 FreeSans 320 0 0 0 Tile_X0Y5_UO_OUT_TT_PROJECT6
port 653 nsew signal input
flabel metal3 s 0 146876 96 146956 0 FreeSans 320 0 0 0 Tile_X0Y5_UO_OUT_TT_PROJECT7
port 654 nsew signal input
flabel metal3 s 0 121004 96 121084 0 FreeSans 320 0 0 0 Tile_X0Y6_CLK_TT_PROJECT
port 655 nsew signal output
flabel metal3 s 0 120500 96 120580 0 FreeSans 320 0 0 0 Tile_X0Y6_ENA_TT_PROJECT
port 656 nsew signal output
flabel metal3 s 0 121508 96 121588 0 FreeSans 320 0 0 0 Tile_X0Y6_RST_N_TT_PROJECT
port 657 nsew signal output
flabel metal3 s 0 116468 96 116548 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_IN_TT_PROJECT0
port 658 nsew signal output
flabel metal3 s 0 116972 96 117052 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_IN_TT_PROJECT1
port 659 nsew signal output
flabel metal3 s 0 117476 96 117556 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_IN_TT_PROJECT2
port 660 nsew signal output
flabel metal3 s 0 117980 96 118060 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_IN_TT_PROJECT3
port 661 nsew signal output
flabel metal3 s 0 118484 96 118564 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_IN_TT_PROJECT4
port 662 nsew signal output
flabel metal3 s 0 118988 96 119068 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_IN_TT_PROJECT5
port 663 nsew signal output
flabel metal3 s 0 119492 96 119572 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_IN_TT_PROJECT6
port 664 nsew signal output
flabel metal3 s 0 119996 96 120076 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_IN_TT_PROJECT7
port 665 nsew signal output
flabel metal3 s 0 108404 96 108484 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OE_TT_PROJECT0
port 666 nsew signal input
flabel metal3 s 0 108908 96 108988 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OE_TT_PROJECT1
port 667 nsew signal input
flabel metal3 s 0 109412 96 109492 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OE_TT_PROJECT2
port 668 nsew signal input
flabel metal3 s 0 109916 96 109996 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OE_TT_PROJECT3
port 669 nsew signal input
flabel metal3 s 0 110420 96 110500 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OE_TT_PROJECT4
port 670 nsew signal input
flabel metal3 s 0 110924 96 111004 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OE_TT_PROJECT5
port 671 nsew signal input
flabel metal3 s 0 111428 96 111508 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OE_TT_PROJECT6
port 672 nsew signal input
flabel metal3 s 0 111932 96 112012 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OE_TT_PROJECT7
port 673 nsew signal input
flabel metal3 s 0 104372 96 104452 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OUT_TT_PROJECT0
port 674 nsew signal input
flabel metal3 s 0 104876 96 104956 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OUT_TT_PROJECT1
port 675 nsew signal input
flabel metal3 s 0 105380 96 105460 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OUT_TT_PROJECT2
port 676 nsew signal input
flabel metal3 s 0 105884 96 105964 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OUT_TT_PROJECT3
port 677 nsew signal input
flabel metal3 s 0 106388 96 106468 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OUT_TT_PROJECT4
port 678 nsew signal input
flabel metal3 s 0 106892 96 106972 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OUT_TT_PROJECT5
port 679 nsew signal input
flabel metal3 s 0 107396 96 107476 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OUT_TT_PROJECT6
port 680 nsew signal input
flabel metal3 s 0 107900 96 107980 0 FreeSans 320 0 0 0 Tile_X0Y6_UIO_OUT_TT_PROJECT7
port 681 nsew signal input
flabel metal3 s 0 112436 96 112516 0 FreeSans 320 0 0 0 Tile_X0Y6_UI_IN_TT_PROJECT0
port 682 nsew signal output
flabel metal3 s 0 112940 96 113020 0 FreeSans 320 0 0 0 Tile_X0Y6_UI_IN_TT_PROJECT1
port 683 nsew signal output
flabel metal3 s 0 113444 96 113524 0 FreeSans 320 0 0 0 Tile_X0Y6_UI_IN_TT_PROJECT2
port 684 nsew signal output
flabel metal3 s 0 113948 96 114028 0 FreeSans 320 0 0 0 Tile_X0Y6_UI_IN_TT_PROJECT3
port 685 nsew signal output
flabel metal3 s 0 114452 96 114532 0 FreeSans 320 0 0 0 Tile_X0Y6_UI_IN_TT_PROJECT4
port 686 nsew signal output
flabel metal3 s 0 114956 96 115036 0 FreeSans 320 0 0 0 Tile_X0Y6_UI_IN_TT_PROJECT5
port 687 nsew signal output
flabel metal3 s 0 115460 96 115540 0 FreeSans 320 0 0 0 Tile_X0Y6_UI_IN_TT_PROJECT6
port 688 nsew signal output
flabel metal3 s 0 115964 96 116044 0 FreeSans 320 0 0 0 Tile_X0Y6_UI_IN_TT_PROJECT7
port 689 nsew signal output
flabel metal3 s 0 100340 96 100420 0 FreeSans 320 0 0 0 Tile_X0Y6_UO_OUT_TT_PROJECT0
port 690 nsew signal input
flabel metal3 s 0 100844 96 100924 0 FreeSans 320 0 0 0 Tile_X0Y6_UO_OUT_TT_PROJECT1
port 691 nsew signal input
flabel metal3 s 0 101348 96 101428 0 FreeSans 320 0 0 0 Tile_X0Y6_UO_OUT_TT_PROJECT2
port 692 nsew signal input
flabel metal3 s 0 101852 96 101932 0 FreeSans 320 0 0 0 Tile_X0Y6_UO_OUT_TT_PROJECT3
port 693 nsew signal input
flabel metal3 s 0 102356 96 102436 0 FreeSans 320 0 0 0 Tile_X0Y6_UO_OUT_TT_PROJECT4
port 694 nsew signal input
flabel metal3 s 0 102860 96 102940 0 FreeSans 320 0 0 0 Tile_X0Y6_UO_OUT_TT_PROJECT5
port 695 nsew signal input
flabel metal3 s 0 103364 96 103444 0 FreeSans 320 0 0 0 Tile_X0Y6_UO_OUT_TT_PROJECT6
port 696 nsew signal input
flabel metal3 s 0 103868 96 103948 0 FreeSans 320 0 0 0 Tile_X0Y6_UO_OUT_TT_PROJECT7
port 697 nsew signal input
flabel metal3 s 0 77996 96 78076 0 FreeSans 320 0 0 0 Tile_X0Y7_CLK_TT_PROJECT
port 698 nsew signal output
flabel metal3 s 0 77492 96 77572 0 FreeSans 320 0 0 0 Tile_X0Y7_ENA_TT_PROJECT
port 699 nsew signal output
flabel metal3 s 0 78500 96 78580 0 FreeSans 320 0 0 0 Tile_X0Y7_RST_N_TT_PROJECT
port 700 nsew signal output
flabel metal3 s 0 73460 96 73540 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_IN_TT_PROJECT0
port 701 nsew signal output
flabel metal3 s 0 73964 96 74044 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_IN_TT_PROJECT1
port 702 nsew signal output
flabel metal3 s 0 74468 96 74548 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_IN_TT_PROJECT2
port 703 nsew signal output
flabel metal3 s 0 74972 96 75052 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_IN_TT_PROJECT3
port 704 nsew signal output
flabel metal3 s 0 75476 96 75556 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_IN_TT_PROJECT4
port 705 nsew signal output
flabel metal3 s 0 75980 96 76060 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_IN_TT_PROJECT5
port 706 nsew signal output
flabel metal3 s 0 76484 96 76564 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_IN_TT_PROJECT6
port 707 nsew signal output
flabel metal3 s 0 76988 96 77068 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_IN_TT_PROJECT7
port 708 nsew signal output
flabel metal3 s 0 65396 96 65476 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OE_TT_PROJECT0
port 709 nsew signal input
flabel metal3 s 0 65900 96 65980 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OE_TT_PROJECT1
port 710 nsew signal input
flabel metal3 s 0 66404 96 66484 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OE_TT_PROJECT2
port 711 nsew signal input
flabel metal3 s 0 66908 96 66988 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OE_TT_PROJECT3
port 712 nsew signal input
flabel metal3 s 0 67412 96 67492 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OE_TT_PROJECT4
port 713 nsew signal input
flabel metal3 s 0 67916 96 67996 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OE_TT_PROJECT5
port 714 nsew signal input
flabel metal3 s 0 68420 96 68500 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OE_TT_PROJECT6
port 715 nsew signal input
flabel metal3 s 0 68924 96 69004 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OE_TT_PROJECT7
port 716 nsew signal input
flabel metal3 s 0 61364 96 61444 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OUT_TT_PROJECT0
port 717 nsew signal input
flabel metal3 s 0 61868 96 61948 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OUT_TT_PROJECT1
port 718 nsew signal input
flabel metal3 s 0 62372 96 62452 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OUT_TT_PROJECT2
port 719 nsew signal input
flabel metal3 s 0 62876 96 62956 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OUT_TT_PROJECT3
port 720 nsew signal input
flabel metal3 s 0 63380 96 63460 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OUT_TT_PROJECT4
port 721 nsew signal input
flabel metal3 s 0 63884 96 63964 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OUT_TT_PROJECT5
port 722 nsew signal input
flabel metal3 s 0 64388 96 64468 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OUT_TT_PROJECT6
port 723 nsew signal input
flabel metal3 s 0 64892 96 64972 0 FreeSans 320 0 0 0 Tile_X0Y7_UIO_OUT_TT_PROJECT7
port 724 nsew signal input
flabel metal3 s 0 69428 96 69508 0 FreeSans 320 0 0 0 Tile_X0Y7_UI_IN_TT_PROJECT0
port 725 nsew signal output
flabel metal3 s 0 69932 96 70012 0 FreeSans 320 0 0 0 Tile_X0Y7_UI_IN_TT_PROJECT1
port 726 nsew signal output
flabel metal3 s 0 70436 96 70516 0 FreeSans 320 0 0 0 Tile_X0Y7_UI_IN_TT_PROJECT2
port 727 nsew signal output
flabel metal3 s 0 70940 96 71020 0 FreeSans 320 0 0 0 Tile_X0Y7_UI_IN_TT_PROJECT3
port 728 nsew signal output
flabel metal3 s 0 71444 96 71524 0 FreeSans 320 0 0 0 Tile_X0Y7_UI_IN_TT_PROJECT4
port 729 nsew signal output
flabel metal3 s 0 71948 96 72028 0 FreeSans 320 0 0 0 Tile_X0Y7_UI_IN_TT_PROJECT5
port 730 nsew signal output
flabel metal3 s 0 72452 96 72532 0 FreeSans 320 0 0 0 Tile_X0Y7_UI_IN_TT_PROJECT6
port 731 nsew signal output
flabel metal3 s 0 72956 96 73036 0 FreeSans 320 0 0 0 Tile_X0Y7_UI_IN_TT_PROJECT7
port 732 nsew signal output
flabel metal3 s 0 57332 96 57412 0 FreeSans 320 0 0 0 Tile_X0Y7_UO_OUT_TT_PROJECT0
port 733 nsew signal input
flabel metal3 s 0 57836 96 57916 0 FreeSans 320 0 0 0 Tile_X0Y7_UO_OUT_TT_PROJECT1
port 734 nsew signal input
flabel metal3 s 0 58340 96 58420 0 FreeSans 320 0 0 0 Tile_X0Y7_UO_OUT_TT_PROJECT2
port 735 nsew signal input
flabel metal3 s 0 58844 96 58924 0 FreeSans 320 0 0 0 Tile_X0Y7_UO_OUT_TT_PROJECT3
port 736 nsew signal input
flabel metal3 s 0 59348 96 59428 0 FreeSans 320 0 0 0 Tile_X0Y7_UO_OUT_TT_PROJECT4
port 737 nsew signal input
flabel metal3 s 0 59852 96 59932 0 FreeSans 320 0 0 0 Tile_X0Y7_UO_OUT_TT_PROJECT5
port 738 nsew signal input
flabel metal3 s 0 60356 96 60436 0 FreeSans 320 0 0 0 Tile_X0Y7_UO_OUT_TT_PROJECT6
port 739 nsew signal input
flabel metal3 s 0 60860 96 60940 0 FreeSans 320 0 0 0 Tile_X0Y7_UO_OUT_TT_PROJECT7
port 740 nsew signal input
flabel metal3 s 0 34988 96 35068 0 FreeSans 320 0 0 0 Tile_X0Y8_CLK_TT_PROJECT
port 741 nsew signal output
flabel metal3 s 0 34484 96 34564 0 FreeSans 320 0 0 0 Tile_X0Y8_ENA_TT_PROJECT
port 742 nsew signal output
flabel metal3 s 0 35492 96 35572 0 FreeSans 320 0 0 0 Tile_X0Y8_RST_N_TT_PROJECT
port 743 nsew signal output
flabel metal3 s 0 30452 96 30532 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_IN_TT_PROJECT0
port 744 nsew signal output
flabel metal3 s 0 30956 96 31036 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_IN_TT_PROJECT1
port 745 nsew signal output
flabel metal3 s 0 31460 96 31540 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_IN_TT_PROJECT2
port 746 nsew signal output
flabel metal3 s 0 31964 96 32044 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_IN_TT_PROJECT3
port 747 nsew signal output
flabel metal3 s 0 32468 96 32548 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_IN_TT_PROJECT4
port 748 nsew signal output
flabel metal3 s 0 32972 96 33052 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_IN_TT_PROJECT5
port 749 nsew signal output
flabel metal3 s 0 33476 96 33556 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_IN_TT_PROJECT6
port 750 nsew signal output
flabel metal3 s 0 33980 96 34060 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_IN_TT_PROJECT7
port 751 nsew signal output
flabel metal3 s 0 22388 96 22468 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OE_TT_PROJECT0
port 752 nsew signal input
flabel metal3 s 0 22892 96 22972 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OE_TT_PROJECT1
port 753 nsew signal input
flabel metal3 s 0 23396 96 23476 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OE_TT_PROJECT2
port 754 nsew signal input
flabel metal3 s 0 23900 96 23980 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OE_TT_PROJECT3
port 755 nsew signal input
flabel metal3 s 0 24404 96 24484 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OE_TT_PROJECT4
port 756 nsew signal input
flabel metal3 s 0 24908 96 24988 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OE_TT_PROJECT5
port 757 nsew signal input
flabel metal3 s 0 25412 96 25492 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OE_TT_PROJECT6
port 758 nsew signal input
flabel metal3 s 0 25916 96 25996 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OE_TT_PROJECT7
port 759 nsew signal input
flabel metal3 s 0 18356 96 18436 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OUT_TT_PROJECT0
port 760 nsew signal input
flabel metal3 s 0 18860 96 18940 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OUT_TT_PROJECT1
port 761 nsew signal input
flabel metal3 s 0 19364 96 19444 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OUT_TT_PROJECT2
port 762 nsew signal input
flabel metal3 s 0 19868 96 19948 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OUT_TT_PROJECT3
port 763 nsew signal input
flabel metal3 s 0 20372 96 20452 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OUT_TT_PROJECT4
port 764 nsew signal input
flabel metal3 s 0 20876 96 20956 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OUT_TT_PROJECT5
port 765 nsew signal input
flabel metal3 s 0 21380 96 21460 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OUT_TT_PROJECT6
port 766 nsew signal input
flabel metal3 s 0 21884 96 21964 0 FreeSans 320 0 0 0 Tile_X0Y8_UIO_OUT_TT_PROJECT7
port 767 nsew signal input
flabel metal3 s 0 26420 96 26500 0 FreeSans 320 0 0 0 Tile_X0Y8_UI_IN_TT_PROJECT0
port 768 nsew signal output
flabel metal3 s 0 26924 96 27004 0 FreeSans 320 0 0 0 Tile_X0Y8_UI_IN_TT_PROJECT1
port 769 nsew signal output
flabel metal3 s 0 27428 96 27508 0 FreeSans 320 0 0 0 Tile_X0Y8_UI_IN_TT_PROJECT2
port 770 nsew signal output
flabel metal3 s 0 27932 96 28012 0 FreeSans 320 0 0 0 Tile_X0Y8_UI_IN_TT_PROJECT3
port 771 nsew signal output
flabel metal3 s 0 28436 96 28516 0 FreeSans 320 0 0 0 Tile_X0Y8_UI_IN_TT_PROJECT4
port 772 nsew signal output
flabel metal3 s 0 28940 96 29020 0 FreeSans 320 0 0 0 Tile_X0Y8_UI_IN_TT_PROJECT5
port 773 nsew signal output
flabel metal3 s 0 29444 96 29524 0 FreeSans 320 0 0 0 Tile_X0Y8_UI_IN_TT_PROJECT6
port 774 nsew signal output
flabel metal3 s 0 29948 96 30028 0 FreeSans 320 0 0 0 Tile_X0Y8_UI_IN_TT_PROJECT7
port 775 nsew signal output
flabel metal3 s 0 14324 96 14404 0 FreeSans 320 0 0 0 Tile_X0Y8_UO_OUT_TT_PROJECT0
port 776 nsew signal input
flabel metal3 s 0 14828 96 14908 0 FreeSans 320 0 0 0 Tile_X0Y8_UO_OUT_TT_PROJECT1
port 777 nsew signal input
flabel metal3 s 0 15332 96 15412 0 FreeSans 320 0 0 0 Tile_X0Y8_UO_OUT_TT_PROJECT2
port 778 nsew signal input
flabel metal3 s 0 15836 96 15916 0 FreeSans 320 0 0 0 Tile_X0Y8_UO_OUT_TT_PROJECT3
port 779 nsew signal input
flabel metal3 s 0 16340 96 16420 0 FreeSans 320 0 0 0 Tile_X0Y8_UO_OUT_TT_PROJECT4
port 780 nsew signal input
flabel metal3 s 0 16844 96 16924 0 FreeSans 320 0 0 0 Tile_X0Y8_UO_OUT_TT_PROJECT5
port 781 nsew signal input
flabel metal3 s 0 17348 96 17428 0 FreeSans 320 0 0 0 Tile_X0Y8_UO_OUT_TT_PROJECT6
port 782 nsew signal input
flabel metal3 s 0 17852 96 17932 0 FreeSans 320 0 0 0 Tile_X0Y8_UO_OUT_TT_PROJECT7
port 783 nsew signal input
flabel metal2 s 25688 366408 25768 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_A_I_top
port 784 nsew signal output
flabel metal2 s 24536 366408 24616 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_A_O_top
port 785 nsew signal input
flabel metal2 s 26840 366408 26920 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_A_T_top
port 786 nsew signal output
flabel metal2 s 29144 366408 29224 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_B_I_top
port 787 nsew signal output
flabel metal2 s 27992 366408 28072 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_B_O_top
port 788 nsew signal input
flabel metal2 s 30296 366408 30376 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_B_T_top
port 789 nsew signal output
flabel metal2 s 32600 366408 32680 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_C_I_top
port 790 nsew signal output
flabel metal2 s 31448 366408 31528 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_C_O_top
port 791 nsew signal input
flabel metal2 s 33752 366408 33832 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_C_T_top
port 792 nsew signal output
flabel metal2 s 36056 366408 36136 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_D_I_top
port 793 nsew signal output
flabel metal2 s 34904 366408 34984 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_D_O_top
port 794 nsew signal input
flabel metal2 s 37208 366408 37288 366504 0 FreeSans 640 0 0 0 Tile_X1Y0_D_T_top
port 795 nsew signal output
flabel metal2 s 25688 0 25768 96 0 FreeSans 640 0 0 0 Tile_X1Y9_A_I_top
port 796 nsew signal output
flabel metal2 s 24536 0 24616 96 0 FreeSans 640 0 0 0 Tile_X1Y9_A_O_top
port 797 nsew signal input
flabel metal2 s 26840 0 26920 96 0 FreeSans 640 0 0 0 Tile_X1Y9_A_T_top
port 798 nsew signal output
flabel metal2 s 29144 0 29224 96 0 FreeSans 640 0 0 0 Tile_X1Y9_B_I_top
port 799 nsew signal output
flabel metal2 s 27992 0 28072 96 0 FreeSans 640 0 0 0 Tile_X1Y9_B_O_top
port 800 nsew signal input
flabel metal2 s 30296 0 30376 96 0 FreeSans 640 0 0 0 Tile_X1Y9_B_T_top
port 801 nsew signal output
flabel metal2 s 32600 0 32680 96 0 FreeSans 640 0 0 0 Tile_X1Y9_C_I_top
port 802 nsew signal output
flabel metal2 s 31448 0 31528 96 0 FreeSans 640 0 0 0 Tile_X1Y9_C_O_top
port 803 nsew signal input
flabel metal2 s 33752 0 33832 96 0 FreeSans 640 0 0 0 Tile_X1Y9_C_T_top
port 804 nsew signal output
flabel metal2 s 36056 0 36136 96 0 FreeSans 640 0 0 0 Tile_X1Y9_D_I_top
port 805 nsew signal output
flabel metal2 s 34904 0 34984 96 0 FreeSans 640 0 0 0 Tile_X1Y9_D_O_top
port 806 nsew signal input
flabel metal2 s 37208 0 37288 96 0 FreeSans 640 0 0 0 Tile_X1Y9_D_T_top
port 807 nsew signal output
flabel metal2 s 68696 366408 68776 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_A_I_top
port 808 nsew signal output
flabel metal2 s 67544 366408 67624 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_A_O_top
port 809 nsew signal input
flabel metal2 s 69848 366408 69928 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_A_T_top
port 810 nsew signal output
flabel metal2 s 72152 366408 72232 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_B_I_top
port 811 nsew signal output
flabel metal2 s 71000 366408 71080 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_B_O_top
port 812 nsew signal input
flabel metal2 s 73304 366408 73384 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_B_T_top
port 813 nsew signal output
flabel metal2 s 75608 366408 75688 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_C_I_top
port 814 nsew signal output
flabel metal2 s 74456 366408 74536 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_C_O_top
port 815 nsew signal input
flabel metal2 s 76760 366408 76840 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_C_T_top
port 816 nsew signal output
flabel metal2 s 79064 366408 79144 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_D_I_top
port 817 nsew signal output
flabel metal2 s 77912 366408 77992 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_D_O_top
port 818 nsew signal input
flabel metal2 s 80216 366408 80296 366504 0 FreeSans 640 0 0 0 Tile_X2Y0_D_T_top
port 819 nsew signal output
flabel metal2 s 68696 0 68776 96 0 FreeSans 640 0 0 0 Tile_X2Y9_A_I_top
port 820 nsew signal output
flabel metal2 s 67544 0 67624 96 0 FreeSans 640 0 0 0 Tile_X2Y9_A_O_top
port 821 nsew signal input
flabel metal2 s 69848 0 69928 96 0 FreeSans 640 0 0 0 Tile_X2Y9_A_T_top
port 822 nsew signal output
flabel metal2 s 72152 0 72232 96 0 FreeSans 640 0 0 0 Tile_X2Y9_B_I_top
port 823 nsew signal output
flabel metal2 s 71000 0 71080 96 0 FreeSans 640 0 0 0 Tile_X2Y9_B_O_top
port 824 nsew signal input
flabel metal2 s 73304 0 73384 96 0 FreeSans 640 0 0 0 Tile_X2Y9_B_T_top
port 825 nsew signal output
flabel metal2 s 75608 0 75688 96 0 FreeSans 640 0 0 0 Tile_X2Y9_C_I_top
port 826 nsew signal output
flabel metal2 s 74456 0 74536 96 0 FreeSans 640 0 0 0 Tile_X2Y9_C_O_top
port 827 nsew signal input
flabel metal2 s 76760 0 76840 96 0 FreeSans 640 0 0 0 Tile_X2Y9_C_T_top
port 828 nsew signal output
flabel metal2 s 79064 0 79144 96 0 FreeSans 640 0 0 0 Tile_X2Y9_D_I_top
port 829 nsew signal output
flabel metal2 s 77912 0 77992 96 0 FreeSans 640 0 0 0 Tile_X2Y9_D_O_top
port 830 nsew signal input
flabel metal2 s 80216 0 80296 96 0 FreeSans 640 0 0 0 Tile_X2Y9_D_T_top
port 831 nsew signal output
flabel metal2 s 111704 366408 111784 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_A_I_top
port 832 nsew signal output
flabel metal2 s 110552 366408 110632 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_A_O_top
port 833 nsew signal input
flabel metal2 s 112856 366408 112936 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_A_T_top
port 834 nsew signal output
flabel metal2 s 115160 366408 115240 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_B_I_top
port 835 nsew signal output
flabel metal2 s 114008 366408 114088 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_B_O_top
port 836 nsew signal input
flabel metal2 s 116312 366408 116392 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_B_T_top
port 837 nsew signal output
flabel metal2 s 118616 366408 118696 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_C_I_top
port 838 nsew signal output
flabel metal2 s 117464 366408 117544 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_C_O_top
port 839 nsew signal input
flabel metal2 s 119768 366408 119848 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_C_T_top
port 840 nsew signal output
flabel metal2 s 122072 366408 122152 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_D_I_top
port 841 nsew signal output
flabel metal2 s 120920 366408 121000 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_D_O_top
port 842 nsew signal input
flabel metal2 s 123224 366408 123304 366504 0 FreeSans 640 0 0 0 Tile_X3Y0_D_T_top
port 843 nsew signal output
flabel metal2 s 111704 0 111784 96 0 FreeSans 640 0 0 0 Tile_X3Y9_A_I_top
port 844 nsew signal output
flabel metal2 s 110552 0 110632 96 0 FreeSans 640 0 0 0 Tile_X3Y9_A_O_top
port 845 nsew signal input
flabel metal2 s 112856 0 112936 96 0 FreeSans 640 0 0 0 Tile_X3Y9_A_T_top
port 846 nsew signal output
flabel metal2 s 115160 0 115240 96 0 FreeSans 640 0 0 0 Tile_X3Y9_B_I_top
port 847 nsew signal output
flabel metal2 s 114008 0 114088 96 0 FreeSans 640 0 0 0 Tile_X3Y9_B_O_top
port 848 nsew signal input
flabel metal2 s 116312 0 116392 96 0 FreeSans 640 0 0 0 Tile_X3Y9_B_T_top
port 849 nsew signal output
flabel metal2 s 118616 0 118696 96 0 FreeSans 640 0 0 0 Tile_X3Y9_C_I_top
port 850 nsew signal output
flabel metal2 s 117464 0 117544 96 0 FreeSans 640 0 0 0 Tile_X3Y9_C_O_top
port 851 nsew signal input
flabel metal2 s 119768 0 119848 96 0 FreeSans 640 0 0 0 Tile_X3Y9_C_T_top
port 852 nsew signal output
flabel metal2 s 122072 0 122152 96 0 FreeSans 640 0 0 0 Tile_X3Y9_D_I_top
port 853 nsew signal output
flabel metal2 s 120920 0 121000 96 0 FreeSans 640 0 0 0 Tile_X3Y9_D_O_top
port 854 nsew signal input
flabel metal2 s 123224 0 123304 96 0 FreeSans 640 0 0 0 Tile_X3Y9_D_T_top
port 855 nsew signal output
flabel metal2 s 154712 366408 154792 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_A_I_top
port 856 nsew signal output
flabel metal2 s 153560 366408 153640 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_A_O_top
port 857 nsew signal input
flabel metal2 s 155864 366408 155944 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_A_T_top
port 858 nsew signal output
flabel metal2 s 158168 366408 158248 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_B_I_top
port 859 nsew signal output
flabel metal2 s 157016 366408 157096 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_B_O_top
port 860 nsew signal input
flabel metal2 s 159320 366408 159400 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_B_T_top
port 861 nsew signal output
flabel metal2 s 161624 366408 161704 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_C_I_top
port 862 nsew signal output
flabel metal2 s 160472 366408 160552 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_C_O_top
port 863 nsew signal input
flabel metal2 s 162776 366408 162856 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_C_T_top
port 864 nsew signal output
flabel metal2 s 165080 366408 165160 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_D_I_top
port 865 nsew signal output
flabel metal2 s 163928 366408 164008 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_D_O_top
port 866 nsew signal input
flabel metal2 s 166232 366408 166312 366504 0 FreeSans 640 0 0 0 Tile_X4Y0_D_T_top
port 867 nsew signal output
flabel metal2 s 154712 0 154792 96 0 FreeSans 640 0 0 0 Tile_X4Y9_A_I_top
port 868 nsew signal output
flabel metal2 s 153560 0 153640 96 0 FreeSans 640 0 0 0 Tile_X4Y9_A_O_top
port 869 nsew signal input
flabel metal2 s 155864 0 155944 96 0 FreeSans 640 0 0 0 Tile_X4Y9_A_T_top
port 870 nsew signal output
flabel metal2 s 158168 0 158248 96 0 FreeSans 640 0 0 0 Tile_X4Y9_B_I_top
port 871 nsew signal output
flabel metal2 s 157016 0 157096 96 0 FreeSans 640 0 0 0 Tile_X4Y9_B_O_top
port 872 nsew signal input
flabel metal2 s 159320 0 159400 96 0 FreeSans 640 0 0 0 Tile_X4Y9_B_T_top
port 873 nsew signal output
flabel metal2 s 161624 0 161704 96 0 FreeSans 640 0 0 0 Tile_X4Y9_C_I_top
port 874 nsew signal output
flabel metal2 s 160472 0 160552 96 0 FreeSans 640 0 0 0 Tile_X4Y9_C_O_top
port 875 nsew signal input
flabel metal2 s 162776 0 162856 96 0 FreeSans 640 0 0 0 Tile_X4Y9_C_T_top
port 876 nsew signal output
flabel metal2 s 165080 0 165160 96 0 FreeSans 640 0 0 0 Tile_X4Y9_D_I_top
port 877 nsew signal output
flabel metal2 s 163928 0 164008 96 0 FreeSans 640 0 0 0 Tile_X4Y9_D_O_top
port 878 nsew signal input
flabel metal2 s 166232 0 166312 96 0 FreeSans 640 0 0 0 Tile_X4Y9_D_T_top
port 879 nsew signal output
flabel metal3 s 215136 294044 215232 294124 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM0
port 880 nsew signal output
flabel metal3 s 215136 294380 215232 294460 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM1
port 881 nsew signal output
flabel metal3 s 215136 294716 215232 294796 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM2
port 882 nsew signal output
flabel metal3 s 215136 295052 215232 295132 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM3
port 883 nsew signal output
flabel metal3 s 215136 295388 215232 295468 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM4
port 884 nsew signal output
flabel metal3 s 215136 295724 215232 295804 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM5
port 885 nsew signal output
flabel metal3 s 215136 296060 215232 296140 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM6
port 886 nsew signal output
flabel metal3 s 215136 296396 215232 296476 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM7
port 887 nsew signal output
flabel metal3 s 215136 296732 215232 296812 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM8
port 888 nsew signal output
flabel metal3 s 215136 297068 215232 297148 0 FreeSans 320 0 0 0 Tile_X5Y2_ADDR_SRAM9
port 889 nsew signal output
flabel metal3 s 215136 308156 215232 308236 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM0
port 890 nsew signal output
flabel metal3 s 215136 308492 215232 308572 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM1
port 891 nsew signal output
flabel metal3 s 215136 311516 215232 311596 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM10
port 892 nsew signal output
flabel metal3 s 215136 311852 215232 311932 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM11
port 893 nsew signal output
flabel metal3 s 215136 312188 215232 312268 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM12
port 894 nsew signal output
flabel metal3 s 215136 312524 215232 312604 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM13
port 895 nsew signal output
flabel metal3 s 215136 312860 215232 312940 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM14
port 896 nsew signal output
flabel metal3 s 215136 313196 215232 313276 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM15
port 897 nsew signal output
flabel metal3 s 215136 313532 215232 313612 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM16
port 898 nsew signal output
flabel metal3 s 215136 313868 215232 313948 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM17
port 899 nsew signal output
flabel metal3 s 215136 314204 215232 314284 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM18
port 900 nsew signal output
flabel metal3 s 215136 314540 215232 314620 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM19
port 901 nsew signal output
flabel metal3 s 215136 308828 215232 308908 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM2
port 902 nsew signal output
flabel metal3 s 215136 314876 215232 314956 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM20
port 903 nsew signal output
flabel metal3 s 215136 315212 215232 315292 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM21
port 904 nsew signal output
flabel metal3 s 215136 315548 215232 315628 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM22
port 905 nsew signal output
flabel metal3 s 215136 315884 215232 315964 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM23
port 906 nsew signal output
flabel metal3 s 215136 316220 215232 316300 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM24
port 907 nsew signal output
flabel metal3 s 215136 316556 215232 316636 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM25
port 908 nsew signal output
flabel metal3 s 215136 316892 215232 316972 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM26
port 909 nsew signal output
flabel metal3 s 215136 317228 215232 317308 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM27
port 910 nsew signal output
flabel metal3 s 215136 317564 215232 317644 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM28
port 911 nsew signal output
flabel metal3 s 215136 317900 215232 317980 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM29
port 912 nsew signal output
flabel metal3 s 215136 309164 215232 309244 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM3
port 913 nsew signal output
flabel metal3 s 215136 318236 215232 318316 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM30
port 914 nsew signal output
flabel metal3 s 215136 318572 215232 318652 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM31
port 915 nsew signal output
flabel metal3 s 215136 309500 215232 309580 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM4
port 916 nsew signal output
flabel metal3 s 215136 309836 215232 309916 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM5
port 917 nsew signal output
flabel metal3 s 215136 310172 215232 310252 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM6
port 918 nsew signal output
flabel metal3 s 215136 310508 215232 310588 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM7
port 919 nsew signal output
flabel metal3 s 215136 310844 215232 310924 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM8
port 920 nsew signal output
flabel metal3 s 215136 311180 215232 311260 0 FreeSans 320 0 0 0 Tile_X5Y2_BM_SRAM9
port 921 nsew signal output
flabel metal3 s 215136 319916 215232 319996 0 FreeSans 320 0 0 0 Tile_X5Y2_CLK_SRAM
port 922 nsew signal output
flabel metal3 s 215136 293708 215232 293788 0 FreeSans 320 0 0 0 Tile_X5Y2_CONFIGURED_top
port 923 nsew signal input
flabel metal3 s 215136 297404 215232 297484 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM0
port 924 nsew signal output
flabel metal3 s 215136 297740 215232 297820 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM1
port 925 nsew signal output
flabel metal3 s 215136 300764 215232 300844 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM10
port 926 nsew signal output
flabel metal3 s 215136 301100 215232 301180 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM11
port 927 nsew signal output
flabel metal3 s 215136 301436 215232 301516 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM12
port 928 nsew signal output
flabel metal3 s 215136 301772 215232 301852 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM13
port 929 nsew signal output
flabel metal3 s 215136 302108 215232 302188 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM14
port 930 nsew signal output
flabel metal3 s 215136 302444 215232 302524 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM15
port 931 nsew signal output
flabel metal3 s 215136 302780 215232 302860 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM16
port 932 nsew signal output
flabel metal3 s 215136 303116 215232 303196 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM17
port 933 nsew signal output
flabel metal3 s 215136 303452 215232 303532 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM18
port 934 nsew signal output
flabel metal3 s 215136 303788 215232 303868 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM19
port 935 nsew signal output
flabel metal3 s 215136 298076 215232 298156 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM2
port 936 nsew signal output
flabel metal3 s 215136 304124 215232 304204 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM20
port 937 nsew signal output
flabel metal3 s 215136 304460 215232 304540 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM21
port 938 nsew signal output
flabel metal3 s 215136 304796 215232 304876 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM22
port 939 nsew signal output
flabel metal3 s 215136 305132 215232 305212 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM23
port 940 nsew signal output
flabel metal3 s 215136 305468 215232 305548 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM24
port 941 nsew signal output
flabel metal3 s 215136 305804 215232 305884 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM25
port 942 nsew signal output
flabel metal3 s 215136 306140 215232 306220 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM26
port 943 nsew signal output
flabel metal3 s 215136 306476 215232 306556 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM27
port 944 nsew signal output
flabel metal3 s 215136 306812 215232 306892 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM28
port 945 nsew signal output
flabel metal3 s 215136 307148 215232 307228 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM29
port 946 nsew signal output
flabel metal3 s 215136 298412 215232 298492 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM3
port 947 nsew signal output
flabel metal3 s 215136 307484 215232 307564 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM30
port 948 nsew signal output
flabel metal3 s 215136 307820 215232 307900 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM31
port 949 nsew signal output
flabel metal3 s 215136 298748 215232 298828 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM4
port 950 nsew signal output
flabel metal3 s 215136 299084 215232 299164 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM5
port 951 nsew signal output
flabel metal3 s 215136 299420 215232 299500 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM6
port 952 nsew signal output
flabel metal3 s 215136 299756 215232 299836 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM7
port 953 nsew signal output
flabel metal3 s 215136 300092 215232 300172 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM8
port 954 nsew signal output
flabel metal3 s 215136 300428 215232 300508 0 FreeSans 320 0 0 0 Tile_X5Y2_DIN_SRAM9
port 955 nsew signal output
flabel metal3 s 215136 282956 215232 283036 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM0
port 956 nsew signal input
flabel metal3 s 215136 283292 215232 283372 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM1
port 957 nsew signal input
flabel metal3 s 215136 286316 215232 286396 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM10
port 958 nsew signal input
flabel metal3 s 215136 286652 215232 286732 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM11
port 959 nsew signal input
flabel metal3 s 215136 286988 215232 287068 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM12
port 960 nsew signal input
flabel metal3 s 215136 287324 215232 287404 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM13
port 961 nsew signal input
flabel metal3 s 215136 287660 215232 287740 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM14
port 962 nsew signal input
flabel metal3 s 215136 287996 215232 288076 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM15
port 963 nsew signal input
flabel metal3 s 215136 288332 215232 288412 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM16
port 964 nsew signal input
flabel metal3 s 215136 288668 215232 288748 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM17
port 965 nsew signal input
flabel metal3 s 215136 289004 215232 289084 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM18
port 966 nsew signal input
flabel metal3 s 215136 289340 215232 289420 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM19
port 967 nsew signal input
flabel metal3 s 215136 283628 215232 283708 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM2
port 968 nsew signal input
flabel metal3 s 215136 289676 215232 289756 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM20
port 969 nsew signal input
flabel metal3 s 215136 290012 215232 290092 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM21
port 970 nsew signal input
flabel metal3 s 215136 290348 215232 290428 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM22
port 971 nsew signal input
flabel metal3 s 215136 290684 215232 290764 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM23
port 972 nsew signal input
flabel metal3 s 215136 291020 215232 291100 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM24
port 973 nsew signal input
flabel metal3 s 215136 291356 215232 291436 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM25
port 974 nsew signal input
flabel metal3 s 215136 291692 215232 291772 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM26
port 975 nsew signal input
flabel metal3 s 215136 292028 215232 292108 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM27
port 976 nsew signal input
flabel metal3 s 215136 292364 215232 292444 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM28
port 977 nsew signal input
flabel metal3 s 215136 292700 215232 292780 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM29
port 978 nsew signal input
flabel metal3 s 215136 283964 215232 284044 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM3
port 979 nsew signal input
flabel metal3 s 215136 293036 215232 293116 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM30
port 980 nsew signal input
flabel metal3 s 215136 293372 215232 293452 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM31
port 981 nsew signal input
flabel metal3 s 215136 284300 215232 284380 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM4
port 982 nsew signal input
flabel metal3 s 215136 284636 215232 284716 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM5
port 983 nsew signal input
flabel metal3 s 215136 284972 215232 285052 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM6
port 984 nsew signal input
flabel metal3 s 215136 285308 215232 285388 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM7
port 985 nsew signal input
flabel metal3 s 215136 285644 215232 285724 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM8
port 986 nsew signal input
flabel metal3 s 215136 285980 215232 286060 0 FreeSans 320 0 0 0 Tile_X5Y2_DOUT_SRAM9
port 987 nsew signal input
flabel metal3 s 215136 319244 215232 319324 0 FreeSans 320 0 0 0 Tile_X5Y2_MEN_SRAM
port 988 nsew signal output
flabel metal3 s 215136 319580 215232 319660 0 FreeSans 320 0 0 0 Tile_X5Y2_REN_SRAM
port 989 nsew signal output
flabel metal3 s 215136 320252 215232 320332 0 FreeSans 320 0 0 0 Tile_X5Y2_TIE_HIGH_SRAM
port 990 nsew signal output
flabel metal3 s 215136 320588 215232 320668 0 FreeSans 320 0 0 0 Tile_X5Y2_TIE_LOW_SRAM
port 991 nsew signal output
flabel metal3 s 215136 318908 215232 318988 0 FreeSans 320 0 0 0 Tile_X5Y2_WEN_SRAM
port 992 nsew signal output
flabel metal3 s 215136 250028 215232 250108 0 FreeSans 320 0 0 0 Tile_X5Y3_CLK_TT_PROJECT
port 993 nsew signal output
flabel metal3 s 215136 249524 215232 249604 0 FreeSans 320 0 0 0 Tile_X5Y3_ENA_TT_PROJECT
port 994 nsew signal output
flabel metal3 s 215136 250532 215232 250612 0 FreeSans 320 0 0 0 Tile_X5Y3_RST_N_TT_PROJECT
port 995 nsew signal output
flabel metal3 s 215136 245492 215232 245572 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_IN_TT_PROJECT0
port 996 nsew signal output
flabel metal3 s 215136 245996 215232 246076 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_IN_TT_PROJECT1
port 997 nsew signal output
flabel metal3 s 215136 246500 215232 246580 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_IN_TT_PROJECT2
port 998 nsew signal output
flabel metal3 s 215136 247004 215232 247084 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_IN_TT_PROJECT3
port 999 nsew signal output
flabel metal3 s 215136 247508 215232 247588 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_IN_TT_PROJECT4
port 1000 nsew signal output
flabel metal3 s 215136 248012 215232 248092 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_IN_TT_PROJECT5
port 1001 nsew signal output
flabel metal3 s 215136 248516 215232 248596 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_IN_TT_PROJECT6
port 1002 nsew signal output
flabel metal3 s 215136 249020 215232 249100 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_IN_TT_PROJECT7
port 1003 nsew signal output
flabel metal3 s 215136 237428 215232 237508 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OE_TT_PROJECT0
port 1004 nsew signal input
flabel metal3 s 215136 237932 215232 238012 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OE_TT_PROJECT1
port 1005 nsew signal input
flabel metal3 s 215136 238436 215232 238516 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OE_TT_PROJECT2
port 1006 nsew signal input
flabel metal3 s 215136 238940 215232 239020 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OE_TT_PROJECT3
port 1007 nsew signal input
flabel metal3 s 215136 239444 215232 239524 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OE_TT_PROJECT4
port 1008 nsew signal input
flabel metal3 s 215136 239948 215232 240028 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OE_TT_PROJECT5
port 1009 nsew signal input
flabel metal3 s 215136 240452 215232 240532 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OE_TT_PROJECT6
port 1010 nsew signal input
flabel metal3 s 215136 240956 215232 241036 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OE_TT_PROJECT7
port 1011 nsew signal input
flabel metal3 s 215136 233396 215232 233476 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OUT_TT_PROJECT0
port 1012 nsew signal input
flabel metal3 s 215136 233900 215232 233980 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OUT_TT_PROJECT1
port 1013 nsew signal input
flabel metal3 s 215136 234404 215232 234484 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OUT_TT_PROJECT2
port 1014 nsew signal input
flabel metal3 s 215136 234908 215232 234988 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OUT_TT_PROJECT3
port 1015 nsew signal input
flabel metal3 s 215136 235412 215232 235492 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OUT_TT_PROJECT4
port 1016 nsew signal input
flabel metal3 s 215136 235916 215232 235996 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OUT_TT_PROJECT5
port 1017 nsew signal input
flabel metal3 s 215136 236420 215232 236500 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OUT_TT_PROJECT6
port 1018 nsew signal input
flabel metal3 s 215136 236924 215232 237004 0 FreeSans 320 0 0 0 Tile_X5Y3_UIO_OUT_TT_PROJECT7
port 1019 nsew signal input
flabel metal3 s 215136 241460 215232 241540 0 FreeSans 320 0 0 0 Tile_X5Y3_UI_IN_TT_PROJECT0
port 1020 nsew signal output
flabel metal3 s 215136 241964 215232 242044 0 FreeSans 320 0 0 0 Tile_X5Y3_UI_IN_TT_PROJECT1
port 1021 nsew signal output
flabel metal3 s 215136 242468 215232 242548 0 FreeSans 320 0 0 0 Tile_X5Y3_UI_IN_TT_PROJECT2
port 1022 nsew signal output
flabel metal3 s 215136 242972 215232 243052 0 FreeSans 320 0 0 0 Tile_X5Y3_UI_IN_TT_PROJECT3
port 1023 nsew signal output
flabel metal3 s 215136 243476 215232 243556 0 FreeSans 320 0 0 0 Tile_X5Y3_UI_IN_TT_PROJECT4
port 1024 nsew signal output
flabel metal3 s 215136 243980 215232 244060 0 FreeSans 320 0 0 0 Tile_X5Y3_UI_IN_TT_PROJECT5
port 1025 nsew signal output
flabel metal3 s 215136 244484 215232 244564 0 FreeSans 320 0 0 0 Tile_X5Y3_UI_IN_TT_PROJECT6
port 1026 nsew signal output
flabel metal3 s 215136 244988 215232 245068 0 FreeSans 320 0 0 0 Tile_X5Y3_UI_IN_TT_PROJECT7
port 1027 nsew signal output
flabel metal3 s 215136 229364 215232 229444 0 FreeSans 320 0 0 0 Tile_X5Y3_UO_OUT_TT_PROJECT0
port 1028 nsew signal input
flabel metal3 s 215136 229868 215232 229948 0 FreeSans 320 0 0 0 Tile_X5Y3_UO_OUT_TT_PROJECT1
port 1029 nsew signal input
flabel metal3 s 215136 230372 215232 230452 0 FreeSans 320 0 0 0 Tile_X5Y3_UO_OUT_TT_PROJECT2
port 1030 nsew signal input
flabel metal3 s 215136 230876 215232 230956 0 FreeSans 320 0 0 0 Tile_X5Y3_UO_OUT_TT_PROJECT3
port 1031 nsew signal input
flabel metal3 s 215136 231380 215232 231460 0 FreeSans 320 0 0 0 Tile_X5Y3_UO_OUT_TT_PROJECT4
port 1032 nsew signal input
flabel metal3 s 215136 231884 215232 231964 0 FreeSans 320 0 0 0 Tile_X5Y3_UO_OUT_TT_PROJECT5
port 1033 nsew signal input
flabel metal3 s 215136 232388 215232 232468 0 FreeSans 320 0 0 0 Tile_X5Y3_UO_OUT_TT_PROJECT6
port 1034 nsew signal input
flabel metal3 s 215136 232892 215232 232972 0 FreeSans 320 0 0 0 Tile_X5Y3_UO_OUT_TT_PROJECT7
port 1035 nsew signal input
flabel metal3 s 215136 207020 215232 207100 0 FreeSans 320 0 0 0 Tile_X5Y4_CLK_TT_PROJECT
port 1036 nsew signal output
flabel metal3 s 215136 206516 215232 206596 0 FreeSans 320 0 0 0 Tile_X5Y4_ENA_TT_PROJECT
port 1037 nsew signal output
flabel metal3 s 215136 207524 215232 207604 0 FreeSans 320 0 0 0 Tile_X5Y4_RST_N_TT_PROJECT
port 1038 nsew signal output
flabel metal3 s 215136 202484 215232 202564 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_IN_TT_PROJECT0
port 1039 nsew signal output
flabel metal3 s 215136 202988 215232 203068 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_IN_TT_PROJECT1
port 1040 nsew signal output
flabel metal3 s 215136 203492 215232 203572 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_IN_TT_PROJECT2
port 1041 nsew signal output
flabel metal3 s 215136 203996 215232 204076 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_IN_TT_PROJECT3
port 1042 nsew signal output
flabel metal3 s 215136 204500 215232 204580 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_IN_TT_PROJECT4
port 1043 nsew signal output
flabel metal3 s 215136 205004 215232 205084 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_IN_TT_PROJECT5
port 1044 nsew signal output
flabel metal3 s 215136 205508 215232 205588 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_IN_TT_PROJECT6
port 1045 nsew signal output
flabel metal3 s 215136 206012 215232 206092 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_IN_TT_PROJECT7
port 1046 nsew signal output
flabel metal3 s 215136 194420 215232 194500 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OE_TT_PROJECT0
port 1047 nsew signal input
flabel metal3 s 215136 194924 215232 195004 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OE_TT_PROJECT1
port 1048 nsew signal input
flabel metal3 s 215136 195428 215232 195508 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OE_TT_PROJECT2
port 1049 nsew signal input
flabel metal3 s 215136 195932 215232 196012 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OE_TT_PROJECT3
port 1050 nsew signal input
flabel metal3 s 215136 196436 215232 196516 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OE_TT_PROJECT4
port 1051 nsew signal input
flabel metal3 s 215136 196940 215232 197020 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OE_TT_PROJECT5
port 1052 nsew signal input
flabel metal3 s 215136 197444 215232 197524 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OE_TT_PROJECT6
port 1053 nsew signal input
flabel metal3 s 215136 197948 215232 198028 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OE_TT_PROJECT7
port 1054 nsew signal input
flabel metal3 s 215136 190388 215232 190468 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OUT_TT_PROJECT0
port 1055 nsew signal input
flabel metal3 s 215136 190892 215232 190972 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OUT_TT_PROJECT1
port 1056 nsew signal input
flabel metal3 s 215136 191396 215232 191476 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OUT_TT_PROJECT2
port 1057 nsew signal input
flabel metal3 s 215136 191900 215232 191980 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OUT_TT_PROJECT3
port 1058 nsew signal input
flabel metal3 s 215136 192404 215232 192484 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OUT_TT_PROJECT4
port 1059 nsew signal input
flabel metal3 s 215136 192908 215232 192988 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OUT_TT_PROJECT5
port 1060 nsew signal input
flabel metal3 s 215136 193412 215232 193492 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OUT_TT_PROJECT6
port 1061 nsew signal input
flabel metal3 s 215136 193916 215232 193996 0 FreeSans 320 0 0 0 Tile_X5Y4_UIO_OUT_TT_PROJECT7
port 1062 nsew signal input
flabel metal3 s 215136 198452 215232 198532 0 FreeSans 320 0 0 0 Tile_X5Y4_UI_IN_TT_PROJECT0
port 1063 nsew signal output
flabel metal3 s 215136 198956 215232 199036 0 FreeSans 320 0 0 0 Tile_X5Y4_UI_IN_TT_PROJECT1
port 1064 nsew signal output
flabel metal3 s 215136 199460 215232 199540 0 FreeSans 320 0 0 0 Tile_X5Y4_UI_IN_TT_PROJECT2
port 1065 nsew signal output
flabel metal3 s 215136 199964 215232 200044 0 FreeSans 320 0 0 0 Tile_X5Y4_UI_IN_TT_PROJECT3
port 1066 nsew signal output
flabel metal3 s 215136 200468 215232 200548 0 FreeSans 320 0 0 0 Tile_X5Y4_UI_IN_TT_PROJECT4
port 1067 nsew signal output
flabel metal3 s 215136 200972 215232 201052 0 FreeSans 320 0 0 0 Tile_X5Y4_UI_IN_TT_PROJECT5
port 1068 nsew signal output
flabel metal3 s 215136 201476 215232 201556 0 FreeSans 320 0 0 0 Tile_X5Y4_UI_IN_TT_PROJECT6
port 1069 nsew signal output
flabel metal3 s 215136 201980 215232 202060 0 FreeSans 320 0 0 0 Tile_X5Y4_UI_IN_TT_PROJECT7
port 1070 nsew signal output
flabel metal3 s 215136 186356 215232 186436 0 FreeSans 320 0 0 0 Tile_X5Y4_UO_OUT_TT_PROJECT0
port 1071 nsew signal input
flabel metal3 s 215136 186860 215232 186940 0 FreeSans 320 0 0 0 Tile_X5Y4_UO_OUT_TT_PROJECT1
port 1072 nsew signal input
flabel metal3 s 215136 187364 215232 187444 0 FreeSans 320 0 0 0 Tile_X5Y4_UO_OUT_TT_PROJECT2
port 1073 nsew signal input
flabel metal3 s 215136 187868 215232 187948 0 FreeSans 320 0 0 0 Tile_X5Y4_UO_OUT_TT_PROJECT3
port 1074 nsew signal input
flabel metal3 s 215136 188372 215232 188452 0 FreeSans 320 0 0 0 Tile_X5Y4_UO_OUT_TT_PROJECT4
port 1075 nsew signal input
flabel metal3 s 215136 188876 215232 188956 0 FreeSans 320 0 0 0 Tile_X5Y4_UO_OUT_TT_PROJECT5
port 1076 nsew signal input
flabel metal3 s 215136 189380 215232 189460 0 FreeSans 320 0 0 0 Tile_X5Y4_UO_OUT_TT_PROJECT6
port 1077 nsew signal input
flabel metal3 s 215136 189884 215232 189964 0 FreeSans 320 0 0 0 Tile_X5Y4_UO_OUT_TT_PROJECT7
port 1078 nsew signal input
flabel metal3 s 215136 164012 215232 164092 0 FreeSans 320 0 0 0 Tile_X5Y5_CLK_TT_PROJECT
port 1079 nsew signal output
flabel metal3 s 215136 163508 215232 163588 0 FreeSans 320 0 0 0 Tile_X5Y5_ENA_TT_PROJECT
port 1080 nsew signal output
flabel metal3 s 215136 164516 215232 164596 0 FreeSans 320 0 0 0 Tile_X5Y5_RST_N_TT_PROJECT
port 1081 nsew signal output
flabel metal3 s 215136 159476 215232 159556 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_IN_TT_PROJECT0
port 1082 nsew signal output
flabel metal3 s 215136 159980 215232 160060 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_IN_TT_PROJECT1
port 1083 nsew signal output
flabel metal3 s 215136 160484 215232 160564 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_IN_TT_PROJECT2
port 1084 nsew signal output
flabel metal3 s 215136 160988 215232 161068 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_IN_TT_PROJECT3
port 1085 nsew signal output
flabel metal3 s 215136 161492 215232 161572 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_IN_TT_PROJECT4
port 1086 nsew signal output
flabel metal3 s 215136 161996 215232 162076 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_IN_TT_PROJECT5
port 1087 nsew signal output
flabel metal3 s 215136 162500 215232 162580 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_IN_TT_PROJECT6
port 1088 nsew signal output
flabel metal3 s 215136 163004 215232 163084 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_IN_TT_PROJECT7
port 1089 nsew signal output
flabel metal3 s 215136 151412 215232 151492 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OE_TT_PROJECT0
port 1090 nsew signal input
flabel metal3 s 215136 151916 215232 151996 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OE_TT_PROJECT1
port 1091 nsew signal input
flabel metal3 s 215136 152420 215232 152500 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OE_TT_PROJECT2
port 1092 nsew signal input
flabel metal3 s 215136 152924 215232 153004 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OE_TT_PROJECT3
port 1093 nsew signal input
flabel metal3 s 215136 153428 215232 153508 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OE_TT_PROJECT4
port 1094 nsew signal input
flabel metal3 s 215136 153932 215232 154012 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OE_TT_PROJECT5
port 1095 nsew signal input
flabel metal3 s 215136 154436 215232 154516 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OE_TT_PROJECT6
port 1096 nsew signal input
flabel metal3 s 215136 154940 215232 155020 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OE_TT_PROJECT7
port 1097 nsew signal input
flabel metal3 s 215136 147380 215232 147460 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OUT_TT_PROJECT0
port 1098 nsew signal input
flabel metal3 s 215136 147884 215232 147964 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OUT_TT_PROJECT1
port 1099 nsew signal input
flabel metal3 s 215136 148388 215232 148468 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OUT_TT_PROJECT2
port 1100 nsew signal input
flabel metal3 s 215136 148892 215232 148972 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OUT_TT_PROJECT3
port 1101 nsew signal input
flabel metal3 s 215136 149396 215232 149476 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OUT_TT_PROJECT4
port 1102 nsew signal input
flabel metal3 s 215136 149900 215232 149980 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OUT_TT_PROJECT5
port 1103 nsew signal input
flabel metal3 s 215136 150404 215232 150484 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OUT_TT_PROJECT6
port 1104 nsew signal input
flabel metal3 s 215136 150908 215232 150988 0 FreeSans 320 0 0 0 Tile_X5Y5_UIO_OUT_TT_PROJECT7
port 1105 nsew signal input
flabel metal3 s 215136 155444 215232 155524 0 FreeSans 320 0 0 0 Tile_X5Y5_UI_IN_TT_PROJECT0
port 1106 nsew signal output
flabel metal3 s 215136 155948 215232 156028 0 FreeSans 320 0 0 0 Tile_X5Y5_UI_IN_TT_PROJECT1
port 1107 nsew signal output
flabel metal3 s 215136 156452 215232 156532 0 FreeSans 320 0 0 0 Tile_X5Y5_UI_IN_TT_PROJECT2
port 1108 nsew signal output
flabel metal3 s 215136 156956 215232 157036 0 FreeSans 320 0 0 0 Tile_X5Y5_UI_IN_TT_PROJECT3
port 1109 nsew signal output
flabel metal3 s 215136 157460 215232 157540 0 FreeSans 320 0 0 0 Tile_X5Y5_UI_IN_TT_PROJECT4
port 1110 nsew signal output
flabel metal3 s 215136 157964 215232 158044 0 FreeSans 320 0 0 0 Tile_X5Y5_UI_IN_TT_PROJECT5
port 1111 nsew signal output
flabel metal3 s 215136 158468 215232 158548 0 FreeSans 320 0 0 0 Tile_X5Y5_UI_IN_TT_PROJECT6
port 1112 nsew signal output
flabel metal3 s 215136 158972 215232 159052 0 FreeSans 320 0 0 0 Tile_X5Y5_UI_IN_TT_PROJECT7
port 1113 nsew signal output
flabel metal3 s 215136 143348 215232 143428 0 FreeSans 320 0 0 0 Tile_X5Y5_UO_OUT_TT_PROJECT0
port 1114 nsew signal input
flabel metal3 s 215136 143852 215232 143932 0 FreeSans 320 0 0 0 Tile_X5Y5_UO_OUT_TT_PROJECT1
port 1115 nsew signal input
flabel metal3 s 215136 144356 215232 144436 0 FreeSans 320 0 0 0 Tile_X5Y5_UO_OUT_TT_PROJECT2
port 1116 nsew signal input
flabel metal3 s 215136 144860 215232 144940 0 FreeSans 320 0 0 0 Tile_X5Y5_UO_OUT_TT_PROJECT3
port 1117 nsew signal input
flabel metal3 s 215136 145364 215232 145444 0 FreeSans 320 0 0 0 Tile_X5Y5_UO_OUT_TT_PROJECT4
port 1118 nsew signal input
flabel metal3 s 215136 145868 215232 145948 0 FreeSans 320 0 0 0 Tile_X5Y5_UO_OUT_TT_PROJECT5
port 1119 nsew signal input
flabel metal3 s 215136 146372 215232 146452 0 FreeSans 320 0 0 0 Tile_X5Y5_UO_OUT_TT_PROJECT6
port 1120 nsew signal input
flabel metal3 s 215136 146876 215232 146956 0 FreeSans 320 0 0 0 Tile_X5Y5_UO_OUT_TT_PROJECT7
port 1121 nsew signal input
flabel metal3 s 215136 121004 215232 121084 0 FreeSans 320 0 0 0 Tile_X5Y6_CLK_TT_PROJECT
port 1122 nsew signal output
flabel metal3 s 215136 120500 215232 120580 0 FreeSans 320 0 0 0 Tile_X5Y6_ENA_TT_PROJECT
port 1123 nsew signal output
flabel metal3 s 215136 121508 215232 121588 0 FreeSans 320 0 0 0 Tile_X5Y6_RST_N_TT_PROJECT
port 1124 nsew signal output
flabel metal3 s 215136 116468 215232 116548 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_IN_TT_PROJECT0
port 1125 nsew signal output
flabel metal3 s 215136 116972 215232 117052 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_IN_TT_PROJECT1
port 1126 nsew signal output
flabel metal3 s 215136 117476 215232 117556 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_IN_TT_PROJECT2
port 1127 nsew signal output
flabel metal3 s 215136 117980 215232 118060 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_IN_TT_PROJECT3
port 1128 nsew signal output
flabel metal3 s 215136 118484 215232 118564 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_IN_TT_PROJECT4
port 1129 nsew signal output
flabel metal3 s 215136 118988 215232 119068 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_IN_TT_PROJECT5
port 1130 nsew signal output
flabel metal3 s 215136 119492 215232 119572 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_IN_TT_PROJECT6
port 1131 nsew signal output
flabel metal3 s 215136 119996 215232 120076 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_IN_TT_PROJECT7
port 1132 nsew signal output
flabel metal3 s 215136 108404 215232 108484 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OE_TT_PROJECT0
port 1133 nsew signal input
flabel metal3 s 215136 108908 215232 108988 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OE_TT_PROJECT1
port 1134 nsew signal input
flabel metal3 s 215136 109412 215232 109492 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OE_TT_PROJECT2
port 1135 nsew signal input
flabel metal3 s 215136 109916 215232 109996 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OE_TT_PROJECT3
port 1136 nsew signal input
flabel metal3 s 215136 110420 215232 110500 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OE_TT_PROJECT4
port 1137 nsew signal input
flabel metal3 s 215136 110924 215232 111004 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OE_TT_PROJECT5
port 1138 nsew signal input
flabel metal3 s 215136 111428 215232 111508 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OE_TT_PROJECT6
port 1139 nsew signal input
flabel metal3 s 215136 111932 215232 112012 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OE_TT_PROJECT7
port 1140 nsew signal input
flabel metal3 s 215136 104372 215232 104452 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OUT_TT_PROJECT0
port 1141 nsew signal input
flabel metal3 s 215136 104876 215232 104956 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OUT_TT_PROJECT1
port 1142 nsew signal input
flabel metal3 s 215136 105380 215232 105460 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OUT_TT_PROJECT2
port 1143 nsew signal input
flabel metal3 s 215136 105884 215232 105964 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OUT_TT_PROJECT3
port 1144 nsew signal input
flabel metal3 s 215136 106388 215232 106468 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OUT_TT_PROJECT4
port 1145 nsew signal input
flabel metal3 s 215136 106892 215232 106972 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OUT_TT_PROJECT5
port 1146 nsew signal input
flabel metal3 s 215136 107396 215232 107476 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OUT_TT_PROJECT6
port 1147 nsew signal input
flabel metal3 s 215136 107900 215232 107980 0 FreeSans 320 0 0 0 Tile_X5Y6_UIO_OUT_TT_PROJECT7
port 1148 nsew signal input
flabel metal3 s 215136 112436 215232 112516 0 FreeSans 320 0 0 0 Tile_X5Y6_UI_IN_TT_PROJECT0
port 1149 nsew signal output
flabel metal3 s 215136 112940 215232 113020 0 FreeSans 320 0 0 0 Tile_X5Y6_UI_IN_TT_PROJECT1
port 1150 nsew signal output
flabel metal3 s 215136 113444 215232 113524 0 FreeSans 320 0 0 0 Tile_X5Y6_UI_IN_TT_PROJECT2
port 1151 nsew signal output
flabel metal3 s 215136 113948 215232 114028 0 FreeSans 320 0 0 0 Tile_X5Y6_UI_IN_TT_PROJECT3
port 1152 nsew signal output
flabel metal3 s 215136 114452 215232 114532 0 FreeSans 320 0 0 0 Tile_X5Y6_UI_IN_TT_PROJECT4
port 1153 nsew signal output
flabel metal3 s 215136 114956 215232 115036 0 FreeSans 320 0 0 0 Tile_X5Y6_UI_IN_TT_PROJECT5
port 1154 nsew signal output
flabel metal3 s 215136 115460 215232 115540 0 FreeSans 320 0 0 0 Tile_X5Y6_UI_IN_TT_PROJECT6
port 1155 nsew signal output
flabel metal3 s 215136 115964 215232 116044 0 FreeSans 320 0 0 0 Tile_X5Y6_UI_IN_TT_PROJECT7
port 1156 nsew signal output
flabel metal3 s 215136 100340 215232 100420 0 FreeSans 320 0 0 0 Tile_X5Y6_UO_OUT_TT_PROJECT0
port 1157 nsew signal input
flabel metal3 s 215136 100844 215232 100924 0 FreeSans 320 0 0 0 Tile_X5Y6_UO_OUT_TT_PROJECT1
port 1158 nsew signal input
flabel metal3 s 215136 101348 215232 101428 0 FreeSans 320 0 0 0 Tile_X5Y6_UO_OUT_TT_PROJECT2
port 1159 nsew signal input
flabel metal3 s 215136 101852 215232 101932 0 FreeSans 320 0 0 0 Tile_X5Y6_UO_OUT_TT_PROJECT3
port 1160 nsew signal input
flabel metal3 s 215136 102356 215232 102436 0 FreeSans 320 0 0 0 Tile_X5Y6_UO_OUT_TT_PROJECT4
port 1161 nsew signal input
flabel metal3 s 215136 102860 215232 102940 0 FreeSans 320 0 0 0 Tile_X5Y6_UO_OUT_TT_PROJECT5
port 1162 nsew signal input
flabel metal3 s 215136 103364 215232 103444 0 FreeSans 320 0 0 0 Tile_X5Y6_UO_OUT_TT_PROJECT6
port 1163 nsew signal input
flabel metal3 s 215136 103868 215232 103948 0 FreeSans 320 0 0 0 Tile_X5Y6_UO_OUT_TT_PROJECT7
port 1164 nsew signal input
flabel metal3 s 215136 77996 215232 78076 0 FreeSans 320 0 0 0 Tile_X5Y7_CLK_TT_PROJECT
port 1165 nsew signal output
flabel metal3 s 215136 77492 215232 77572 0 FreeSans 320 0 0 0 Tile_X5Y7_ENA_TT_PROJECT
port 1166 nsew signal output
flabel metal3 s 215136 78500 215232 78580 0 FreeSans 320 0 0 0 Tile_X5Y7_RST_N_TT_PROJECT
port 1167 nsew signal output
flabel metal3 s 215136 73460 215232 73540 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_IN_TT_PROJECT0
port 1168 nsew signal output
flabel metal3 s 215136 73964 215232 74044 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_IN_TT_PROJECT1
port 1169 nsew signal output
flabel metal3 s 215136 74468 215232 74548 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_IN_TT_PROJECT2
port 1170 nsew signal output
flabel metal3 s 215136 74972 215232 75052 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_IN_TT_PROJECT3
port 1171 nsew signal output
flabel metal3 s 215136 75476 215232 75556 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_IN_TT_PROJECT4
port 1172 nsew signal output
flabel metal3 s 215136 75980 215232 76060 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_IN_TT_PROJECT5
port 1173 nsew signal output
flabel metal3 s 215136 76484 215232 76564 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_IN_TT_PROJECT6
port 1174 nsew signal output
flabel metal3 s 215136 76988 215232 77068 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_IN_TT_PROJECT7
port 1175 nsew signal output
flabel metal3 s 215136 65396 215232 65476 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OE_TT_PROJECT0
port 1176 nsew signal input
flabel metal3 s 215136 65900 215232 65980 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OE_TT_PROJECT1
port 1177 nsew signal input
flabel metal3 s 215136 66404 215232 66484 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OE_TT_PROJECT2
port 1178 nsew signal input
flabel metal3 s 215136 66908 215232 66988 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OE_TT_PROJECT3
port 1179 nsew signal input
flabel metal3 s 215136 67412 215232 67492 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OE_TT_PROJECT4
port 1180 nsew signal input
flabel metal3 s 215136 67916 215232 67996 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OE_TT_PROJECT5
port 1181 nsew signal input
flabel metal3 s 215136 68420 215232 68500 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OE_TT_PROJECT6
port 1182 nsew signal input
flabel metal3 s 215136 68924 215232 69004 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OE_TT_PROJECT7
port 1183 nsew signal input
flabel metal3 s 215136 61364 215232 61444 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OUT_TT_PROJECT0
port 1184 nsew signal input
flabel metal3 s 215136 61868 215232 61948 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OUT_TT_PROJECT1
port 1185 nsew signal input
flabel metal3 s 215136 62372 215232 62452 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OUT_TT_PROJECT2
port 1186 nsew signal input
flabel metal3 s 215136 62876 215232 62956 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OUT_TT_PROJECT3
port 1187 nsew signal input
flabel metal3 s 215136 63380 215232 63460 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OUT_TT_PROJECT4
port 1188 nsew signal input
flabel metal3 s 215136 63884 215232 63964 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OUT_TT_PROJECT5
port 1189 nsew signal input
flabel metal3 s 215136 64388 215232 64468 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OUT_TT_PROJECT6
port 1190 nsew signal input
flabel metal3 s 215136 64892 215232 64972 0 FreeSans 320 0 0 0 Tile_X5Y7_UIO_OUT_TT_PROJECT7
port 1191 nsew signal input
flabel metal3 s 215136 69428 215232 69508 0 FreeSans 320 0 0 0 Tile_X5Y7_UI_IN_TT_PROJECT0
port 1192 nsew signal output
flabel metal3 s 215136 69932 215232 70012 0 FreeSans 320 0 0 0 Tile_X5Y7_UI_IN_TT_PROJECT1
port 1193 nsew signal output
flabel metal3 s 215136 70436 215232 70516 0 FreeSans 320 0 0 0 Tile_X5Y7_UI_IN_TT_PROJECT2
port 1194 nsew signal output
flabel metal3 s 215136 70940 215232 71020 0 FreeSans 320 0 0 0 Tile_X5Y7_UI_IN_TT_PROJECT3
port 1195 nsew signal output
flabel metal3 s 215136 71444 215232 71524 0 FreeSans 320 0 0 0 Tile_X5Y7_UI_IN_TT_PROJECT4
port 1196 nsew signal output
flabel metal3 s 215136 71948 215232 72028 0 FreeSans 320 0 0 0 Tile_X5Y7_UI_IN_TT_PROJECT5
port 1197 nsew signal output
flabel metal3 s 215136 72452 215232 72532 0 FreeSans 320 0 0 0 Tile_X5Y7_UI_IN_TT_PROJECT6
port 1198 nsew signal output
flabel metal3 s 215136 72956 215232 73036 0 FreeSans 320 0 0 0 Tile_X5Y7_UI_IN_TT_PROJECT7
port 1199 nsew signal output
flabel metal3 s 215136 57332 215232 57412 0 FreeSans 320 0 0 0 Tile_X5Y7_UO_OUT_TT_PROJECT0
port 1200 nsew signal input
flabel metal3 s 215136 57836 215232 57916 0 FreeSans 320 0 0 0 Tile_X5Y7_UO_OUT_TT_PROJECT1
port 1201 nsew signal input
flabel metal3 s 215136 58340 215232 58420 0 FreeSans 320 0 0 0 Tile_X5Y7_UO_OUT_TT_PROJECT2
port 1202 nsew signal input
flabel metal3 s 215136 58844 215232 58924 0 FreeSans 320 0 0 0 Tile_X5Y7_UO_OUT_TT_PROJECT3
port 1203 nsew signal input
flabel metal3 s 215136 59348 215232 59428 0 FreeSans 320 0 0 0 Tile_X5Y7_UO_OUT_TT_PROJECT4
port 1204 nsew signal input
flabel metal3 s 215136 59852 215232 59932 0 FreeSans 320 0 0 0 Tile_X5Y7_UO_OUT_TT_PROJECT5
port 1205 nsew signal input
flabel metal3 s 215136 60356 215232 60436 0 FreeSans 320 0 0 0 Tile_X5Y7_UO_OUT_TT_PROJECT6
port 1206 nsew signal input
flabel metal3 s 215136 60860 215232 60940 0 FreeSans 320 0 0 0 Tile_X5Y7_UO_OUT_TT_PROJECT7
port 1207 nsew signal input
flabel metal3 s 215136 34988 215232 35068 0 FreeSans 320 0 0 0 Tile_X5Y8_CLK_TT_PROJECT
port 1208 nsew signal output
flabel metal3 s 215136 34484 215232 34564 0 FreeSans 320 0 0 0 Tile_X5Y8_ENA_TT_PROJECT
port 1209 nsew signal output
flabel metal3 s 215136 35492 215232 35572 0 FreeSans 320 0 0 0 Tile_X5Y8_RST_N_TT_PROJECT
port 1210 nsew signal output
flabel metal3 s 215136 30452 215232 30532 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_IN_TT_PROJECT0
port 1211 nsew signal output
flabel metal3 s 215136 30956 215232 31036 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_IN_TT_PROJECT1
port 1212 nsew signal output
flabel metal3 s 215136 31460 215232 31540 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_IN_TT_PROJECT2
port 1213 nsew signal output
flabel metal3 s 215136 31964 215232 32044 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_IN_TT_PROJECT3
port 1214 nsew signal output
flabel metal3 s 215136 32468 215232 32548 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_IN_TT_PROJECT4
port 1215 nsew signal output
flabel metal3 s 215136 32972 215232 33052 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_IN_TT_PROJECT5
port 1216 nsew signal output
flabel metal3 s 215136 33476 215232 33556 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_IN_TT_PROJECT6
port 1217 nsew signal output
flabel metal3 s 215136 33980 215232 34060 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_IN_TT_PROJECT7
port 1218 nsew signal output
flabel metal3 s 215136 22388 215232 22468 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OE_TT_PROJECT0
port 1219 nsew signal input
flabel metal3 s 215136 22892 215232 22972 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OE_TT_PROJECT1
port 1220 nsew signal input
flabel metal3 s 215136 23396 215232 23476 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OE_TT_PROJECT2
port 1221 nsew signal input
flabel metal3 s 215136 23900 215232 23980 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OE_TT_PROJECT3
port 1222 nsew signal input
flabel metal3 s 215136 24404 215232 24484 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OE_TT_PROJECT4
port 1223 nsew signal input
flabel metal3 s 215136 24908 215232 24988 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OE_TT_PROJECT5
port 1224 nsew signal input
flabel metal3 s 215136 25412 215232 25492 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OE_TT_PROJECT6
port 1225 nsew signal input
flabel metal3 s 215136 25916 215232 25996 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OE_TT_PROJECT7
port 1226 nsew signal input
flabel metal3 s 215136 18356 215232 18436 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OUT_TT_PROJECT0
port 1227 nsew signal input
flabel metal3 s 215136 18860 215232 18940 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OUT_TT_PROJECT1
port 1228 nsew signal input
flabel metal3 s 215136 19364 215232 19444 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OUT_TT_PROJECT2
port 1229 nsew signal input
flabel metal3 s 215136 19868 215232 19948 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OUT_TT_PROJECT3
port 1230 nsew signal input
flabel metal3 s 215136 20372 215232 20452 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OUT_TT_PROJECT4
port 1231 nsew signal input
flabel metal3 s 215136 20876 215232 20956 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OUT_TT_PROJECT5
port 1232 nsew signal input
flabel metal3 s 215136 21380 215232 21460 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OUT_TT_PROJECT6
port 1233 nsew signal input
flabel metal3 s 215136 21884 215232 21964 0 FreeSans 320 0 0 0 Tile_X5Y8_UIO_OUT_TT_PROJECT7
port 1234 nsew signal input
flabel metal3 s 215136 26420 215232 26500 0 FreeSans 320 0 0 0 Tile_X5Y8_UI_IN_TT_PROJECT0
port 1235 nsew signal output
flabel metal3 s 215136 26924 215232 27004 0 FreeSans 320 0 0 0 Tile_X5Y8_UI_IN_TT_PROJECT1
port 1236 nsew signal output
flabel metal3 s 215136 27428 215232 27508 0 FreeSans 320 0 0 0 Tile_X5Y8_UI_IN_TT_PROJECT2
port 1237 nsew signal output
flabel metal3 s 215136 27932 215232 28012 0 FreeSans 320 0 0 0 Tile_X5Y8_UI_IN_TT_PROJECT3
port 1238 nsew signal output
flabel metal3 s 215136 28436 215232 28516 0 FreeSans 320 0 0 0 Tile_X5Y8_UI_IN_TT_PROJECT4
port 1239 nsew signal output
flabel metal3 s 215136 28940 215232 29020 0 FreeSans 320 0 0 0 Tile_X5Y8_UI_IN_TT_PROJECT5
port 1240 nsew signal output
flabel metal3 s 215136 29444 215232 29524 0 FreeSans 320 0 0 0 Tile_X5Y8_UI_IN_TT_PROJECT6
port 1241 nsew signal output
flabel metal3 s 215136 29948 215232 30028 0 FreeSans 320 0 0 0 Tile_X5Y8_UI_IN_TT_PROJECT7
port 1242 nsew signal output
flabel metal3 s 215136 14324 215232 14404 0 FreeSans 320 0 0 0 Tile_X5Y8_UO_OUT_TT_PROJECT0
port 1243 nsew signal input
flabel metal3 s 215136 14828 215232 14908 0 FreeSans 320 0 0 0 Tile_X5Y8_UO_OUT_TT_PROJECT1
port 1244 nsew signal input
flabel metal3 s 215136 15332 215232 15412 0 FreeSans 320 0 0 0 Tile_X5Y8_UO_OUT_TT_PROJECT2
port 1245 nsew signal input
flabel metal3 s 215136 15836 215232 15916 0 FreeSans 320 0 0 0 Tile_X5Y8_UO_OUT_TT_PROJECT3
port 1246 nsew signal input
flabel metal3 s 215136 16340 215232 16420 0 FreeSans 320 0 0 0 Tile_X5Y8_UO_OUT_TT_PROJECT4
port 1247 nsew signal input
flabel metal3 s 215136 16844 215232 16924 0 FreeSans 320 0 0 0 Tile_X5Y8_UO_OUT_TT_PROJECT5
port 1248 nsew signal input
flabel metal3 s 215136 17348 215232 17428 0 FreeSans 320 0 0 0 Tile_X5Y8_UO_OUT_TT_PROJECT6
port 1249 nsew signal input
flabel metal3 s 215136 17852 215232 17932 0 FreeSans 320 0 0 0 Tile_X5Y8_UO_OUT_TT_PROJECT7
port 1250 nsew signal input
flabel metal2 s 1112 0 1192 96 0 FreeSans 640 0 0 0 UserCLK
port 1251 nsew signal input
flabel metal6 s 4988 840 5428 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 26492 840 26932 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 41612 840 42052 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 56732 840 57172 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 69500 840 69940 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 84620 840 85060 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 99740 840 100180 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 112508 840 112948 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 127628 840 128068 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 142748 840 143188 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 155516 840 155956 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 170636 840 171076 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 185756 840 186196 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 198524 840 198964 366408 0 FreeSans 2624 90 0 0 VGND
port 1252 nsew ground bidirectional
flabel metal6 s 3748 840 4188 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 18868 840 19308 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 25252 840 25692 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 40372 840 40812 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 55492 840 55932 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 68260 840 68700 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 83380 840 83820 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 98500 840 98940 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 111268 840 111708 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 126388 840 126828 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 141508 840 141948 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 154276 840 154716 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 169396 840 169836 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 184516 840 184956 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 197284 840 197724 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
flabel metal6 s 212404 840 212844 366408 0 FreeSans 2624 90 0 0 VPWR
port 1253 nsew power bidirectional
rlabel metal6 198744 183624 198744 183624 0 VGND
rlabel metal6 212624 183624 212624 183624 0 VPWR
rlabel metal3 82 355740 82 355740 0 FrameData[0]
rlabel metal3 82 253092 82 253092 0 FrameData[100]
rlabel metal3 82 253596 82 253596 0 FrameData[101]
rlabel metal3 82 254100 82 254100 0 FrameData[102]
rlabel metal3 82 254604 82 254604 0 FrameData[103]
rlabel metal3 82 255108 82 255108 0 FrameData[104]
rlabel metal3 82 255612 82 255612 0 FrameData[105]
rlabel metal3 82 256116 82 256116 0 FrameData[106]
rlabel metal3 82 256620 82 256620 0 FrameData[107]
rlabel metal3 82 257124 82 257124 0 FrameData[108]
rlabel metal3 82 257628 82 257628 0 FrameData[109]
rlabel metal3 82 359100 82 359100 0 FrameData[10]
rlabel metal3 82 258132 82 258132 0 FrameData[110]
rlabel metal3 82 258636 82 258636 0 FrameData[111]
rlabel metal3 82 259140 82 259140 0 FrameData[112]
rlabel metal3 82 259644 82 259644 0 FrameData[113]
rlabel metal3 82 260148 82 260148 0 FrameData[114]
rlabel metal3 82 260652 82 260652 0 FrameData[115]
rlabel metal3 82 261156 82 261156 0 FrameData[116]
rlabel metal3 82 261660 82 261660 0 FrameData[117]
rlabel metal3 82 262164 82 262164 0 FrameData[118]
rlabel metal3 82 262668 82 262668 0 FrameData[119]
rlabel metal3 82 359436 82 359436 0 FrameData[11]
rlabel metal3 82 263172 82 263172 0 FrameData[120]
rlabel metal3 82 263676 82 263676 0 FrameData[121]
rlabel metal3 82 264180 82 264180 0 FrameData[122]
rlabel metal3 82 264684 82 264684 0 FrameData[123]
rlabel metal3 82 265188 82 265188 0 FrameData[124]
rlabel metal3 82 265692 82 265692 0 FrameData[125]
rlabel metal3 82 266196 82 266196 0 FrameData[126]
rlabel metal3 82 266700 82 266700 0 FrameData[127]
rlabel metal3 82 208068 82 208068 0 FrameData[128]
rlabel metal3 82 208572 82 208572 0 FrameData[129]
rlabel metal3 82 359772 82 359772 0 FrameData[12]
rlabel metal3 82 209076 82 209076 0 FrameData[130]
rlabel metal3 82 209580 82 209580 0 FrameData[131]
rlabel metal3 82 210084 82 210084 0 FrameData[132]
rlabel metal3 82 210588 82 210588 0 FrameData[133]
rlabel metal3 82 211092 82 211092 0 FrameData[134]
rlabel metal3 82 211596 82 211596 0 FrameData[135]
rlabel metal3 82 212100 82 212100 0 FrameData[136]
rlabel metal3 82 212604 82 212604 0 FrameData[137]
rlabel metal3 82 213108 82 213108 0 FrameData[138]
rlabel metal3 82 213612 82 213612 0 FrameData[139]
rlabel metal3 82 360108 82 360108 0 FrameData[13]
rlabel metal3 82 214116 82 214116 0 FrameData[140]
rlabel metal3 82 214620 82 214620 0 FrameData[141]
rlabel metal3 82 215124 82 215124 0 FrameData[142]
rlabel metal3 82 215628 82 215628 0 FrameData[143]
rlabel metal3 82 216132 82 216132 0 FrameData[144]
rlabel metal3 82 216636 82 216636 0 FrameData[145]
rlabel metal3 82 217140 82 217140 0 FrameData[146]
rlabel metal3 82 217644 82 217644 0 FrameData[147]
rlabel metal3 82 218148 82 218148 0 FrameData[148]
rlabel metal3 82 218652 82 218652 0 FrameData[149]
rlabel metal3 82 360444 82 360444 0 FrameData[14]
rlabel metal3 82 219156 82 219156 0 FrameData[150]
rlabel metal3 82 219660 82 219660 0 FrameData[151]
rlabel metal3 82 220164 82 220164 0 FrameData[152]
rlabel metal3 82 220668 82 220668 0 FrameData[153]
rlabel metal3 82 221172 82 221172 0 FrameData[154]
rlabel metal3 82 221676 82 221676 0 FrameData[155]
rlabel metal3 82 222180 82 222180 0 FrameData[156]
rlabel metal3 82 222684 82 222684 0 FrameData[157]
rlabel metal3 82 223188 82 223188 0 FrameData[158]
rlabel metal3 82 223692 82 223692 0 FrameData[159]
rlabel metal3 82 360780 82 360780 0 FrameData[15]
rlabel metal3 82 165060 82 165060 0 FrameData[160]
rlabel metal3 82 165564 82 165564 0 FrameData[161]
rlabel metal3 82 166068 82 166068 0 FrameData[162]
rlabel metal3 82 166572 82 166572 0 FrameData[163]
rlabel metal3 82 167076 82 167076 0 FrameData[164]
rlabel metal3 82 167580 82 167580 0 FrameData[165]
rlabel metal3 82 168084 82 168084 0 FrameData[166]
rlabel metal3 82 168588 82 168588 0 FrameData[167]
rlabel metal3 82 169092 82 169092 0 FrameData[168]
rlabel metal3 82 169596 82 169596 0 FrameData[169]
rlabel metal3 82 361116 82 361116 0 FrameData[16]
rlabel metal3 82 170100 82 170100 0 FrameData[170]
rlabel metal3 82 170604 82 170604 0 FrameData[171]
rlabel metal3 82 171108 82 171108 0 FrameData[172]
rlabel metal3 82 171612 82 171612 0 FrameData[173]
rlabel metal3 82 172116 82 172116 0 FrameData[174]
rlabel metal3 82 172620 82 172620 0 FrameData[175]
rlabel metal3 82 173124 82 173124 0 FrameData[176]
rlabel metal3 82 173628 82 173628 0 FrameData[177]
rlabel metal3 82 174132 82 174132 0 FrameData[178]
rlabel metal3 82 174636 82 174636 0 FrameData[179]
rlabel metal3 82 361452 82 361452 0 FrameData[17]
rlabel metal3 82 175140 82 175140 0 FrameData[180]
rlabel metal3 82 175644 82 175644 0 FrameData[181]
rlabel metal3 82 176148 82 176148 0 FrameData[182]
rlabel metal3 82 176652 82 176652 0 FrameData[183]
rlabel metal3 82 177156 82 177156 0 FrameData[184]
rlabel metal3 82 177660 82 177660 0 FrameData[185]
rlabel metal3 82 178164 82 178164 0 FrameData[186]
rlabel metal3 82 178668 82 178668 0 FrameData[187]
rlabel metal3 82 179172 82 179172 0 FrameData[188]
rlabel metal3 82 179676 82 179676 0 FrameData[189]
rlabel metal3 82 361788 82 361788 0 FrameData[18]
rlabel metal3 82 180180 82 180180 0 FrameData[190]
rlabel metal3 82 180684 82 180684 0 FrameData[191]
rlabel metal3 82 122052 82 122052 0 FrameData[192]
rlabel metal3 82 122556 82 122556 0 FrameData[193]
rlabel metal3 82 123060 82 123060 0 FrameData[194]
rlabel metal3 82 123564 82 123564 0 FrameData[195]
rlabel metal3 82 124068 82 124068 0 FrameData[196]
rlabel metal3 82 124572 82 124572 0 FrameData[197]
rlabel metal3 82 125076 82 125076 0 FrameData[198]
rlabel metal3 82 125580 82 125580 0 FrameData[199]
rlabel metal3 82 362124 82 362124 0 FrameData[19]
rlabel metal3 82 356076 82 356076 0 FrameData[1]
rlabel metal3 82 126084 82 126084 0 FrameData[200]
rlabel metal3 82 126588 82 126588 0 FrameData[201]
rlabel metal3 82 127092 82 127092 0 FrameData[202]
rlabel metal3 82 127596 82 127596 0 FrameData[203]
rlabel metal3 82 128100 82 128100 0 FrameData[204]
rlabel metal3 82 128604 82 128604 0 FrameData[205]
rlabel metal3 82 129108 82 129108 0 FrameData[206]
rlabel metal3 82 129612 82 129612 0 FrameData[207]
rlabel metal3 82 130116 82 130116 0 FrameData[208]
rlabel metal3 82 130620 82 130620 0 FrameData[209]
rlabel metal3 82 362460 82 362460 0 FrameData[20]
rlabel metal3 82 131124 82 131124 0 FrameData[210]
rlabel metal3 82 131628 82 131628 0 FrameData[211]
rlabel metal3 82 132132 82 132132 0 FrameData[212]
rlabel metal3 82 132636 82 132636 0 FrameData[213]
rlabel metal3 82 133140 82 133140 0 FrameData[214]
rlabel metal3 82 133644 82 133644 0 FrameData[215]
rlabel metal3 82 134148 82 134148 0 FrameData[216]
rlabel metal3 82 134652 82 134652 0 FrameData[217]
rlabel metal3 82 135156 82 135156 0 FrameData[218]
rlabel metal3 82 135660 82 135660 0 FrameData[219]
rlabel metal3 82 362796 82 362796 0 FrameData[21]
rlabel metal3 82 136164 82 136164 0 FrameData[220]
rlabel metal3 82 136668 82 136668 0 FrameData[221]
rlabel metal3 82 137172 82 137172 0 FrameData[222]
rlabel metal3 82 137676 82 137676 0 FrameData[223]
rlabel metal3 82 79044 82 79044 0 FrameData[224]
rlabel metal3 82 79548 82 79548 0 FrameData[225]
rlabel metal3 82 80052 82 80052 0 FrameData[226]
rlabel metal3 82 80556 82 80556 0 FrameData[227]
rlabel metal3 82 81060 82 81060 0 FrameData[228]
rlabel metal3 82 81564 82 81564 0 FrameData[229]
rlabel metal3 82 363132 82 363132 0 FrameData[22]
rlabel metal3 82 82068 82 82068 0 FrameData[230]
rlabel metal3 82 82572 82 82572 0 FrameData[231]
rlabel metal3 82 83076 82 83076 0 FrameData[232]
rlabel metal3 82 83580 82 83580 0 FrameData[233]
rlabel metal3 82 84084 82 84084 0 FrameData[234]
rlabel metal3 82 84588 82 84588 0 FrameData[235]
rlabel metal3 82 85092 82 85092 0 FrameData[236]
rlabel metal3 82 85596 82 85596 0 FrameData[237]
rlabel metal3 82 86100 82 86100 0 FrameData[238]
rlabel metal3 82 86604 82 86604 0 FrameData[239]
rlabel metal3 82 363468 82 363468 0 FrameData[23]
rlabel metal3 82 87108 82 87108 0 FrameData[240]
rlabel metal3 82 87612 82 87612 0 FrameData[241]
rlabel metal3 82 88116 82 88116 0 FrameData[242]
rlabel metal3 82 88620 82 88620 0 FrameData[243]
rlabel metal3 82 89124 82 89124 0 FrameData[244]
rlabel metal3 82 89628 82 89628 0 FrameData[245]
rlabel metal3 82 90132 82 90132 0 FrameData[246]
rlabel metal3 82 90636 82 90636 0 FrameData[247]
rlabel metal3 82 91140 82 91140 0 FrameData[248]
rlabel metal3 82 91644 82 91644 0 FrameData[249]
rlabel metal3 82 363804 82 363804 0 FrameData[24]
rlabel metal3 82 92148 82 92148 0 FrameData[250]
rlabel metal3 82 92652 82 92652 0 FrameData[251]
rlabel metal3 82 93156 82 93156 0 FrameData[252]
rlabel metal3 82 93660 82 93660 0 FrameData[253]
rlabel metal3 82 94164 82 94164 0 FrameData[254]
rlabel metal3 82 94668 82 94668 0 FrameData[255]
rlabel metal3 82 36036 82 36036 0 FrameData[256]
rlabel metal3 82 36540 82 36540 0 FrameData[257]
rlabel metal3 82 37044 82 37044 0 FrameData[258]
rlabel metal3 82 37548 82 37548 0 FrameData[259]
rlabel metal3 82 364140 82 364140 0 FrameData[25]
rlabel metal3 82 38052 82 38052 0 FrameData[260]
rlabel metal3 82 38556 82 38556 0 FrameData[261]
rlabel metal3 82 39060 82 39060 0 FrameData[262]
rlabel metal3 82 39564 82 39564 0 FrameData[263]
rlabel metal3 82 40068 82 40068 0 FrameData[264]
rlabel metal3 82 40572 82 40572 0 FrameData[265]
rlabel metal3 82 41076 82 41076 0 FrameData[266]
rlabel metal3 82 41580 82 41580 0 FrameData[267]
rlabel metal3 82 42084 82 42084 0 FrameData[268]
rlabel metal3 82 42588 82 42588 0 FrameData[269]
rlabel metal3 82 364476 82 364476 0 FrameData[26]
rlabel metal3 82 43092 82 43092 0 FrameData[270]
rlabel metal3 82 43596 82 43596 0 FrameData[271]
rlabel metal3 82 44100 82 44100 0 FrameData[272]
rlabel metal3 82 44604 82 44604 0 FrameData[273]
rlabel metal3 82 45108 82 45108 0 FrameData[274]
rlabel metal3 82 45612 82 45612 0 FrameData[275]
rlabel metal3 82 46116 82 46116 0 FrameData[276]
rlabel metal3 82 46620 82 46620 0 FrameData[277]
rlabel metal3 82 47124 82 47124 0 FrameData[278]
rlabel metal3 82 47628 82 47628 0 FrameData[279]
rlabel metal3 82 364812 82 364812 0 FrameData[27]
rlabel metal3 82 48132 82 48132 0 FrameData[280]
rlabel metal3 82 48636 82 48636 0 FrameData[281]
rlabel metal3 82 49140 82 49140 0 FrameData[282]
rlabel metal3 82 49644 82 49644 0 FrameData[283]
rlabel metal3 82 50148 82 50148 0 FrameData[284]
rlabel metal3 82 50652 82 50652 0 FrameData[285]
rlabel metal3 82 51156 82 51156 0 FrameData[286]
rlabel metal3 82 51660 82 51660 0 FrameData[287]
rlabel metal3 82 924 82 924 0 FrameData[288]
rlabel metal3 82 1260 82 1260 0 FrameData[289]
rlabel metal3 82 365148 82 365148 0 FrameData[28]
rlabel metal3 82 1596 82 1596 0 FrameData[290]
rlabel metal3 82 1932 82 1932 0 FrameData[291]
rlabel metal3 82 2268 82 2268 0 FrameData[292]
rlabel metal3 82 2604 82 2604 0 FrameData[293]
rlabel metal3 82 2940 82 2940 0 FrameData[294]
rlabel metal3 82 3276 82 3276 0 FrameData[295]
rlabel metal3 82 3612 82 3612 0 FrameData[296]
rlabel metal3 82 3948 82 3948 0 FrameData[297]
rlabel metal3 82 4284 82 4284 0 FrameData[298]
rlabel metal3 82 4620 82 4620 0 FrameData[299]
rlabel metal3 82 365484 82 365484 0 FrameData[29]
rlabel metal3 82 356412 82 356412 0 FrameData[2]
rlabel metal3 82 4956 82 4956 0 FrameData[300]
rlabel metal3 82 5292 82 5292 0 FrameData[301]
rlabel metal3 82 5628 82 5628 0 FrameData[302]
rlabel metal3 82 5964 82 5964 0 FrameData[303]
rlabel metal3 82 6300 82 6300 0 FrameData[304]
rlabel metal3 82 6636 82 6636 0 FrameData[305]
rlabel metal3 82 6972 82 6972 0 FrameData[306]
rlabel metal3 82 7308 82 7308 0 FrameData[307]
rlabel metal3 82 7644 82 7644 0 FrameData[308]
rlabel metal3 82 7980 82 7980 0 FrameData[309]
rlabel metal3 82 365820 82 365820 0 FrameData[30]
rlabel metal3 82 8316 82 8316 0 FrameData[310]
rlabel metal3 82 8652 82 8652 0 FrameData[311]
rlabel metal3 82 8988 82 8988 0 FrameData[312]
rlabel metal3 82 9324 82 9324 0 FrameData[313]
rlabel metal3 82 9660 82 9660 0 FrameData[314]
rlabel metal3 82 9996 82 9996 0 FrameData[315]
rlabel metal3 82 10332 82 10332 0 FrameData[316]
rlabel metal3 82 10668 82 10668 0 FrameData[317]
rlabel metal3 82 11004 82 11004 0 FrameData[318]
rlabel metal3 82 11340 82 11340 0 FrameData[319]
rlabel metal3 82 366156 82 366156 0 FrameData[31]
rlabel metal3 82 337092 82 337092 0 FrameData[32]
rlabel metal3 82 337596 82 337596 0 FrameData[33]
rlabel metal3 82 338100 82 338100 0 FrameData[34]
rlabel metal3 82 338604 82 338604 0 FrameData[35]
rlabel metal3 82 339108 82 339108 0 FrameData[36]
rlabel metal3 82 339612 82 339612 0 FrameData[37]
rlabel metal3 82 340116 82 340116 0 FrameData[38]
rlabel metal3 82 340620 82 340620 0 FrameData[39]
rlabel metal3 82 356748 82 356748 0 FrameData[3]
rlabel metal3 82 341124 82 341124 0 FrameData[40]
rlabel metal3 82 341628 82 341628 0 FrameData[41]
rlabel metal3 82 342132 82 342132 0 FrameData[42]
rlabel metal3 82 342636 82 342636 0 FrameData[43]
rlabel metal3 82 343140 82 343140 0 FrameData[44]
rlabel metal3 82 343644 82 343644 0 FrameData[45]
rlabel metal3 82 344148 82 344148 0 FrameData[46]
rlabel metal3 82 344652 82 344652 0 FrameData[47]
rlabel metal3 82 345156 82 345156 0 FrameData[48]
rlabel metal3 82 345660 82 345660 0 FrameData[49]
rlabel metal3 82 357084 82 357084 0 FrameData[4]
rlabel metal3 82 346164 82 346164 0 FrameData[50]
rlabel metal3 82 346668 82 346668 0 FrameData[51]
rlabel metal3 82 347172 82 347172 0 FrameData[52]
rlabel metal3 82 347676 82 347676 0 FrameData[53]
rlabel metal3 82 348180 82 348180 0 FrameData[54]
rlabel metal3 82 348684 82 348684 0 FrameData[55]
rlabel metal3 82 349188 82 349188 0 FrameData[56]
rlabel metal3 82 349692 82 349692 0 FrameData[57]
rlabel metal3 82 350196 82 350196 0 FrameData[58]
rlabel metal3 82 350700 82 350700 0 FrameData[59]
rlabel metal3 82 357420 82 357420 0 FrameData[5]
rlabel metal3 82 351204 82 351204 0 FrameData[60]
rlabel metal3 82 351708 82 351708 0 FrameData[61]
rlabel metal3 82 352212 82 352212 0 FrameData[62]
rlabel metal3 82 352716 82 352716 0 FrameData[63]
rlabel metal3 82 294084 82 294084 0 FrameData[64]
rlabel metal3 82 294588 82 294588 0 FrameData[65]
rlabel metal3 82 295092 82 295092 0 FrameData[66]
rlabel metal3 82 295596 82 295596 0 FrameData[67]
rlabel metal3 82 296100 82 296100 0 FrameData[68]
rlabel metal3 82 296604 82 296604 0 FrameData[69]
rlabel metal3 82 357756 82 357756 0 FrameData[6]
rlabel metal3 82 297108 82 297108 0 FrameData[70]
rlabel metal3 82 297612 82 297612 0 FrameData[71]
rlabel metal3 82 298116 82 298116 0 FrameData[72]
rlabel metal3 82 298620 82 298620 0 FrameData[73]
rlabel metal3 82 299124 82 299124 0 FrameData[74]
rlabel metal3 82 299628 82 299628 0 FrameData[75]
rlabel metal3 82 300132 82 300132 0 FrameData[76]
rlabel metal3 82 300636 82 300636 0 FrameData[77]
rlabel metal3 82 301140 82 301140 0 FrameData[78]
rlabel metal3 82 301644 82 301644 0 FrameData[79]
rlabel metal3 82 358092 82 358092 0 FrameData[7]
rlabel metal3 82 302148 82 302148 0 FrameData[80]
rlabel metal3 82 302652 82 302652 0 FrameData[81]
rlabel metal3 82 303156 82 303156 0 FrameData[82]
rlabel metal3 82 303660 82 303660 0 FrameData[83]
rlabel metal3 82 304164 82 304164 0 FrameData[84]
rlabel metal3 82 304668 82 304668 0 FrameData[85]
rlabel metal3 82 305172 82 305172 0 FrameData[86]
rlabel metal3 82 305676 82 305676 0 FrameData[87]
rlabel metal3 82 306180 82 306180 0 FrameData[88]
rlabel metal3 82 306684 82 306684 0 FrameData[89]
rlabel metal3 82 358428 82 358428 0 FrameData[8]
rlabel metal3 82 307188 82 307188 0 FrameData[90]
rlabel metal3 82 307692 82 307692 0 FrameData[91]
rlabel metal3 82 308196 82 308196 0 FrameData[92]
rlabel metal3 82 308700 82 308700 0 FrameData[93]
rlabel metal3 82 309204 82 309204 0 FrameData[94]
rlabel metal3 82 309708 82 309708 0 FrameData[95]
rlabel metal3 82 251076 82 251076 0 FrameData[96]
rlabel metal3 82 251580 82 251580 0 FrameData[97]
rlabel metal3 82 252084 82 252084 0 FrameData[98]
rlabel metal3 82 252588 82 252588 0 FrameData[99]
rlabel metal3 82 358764 82 358764 0 FrameData[9]
rlabel metal2 2112 454 2112 454 0 FrameStrobe[0]
rlabel metal2 195648 454 195648 454 0 FrameStrobe[100]
rlabel metal2 196608 454 196608 454 0 FrameStrobe[101]
rlabel metal2 197568 454 197568 454 0 FrameStrobe[102]
rlabel metal2 198528 454 198528 454 0 FrameStrobe[103]
rlabel metal2 199488 454 199488 454 0 FrameStrobe[104]
rlabel metal2 200448 454 200448 454 0 FrameStrobe[105]
rlabel metal2 201408 454 201408 454 0 FrameStrobe[106]
rlabel metal2 202368 454 202368 454 0 FrameStrobe[107]
rlabel metal2 203328 454 203328 454 0 FrameStrobe[108]
rlabel metal2 204288 454 204288 454 0 FrameStrobe[109]
rlabel metal2 11712 454 11712 454 0 FrameStrobe[10]
rlabel metal2 205248 454 205248 454 0 FrameStrobe[110]
rlabel metal2 206208 454 206208 454 0 FrameStrobe[111]
rlabel metal2 207168 454 207168 454 0 FrameStrobe[112]
rlabel metal2 208128 454 208128 454 0 FrameStrobe[113]
rlabel metal2 209088 454 209088 454 0 FrameStrobe[114]
rlabel metal2 210048 454 210048 454 0 FrameStrobe[115]
rlabel metal2 211008 454 211008 454 0 FrameStrobe[116]
rlabel metal2 211968 454 211968 454 0 FrameStrobe[117]
rlabel metal2 212928 454 212928 454 0 FrameStrobe[118]
rlabel metal2 213888 454 213888 454 0 FrameStrobe[119]
rlabel metal2 12672 454 12672 454 0 FrameStrobe[11]
rlabel metal2 13632 454 13632 454 0 FrameStrobe[12]
rlabel metal2 14592 454 14592 454 0 FrameStrobe[13]
rlabel metal2 15552 454 15552 454 0 FrameStrobe[14]
rlabel metal2 16512 454 16512 454 0 FrameStrobe[15]
rlabel metal2 17472 454 17472 454 0 FrameStrobe[16]
rlabel metal2 18432 454 18432 454 0 FrameStrobe[17]
rlabel metal2 19392 454 19392 454 0 FrameStrobe[18]
rlabel metal2 20352 454 20352 454 0 FrameStrobe[19]
rlabel metal2 3072 454 3072 454 0 FrameStrobe[1]
rlabel metal2 39552 454 39552 454 0 FrameStrobe[20]
rlabel metal2 40704 454 40704 454 0 FrameStrobe[21]
rlabel metal2 41856 454 41856 454 0 FrameStrobe[22]
rlabel metal2 43008 454 43008 454 0 FrameStrobe[23]
rlabel metal2 44160 454 44160 454 0 FrameStrobe[24]
rlabel metal2 45312 454 45312 454 0 FrameStrobe[25]
rlabel metal2 46464 454 46464 454 0 FrameStrobe[26]
rlabel metal2 47616 454 47616 454 0 FrameStrobe[27]
rlabel metal2 48768 454 48768 454 0 FrameStrobe[28]
rlabel metal2 49920 454 49920 454 0 FrameStrobe[29]
rlabel metal2 4032 454 4032 454 0 FrameStrobe[2]
rlabel metal2 51072 454 51072 454 0 FrameStrobe[30]
rlabel metal2 52224 454 52224 454 0 FrameStrobe[31]
rlabel metal2 53376 454 53376 454 0 FrameStrobe[32]
rlabel metal2 54528 454 54528 454 0 FrameStrobe[33]
rlabel metal2 55680 454 55680 454 0 FrameStrobe[34]
rlabel metal2 56832 454 56832 454 0 FrameStrobe[35]
rlabel metal2 57984 454 57984 454 0 FrameStrobe[36]
rlabel metal2 59136 454 59136 454 0 FrameStrobe[37]
rlabel metal2 60288 454 60288 454 0 FrameStrobe[38]
rlabel metal2 61440 454 61440 454 0 FrameStrobe[39]
rlabel metal2 4992 454 4992 454 0 FrameStrobe[3]
rlabel metal2 82560 454 82560 454 0 FrameStrobe[40]
rlabel metal2 83712 454 83712 454 0 FrameStrobe[41]
rlabel metal2 84864 454 84864 454 0 FrameStrobe[42]
rlabel metal2 86016 454 86016 454 0 FrameStrobe[43]
rlabel metal2 87168 454 87168 454 0 FrameStrobe[44]
rlabel metal2 88320 454 88320 454 0 FrameStrobe[45]
rlabel metal2 89472 454 89472 454 0 FrameStrobe[46]
rlabel metal2 90624 454 90624 454 0 FrameStrobe[47]
rlabel metal2 91776 454 91776 454 0 FrameStrobe[48]
rlabel metal2 92928 454 92928 454 0 FrameStrobe[49]
rlabel metal2 5952 454 5952 454 0 FrameStrobe[4]
rlabel metal2 94080 454 94080 454 0 FrameStrobe[50]
rlabel metal2 95232 454 95232 454 0 FrameStrobe[51]
rlabel metal2 96384 454 96384 454 0 FrameStrobe[52]
rlabel metal2 97536 454 97536 454 0 FrameStrobe[53]
rlabel metal2 98688 454 98688 454 0 FrameStrobe[54]
rlabel metal2 99840 454 99840 454 0 FrameStrobe[55]
rlabel metal2 100992 454 100992 454 0 FrameStrobe[56]
rlabel metal2 102144 454 102144 454 0 FrameStrobe[57]
rlabel metal2 103296 454 103296 454 0 FrameStrobe[58]
rlabel metal2 104448 454 104448 454 0 FrameStrobe[59]
rlabel metal2 6912 454 6912 454 0 FrameStrobe[5]
rlabel metal2 125568 454 125568 454 0 FrameStrobe[60]
rlabel metal2 126720 454 126720 454 0 FrameStrobe[61]
rlabel metal2 127872 454 127872 454 0 FrameStrobe[62]
rlabel metal2 129024 454 129024 454 0 FrameStrobe[63]
rlabel metal2 130176 454 130176 454 0 FrameStrobe[64]
rlabel metal2 131328 454 131328 454 0 FrameStrobe[65]
rlabel metal2 132480 454 132480 454 0 FrameStrobe[66]
rlabel metal2 133632 454 133632 454 0 FrameStrobe[67]
rlabel metal2 134784 454 134784 454 0 FrameStrobe[68]
rlabel metal2 135936 454 135936 454 0 FrameStrobe[69]
rlabel metal2 7872 454 7872 454 0 FrameStrobe[6]
rlabel metal2 137088 454 137088 454 0 FrameStrobe[70]
rlabel metal2 138240 454 138240 454 0 FrameStrobe[71]
rlabel metal2 139392 454 139392 454 0 FrameStrobe[72]
rlabel metal2 140544 454 140544 454 0 FrameStrobe[73]
rlabel metal2 141696 454 141696 454 0 FrameStrobe[74]
rlabel metal2 142848 454 142848 454 0 FrameStrobe[75]
rlabel metal2 144000 454 144000 454 0 FrameStrobe[76]
rlabel metal2 145152 454 145152 454 0 FrameStrobe[77]
rlabel metal2 146304 454 146304 454 0 FrameStrobe[78]
rlabel metal2 147456 454 147456 454 0 FrameStrobe[79]
rlabel metal2 8832 454 8832 454 0 FrameStrobe[7]
rlabel metal2 168576 454 168576 454 0 FrameStrobe[80]
rlabel metal2 169728 454 169728 454 0 FrameStrobe[81]
rlabel metal2 170880 454 170880 454 0 FrameStrobe[82]
rlabel metal2 172032 454 172032 454 0 FrameStrobe[83]
rlabel metal2 173184 454 173184 454 0 FrameStrobe[84]
rlabel metal2 174336 454 174336 454 0 FrameStrobe[85]
rlabel metal2 175488 454 175488 454 0 FrameStrobe[86]
rlabel metal2 176640 454 176640 454 0 FrameStrobe[87]
rlabel metal2 177792 454 177792 454 0 FrameStrobe[88]
rlabel metal2 178944 454 178944 454 0 FrameStrobe[89]
rlabel metal2 9792 454 9792 454 0 FrameStrobe[8]
rlabel metal2 180096 454 180096 454 0 FrameStrobe[90]
rlabel metal2 181248 454 181248 454 0 FrameStrobe[91]
rlabel metal2 182400 454 182400 454 0 FrameStrobe[92]
rlabel metal2 183552 454 183552 454 0 FrameStrobe[93]
rlabel metal2 184704 454 184704 454 0 FrameStrobe[94]
rlabel metal2 185856 454 185856 454 0 FrameStrobe[95]
rlabel metal2 187008 454 187008 454 0 FrameStrobe[96]
rlabel metal2 188160 454 188160 454 0 FrameStrobe[97]
rlabel metal2 189312 454 189312 454 0 FrameStrobe[98]
rlabel metal2 190464 454 190464 454 0 FrameStrobe[99]
rlabel metal2 10752 454 10752 454 0 FrameStrobe[9]
rlabel metal3 82 336084 82 336084 0 Tile_X0Y1_CLK_TT_PROJECT
rlabel metal3 82 335580 82 335580 0 Tile_X0Y1_ENA_TT_PROJECT
rlabel metal3 82 336588 82 336588 0 Tile_X0Y1_RST_N_TT_PROJECT
rlabel metal3 82 331548 82 331548 0 Tile_X0Y1_UIO_IN_TT_PROJECT0
rlabel metal3 82 332052 82 332052 0 Tile_X0Y1_UIO_IN_TT_PROJECT1
rlabel metal3 82 332556 82 332556 0 Tile_X0Y1_UIO_IN_TT_PROJECT2
rlabel metal3 82 333060 82 333060 0 Tile_X0Y1_UIO_IN_TT_PROJECT3
rlabel metal3 82 333564 82 333564 0 Tile_X0Y1_UIO_IN_TT_PROJECT4
rlabel metal3 82 334068 82 334068 0 Tile_X0Y1_UIO_IN_TT_PROJECT5
rlabel metal3 82 334572 82 334572 0 Tile_X0Y1_UIO_IN_TT_PROJECT6
rlabel metal3 82 335076 82 335076 0 Tile_X0Y1_UIO_IN_TT_PROJECT7
rlabel metal3 82 323484 82 323484 0 Tile_X0Y1_UIO_OE_TT_PROJECT0
rlabel metal3 82 323988 82 323988 0 Tile_X0Y1_UIO_OE_TT_PROJECT1
rlabel metal3 82 324492 82 324492 0 Tile_X0Y1_UIO_OE_TT_PROJECT2
rlabel metal3 82 324996 82 324996 0 Tile_X0Y1_UIO_OE_TT_PROJECT3
rlabel metal3 82 325500 82 325500 0 Tile_X0Y1_UIO_OE_TT_PROJECT4
rlabel metal3 82 326004 82 326004 0 Tile_X0Y1_UIO_OE_TT_PROJECT5
rlabel metal3 82 326508 82 326508 0 Tile_X0Y1_UIO_OE_TT_PROJECT6
rlabel metal3 82 327012 82 327012 0 Tile_X0Y1_UIO_OE_TT_PROJECT7
rlabel metal3 82 319452 82 319452 0 Tile_X0Y1_UIO_OUT_TT_PROJECT0
rlabel metal3 82 319956 82 319956 0 Tile_X0Y1_UIO_OUT_TT_PROJECT1
rlabel metal3 82 320460 82 320460 0 Tile_X0Y1_UIO_OUT_TT_PROJECT2
rlabel metal3 82 320964 82 320964 0 Tile_X0Y1_UIO_OUT_TT_PROJECT3
rlabel metal3 82 321468 82 321468 0 Tile_X0Y1_UIO_OUT_TT_PROJECT4
rlabel metal3 82 321972 82 321972 0 Tile_X0Y1_UIO_OUT_TT_PROJECT5
rlabel metal3 82 322476 82 322476 0 Tile_X0Y1_UIO_OUT_TT_PROJECT6
rlabel metal3 82 322980 82 322980 0 Tile_X0Y1_UIO_OUT_TT_PROJECT7
rlabel metal3 82 327516 82 327516 0 Tile_X0Y1_UI_IN_TT_PROJECT0
rlabel metal3 82 328020 82 328020 0 Tile_X0Y1_UI_IN_TT_PROJECT1
rlabel metal3 82 328524 82 328524 0 Tile_X0Y1_UI_IN_TT_PROJECT2
rlabel metal3 82 329028 82 329028 0 Tile_X0Y1_UI_IN_TT_PROJECT3
rlabel metal3 82 329532 82 329532 0 Tile_X0Y1_UI_IN_TT_PROJECT4
rlabel metal3 82 330036 82 330036 0 Tile_X0Y1_UI_IN_TT_PROJECT5
rlabel metal3 82 330540 82 330540 0 Tile_X0Y1_UI_IN_TT_PROJECT6
rlabel metal3 82 331044 82 331044 0 Tile_X0Y1_UI_IN_TT_PROJECT7
rlabel metal3 82 315420 82 315420 0 Tile_X0Y1_UO_OUT_TT_PROJECT0
rlabel metal3 82 315924 82 315924 0 Tile_X0Y1_UO_OUT_TT_PROJECT1
rlabel metal3 82 316428 82 316428 0 Tile_X0Y1_UO_OUT_TT_PROJECT2
rlabel metal3 82 316932 82 316932 0 Tile_X0Y1_UO_OUT_TT_PROJECT3
rlabel metal3 82 317436 82 317436 0 Tile_X0Y1_UO_OUT_TT_PROJECT4
rlabel metal3 82 317940 82 317940 0 Tile_X0Y1_UO_OUT_TT_PROJECT5
rlabel metal3 82 318444 82 318444 0 Tile_X0Y1_UO_OUT_TT_PROJECT6
rlabel metal3 82 318948 82 318948 0 Tile_X0Y1_UO_OUT_TT_PROJECT7
rlabel metal3 82 293076 82 293076 0 Tile_X0Y2_CLK_TT_PROJECT
rlabel metal3 82 292572 82 292572 0 Tile_X0Y2_ENA_TT_PROJECT
rlabel metal3 82 293580 82 293580 0 Tile_X0Y2_RST_N_TT_PROJECT
rlabel metal3 82 288540 82 288540 0 Tile_X0Y2_UIO_IN_TT_PROJECT0
rlabel metal3 82 289044 82 289044 0 Tile_X0Y2_UIO_IN_TT_PROJECT1
rlabel metal3 82 289548 82 289548 0 Tile_X0Y2_UIO_IN_TT_PROJECT2
rlabel metal3 82 290052 82 290052 0 Tile_X0Y2_UIO_IN_TT_PROJECT3
rlabel metal3 82 290556 82 290556 0 Tile_X0Y2_UIO_IN_TT_PROJECT4
rlabel metal3 82 291060 82 291060 0 Tile_X0Y2_UIO_IN_TT_PROJECT5
rlabel metal3 82 291564 82 291564 0 Tile_X0Y2_UIO_IN_TT_PROJECT6
rlabel metal3 82 292068 82 292068 0 Tile_X0Y2_UIO_IN_TT_PROJECT7
rlabel metal3 82 280476 82 280476 0 Tile_X0Y2_UIO_OE_TT_PROJECT0
rlabel metal3 82 280980 82 280980 0 Tile_X0Y2_UIO_OE_TT_PROJECT1
rlabel metal3 82 281484 82 281484 0 Tile_X0Y2_UIO_OE_TT_PROJECT2
rlabel metal3 82 281988 82 281988 0 Tile_X0Y2_UIO_OE_TT_PROJECT3
rlabel metal3 82 282492 82 282492 0 Tile_X0Y2_UIO_OE_TT_PROJECT4
rlabel metal3 82 282996 82 282996 0 Tile_X0Y2_UIO_OE_TT_PROJECT5
rlabel metal3 82 283500 82 283500 0 Tile_X0Y2_UIO_OE_TT_PROJECT6
rlabel metal3 82 284004 82 284004 0 Tile_X0Y2_UIO_OE_TT_PROJECT7
rlabel metal3 82 276444 82 276444 0 Tile_X0Y2_UIO_OUT_TT_PROJECT0
rlabel metal3 82 276948 82 276948 0 Tile_X0Y2_UIO_OUT_TT_PROJECT1
rlabel metal3 82 277452 82 277452 0 Tile_X0Y2_UIO_OUT_TT_PROJECT2
rlabel metal3 82 277956 82 277956 0 Tile_X0Y2_UIO_OUT_TT_PROJECT3
rlabel metal3 82 278460 82 278460 0 Tile_X0Y2_UIO_OUT_TT_PROJECT4
rlabel metal3 82 278964 82 278964 0 Tile_X0Y2_UIO_OUT_TT_PROJECT5
rlabel metal3 82 279468 82 279468 0 Tile_X0Y2_UIO_OUT_TT_PROJECT6
rlabel metal3 82 279972 82 279972 0 Tile_X0Y2_UIO_OUT_TT_PROJECT7
rlabel metal3 82 284508 82 284508 0 Tile_X0Y2_UI_IN_TT_PROJECT0
rlabel metal3 82 285012 82 285012 0 Tile_X0Y2_UI_IN_TT_PROJECT1
rlabel metal3 82 285516 82 285516 0 Tile_X0Y2_UI_IN_TT_PROJECT2
rlabel metal3 82 286020 82 286020 0 Tile_X0Y2_UI_IN_TT_PROJECT3
rlabel metal3 82 286524 82 286524 0 Tile_X0Y2_UI_IN_TT_PROJECT4
rlabel metal3 82 287028 82 287028 0 Tile_X0Y2_UI_IN_TT_PROJECT5
rlabel metal3 82 287532 82 287532 0 Tile_X0Y2_UI_IN_TT_PROJECT6
rlabel metal3 82 288036 82 288036 0 Tile_X0Y2_UI_IN_TT_PROJECT7
rlabel metal3 82 272412 82 272412 0 Tile_X0Y2_UO_OUT_TT_PROJECT0
rlabel metal3 82 272916 82 272916 0 Tile_X0Y2_UO_OUT_TT_PROJECT1
rlabel metal3 82 273420 82 273420 0 Tile_X0Y2_UO_OUT_TT_PROJECT2
rlabel metal3 82 273924 82 273924 0 Tile_X0Y2_UO_OUT_TT_PROJECT3
rlabel metal3 82 274428 82 274428 0 Tile_X0Y2_UO_OUT_TT_PROJECT4
rlabel metal3 82 274932 82 274932 0 Tile_X0Y2_UO_OUT_TT_PROJECT5
rlabel metal3 82 275436 82 275436 0 Tile_X0Y2_UO_OUT_TT_PROJECT6
rlabel metal3 82 275940 82 275940 0 Tile_X0Y2_UO_OUT_TT_PROJECT7
rlabel metal3 82 250068 82 250068 0 Tile_X0Y3_CLK_TT_PROJECT
rlabel metal3 82 249564 82 249564 0 Tile_X0Y3_ENA_TT_PROJECT
rlabel metal3 82 250572 82 250572 0 Tile_X0Y3_RST_N_TT_PROJECT
rlabel metal3 82 245532 82 245532 0 Tile_X0Y3_UIO_IN_TT_PROJECT0
rlabel metal3 82 246036 82 246036 0 Tile_X0Y3_UIO_IN_TT_PROJECT1
rlabel metal3 82 246540 82 246540 0 Tile_X0Y3_UIO_IN_TT_PROJECT2
rlabel metal3 82 247044 82 247044 0 Tile_X0Y3_UIO_IN_TT_PROJECT3
rlabel metal3 82 247548 82 247548 0 Tile_X0Y3_UIO_IN_TT_PROJECT4
rlabel metal3 82 248052 82 248052 0 Tile_X0Y3_UIO_IN_TT_PROJECT5
rlabel metal3 82 248556 82 248556 0 Tile_X0Y3_UIO_IN_TT_PROJECT6
rlabel metal3 82 249060 82 249060 0 Tile_X0Y3_UIO_IN_TT_PROJECT7
rlabel metal3 82 237468 82 237468 0 Tile_X0Y3_UIO_OE_TT_PROJECT0
rlabel metal3 82 237972 82 237972 0 Tile_X0Y3_UIO_OE_TT_PROJECT1
rlabel metal3 82 238476 82 238476 0 Tile_X0Y3_UIO_OE_TT_PROJECT2
rlabel metal3 82 238980 82 238980 0 Tile_X0Y3_UIO_OE_TT_PROJECT3
rlabel metal3 82 239484 82 239484 0 Tile_X0Y3_UIO_OE_TT_PROJECT4
rlabel metal3 82 239988 82 239988 0 Tile_X0Y3_UIO_OE_TT_PROJECT5
rlabel metal3 82 240492 82 240492 0 Tile_X0Y3_UIO_OE_TT_PROJECT6
rlabel metal3 82 240996 82 240996 0 Tile_X0Y3_UIO_OE_TT_PROJECT7
rlabel metal3 82 233436 82 233436 0 Tile_X0Y3_UIO_OUT_TT_PROJECT0
rlabel metal3 82 233940 82 233940 0 Tile_X0Y3_UIO_OUT_TT_PROJECT1
rlabel metal3 82 234444 82 234444 0 Tile_X0Y3_UIO_OUT_TT_PROJECT2
rlabel metal3 82 234948 82 234948 0 Tile_X0Y3_UIO_OUT_TT_PROJECT3
rlabel metal3 82 235452 82 235452 0 Tile_X0Y3_UIO_OUT_TT_PROJECT4
rlabel metal3 82 235956 82 235956 0 Tile_X0Y3_UIO_OUT_TT_PROJECT5
rlabel metal3 82 236460 82 236460 0 Tile_X0Y3_UIO_OUT_TT_PROJECT6
rlabel metal3 82 236964 82 236964 0 Tile_X0Y3_UIO_OUT_TT_PROJECT7
rlabel metal3 82 241500 82 241500 0 Tile_X0Y3_UI_IN_TT_PROJECT0
rlabel metal3 82 242004 82 242004 0 Tile_X0Y3_UI_IN_TT_PROJECT1
rlabel metal3 82 242508 82 242508 0 Tile_X0Y3_UI_IN_TT_PROJECT2
rlabel metal3 82 243012 82 243012 0 Tile_X0Y3_UI_IN_TT_PROJECT3
rlabel metal3 82 243516 82 243516 0 Tile_X0Y3_UI_IN_TT_PROJECT4
rlabel metal3 82 244020 82 244020 0 Tile_X0Y3_UI_IN_TT_PROJECT5
rlabel metal3 82 244524 82 244524 0 Tile_X0Y3_UI_IN_TT_PROJECT6
rlabel metal3 82 245028 82 245028 0 Tile_X0Y3_UI_IN_TT_PROJECT7
rlabel metal3 82 229404 82 229404 0 Tile_X0Y3_UO_OUT_TT_PROJECT0
rlabel metal3 82 229908 82 229908 0 Tile_X0Y3_UO_OUT_TT_PROJECT1
rlabel metal3 82 230412 82 230412 0 Tile_X0Y3_UO_OUT_TT_PROJECT2
rlabel metal3 82 230916 82 230916 0 Tile_X0Y3_UO_OUT_TT_PROJECT3
rlabel metal3 82 231420 82 231420 0 Tile_X0Y3_UO_OUT_TT_PROJECT4
rlabel metal3 82 231924 82 231924 0 Tile_X0Y3_UO_OUT_TT_PROJECT5
rlabel metal3 82 232428 82 232428 0 Tile_X0Y3_UO_OUT_TT_PROJECT6
rlabel metal3 82 232932 82 232932 0 Tile_X0Y3_UO_OUT_TT_PROJECT7
rlabel metal3 82 207060 82 207060 0 Tile_X0Y4_CLK_TT_PROJECT
rlabel metal3 82 206556 82 206556 0 Tile_X0Y4_ENA_TT_PROJECT
rlabel metal3 82 207564 82 207564 0 Tile_X0Y4_RST_N_TT_PROJECT
rlabel metal3 82 202524 82 202524 0 Tile_X0Y4_UIO_IN_TT_PROJECT0
rlabel metal3 82 203028 82 203028 0 Tile_X0Y4_UIO_IN_TT_PROJECT1
rlabel metal3 82 203532 82 203532 0 Tile_X0Y4_UIO_IN_TT_PROJECT2
rlabel metal3 82 204036 82 204036 0 Tile_X0Y4_UIO_IN_TT_PROJECT3
rlabel metal3 82 204540 82 204540 0 Tile_X0Y4_UIO_IN_TT_PROJECT4
rlabel metal3 82 205044 82 205044 0 Tile_X0Y4_UIO_IN_TT_PROJECT5
rlabel metal3 82 205548 82 205548 0 Tile_X0Y4_UIO_IN_TT_PROJECT6
rlabel metal3 82 206052 82 206052 0 Tile_X0Y4_UIO_IN_TT_PROJECT7
rlabel metal3 82 194460 82 194460 0 Tile_X0Y4_UIO_OE_TT_PROJECT0
rlabel metal3 82 194964 82 194964 0 Tile_X0Y4_UIO_OE_TT_PROJECT1
rlabel metal3 82 195468 82 195468 0 Tile_X0Y4_UIO_OE_TT_PROJECT2
rlabel metal3 82 195972 82 195972 0 Tile_X0Y4_UIO_OE_TT_PROJECT3
rlabel metal3 82 196476 82 196476 0 Tile_X0Y4_UIO_OE_TT_PROJECT4
rlabel metal3 82 196980 82 196980 0 Tile_X0Y4_UIO_OE_TT_PROJECT5
rlabel metal3 82 197484 82 197484 0 Tile_X0Y4_UIO_OE_TT_PROJECT6
rlabel metal3 82 197988 82 197988 0 Tile_X0Y4_UIO_OE_TT_PROJECT7
rlabel metal3 82 190428 82 190428 0 Tile_X0Y4_UIO_OUT_TT_PROJECT0
rlabel metal3 82 190932 82 190932 0 Tile_X0Y4_UIO_OUT_TT_PROJECT1
rlabel metal3 82 191436 82 191436 0 Tile_X0Y4_UIO_OUT_TT_PROJECT2
rlabel metal3 82 191940 82 191940 0 Tile_X0Y4_UIO_OUT_TT_PROJECT3
rlabel metal3 82 192444 82 192444 0 Tile_X0Y4_UIO_OUT_TT_PROJECT4
rlabel metal3 82 192948 82 192948 0 Tile_X0Y4_UIO_OUT_TT_PROJECT5
rlabel metal3 82 193452 82 193452 0 Tile_X0Y4_UIO_OUT_TT_PROJECT6
rlabel metal3 82 193956 82 193956 0 Tile_X0Y4_UIO_OUT_TT_PROJECT7
rlabel metal3 82 198492 82 198492 0 Tile_X0Y4_UI_IN_TT_PROJECT0
rlabel metal3 82 198996 82 198996 0 Tile_X0Y4_UI_IN_TT_PROJECT1
rlabel metal3 82 199500 82 199500 0 Tile_X0Y4_UI_IN_TT_PROJECT2
rlabel metal3 82 200004 82 200004 0 Tile_X0Y4_UI_IN_TT_PROJECT3
rlabel metal3 82 200508 82 200508 0 Tile_X0Y4_UI_IN_TT_PROJECT4
rlabel metal3 82 201012 82 201012 0 Tile_X0Y4_UI_IN_TT_PROJECT5
rlabel metal3 82 201516 82 201516 0 Tile_X0Y4_UI_IN_TT_PROJECT6
rlabel metal3 82 202020 82 202020 0 Tile_X0Y4_UI_IN_TT_PROJECT7
rlabel metal3 82 186396 82 186396 0 Tile_X0Y4_UO_OUT_TT_PROJECT0
rlabel metal3 82 186900 82 186900 0 Tile_X0Y4_UO_OUT_TT_PROJECT1
rlabel metal3 82 187404 82 187404 0 Tile_X0Y4_UO_OUT_TT_PROJECT2
rlabel metal3 82 187908 82 187908 0 Tile_X0Y4_UO_OUT_TT_PROJECT3
rlabel metal3 82 188412 82 188412 0 Tile_X0Y4_UO_OUT_TT_PROJECT4
rlabel metal3 82 188916 82 188916 0 Tile_X0Y4_UO_OUT_TT_PROJECT5
rlabel metal3 82 189420 82 189420 0 Tile_X0Y4_UO_OUT_TT_PROJECT6
rlabel metal3 82 189924 82 189924 0 Tile_X0Y4_UO_OUT_TT_PROJECT7
rlabel metal3 82 164052 82 164052 0 Tile_X0Y5_CLK_TT_PROJECT
rlabel metal3 82 163548 82 163548 0 Tile_X0Y5_ENA_TT_PROJECT
rlabel metal3 82 164556 82 164556 0 Tile_X0Y5_RST_N_TT_PROJECT
rlabel metal3 82 159516 82 159516 0 Tile_X0Y5_UIO_IN_TT_PROJECT0
rlabel metal3 82 160020 82 160020 0 Tile_X0Y5_UIO_IN_TT_PROJECT1
rlabel metal3 82 160524 82 160524 0 Tile_X0Y5_UIO_IN_TT_PROJECT2
rlabel metal3 82 161028 82 161028 0 Tile_X0Y5_UIO_IN_TT_PROJECT3
rlabel metal3 82 161532 82 161532 0 Tile_X0Y5_UIO_IN_TT_PROJECT4
rlabel metal3 82 162036 82 162036 0 Tile_X0Y5_UIO_IN_TT_PROJECT5
rlabel metal3 82 162540 82 162540 0 Tile_X0Y5_UIO_IN_TT_PROJECT6
rlabel metal3 82 163044 82 163044 0 Tile_X0Y5_UIO_IN_TT_PROJECT7
rlabel metal3 82 151452 82 151452 0 Tile_X0Y5_UIO_OE_TT_PROJECT0
rlabel metal3 82 151956 82 151956 0 Tile_X0Y5_UIO_OE_TT_PROJECT1
rlabel metal3 82 152460 82 152460 0 Tile_X0Y5_UIO_OE_TT_PROJECT2
rlabel metal3 82 152964 82 152964 0 Tile_X0Y5_UIO_OE_TT_PROJECT3
rlabel metal3 82 153468 82 153468 0 Tile_X0Y5_UIO_OE_TT_PROJECT4
rlabel metal3 82 153972 82 153972 0 Tile_X0Y5_UIO_OE_TT_PROJECT5
rlabel metal3 82 154476 82 154476 0 Tile_X0Y5_UIO_OE_TT_PROJECT6
rlabel metal3 82 154980 82 154980 0 Tile_X0Y5_UIO_OE_TT_PROJECT7
rlabel metal3 82 147420 82 147420 0 Tile_X0Y5_UIO_OUT_TT_PROJECT0
rlabel metal3 82 147924 82 147924 0 Tile_X0Y5_UIO_OUT_TT_PROJECT1
rlabel metal3 82 148428 82 148428 0 Tile_X0Y5_UIO_OUT_TT_PROJECT2
rlabel metal3 82 148932 82 148932 0 Tile_X0Y5_UIO_OUT_TT_PROJECT3
rlabel metal3 82 149436 82 149436 0 Tile_X0Y5_UIO_OUT_TT_PROJECT4
rlabel metal3 82 149940 82 149940 0 Tile_X0Y5_UIO_OUT_TT_PROJECT5
rlabel metal3 82 150444 82 150444 0 Tile_X0Y5_UIO_OUT_TT_PROJECT6
rlabel metal3 82 150948 82 150948 0 Tile_X0Y5_UIO_OUT_TT_PROJECT7
rlabel metal3 82 155484 82 155484 0 Tile_X0Y5_UI_IN_TT_PROJECT0
rlabel metal3 82 155988 82 155988 0 Tile_X0Y5_UI_IN_TT_PROJECT1
rlabel metal3 82 156492 82 156492 0 Tile_X0Y5_UI_IN_TT_PROJECT2
rlabel metal3 82 156996 82 156996 0 Tile_X0Y5_UI_IN_TT_PROJECT3
rlabel metal3 82 157500 82 157500 0 Tile_X0Y5_UI_IN_TT_PROJECT4
rlabel metal3 82 158004 82 158004 0 Tile_X0Y5_UI_IN_TT_PROJECT5
rlabel metal3 82 158508 82 158508 0 Tile_X0Y5_UI_IN_TT_PROJECT6
rlabel metal3 82 159012 82 159012 0 Tile_X0Y5_UI_IN_TT_PROJECT7
rlabel metal3 82 143388 82 143388 0 Tile_X0Y5_UO_OUT_TT_PROJECT0
rlabel metal3 82 143892 82 143892 0 Tile_X0Y5_UO_OUT_TT_PROJECT1
rlabel metal3 82 144396 82 144396 0 Tile_X0Y5_UO_OUT_TT_PROJECT2
rlabel metal3 82 144900 82 144900 0 Tile_X0Y5_UO_OUT_TT_PROJECT3
rlabel metal3 82 145404 82 145404 0 Tile_X0Y5_UO_OUT_TT_PROJECT4
rlabel metal3 82 145908 82 145908 0 Tile_X0Y5_UO_OUT_TT_PROJECT5
rlabel metal3 82 146412 82 146412 0 Tile_X0Y5_UO_OUT_TT_PROJECT6
rlabel metal3 82 146916 82 146916 0 Tile_X0Y5_UO_OUT_TT_PROJECT7
rlabel metal3 82 121044 82 121044 0 Tile_X0Y6_CLK_TT_PROJECT
rlabel metal3 82 120540 82 120540 0 Tile_X0Y6_ENA_TT_PROJECT
rlabel metal3 82 121548 82 121548 0 Tile_X0Y6_RST_N_TT_PROJECT
rlabel metal3 82 116508 82 116508 0 Tile_X0Y6_UIO_IN_TT_PROJECT0
rlabel metal3 82 117012 82 117012 0 Tile_X0Y6_UIO_IN_TT_PROJECT1
rlabel metal3 82 117516 82 117516 0 Tile_X0Y6_UIO_IN_TT_PROJECT2
rlabel metal3 82 118020 82 118020 0 Tile_X0Y6_UIO_IN_TT_PROJECT3
rlabel metal3 82 118524 82 118524 0 Tile_X0Y6_UIO_IN_TT_PROJECT4
rlabel metal3 82 119028 82 119028 0 Tile_X0Y6_UIO_IN_TT_PROJECT5
rlabel metal3 82 119532 82 119532 0 Tile_X0Y6_UIO_IN_TT_PROJECT6
rlabel metal3 82 120036 82 120036 0 Tile_X0Y6_UIO_IN_TT_PROJECT7
rlabel metal3 82 108444 82 108444 0 Tile_X0Y6_UIO_OE_TT_PROJECT0
rlabel metal3 82 108948 82 108948 0 Tile_X0Y6_UIO_OE_TT_PROJECT1
rlabel metal3 82 109452 82 109452 0 Tile_X0Y6_UIO_OE_TT_PROJECT2
rlabel metal3 82 109956 82 109956 0 Tile_X0Y6_UIO_OE_TT_PROJECT3
rlabel metal3 82 110460 82 110460 0 Tile_X0Y6_UIO_OE_TT_PROJECT4
rlabel metal3 82 110964 82 110964 0 Tile_X0Y6_UIO_OE_TT_PROJECT5
rlabel metal3 82 111468 82 111468 0 Tile_X0Y6_UIO_OE_TT_PROJECT6
rlabel metal3 82 111972 82 111972 0 Tile_X0Y6_UIO_OE_TT_PROJECT7
rlabel metal3 82 104412 82 104412 0 Tile_X0Y6_UIO_OUT_TT_PROJECT0
rlabel metal3 82 104916 82 104916 0 Tile_X0Y6_UIO_OUT_TT_PROJECT1
rlabel metal3 82 105420 82 105420 0 Tile_X0Y6_UIO_OUT_TT_PROJECT2
rlabel metal3 82 105924 82 105924 0 Tile_X0Y6_UIO_OUT_TT_PROJECT3
rlabel metal3 82 106428 82 106428 0 Tile_X0Y6_UIO_OUT_TT_PROJECT4
rlabel metal3 82 106932 82 106932 0 Tile_X0Y6_UIO_OUT_TT_PROJECT5
rlabel metal3 82 107436 82 107436 0 Tile_X0Y6_UIO_OUT_TT_PROJECT6
rlabel metal3 82 107940 82 107940 0 Tile_X0Y6_UIO_OUT_TT_PROJECT7
rlabel metal3 82 112476 82 112476 0 Tile_X0Y6_UI_IN_TT_PROJECT0
rlabel metal3 82 112980 82 112980 0 Tile_X0Y6_UI_IN_TT_PROJECT1
rlabel metal3 82 113484 82 113484 0 Tile_X0Y6_UI_IN_TT_PROJECT2
rlabel metal3 82 113988 82 113988 0 Tile_X0Y6_UI_IN_TT_PROJECT3
rlabel metal3 82 114492 82 114492 0 Tile_X0Y6_UI_IN_TT_PROJECT4
rlabel metal3 82 114996 82 114996 0 Tile_X0Y6_UI_IN_TT_PROJECT5
rlabel metal3 82 115500 82 115500 0 Tile_X0Y6_UI_IN_TT_PROJECT6
rlabel metal3 82 116004 82 116004 0 Tile_X0Y6_UI_IN_TT_PROJECT7
rlabel metal3 82 100380 82 100380 0 Tile_X0Y6_UO_OUT_TT_PROJECT0
rlabel metal3 82 100884 82 100884 0 Tile_X0Y6_UO_OUT_TT_PROJECT1
rlabel metal3 82 101388 82 101388 0 Tile_X0Y6_UO_OUT_TT_PROJECT2
rlabel metal3 82 101892 82 101892 0 Tile_X0Y6_UO_OUT_TT_PROJECT3
rlabel metal3 82 102396 82 102396 0 Tile_X0Y6_UO_OUT_TT_PROJECT4
rlabel metal3 82 102900 82 102900 0 Tile_X0Y6_UO_OUT_TT_PROJECT5
rlabel metal3 82 103404 82 103404 0 Tile_X0Y6_UO_OUT_TT_PROJECT6
rlabel metal3 82 103908 82 103908 0 Tile_X0Y6_UO_OUT_TT_PROJECT7
rlabel metal3 82 78036 82 78036 0 Tile_X0Y7_CLK_TT_PROJECT
rlabel metal3 82 77532 82 77532 0 Tile_X0Y7_ENA_TT_PROJECT
rlabel metal3 82 78540 82 78540 0 Tile_X0Y7_RST_N_TT_PROJECT
rlabel metal3 82 73500 82 73500 0 Tile_X0Y7_UIO_IN_TT_PROJECT0
rlabel metal3 82 74004 82 74004 0 Tile_X0Y7_UIO_IN_TT_PROJECT1
rlabel metal3 82 74508 82 74508 0 Tile_X0Y7_UIO_IN_TT_PROJECT2
rlabel metal3 82 75012 82 75012 0 Tile_X0Y7_UIO_IN_TT_PROJECT3
rlabel metal3 82 75516 82 75516 0 Tile_X0Y7_UIO_IN_TT_PROJECT4
rlabel metal3 82 76020 82 76020 0 Tile_X0Y7_UIO_IN_TT_PROJECT5
rlabel metal3 82 76524 82 76524 0 Tile_X0Y7_UIO_IN_TT_PROJECT6
rlabel metal3 82 77028 82 77028 0 Tile_X0Y7_UIO_IN_TT_PROJECT7
rlabel metal3 82 65436 82 65436 0 Tile_X0Y7_UIO_OE_TT_PROJECT0
rlabel metal3 82 65940 82 65940 0 Tile_X0Y7_UIO_OE_TT_PROJECT1
rlabel metal3 82 66444 82 66444 0 Tile_X0Y7_UIO_OE_TT_PROJECT2
rlabel metal3 82 66948 82 66948 0 Tile_X0Y7_UIO_OE_TT_PROJECT3
rlabel metal3 82 67452 82 67452 0 Tile_X0Y7_UIO_OE_TT_PROJECT4
rlabel metal3 82 67956 82 67956 0 Tile_X0Y7_UIO_OE_TT_PROJECT5
rlabel metal3 82 68460 82 68460 0 Tile_X0Y7_UIO_OE_TT_PROJECT6
rlabel metal3 82 68964 82 68964 0 Tile_X0Y7_UIO_OE_TT_PROJECT7
rlabel metal3 82 61404 82 61404 0 Tile_X0Y7_UIO_OUT_TT_PROJECT0
rlabel metal3 82 61908 82 61908 0 Tile_X0Y7_UIO_OUT_TT_PROJECT1
rlabel metal3 82 62412 82 62412 0 Tile_X0Y7_UIO_OUT_TT_PROJECT2
rlabel metal3 82 62916 82 62916 0 Tile_X0Y7_UIO_OUT_TT_PROJECT3
rlabel metal3 82 63420 82 63420 0 Tile_X0Y7_UIO_OUT_TT_PROJECT4
rlabel metal3 82 63924 82 63924 0 Tile_X0Y7_UIO_OUT_TT_PROJECT5
rlabel metal3 82 64428 82 64428 0 Tile_X0Y7_UIO_OUT_TT_PROJECT6
rlabel metal3 82 64932 82 64932 0 Tile_X0Y7_UIO_OUT_TT_PROJECT7
rlabel metal3 82 69468 82 69468 0 Tile_X0Y7_UI_IN_TT_PROJECT0
rlabel metal3 82 69972 82 69972 0 Tile_X0Y7_UI_IN_TT_PROJECT1
rlabel metal3 82 70476 82 70476 0 Tile_X0Y7_UI_IN_TT_PROJECT2
rlabel metal3 82 70980 82 70980 0 Tile_X0Y7_UI_IN_TT_PROJECT3
rlabel metal3 82 71484 82 71484 0 Tile_X0Y7_UI_IN_TT_PROJECT4
rlabel metal3 82 71988 82 71988 0 Tile_X0Y7_UI_IN_TT_PROJECT5
rlabel metal3 82 72492 82 72492 0 Tile_X0Y7_UI_IN_TT_PROJECT6
rlabel metal3 82 72996 82 72996 0 Tile_X0Y7_UI_IN_TT_PROJECT7
rlabel metal3 82 57372 82 57372 0 Tile_X0Y7_UO_OUT_TT_PROJECT0
rlabel metal3 82 57876 82 57876 0 Tile_X0Y7_UO_OUT_TT_PROJECT1
rlabel metal3 82 58380 82 58380 0 Tile_X0Y7_UO_OUT_TT_PROJECT2
rlabel metal3 82 58884 82 58884 0 Tile_X0Y7_UO_OUT_TT_PROJECT3
rlabel metal3 82 59388 82 59388 0 Tile_X0Y7_UO_OUT_TT_PROJECT4
rlabel metal3 82 59892 82 59892 0 Tile_X0Y7_UO_OUT_TT_PROJECT5
rlabel metal3 82 60396 82 60396 0 Tile_X0Y7_UO_OUT_TT_PROJECT6
rlabel metal3 82 60900 82 60900 0 Tile_X0Y7_UO_OUT_TT_PROJECT7
rlabel metal3 82 35028 82 35028 0 Tile_X0Y8_CLK_TT_PROJECT
rlabel metal3 82 34524 82 34524 0 Tile_X0Y8_ENA_TT_PROJECT
rlabel metal3 82 35532 82 35532 0 Tile_X0Y8_RST_N_TT_PROJECT
rlabel metal3 82 30492 82 30492 0 Tile_X0Y8_UIO_IN_TT_PROJECT0
rlabel metal3 82 30996 82 30996 0 Tile_X0Y8_UIO_IN_TT_PROJECT1
rlabel metal3 82 31500 82 31500 0 Tile_X0Y8_UIO_IN_TT_PROJECT2
rlabel metal3 82 32004 82 32004 0 Tile_X0Y8_UIO_IN_TT_PROJECT3
rlabel metal3 82 32508 82 32508 0 Tile_X0Y8_UIO_IN_TT_PROJECT4
rlabel metal3 82 33012 82 33012 0 Tile_X0Y8_UIO_IN_TT_PROJECT5
rlabel metal3 82 33516 82 33516 0 Tile_X0Y8_UIO_IN_TT_PROJECT6
rlabel metal3 82 34020 82 34020 0 Tile_X0Y8_UIO_IN_TT_PROJECT7
rlabel metal3 82 22428 82 22428 0 Tile_X0Y8_UIO_OE_TT_PROJECT0
rlabel metal3 82 22932 82 22932 0 Tile_X0Y8_UIO_OE_TT_PROJECT1
rlabel metal3 82 23436 82 23436 0 Tile_X0Y8_UIO_OE_TT_PROJECT2
rlabel metal3 82 23940 82 23940 0 Tile_X0Y8_UIO_OE_TT_PROJECT3
rlabel metal3 82 24444 82 24444 0 Tile_X0Y8_UIO_OE_TT_PROJECT4
rlabel metal3 82 24948 82 24948 0 Tile_X0Y8_UIO_OE_TT_PROJECT5
rlabel metal3 82 25452 82 25452 0 Tile_X0Y8_UIO_OE_TT_PROJECT6
rlabel metal3 82 25956 82 25956 0 Tile_X0Y8_UIO_OE_TT_PROJECT7
rlabel metal3 82 18396 82 18396 0 Tile_X0Y8_UIO_OUT_TT_PROJECT0
rlabel metal3 82 18900 82 18900 0 Tile_X0Y8_UIO_OUT_TT_PROJECT1
rlabel metal3 82 19404 82 19404 0 Tile_X0Y8_UIO_OUT_TT_PROJECT2
rlabel metal3 82 19908 82 19908 0 Tile_X0Y8_UIO_OUT_TT_PROJECT3
rlabel metal3 82 20412 82 20412 0 Tile_X0Y8_UIO_OUT_TT_PROJECT4
rlabel metal3 82 20916 82 20916 0 Tile_X0Y8_UIO_OUT_TT_PROJECT5
rlabel metal3 82 21420 82 21420 0 Tile_X0Y8_UIO_OUT_TT_PROJECT6
rlabel metal3 82 21924 82 21924 0 Tile_X0Y8_UIO_OUT_TT_PROJECT7
rlabel metal3 82 26460 82 26460 0 Tile_X0Y8_UI_IN_TT_PROJECT0
rlabel metal3 82 26964 82 26964 0 Tile_X0Y8_UI_IN_TT_PROJECT1
rlabel metal3 82 27468 82 27468 0 Tile_X0Y8_UI_IN_TT_PROJECT2
rlabel metal3 82 27972 82 27972 0 Tile_X0Y8_UI_IN_TT_PROJECT3
rlabel metal3 82 28476 82 28476 0 Tile_X0Y8_UI_IN_TT_PROJECT4
rlabel metal3 82 28980 82 28980 0 Tile_X0Y8_UI_IN_TT_PROJECT5
rlabel metal3 82 29484 82 29484 0 Tile_X0Y8_UI_IN_TT_PROJECT6
rlabel metal3 82 29988 82 29988 0 Tile_X0Y8_UI_IN_TT_PROJECT7
rlabel metal3 82 14364 82 14364 0 Tile_X0Y8_UO_OUT_TT_PROJECT0
rlabel metal3 82 14868 82 14868 0 Tile_X0Y8_UO_OUT_TT_PROJECT1
rlabel metal3 82 15372 82 15372 0 Tile_X0Y8_UO_OUT_TT_PROJECT2
rlabel metal3 82 15876 82 15876 0 Tile_X0Y8_UO_OUT_TT_PROJECT3
rlabel metal3 82 16380 82 16380 0 Tile_X0Y8_UO_OUT_TT_PROJECT4
rlabel metal3 82 16884 82 16884 0 Tile_X0Y8_UO_OUT_TT_PROJECT5
rlabel metal3 82 17388 82 17388 0 Tile_X0Y8_UO_OUT_TT_PROJECT6
rlabel metal3 82 17892 82 17892 0 Tile_X0Y8_UO_OUT_TT_PROJECT7
rlabel metal2 25728 366421 25728 366421 0 Tile_X1Y0_A_I_top
rlabel metal2 24576 366421 24576 366421 0 Tile_X1Y0_A_O_top
rlabel metal2 26880 366421 26880 366421 0 Tile_X1Y0_A_T_top
rlabel metal2 29184 366421 29184 366421 0 Tile_X1Y0_B_I_top
rlabel metal2 28032 366421 28032 366421 0 Tile_X1Y0_B_O_top
rlabel metal2 30336 366421 30336 366421 0 Tile_X1Y0_B_T_top
rlabel metal2 32640 366421 32640 366421 0 Tile_X1Y0_C_I_top
rlabel metal2 31488 366421 31488 366421 0 Tile_X1Y0_C_O_top
rlabel metal2 33792 366421 33792 366421 0 Tile_X1Y0_C_T_top
rlabel metal2 36096 366421 36096 366421 0 Tile_X1Y0_D_I_top
rlabel metal2 34944 366421 34944 366421 0 Tile_X1Y0_D_O_top
rlabel metal2 37248 366421 37248 366421 0 Tile_X1Y0_D_T_top
rlabel metal2 25728 454 25728 454 0 Tile_X1Y9_A_I_top
rlabel metal2 24576 454 24576 454 0 Tile_X1Y9_A_O_top
rlabel metal2 26880 454 26880 454 0 Tile_X1Y9_A_T_top
rlabel metal2 29184 454 29184 454 0 Tile_X1Y9_B_I_top
rlabel metal2 28032 454 28032 454 0 Tile_X1Y9_B_O_top
rlabel metal2 30336 454 30336 454 0 Tile_X1Y9_B_T_top
rlabel metal2 32640 454 32640 454 0 Tile_X1Y9_C_I_top
rlabel metal2 31488 454 31488 454 0 Tile_X1Y9_C_O_top
rlabel metal2 33792 454 33792 454 0 Tile_X1Y9_C_T_top
rlabel metal2 36096 454 36096 454 0 Tile_X1Y9_D_I_top
rlabel metal2 34944 454 34944 454 0 Tile_X1Y9_D_O_top
rlabel metal2 37248 454 37248 454 0 Tile_X1Y9_D_T_top
rlabel metal2 68736 366421 68736 366421 0 Tile_X2Y0_A_I_top
rlabel metal2 67584 366421 67584 366421 0 Tile_X2Y0_A_O_top
rlabel metal2 69888 366421 69888 366421 0 Tile_X2Y0_A_T_top
rlabel metal2 72192 366421 72192 366421 0 Tile_X2Y0_B_I_top
rlabel metal2 71040 366421 71040 366421 0 Tile_X2Y0_B_O_top
rlabel metal2 73344 366421 73344 366421 0 Tile_X2Y0_B_T_top
rlabel metal2 75648 366421 75648 366421 0 Tile_X2Y0_C_I_top
rlabel metal2 74496 366421 74496 366421 0 Tile_X2Y0_C_O_top
rlabel metal2 76800 366421 76800 366421 0 Tile_X2Y0_C_T_top
rlabel metal2 79104 366421 79104 366421 0 Tile_X2Y0_D_I_top
rlabel metal2 77952 366421 77952 366421 0 Tile_X2Y0_D_O_top
rlabel metal2 80256 366421 80256 366421 0 Tile_X2Y0_D_T_top
rlabel metal2 68736 454 68736 454 0 Tile_X2Y9_A_I_top
rlabel metal2 67584 454 67584 454 0 Tile_X2Y9_A_O_top
rlabel metal2 69888 454 69888 454 0 Tile_X2Y9_A_T_top
rlabel metal2 72192 454 72192 454 0 Tile_X2Y9_B_I_top
rlabel metal2 71040 454 71040 454 0 Tile_X2Y9_B_O_top
rlabel metal2 73344 454 73344 454 0 Tile_X2Y9_B_T_top
rlabel metal2 75648 454 75648 454 0 Tile_X2Y9_C_I_top
rlabel metal2 74496 454 74496 454 0 Tile_X2Y9_C_O_top
rlabel metal2 76800 454 76800 454 0 Tile_X2Y9_C_T_top
rlabel metal2 79104 454 79104 454 0 Tile_X2Y9_D_I_top
rlabel metal2 77952 454 77952 454 0 Tile_X2Y9_D_O_top
rlabel metal2 80256 454 80256 454 0 Tile_X2Y9_D_T_top
rlabel metal2 111744 366421 111744 366421 0 Tile_X3Y0_A_I_top
rlabel metal2 110592 366421 110592 366421 0 Tile_X3Y0_A_O_top
rlabel metal2 112896 366421 112896 366421 0 Tile_X3Y0_A_T_top
rlabel metal2 115200 366421 115200 366421 0 Tile_X3Y0_B_I_top
rlabel metal2 114048 366421 114048 366421 0 Tile_X3Y0_B_O_top
rlabel metal2 116352 366421 116352 366421 0 Tile_X3Y0_B_T_top
rlabel metal2 118656 366421 118656 366421 0 Tile_X3Y0_C_I_top
rlabel metal2 117504 366421 117504 366421 0 Tile_X3Y0_C_O_top
rlabel metal2 119808 366421 119808 366421 0 Tile_X3Y0_C_T_top
rlabel metal2 122112 366421 122112 366421 0 Tile_X3Y0_D_I_top
rlabel metal2 120960 366421 120960 366421 0 Tile_X3Y0_D_O_top
rlabel metal2 123264 366421 123264 366421 0 Tile_X3Y0_D_T_top
rlabel metal2 111744 454 111744 454 0 Tile_X3Y9_A_I_top
rlabel metal2 110592 454 110592 454 0 Tile_X3Y9_A_O_top
rlabel metal2 112896 454 112896 454 0 Tile_X3Y9_A_T_top
rlabel metal2 115200 454 115200 454 0 Tile_X3Y9_B_I_top
rlabel metal2 114048 454 114048 454 0 Tile_X3Y9_B_O_top
rlabel metal2 116352 454 116352 454 0 Tile_X3Y9_B_T_top
rlabel metal2 118656 454 118656 454 0 Tile_X3Y9_C_I_top
rlabel metal2 117504 454 117504 454 0 Tile_X3Y9_C_O_top
rlabel metal2 119808 454 119808 454 0 Tile_X3Y9_C_T_top
rlabel metal2 122112 454 122112 454 0 Tile_X3Y9_D_I_top
rlabel metal2 120960 454 120960 454 0 Tile_X3Y9_D_O_top
rlabel metal2 123264 454 123264 454 0 Tile_X3Y9_D_T_top
rlabel metal2 154752 366421 154752 366421 0 Tile_X4Y0_A_I_top
rlabel metal2 153600 366421 153600 366421 0 Tile_X4Y0_A_O_top
rlabel metal2 155904 366421 155904 366421 0 Tile_X4Y0_A_T_top
rlabel metal2 158208 366421 158208 366421 0 Tile_X4Y0_B_I_top
rlabel metal2 157056 366421 157056 366421 0 Tile_X4Y0_B_O_top
rlabel metal2 159360 366421 159360 366421 0 Tile_X4Y0_B_T_top
rlabel metal2 161664 366421 161664 366421 0 Tile_X4Y0_C_I_top
rlabel metal2 160512 366421 160512 366421 0 Tile_X4Y0_C_O_top
rlabel metal2 162816 366421 162816 366421 0 Tile_X4Y0_C_T_top
rlabel metal2 165120 366421 165120 366421 0 Tile_X4Y0_D_I_top
rlabel metal2 163968 366421 163968 366421 0 Tile_X4Y0_D_O_top
rlabel metal2 166272 366421 166272 366421 0 Tile_X4Y0_D_T_top
rlabel metal2 154752 454 154752 454 0 Tile_X4Y9_A_I_top
rlabel metal2 153600 454 153600 454 0 Tile_X4Y9_A_O_top
rlabel metal2 155904 454 155904 454 0 Tile_X4Y9_A_T_top
rlabel metal2 158208 454 158208 454 0 Tile_X4Y9_B_I_top
rlabel metal2 157056 454 157056 454 0 Tile_X4Y9_B_O_top
rlabel metal2 159360 454 159360 454 0 Tile_X4Y9_B_T_top
rlabel metal2 161664 454 161664 454 0 Tile_X4Y9_C_I_top
rlabel metal2 160512 454 160512 454 0 Tile_X4Y9_C_O_top
rlabel metal2 162816 454 162816 454 0 Tile_X4Y9_C_T_top
rlabel metal2 165120 454 165120 454 0 Tile_X4Y9_D_I_top
rlabel metal2 163968 454 163968 454 0 Tile_X4Y9_D_O_top
rlabel metal2 166272 454 166272 454 0 Tile_X4Y9_D_T_top
rlabel metal3 215149 294084 215149 294084 0 Tile_X5Y2_ADDR_SRAM0
rlabel metal3 215149 294420 215149 294420 0 Tile_X5Y2_ADDR_SRAM1
rlabel metal3 215149 294756 215149 294756 0 Tile_X5Y2_ADDR_SRAM2
rlabel metal3 215149 295092 215149 295092 0 Tile_X5Y2_ADDR_SRAM3
rlabel metal3 215149 295428 215149 295428 0 Tile_X5Y2_ADDR_SRAM4
rlabel metal3 215149 295764 215149 295764 0 Tile_X5Y2_ADDR_SRAM5
rlabel metal3 215149 296100 215149 296100 0 Tile_X5Y2_ADDR_SRAM6
rlabel metal3 215149 296436 215149 296436 0 Tile_X5Y2_ADDR_SRAM7
rlabel metal3 215149 296772 215149 296772 0 Tile_X5Y2_ADDR_SRAM8
rlabel metal3 215149 297108 215149 297108 0 Tile_X5Y2_ADDR_SRAM9
rlabel metal3 215149 308196 215149 308196 0 Tile_X5Y2_BM_SRAM0
rlabel metal3 215149 308532 215149 308532 0 Tile_X5Y2_BM_SRAM1
rlabel metal3 215149 311556 215149 311556 0 Tile_X5Y2_BM_SRAM10
rlabel metal3 215149 311892 215149 311892 0 Tile_X5Y2_BM_SRAM11
rlabel metal3 215149 312228 215149 312228 0 Tile_X5Y2_BM_SRAM12
rlabel metal3 215149 312564 215149 312564 0 Tile_X5Y2_BM_SRAM13
rlabel metal3 215149 312900 215149 312900 0 Tile_X5Y2_BM_SRAM14
rlabel metal3 215149 313236 215149 313236 0 Tile_X5Y2_BM_SRAM15
rlabel metal3 215149 313572 215149 313572 0 Tile_X5Y2_BM_SRAM16
rlabel metal3 215149 313908 215149 313908 0 Tile_X5Y2_BM_SRAM17
rlabel metal3 215149 314244 215149 314244 0 Tile_X5Y2_BM_SRAM18
rlabel metal3 215149 314580 215149 314580 0 Tile_X5Y2_BM_SRAM19
rlabel metal3 215149 308868 215149 308868 0 Tile_X5Y2_BM_SRAM2
rlabel metal3 215149 314916 215149 314916 0 Tile_X5Y2_BM_SRAM20
rlabel metal3 215149 315252 215149 315252 0 Tile_X5Y2_BM_SRAM21
rlabel metal3 215149 315588 215149 315588 0 Tile_X5Y2_BM_SRAM22
rlabel metal3 215149 315924 215149 315924 0 Tile_X5Y2_BM_SRAM23
rlabel metal3 215149 316260 215149 316260 0 Tile_X5Y2_BM_SRAM24
rlabel metal3 215149 316596 215149 316596 0 Tile_X5Y2_BM_SRAM25
rlabel metal3 215149 316932 215149 316932 0 Tile_X5Y2_BM_SRAM26
rlabel metal3 215149 317268 215149 317268 0 Tile_X5Y2_BM_SRAM27
rlabel metal3 215149 317604 215149 317604 0 Tile_X5Y2_BM_SRAM28
rlabel metal3 215149 317940 215149 317940 0 Tile_X5Y2_BM_SRAM29
rlabel metal3 215149 309204 215149 309204 0 Tile_X5Y2_BM_SRAM3
rlabel metal3 215149 318276 215149 318276 0 Tile_X5Y2_BM_SRAM30
rlabel metal3 215149 318612 215149 318612 0 Tile_X5Y2_BM_SRAM31
rlabel metal3 215149 309540 215149 309540 0 Tile_X5Y2_BM_SRAM4
rlabel metal3 215149 309876 215149 309876 0 Tile_X5Y2_BM_SRAM5
rlabel metal3 215149 310212 215149 310212 0 Tile_X5Y2_BM_SRAM6
rlabel metal3 215149 310548 215149 310548 0 Tile_X5Y2_BM_SRAM7
rlabel metal3 215149 310884 215149 310884 0 Tile_X5Y2_BM_SRAM8
rlabel metal3 215149 311220 215149 311220 0 Tile_X5Y2_BM_SRAM9
rlabel metal3 215149 319956 215149 319956 0 Tile_X5Y2_CLK_SRAM
rlabel metal3 215149 293748 215149 293748 0 Tile_X5Y2_CONFIGURED_top
rlabel metal3 215149 297444 215149 297444 0 Tile_X5Y2_DIN_SRAM0
rlabel metal3 215149 297780 215149 297780 0 Tile_X5Y2_DIN_SRAM1
rlabel metal3 215149 300804 215149 300804 0 Tile_X5Y2_DIN_SRAM10
rlabel metal3 215149 301140 215149 301140 0 Tile_X5Y2_DIN_SRAM11
rlabel metal3 215149 301476 215149 301476 0 Tile_X5Y2_DIN_SRAM12
rlabel metal3 215149 301812 215149 301812 0 Tile_X5Y2_DIN_SRAM13
rlabel metal3 215149 302148 215149 302148 0 Tile_X5Y2_DIN_SRAM14
rlabel metal3 215149 302484 215149 302484 0 Tile_X5Y2_DIN_SRAM15
rlabel metal3 215149 302820 215149 302820 0 Tile_X5Y2_DIN_SRAM16
rlabel metal3 215149 303156 215149 303156 0 Tile_X5Y2_DIN_SRAM17
rlabel metal3 215149 303492 215149 303492 0 Tile_X5Y2_DIN_SRAM18
rlabel metal3 215149 303828 215149 303828 0 Tile_X5Y2_DIN_SRAM19
rlabel metal3 215149 298116 215149 298116 0 Tile_X5Y2_DIN_SRAM2
rlabel metal3 215149 304164 215149 304164 0 Tile_X5Y2_DIN_SRAM20
rlabel metal3 215149 304500 215149 304500 0 Tile_X5Y2_DIN_SRAM21
rlabel metal3 215149 304836 215149 304836 0 Tile_X5Y2_DIN_SRAM22
rlabel metal3 215149 305172 215149 305172 0 Tile_X5Y2_DIN_SRAM23
rlabel metal3 215149 305508 215149 305508 0 Tile_X5Y2_DIN_SRAM24
rlabel metal3 215149 305844 215149 305844 0 Tile_X5Y2_DIN_SRAM25
rlabel metal3 215149 306180 215149 306180 0 Tile_X5Y2_DIN_SRAM26
rlabel metal3 215149 306516 215149 306516 0 Tile_X5Y2_DIN_SRAM27
rlabel metal3 215149 306852 215149 306852 0 Tile_X5Y2_DIN_SRAM28
rlabel metal3 215149 307188 215149 307188 0 Tile_X5Y2_DIN_SRAM29
rlabel metal3 215149 298452 215149 298452 0 Tile_X5Y2_DIN_SRAM3
rlabel metal3 215149 307524 215149 307524 0 Tile_X5Y2_DIN_SRAM30
rlabel metal3 215149 307860 215149 307860 0 Tile_X5Y2_DIN_SRAM31
rlabel metal3 215149 298788 215149 298788 0 Tile_X5Y2_DIN_SRAM4
rlabel metal3 215149 299124 215149 299124 0 Tile_X5Y2_DIN_SRAM5
rlabel metal3 215149 299460 215149 299460 0 Tile_X5Y2_DIN_SRAM6
rlabel metal3 215149 299796 215149 299796 0 Tile_X5Y2_DIN_SRAM7
rlabel metal3 215149 300132 215149 300132 0 Tile_X5Y2_DIN_SRAM8
rlabel metal3 215149 300468 215149 300468 0 Tile_X5Y2_DIN_SRAM9
rlabel metal3 215149 282996 215149 282996 0 Tile_X5Y2_DOUT_SRAM0
rlabel metal3 215149 283332 215149 283332 0 Tile_X5Y2_DOUT_SRAM1
rlabel metal3 215149 286356 215149 286356 0 Tile_X5Y2_DOUT_SRAM10
rlabel metal3 215149 286692 215149 286692 0 Tile_X5Y2_DOUT_SRAM11
rlabel metal3 215149 287028 215149 287028 0 Tile_X5Y2_DOUT_SRAM12
rlabel metal3 215149 287364 215149 287364 0 Tile_X5Y2_DOUT_SRAM13
rlabel metal3 215149 287700 215149 287700 0 Tile_X5Y2_DOUT_SRAM14
rlabel metal3 215149 288036 215149 288036 0 Tile_X5Y2_DOUT_SRAM15
rlabel metal3 215149 288372 215149 288372 0 Tile_X5Y2_DOUT_SRAM16
rlabel metal3 215149 288708 215149 288708 0 Tile_X5Y2_DOUT_SRAM17
rlabel metal3 215149 289044 215149 289044 0 Tile_X5Y2_DOUT_SRAM18
rlabel metal3 215149 289380 215149 289380 0 Tile_X5Y2_DOUT_SRAM19
rlabel metal3 215149 283668 215149 283668 0 Tile_X5Y2_DOUT_SRAM2
rlabel metal3 215149 289716 215149 289716 0 Tile_X5Y2_DOUT_SRAM20
rlabel metal3 215149 290052 215149 290052 0 Tile_X5Y2_DOUT_SRAM21
rlabel metal3 215149 290388 215149 290388 0 Tile_X5Y2_DOUT_SRAM22
rlabel metal3 215149 290724 215149 290724 0 Tile_X5Y2_DOUT_SRAM23
rlabel metal3 215149 291060 215149 291060 0 Tile_X5Y2_DOUT_SRAM24
rlabel metal3 215149 291396 215149 291396 0 Tile_X5Y2_DOUT_SRAM25
rlabel metal3 215149 291732 215149 291732 0 Tile_X5Y2_DOUT_SRAM26
rlabel metal3 215149 292068 215149 292068 0 Tile_X5Y2_DOUT_SRAM27
rlabel metal3 215149 292404 215149 292404 0 Tile_X5Y2_DOUT_SRAM28
rlabel metal3 215149 292740 215149 292740 0 Tile_X5Y2_DOUT_SRAM29
rlabel metal3 215149 284004 215149 284004 0 Tile_X5Y2_DOUT_SRAM3
rlabel metal3 215149 293076 215149 293076 0 Tile_X5Y2_DOUT_SRAM30
rlabel metal3 215149 293412 215149 293412 0 Tile_X5Y2_DOUT_SRAM31
rlabel metal3 215149 284340 215149 284340 0 Tile_X5Y2_DOUT_SRAM4
rlabel metal3 215149 284676 215149 284676 0 Tile_X5Y2_DOUT_SRAM5
rlabel metal3 215149 285012 215149 285012 0 Tile_X5Y2_DOUT_SRAM6
rlabel metal3 215149 285348 215149 285348 0 Tile_X5Y2_DOUT_SRAM7
rlabel metal3 215149 285684 215149 285684 0 Tile_X5Y2_DOUT_SRAM8
rlabel metal3 215149 286020 215149 286020 0 Tile_X5Y2_DOUT_SRAM9
rlabel metal3 215149 319284 215149 319284 0 Tile_X5Y2_MEN_SRAM
rlabel metal3 215149 319620 215149 319620 0 Tile_X5Y2_REN_SRAM
rlabel metal3 215149 320292 215149 320292 0 Tile_X5Y2_TIE_HIGH_SRAM
rlabel metal3 215149 320628 215149 320628 0 Tile_X5Y2_TIE_LOW_SRAM
rlabel metal3 215149 318948 215149 318948 0 Tile_X5Y2_WEN_SRAM
rlabel metal3 215149 250068 215149 250068 0 Tile_X5Y3_CLK_TT_PROJECT
rlabel metal3 215149 249564 215149 249564 0 Tile_X5Y3_ENA_TT_PROJECT
rlabel metal3 215149 250572 215149 250572 0 Tile_X5Y3_RST_N_TT_PROJECT
rlabel metal3 215149 245532 215149 245532 0 Tile_X5Y3_UIO_IN_TT_PROJECT0
rlabel metal3 215149 246036 215149 246036 0 Tile_X5Y3_UIO_IN_TT_PROJECT1
rlabel metal3 215149 246540 215149 246540 0 Tile_X5Y3_UIO_IN_TT_PROJECT2
rlabel metal3 215149 247044 215149 247044 0 Tile_X5Y3_UIO_IN_TT_PROJECT3
rlabel metal3 215149 247548 215149 247548 0 Tile_X5Y3_UIO_IN_TT_PROJECT4
rlabel metal3 215149 248052 215149 248052 0 Tile_X5Y3_UIO_IN_TT_PROJECT5
rlabel metal3 215149 248556 215149 248556 0 Tile_X5Y3_UIO_IN_TT_PROJECT6
rlabel metal3 215149 249060 215149 249060 0 Tile_X5Y3_UIO_IN_TT_PROJECT7
rlabel metal3 215149 237468 215149 237468 0 Tile_X5Y3_UIO_OE_TT_PROJECT0
rlabel metal3 215149 237972 215149 237972 0 Tile_X5Y3_UIO_OE_TT_PROJECT1
rlabel metal3 215149 238476 215149 238476 0 Tile_X5Y3_UIO_OE_TT_PROJECT2
rlabel metal3 215149 238980 215149 238980 0 Tile_X5Y3_UIO_OE_TT_PROJECT3
rlabel metal3 215149 239484 215149 239484 0 Tile_X5Y3_UIO_OE_TT_PROJECT4
rlabel metal3 215149 239988 215149 239988 0 Tile_X5Y3_UIO_OE_TT_PROJECT5
rlabel metal3 215149 240492 215149 240492 0 Tile_X5Y3_UIO_OE_TT_PROJECT6
rlabel metal3 215149 240996 215149 240996 0 Tile_X5Y3_UIO_OE_TT_PROJECT7
rlabel metal3 215149 233436 215149 233436 0 Tile_X5Y3_UIO_OUT_TT_PROJECT0
rlabel metal3 215149 233940 215149 233940 0 Tile_X5Y3_UIO_OUT_TT_PROJECT1
rlabel metal3 215149 234444 215149 234444 0 Tile_X5Y3_UIO_OUT_TT_PROJECT2
rlabel metal3 215149 234948 215149 234948 0 Tile_X5Y3_UIO_OUT_TT_PROJECT3
rlabel metal3 215149 235452 215149 235452 0 Tile_X5Y3_UIO_OUT_TT_PROJECT4
rlabel metal3 215149 235956 215149 235956 0 Tile_X5Y3_UIO_OUT_TT_PROJECT5
rlabel metal3 215149 236460 215149 236460 0 Tile_X5Y3_UIO_OUT_TT_PROJECT6
rlabel metal3 215149 236964 215149 236964 0 Tile_X5Y3_UIO_OUT_TT_PROJECT7
rlabel metal3 215149 241500 215149 241500 0 Tile_X5Y3_UI_IN_TT_PROJECT0
rlabel metal3 215149 242004 215149 242004 0 Tile_X5Y3_UI_IN_TT_PROJECT1
rlabel metal3 215149 242508 215149 242508 0 Tile_X5Y3_UI_IN_TT_PROJECT2
rlabel metal3 215149 243012 215149 243012 0 Tile_X5Y3_UI_IN_TT_PROJECT3
rlabel metal3 215149 243516 215149 243516 0 Tile_X5Y3_UI_IN_TT_PROJECT4
rlabel metal3 215149 244020 215149 244020 0 Tile_X5Y3_UI_IN_TT_PROJECT5
rlabel metal3 215149 244524 215149 244524 0 Tile_X5Y3_UI_IN_TT_PROJECT6
rlabel metal3 215149 245028 215149 245028 0 Tile_X5Y3_UI_IN_TT_PROJECT7
rlabel metal3 215149 229404 215149 229404 0 Tile_X5Y3_UO_OUT_TT_PROJECT0
rlabel metal3 215149 229908 215149 229908 0 Tile_X5Y3_UO_OUT_TT_PROJECT1
rlabel metal3 215149 230412 215149 230412 0 Tile_X5Y3_UO_OUT_TT_PROJECT2
rlabel metal3 215149 230916 215149 230916 0 Tile_X5Y3_UO_OUT_TT_PROJECT3
rlabel metal3 215149 231420 215149 231420 0 Tile_X5Y3_UO_OUT_TT_PROJECT4
rlabel metal3 215149 231924 215149 231924 0 Tile_X5Y3_UO_OUT_TT_PROJECT5
rlabel metal3 215149 232428 215149 232428 0 Tile_X5Y3_UO_OUT_TT_PROJECT6
rlabel metal3 215149 232932 215149 232932 0 Tile_X5Y3_UO_OUT_TT_PROJECT7
rlabel metal3 215149 207060 215149 207060 0 Tile_X5Y4_CLK_TT_PROJECT
rlabel metal3 215149 206556 215149 206556 0 Tile_X5Y4_ENA_TT_PROJECT
rlabel metal3 215149 207564 215149 207564 0 Tile_X5Y4_RST_N_TT_PROJECT
rlabel metal3 215149 202524 215149 202524 0 Tile_X5Y4_UIO_IN_TT_PROJECT0
rlabel metal3 215149 203028 215149 203028 0 Tile_X5Y4_UIO_IN_TT_PROJECT1
rlabel metal3 215149 203532 215149 203532 0 Tile_X5Y4_UIO_IN_TT_PROJECT2
rlabel metal3 215149 204036 215149 204036 0 Tile_X5Y4_UIO_IN_TT_PROJECT3
rlabel metal3 215149 204540 215149 204540 0 Tile_X5Y4_UIO_IN_TT_PROJECT4
rlabel metal3 215149 205044 215149 205044 0 Tile_X5Y4_UIO_IN_TT_PROJECT5
rlabel metal3 215149 205548 215149 205548 0 Tile_X5Y4_UIO_IN_TT_PROJECT6
rlabel metal3 215149 206052 215149 206052 0 Tile_X5Y4_UIO_IN_TT_PROJECT7
rlabel metal3 215149 194460 215149 194460 0 Tile_X5Y4_UIO_OE_TT_PROJECT0
rlabel metal3 215149 194964 215149 194964 0 Tile_X5Y4_UIO_OE_TT_PROJECT1
rlabel metal3 215149 195468 215149 195468 0 Tile_X5Y4_UIO_OE_TT_PROJECT2
rlabel metal3 215149 195972 215149 195972 0 Tile_X5Y4_UIO_OE_TT_PROJECT3
rlabel metal3 215149 196476 215149 196476 0 Tile_X5Y4_UIO_OE_TT_PROJECT4
rlabel metal3 215149 196980 215149 196980 0 Tile_X5Y4_UIO_OE_TT_PROJECT5
rlabel metal3 215149 197484 215149 197484 0 Tile_X5Y4_UIO_OE_TT_PROJECT6
rlabel metal3 215149 197988 215149 197988 0 Tile_X5Y4_UIO_OE_TT_PROJECT7
rlabel metal3 215149 190428 215149 190428 0 Tile_X5Y4_UIO_OUT_TT_PROJECT0
rlabel metal3 215149 190932 215149 190932 0 Tile_X5Y4_UIO_OUT_TT_PROJECT1
rlabel metal3 215149 191436 215149 191436 0 Tile_X5Y4_UIO_OUT_TT_PROJECT2
rlabel metal3 215149 191940 215149 191940 0 Tile_X5Y4_UIO_OUT_TT_PROJECT3
rlabel metal3 215149 192444 215149 192444 0 Tile_X5Y4_UIO_OUT_TT_PROJECT4
rlabel metal3 215149 192948 215149 192948 0 Tile_X5Y4_UIO_OUT_TT_PROJECT5
rlabel metal3 215149 193452 215149 193452 0 Tile_X5Y4_UIO_OUT_TT_PROJECT6
rlabel metal3 215149 193956 215149 193956 0 Tile_X5Y4_UIO_OUT_TT_PROJECT7
rlabel metal3 215149 198492 215149 198492 0 Tile_X5Y4_UI_IN_TT_PROJECT0
rlabel metal3 215149 198996 215149 198996 0 Tile_X5Y4_UI_IN_TT_PROJECT1
rlabel metal3 215149 199500 215149 199500 0 Tile_X5Y4_UI_IN_TT_PROJECT2
rlabel metal3 215149 200004 215149 200004 0 Tile_X5Y4_UI_IN_TT_PROJECT3
rlabel metal3 215149 200508 215149 200508 0 Tile_X5Y4_UI_IN_TT_PROJECT4
rlabel metal3 215149 201012 215149 201012 0 Tile_X5Y4_UI_IN_TT_PROJECT5
rlabel metal3 215149 201516 215149 201516 0 Tile_X5Y4_UI_IN_TT_PROJECT6
rlabel metal3 215149 202020 215149 202020 0 Tile_X5Y4_UI_IN_TT_PROJECT7
rlabel metal3 215149 186396 215149 186396 0 Tile_X5Y4_UO_OUT_TT_PROJECT0
rlabel metal3 215149 186900 215149 186900 0 Tile_X5Y4_UO_OUT_TT_PROJECT1
rlabel metal3 215149 187404 215149 187404 0 Tile_X5Y4_UO_OUT_TT_PROJECT2
rlabel metal3 215149 187908 215149 187908 0 Tile_X5Y4_UO_OUT_TT_PROJECT3
rlabel metal3 215149 188412 215149 188412 0 Tile_X5Y4_UO_OUT_TT_PROJECT4
rlabel metal3 215149 188916 215149 188916 0 Tile_X5Y4_UO_OUT_TT_PROJECT5
rlabel metal3 215149 189420 215149 189420 0 Tile_X5Y4_UO_OUT_TT_PROJECT6
rlabel metal3 215149 189924 215149 189924 0 Tile_X5Y4_UO_OUT_TT_PROJECT7
rlabel metal3 215149 164052 215149 164052 0 Tile_X5Y5_CLK_TT_PROJECT
rlabel metal3 215149 163548 215149 163548 0 Tile_X5Y5_ENA_TT_PROJECT
rlabel metal3 215149 164556 215149 164556 0 Tile_X5Y5_RST_N_TT_PROJECT
rlabel metal3 215149 159516 215149 159516 0 Tile_X5Y5_UIO_IN_TT_PROJECT0
rlabel metal3 215149 160020 215149 160020 0 Tile_X5Y5_UIO_IN_TT_PROJECT1
rlabel metal3 215149 160524 215149 160524 0 Tile_X5Y5_UIO_IN_TT_PROJECT2
rlabel metal3 215149 161028 215149 161028 0 Tile_X5Y5_UIO_IN_TT_PROJECT3
rlabel metal3 215149 161532 215149 161532 0 Tile_X5Y5_UIO_IN_TT_PROJECT4
rlabel metal3 215149 162036 215149 162036 0 Tile_X5Y5_UIO_IN_TT_PROJECT5
rlabel metal3 215149 162540 215149 162540 0 Tile_X5Y5_UIO_IN_TT_PROJECT6
rlabel metal3 215149 163044 215149 163044 0 Tile_X5Y5_UIO_IN_TT_PROJECT7
rlabel metal3 215149 151452 215149 151452 0 Tile_X5Y5_UIO_OE_TT_PROJECT0
rlabel metal3 215149 151956 215149 151956 0 Tile_X5Y5_UIO_OE_TT_PROJECT1
rlabel metal3 215149 152460 215149 152460 0 Tile_X5Y5_UIO_OE_TT_PROJECT2
rlabel metal3 215149 152964 215149 152964 0 Tile_X5Y5_UIO_OE_TT_PROJECT3
rlabel metal3 215149 153468 215149 153468 0 Tile_X5Y5_UIO_OE_TT_PROJECT4
rlabel metal3 215149 153972 215149 153972 0 Tile_X5Y5_UIO_OE_TT_PROJECT5
rlabel metal3 215149 154476 215149 154476 0 Tile_X5Y5_UIO_OE_TT_PROJECT6
rlabel metal3 215149 154980 215149 154980 0 Tile_X5Y5_UIO_OE_TT_PROJECT7
rlabel metal3 215149 147420 215149 147420 0 Tile_X5Y5_UIO_OUT_TT_PROJECT0
rlabel metal3 215149 147924 215149 147924 0 Tile_X5Y5_UIO_OUT_TT_PROJECT1
rlabel metal3 215149 148428 215149 148428 0 Tile_X5Y5_UIO_OUT_TT_PROJECT2
rlabel metal3 215149 148932 215149 148932 0 Tile_X5Y5_UIO_OUT_TT_PROJECT3
rlabel metal3 215149 149436 215149 149436 0 Tile_X5Y5_UIO_OUT_TT_PROJECT4
rlabel metal3 215149 149940 215149 149940 0 Tile_X5Y5_UIO_OUT_TT_PROJECT5
rlabel metal3 215149 150444 215149 150444 0 Tile_X5Y5_UIO_OUT_TT_PROJECT6
rlabel metal3 215149 150948 215149 150948 0 Tile_X5Y5_UIO_OUT_TT_PROJECT7
rlabel metal3 215149 155484 215149 155484 0 Tile_X5Y5_UI_IN_TT_PROJECT0
rlabel metal3 215149 155988 215149 155988 0 Tile_X5Y5_UI_IN_TT_PROJECT1
rlabel metal3 215149 156492 215149 156492 0 Tile_X5Y5_UI_IN_TT_PROJECT2
rlabel metal3 215149 156996 215149 156996 0 Tile_X5Y5_UI_IN_TT_PROJECT3
rlabel metal3 215149 157500 215149 157500 0 Tile_X5Y5_UI_IN_TT_PROJECT4
rlabel metal3 215149 158004 215149 158004 0 Tile_X5Y5_UI_IN_TT_PROJECT5
rlabel metal3 215149 158508 215149 158508 0 Tile_X5Y5_UI_IN_TT_PROJECT6
rlabel metal3 215149 159012 215149 159012 0 Tile_X5Y5_UI_IN_TT_PROJECT7
rlabel metal3 215149 143388 215149 143388 0 Tile_X5Y5_UO_OUT_TT_PROJECT0
rlabel metal3 215149 143892 215149 143892 0 Tile_X5Y5_UO_OUT_TT_PROJECT1
rlabel metal3 215149 144396 215149 144396 0 Tile_X5Y5_UO_OUT_TT_PROJECT2
rlabel metal3 215149 144900 215149 144900 0 Tile_X5Y5_UO_OUT_TT_PROJECT3
rlabel metal3 215149 145404 215149 145404 0 Tile_X5Y5_UO_OUT_TT_PROJECT4
rlabel metal3 215149 145908 215149 145908 0 Tile_X5Y5_UO_OUT_TT_PROJECT5
rlabel metal3 215149 146412 215149 146412 0 Tile_X5Y5_UO_OUT_TT_PROJECT6
rlabel metal3 215149 146916 215149 146916 0 Tile_X5Y5_UO_OUT_TT_PROJECT7
rlabel metal3 215149 121044 215149 121044 0 Tile_X5Y6_CLK_TT_PROJECT
rlabel metal3 215149 120540 215149 120540 0 Tile_X5Y6_ENA_TT_PROJECT
rlabel metal3 215149 121548 215149 121548 0 Tile_X5Y6_RST_N_TT_PROJECT
rlabel metal3 215149 116508 215149 116508 0 Tile_X5Y6_UIO_IN_TT_PROJECT0
rlabel metal3 215149 117012 215149 117012 0 Tile_X5Y6_UIO_IN_TT_PROJECT1
rlabel metal3 215149 117516 215149 117516 0 Tile_X5Y6_UIO_IN_TT_PROJECT2
rlabel metal3 215149 118020 215149 118020 0 Tile_X5Y6_UIO_IN_TT_PROJECT3
rlabel metal3 215149 118524 215149 118524 0 Tile_X5Y6_UIO_IN_TT_PROJECT4
rlabel metal3 215149 119028 215149 119028 0 Tile_X5Y6_UIO_IN_TT_PROJECT5
rlabel metal3 215149 119532 215149 119532 0 Tile_X5Y6_UIO_IN_TT_PROJECT6
rlabel metal3 215149 120036 215149 120036 0 Tile_X5Y6_UIO_IN_TT_PROJECT7
rlabel metal3 215149 108444 215149 108444 0 Tile_X5Y6_UIO_OE_TT_PROJECT0
rlabel metal3 215149 108948 215149 108948 0 Tile_X5Y6_UIO_OE_TT_PROJECT1
rlabel metal3 215149 109452 215149 109452 0 Tile_X5Y6_UIO_OE_TT_PROJECT2
rlabel metal3 215149 109956 215149 109956 0 Tile_X5Y6_UIO_OE_TT_PROJECT3
rlabel metal3 215149 110460 215149 110460 0 Tile_X5Y6_UIO_OE_TT_PROJECT4
rlabel metal3 215149 110964 215149 110964 0 Tile_X5Y6_UIO_OE_TT_PROJECT5
rlabel metal3 215149 111468 215149 111468 0 Tile_X5Y6_UIO_OE_TT_PROJECT6
rlabel metal3 215149 111972 215149 111972 0 Tile_X5Y6_UIO_OE_TT_PROJECT7
rlabel metal3 215149 104412 215149 104412 0 Tile_X5Y6_UIO_OUT_TT_PROJECT0
rlabel metal3 215149 104916 215149 104916 0 Tile_X5Y6_UIO_OUT_TT_PROJECT1
rlabel metal3 215149 105420 215149 105420 0 Tile_X5Y6_UIO_OUT_TT_PROJECT2
rlabel metal3 215149 105924 215149 105924 0 Tile_X5Y6_UIO_OUT_TT_PROJECT3
rlabel metal3 215149 106428 215149 106428 0 Tile_X5Y6_UIO_OUT_TT_PROJECT4
rlabel metal3 215149 106932 215149 106932 0 Tile_X5Y6_UIO_OUT_TT_PROJECT5
rlabel metal3 215149 107436 215149 107436 0 Tile_X5Y6_UIO_OUT_TT_PROJECT6
rlabel metal3 215149 107940 215149 107940 0 Tile_X5Y6_UIO_OUT_TT_PROJECT7
rlabel metal3 215149 112476 215149 112476 0 Tile_X5Y6_UI_IN_TT_PROJECT0
rlabel metal3 215149 112980 215149 112980 0 Tile_X5Y6_UI_IN_TT_PROJECT1
rlabel metal3 215149 113484 215149 113484 0 Tile_X5Y6_UI_IN_TT_PROJECT2
rlabel metal3 215149 113988 215149 113988 0 Tile_X5Y6_UI_IN_TT_PROJECT3
rlabel metal3 215149 114492 215149 114492 0 Tile_X5Y6_UI_IN_TT_PROJECT4
rlabel metal3 215149 114996 215149 114996 0 Tile_X5Y6_UI_IN_TT_PROJECT5
rlabel metal3 215149 115500 215149 115500 0 Tile_X5Y6_UI_IN_TT_PROJECT6
rlabel metal3 215149 116004 215149 116004 0 Tile_X5Y6_UI_IN_TT_PROJECT7
rlabel metal3 215149 100380 215149 100380 0 Tile_X5Y6_UO_OUT_TT_PROJECT0
rlabel metal3 215149 100884 215149 100884 0 Tile_X5Y6_UO_OUT_TT_PROJECT1
rlabel metal3 215149 101388 215149 101388 0 Tile_X5Y6_UO_OUT_TT_PROJECT2
rlabel metal3 215149 101892 215149 101892 0 Tile_X5Y6_UO_OUT_TT_PROJECT3
rlabel metal3 215149 102396 215149 102396 0 Tile_X5Y6_UO_OUT_TT_PROJECT4
rlabel metal3 215149 102900 215149 102900 0 Tile_X5Y6_UO_OUT_TT_PROJECT5
rlabel metal3 215149 103404 215149 103404 0 Tile_X5Y6_UO_OUT_TT_PROJECT6
rlabel metal3 215149 103908 215149 103908 0 Tile_X5Y6_UO_OUT_TT_PROJECT7
rlabel metal3 215149 78036 215149 78036 0 Tile_X5Y7_CLK_TT_PROJECT
rlabel metal3 215149 77532 215149 77532 0 Tile_X5Y7_ENA_TT_PROJECT
rlabel metal3 215149 78540 215149 78540 0 Tile_X5Y7_RST_N_TT_PROJECT
rlabel metal3 215149 73500 215149 73500 0 Tile_X5Y7_UIO_IN_TT_PROJECT0
rlabel metal3 215149 74004 215149 74004 0 Tile_X5Y7_UIO_IN_TT_PROJECT1
rlabel metal3 215149 74508 215149 74508 0 Tile_X5Y7_UIO_IN_TT_PROJECT2
rlabel metal3 215149 75012 215149 75012 0 Tile_X5Y7_UIO_IN_TT_PROJECT3
rlabel metal3 215149 75516 215149 75516 0 Tile_X5Y7_UIO_IN_TT_PROJECT4
rlabel metal3 215149 76020 215149 76020 0 Tile_X5Y7_UIO_IN_TT_PROJECT5
rlabel metal3 215149 76524 215149 76524 0 Tile_X5Y7_UIO_IN_TT_PROJECT6
rlabel metal3 215149 77028 215149 77028 0 Tile_X5Y7_UIO_IN_TT_PROJECT7
rlabel metal3 215149 65436 215149 65436 0 Tile_X5Y7_UIO_OE_TT_PROJECT0
rlabel metal3 215149 65940 215149 65940 0 Tile_X5Y7_UIO_OE_TT_PROJECT1
rlabel metal3 215149 66444 215149 66444 0 Tile_X5Y7_UIO_OE_TT_PROJECT2
rlabel metal3 215149 66948 215149 66948 0 Tile_X5Y7_UIO_OE_TT_PROJECT3
rlabel metal3 215149 67452 215149 67452 0 Tile_X5Y7_UIO_OE_TT_PROJECT4
rlabel metal3 215149 67956 215149 67956 0 Tile_X5Y7_UIO_OE_TT_PROJECT5
rlabel metal3 215149 68460 215149 68460 0 Tile_X5Y7_UIO_OE_TT_PROJECT6
rlabel metal3 215149 68964 215149 68964 0 Tile_X5Y7_UIO_OE_TT_PROJECT7
rlabel metal3 215149 61404 215149 61404 0 Tile_X5Y7_UIO_OUT_TT_PROJECT0
rlabel metal3 215149 61908 215149 61908 0 Tile_X5Y7_UIO_OUT_TT_PROJECT1
rlabel metal3 215149 62412 215149 62412 0 Tile_X5Y7_UIO_OUT_TT_PROJECT2
rlabel metal3 215149 62916 215149 62916 0 Tile_X5Y7_UIO_OUT_TT_PROJECT3
rlabel metal3 215149 63420 215149 63420 0 Tile_X5Y7_UIO_OUT_TT_PROJECT4
rlabel metal3 215149 63924 215149 63924 0 Tile_X5Y7_UIO_OUT_TT_PROJECT5
rlabel metal3 215149 64428 215149 64428 0 Tile_X5Y7_UIO_OUT_TT_PROJECT6
rlabel metal3 215149 64932 215149 64932 0 Tile_X5Y7_UIO_OUT_TT_PROJECT7
rlabel metal3 215149 69468 215149 69468 0 Tile_X5Y7_UI_IN_TT_PROJECT0
rlabel metal3 215149 69972 215149 69972 0 Tile_X5Y7_UI_IN_TT_PROJECT1
rlabel metal3 215149 70476 215149 70476 0 Tile_X5Y7_UI_IN_TT_PROJECT2
rlabel metal3 215149 70980 215149 70980 0 Tile_X5Y7_UI_IN_TT_PROJECT3
rlabel metal3 215149 71484 215149 71484 0 Tile_X5Y7_UI_IN_TT_PROJECT4
rlabel metal3 215149 71988 215149 71988 0 Tile_X5Y7_UI_IN_TT_PROJECT5
rlabel metal3 215149 72492 215149 72492 0 Tile_X5Y7_UI_IN_TT_PROJECT6
rlabel metal3 215149 72996 215149 72996 0 Tile_X5Y7_UI_IN_TT_PROJECT7
rlabel metal3 215149 57372 215149 57372 0 Tile_X5Y7_UO_OUT_TT_PROJECT0
rlabel metal3 215149 57876 215149 57876 0 Tile_X5Y7_UO_OUT_TT_PROJECT1
rlabel metal3 215149 58380 215149 58380 0 Tile_X5Y7_UO_OUT_TT_PROJECT2
rlabel metal3 215149 58884 215149 58884 0 Tile_X5Y7_UO_OUT_TT_PROJECT3
rlabel metal3 215149 59388 215149 59388 0 Tile_X5Y7_UO_OUT_TT_PROJECT4
rlabel metal3 215149 59892 215149 59892 0 Tile_X5Y7_UO_OUT_TT_PROJECT5
rlabel metal3 215149 60396 215149 60396 0 Tile_X5Y7_UO_OUT_TT_PROJECT6
rlabel metal3 215149 60900 215149 60900 0 Tile_X5Y7_UO_OUT_TT_PROJECT7
rlabel metal3 215149 35028 215149 35028 0 Tile_X5Y8_CLK_TT_PROJECT
rlabel metal3 215149 34524 215149 34524 0 Tile_X5Y8_ENA_TT_PROJECT
rlabel metal3 215149 35532 215149 35532 0 Tile_X5Y8_RST_N_TT_PROJECT
rlabel metal3 215149 30492 215149 30492 0 Tile_X5Y8_UIO_IN_TT_PROJECT0
rlabel metal3 215149 30996 215149 30996 0 Tile_X5Y8_UIO_IN_TT_PROJECT1
rlabel metal3 215149 31500 215149 31500 0 Tile_X5Y8_UIO_IN_TT_PROJECT2
rlabel metal3 215149 32004 215149 32004 0 Tile_X5Y8_UIO_IN_TT_PROJECT3
rlabel metal3 215149 32508 215149 32508 0 Tile_X5Y8_UIO_IN_TT_PROJECT4
rlabel metal3 215149 33012 215149 33012 0 Tile_X5Y8_UIO_IN_TT_PROJECT5
rlabel metal3 215149 33516 215149 33516 0 Tile_X5Y8_UIO_IN_TT_PROJECT6
rlabel metal3 215149 34020 215149 34020 0 Tile_X5Y8_UIO_IN_TT_PROJECT7
rlabel metal3 215149 22428 215149 22428 0 Tile_X5Y8_UIO_OE_TT_PROJECT0
rlabel metal3 215149 22932 215149 22932 0 Tile_X5Y8_UIO_OE_TT_PROJECT1
rlabel metal3 215149 23436 215149 23436 0 Tile_X5Y8_UIO_OE_TT_PROJECT2
rlabel metal3 215149 23940 215149 23940 0 Tile_X5Y8_UIO_OE_TT_PROJECT3
rlabel metal3 215149 24444 215149 24444 0 Tile_X5Y8_UIO_OE_TT_PROJECT4
rlabel metal3 215149 24948 215149 24948 0 Tile_X5Y8_UIO_OE_TT_PROJECT5
rlabel metal3 215149 25452 215149 25452 0 Tile_X5Y8_UIO_OE_TT_PROJECT6
rlabel metal3 215149 25956 215149 25956 0 Tile_X5Y8_UIO_OE_TT_PROJECT7
rlabel metal3 215149 18396 215149 18396 0 Tile_X5Y8_UIO_OUT_TT_PROJECT0
rlabel metal3 215149 18900 215149 18900 0 Tile_X5Y8_UIO_OUT_TT_PROJECT1
rlabel metal3 215149 19404 215149 19404 0 Tile_X5Y8_UIO_OUT_TT_PROJECT2
rlabel metal3 215149 19908 215149 19908 0 Tile_X5Y8_UIO_OUT_TT_PROJECT3
rlabel metal3 215149 20412 215149 20412 0 Tile_X5Y8_UIO_OUT_TT_PROJECT4
rlabel metal3 215149 20916 215149 20916 0 Tile_X5Y8_UIO_OUT_TT_PROJECT5
rlabel metal3 215149 21420 215149 21420 0 Tile_X5Y8_UIO_OUT_TT_PROJECT6
rlabel metal3 215149 21924 215149 21924 0 Tile_X5Y8_UIO_OUT_TT_PROJECT7
rlabel metal3 215149 26460 215149 26460 0 Tile_X5Y8_UI_IN_TT_PROJECT0
rlabel metal3 215149 26964 215149 26964 0 Tile_X5Y8_UI_IN_TT_PROJECT1
rlabel metal3 215149 27468 215149 27468 0 Tile_X5Y8_UI_IN_TT_PROJECT2
rlabel metal3 215149 27972 215149 27972 0 Tile_X5Y8_UI_IN_TT_PROJECT3
rlabel metal3 215149 28476 215149 28476 0 Tile_X5Y8_UI_IN_TT_PROJECT4
rlabel metal3 215149 28980 215149 28980 0 Tile_X5Y8_UI_IN_TT_PROJECT5
rlabel metal3 215149 29484 215149 29484 0 Tile_X5Y8_UI_IN_TT_PROJECT6
rlabel metal3 215149 29988 215149 29988 0 Tile_X5Y8_UI_IN_TT_PROJECT7
rlabel metal3 215149 14364 215149 14364 0 Tile_X5Y8_UO_OUT_TT_PROJECT0
rlabel metal3 215149 14868 215149 14868 0 Tile_X5Y8_UO_OUT_TT_PROJECT1
rlabel metal3 215149 15372 215149 15372 0 Tile_X5Y8_UO_OUT_TT_PROJECT2
rlabel metal3 215149 15876 215149 15876 0 Tile_X5Y8_UO_OUT_TT_PROJECT3
rlabel metal3 215149 16380 215149 16380 0 Tile_X5Y8_UO_OUT_TT_PROJECT4
rlabel metal3 215149 16884 215149 16884 0 Tile_X5Y8_UO_OUT_TT_PROJECT5
rlabel metal3 215149 17388 215149 17388 0 Tile_X5Y8_UO_OUT_TT_PROJECT6
rlabel metal3 215149 17892 215149 17892 0 Tile_X5Y8_UO_OUT_TT_PROJECT7
rlabel metal2 1152 118 1152 118 0 UserCLK
<< properties >>
string FIXED_BBOX 0 0 215232 366504
<< end >>
