* NGSPICE file created from IHP_SRAM.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand4_1 abstract view
.subckt sg13g2_nand4_1 B C A Y VDD VSS D
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

.subckt IHP_SRAM ADDR_SRAM0 ADDR_SRAM1 ADDR_SRAM2 ADDR_SRAM3 ADDR_SRAM4 ADDR_SRAM5
+ ADDR_SRAM6 ADDR_SRAM7 ADDR_SRAM8 ADDR_SRAM9 BM_SRAM0 BM_SRAM1 BM_SRAM10 BM_SRAM11
+ BM_SRAM12 BM_SRAM13 BM_SRAM14 BM_SRAM15 BM_SRAM16 BM_SRAM17 BM_SRAM18 BM_SRAM19
+ BM_SRAM2 BM_SRAM20 BM_SRAM21 BM_SRAM22 BM_SRAM23 BM_SRAM24 BM_SRAM25 BM_SRAM26 BM_SRAM27
+ BM_SRAM28 BM_SRAM29 BM_SRAM3 BM_SRAM30 BM_SRAM31 BM_SRAM4 BM_SRAM5 BM_SRAM6 BM_SRAM7
+ BM_SRAM8 BM_SRAM9 CLK_SRAM CONFIGURED_top DIN_SRAM0 DIN_SRAM1 DIN_SRAM10 DIN_SRAM11
+ DIN_SRAM12 DIN_SRAM13 DIN_SRAM14 DIN_SRAM15 DIN_SRAM16 DIN_SRAM17 DIN_SRAM18 DIN_SRAM19
+ DIN_SRAM2 DIN_SRAM20 DIN_SRAM21 DIN_SRAM22 DIN_SRAM23 DIN_SRAM24 DIN_SRAM25 DIN_SRAM26
+ DIN_SRAM27 DIN_SRAM28 DIN_SRAM29 DIN_SRAM3 DIN_SRAM30 DIN_SRAM31 DIN_SRAM4 DIN_SRAM5
+ DIN_SRAM6 DIN_SRAM7 DIN_SRAM8 DIN_SRAM9 DOUT_SRAM0 DOUT_SRAM1 DOUT_SRAM10 DOUT_SRAM11
+ DOUT_SRAM12 DOUT_SRAM13 DOUT_SRAM14 DOUT_SRAM15 DOUT_SRAM16 DOUT_SRAM17 DOUT_SRAM18
+ DOUT_SRAM19 DOUT_SRAM2 DOUT_SRAM20 DOUT_SRAM21 DOUT_SRAM22 DOUT_SRAM23 DOUT_SRAM24
+ DOUT_SRAM25 DOUT_SRAM26 DOUT_SRAM27 DOUT_SRAM28 DOUT_SRAM29 DOUT_SRAM3 DOUT_SRAM30
+ DOUT_SRAM31 DOUT_SRAM4 DOUT_SRAM5 DOUT_SRAM6 DOUT_SRAM7 DOUT_SRAM8 DOUT_SRAM9 MEN_SRAM
+ REN_SRAM TIE_HIGH_SRAM TIE_LOW_SRAM Tile_X0Y0_E1END[0] Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E1END[3] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1] Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6] Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3] Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6END[0] Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11]
+ Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3] Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5]
+ Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8] Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11] Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13]
+ Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15] Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6]
+ Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8] Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0]
+ Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11] Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13]
+ Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15] Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17]
+ Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19] Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20]
+ Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22] Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24]
+ Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26] Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28]
+ Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2] Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31]
+ Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4] Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6]
+ Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8] Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0]
+ Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11] Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13]
+ Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15] Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17]
+ Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19] Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20]
+ Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22] Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24]
+ Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26] Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28]
+ Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2] Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31]
+ Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4] Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6]
+ Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8] Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0]
+ Tile_X0Y0_FrameStrobe_O[10] Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12]
+ Tile_X0Y0_FrameStrobe_O[13] Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15]
+ Tile_X0Y0_FrameStrobe_O[16] Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18]
+ Tile_X0Y0_FrameStrobe_O[19] Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2]
+ Tile_X0Y0_FrameStrobe_O[3] Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5]
+ Tile_X0Y0_FrameStrobe_O[6] Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8]
+ Tile_X0Y0_FrameStrobe_O[9] Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2]
+ Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0] Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3]
+ Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5] Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0]
+ Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2] Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4]
+ Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6] Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10]
+ Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12] Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14]
+ Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2] Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4]
+ Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7] Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9]
+ Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2] Tile_X0Y0_S1END[3] Tile_X0Y0_S2END[0]
+ Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3] Tile_X0Y0_S2END[4] Tile_X0Y0_S2END[5]
+ Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0] Tile_X0Y0_S2MID[1] Tile_X0Y0_S2MID[2]
+ Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5] Tile_X0Y0_S2MID[6] Tile_X0Y0_S2MID[7]
+ Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11] Tile_X0Y0_S4END[12] Tile_X0Y0_S4END[13]
+ Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15] Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2] Tile_X0Y0_S4END[3]
+ Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5] Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7] Tile_X0Y0_S4END[8]
+ Tile_X0Y0_S4END[9] Tile_X0Y0_UserCLKo Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2]
+ Tile_X0Y0_W1BEG[3] Tile_X0Y0_W2BEG[0] Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3]
+ Tile_X0Y0_W2BEG[4] Tile_X0Y0_W2BEG[5] Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0]
+ Tile_X0Y0_W2BEGb[1] Tile_X0Y0_W2BEGb[2] Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4]
+ Tile_X0Y0_W2BEGb[5] Tile_X0Y0_W2BEGb[6] Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10]
+ Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1] Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4]
+ Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6] Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9]
+ Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10] Tile_X0Y0_WW4BEG[11] Tile_X0Y0_WW4BEG[12]
+ Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14] Tile_X0Y0_WW4BEG[15] Tile_X0Y0_WW4BEG[1]
+ Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3] Tile_X0Y0_WW4BEG[4] Tile_X0Y0_WW4BEG[5]
+ Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7] Tile_X0Y0_WW4BEG[8] Tile_X0Y0_WW4BEG[9]
+ Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2] Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[0]
+ Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3] Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5]
+ Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0] Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2]
+ Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5] Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7]
+ Tile_X0Y1_E6END[0] Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2]
+ Tile_X0Y1_E6END[3] Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5] Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7]
+ Tile_X0Y1_E6END[8] Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[0] Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15]
+ Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2] Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11]
+ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15]
+ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19]
+ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22]
+ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26]
+ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2]
+ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4]
+ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8]
+ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0] Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11]
+ Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13] Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15]
+ Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17] Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19]
+ Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20] Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22]
+ Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24] Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26]
+ Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28] Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2]
+ Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31] Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4]
+ Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6] Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8]
+ Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11]
+ Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13] Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15]
+ Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17] Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19]
+ Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4]
+ Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8]
+ Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0] Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1] Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3]
+ Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6] Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3] Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0] Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11]
+ Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13] Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15]
+ Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3] Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5]
+ Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8] Tile_X0Y1_N4END[9] Tile_X0Y1_S1BEG[0]
+ Tile_X0Y1_S1BEG[1] Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3] Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1]
+ Tile_X0Y1_S2BEG[2] Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4] Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6]
+ Tile_X0Y1_S2BEG[7] Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1] Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3]
+ Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5] Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7]
+ Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11] Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13]
+ Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15] Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3]
+ Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5] Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8]
+ Tile_X0Y1_S4BEG[9] Tile_X0Y1_UserCLK Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2]
+ Tile_X0Y1_W1BEG[3] Tile_X0Y1_W2BEG[0] Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3]
+ Tile_X0Y1_W2BEG[4] Tile_X0Y1_W2BEG[5] Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0]
+ Tile_X0Y1_W2BEGb[1] Tile_X0Y1_W2BEGb[2] Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4]
+ Tile_X0Y1_W2BEGb[5] Tile_X0Y1_W2BEGb[6] Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10]
+ Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1] Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4]
+ Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6] Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9]
+ Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10] Tile_X0Y1_WW4BEG[11] Tile_X0Y1_WW4BEG[12]
+ Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14] Tile_X0Y1_WW4BEG[15] Tile_X0Y1_WW4BEG[1]
+ Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3] Tile_X0Y1_WW4BEG[4] Tile_X0Y1_WW4BEG[5]
+ Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7] Tile_X0Y1_WW4BEG[8] Tile_X0Y1_WW4BEG[9]
+ VGND VPWR WEN_SRAM
XFILLER_100_138 VPWR VGND sg13g2_fill_1
XFILLER_100_127 VPWR VGND sg13g2_decap_8
X_0367_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_E6END[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13
+ _0059_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1
+ VPWR VGND sg13g2_mux4_1
X_0298_ VPWR _0001_ Tile_X0Y1_E2END[5] VGND sg13g2_inv_1
XFILLER_22_144 VPWR VGND sg13g2_decap_4
XFILLER_22_199 VPWR VGND sg13g2_fill_1
XFILLER_89_177 VPWR VGND sg13g2_fill_2
XFILLER_26_74 VPWR VGND sg13g2_fill_1
XFILLER_13_199 VPWR VGND sg13g2_fill_1
XFILLER_9_115 VPWR VGND sg13g2_fill_2
XFILLER_3_67 VPWR VGND sg13g2_fill_1
X_1270_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0985_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1606_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11 Tile_X0Y0_WW4BEG[11]
+ VPWR VGND sg13g2_buf_1
X_1537_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7 Tile_X0Y0_N2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_0419_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E2MID[0] Tile_X0Y0_E2END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7
+ VPWR VGND sg13g2_mux4_1
X_1399_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1468_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_12_21 VPWR VGND sg13g2_fill_2
XFILLER_10_136 VPWR VGND sg13g2_decap_4
XFILLER_92_106 VPWR VGND sg13g2_decap_4
X_0770_ VGND VPWR _0026_ _0210_ _0211_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q
+ sg13g2_a21oi_1
X_1322_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1253_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1184_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0968_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0899_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_147 VPWR VGND sg13g2_decap_4
XFILLER_2_143 VPWR VGND sg13g2_fill_1
X_0822_ _0258_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q VPWR VGND
+ sg13g2_nand2b_1
X_0684_ _0162_ VPWR ADDR_SRAM0 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
+ _0164_ sg13g2_o21ai_1
X_0753_ VGND VPWR _0022_ _0194_ _0196_ _0195_ sg13g2_a21oi_1
X_1305_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1236_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_128 VPWR VGND sg13g2_fill_2
X_1098_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_109 VPWR VGND sg13g2_fill_1
X_1167_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_29 VPWR VGND sg13g2_fill_1
XFILLER_69_49 VPWR VGND sg13g2_decap_8
XFILLER_85_37 VPWR VGND sg13g2_decap_8
XFILLER_47_117 VPWR VGND sg13g2_fill_2
XFILLER_34_74 VPWR VGND sg13g2_fill_2
XFILLER_59_71 VPWR VGND sg13g2_decap_8
XFILLER_75_92 VPWR VGND sg13g2_fill_1
X_1021_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_46_161 VPWR VGND sg13g2_fill_2
XFILLER_61_175 VPWR VGND sg13g2_fill_2
X_0805_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q VPWR
+ _0243_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
X_0598_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q VPWR
+ _0153_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
X_0667_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0088_ Tile_X0Y0_S4END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
+ _0161_ VPWR VGND sg13g2_mux4_1
X_0736_ Tile_X0Y1_E1END[0] Tile_X0Y1_EE4END[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ _0180_ VPWR VGND sg13g2_mux2_1
XFILLER_29_139 VPWR VGND sg13g2_fill_2
X_1219_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_194 VPWR VGND sg13g2_decap_4
XFILLER_52_131 VPWR VGND sg13g2_fill_2
XFILLER_52_175 VPWR VGND sg13g2_fill_2
XFILLER_29_74 VPWR VGND sg13g2_fill_1
XFILLER_61_72 VPWR VGND sg13g2_decap_4
XANTENNA_5 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
X_0521_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[12] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q BM_SRAM28
+ VPWR VGND sg13g2_mux4_1
X_0452_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q DOUT_SRAM16
+ DOUT_SRAM28 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0
+ VPWR VGND sg13g2_mux4_1
XFILLER_6_78 VPWR VGND sg13g2_fill_2
X_1570_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3 Tile_X0Y0_W2BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_20_4 VPWR VGND sg13g2_decap_8
X_0383_ _0076_ _0074_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_96_0 VPWR VGND sg13g2_fill_2
X_1004_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_120 VPWR VGND sg13g2_decap_4
X_1699_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 Tile_X0Y1_W6BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0719_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y1_EE4END[2]
+ Tile_X0Y1_EE4END[10] Tile_X0Y1_E6END[2] _0159_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
+ BM_SRAM2 VPWR VGND sg13g2_mux4_1
XFILLER_56_83 VPWR VGND sg13g2_fill_1
XFILLER_72_93 VPWR VGND sg13g2_decap_8
XFILLER_16_120 VPWR VGND sg13g2_decap_4
XFILLER_56_94 VPWR VGND sg13g2_decap_8
X_1622_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameData_O[11] VPWR VGND sg13g2_buf_1
X_0504_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y0_EE4END[3]
+ Tile_X0Y0_EE4END[11] Tile_X0Y0_E6END[11] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q DIN_SRAM27
+ VPWR VGND sg13g2_mux4_1
XFILLER_98_145 VPWR VGND sg13g2_fill_1
X_1484_ Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData_O[10] VPWR VGND sg13g2_buf_1
X_0435_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ DOUT_SRAM17 Tile_X0Y0_S1END[3] DOUT_SRAM20 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 VPWR VGND sg13g2_mux4_1
X_1553_ Tile_X0Y1_N4END[15] Tile_X0Y0_N4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_0297_ VPWR _0000_ Tile_X0Y1_E2MID[3] VGND sg13g2_inv_1
X_0366_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_mux4_1
XFILLER_13_178 VPWR VGND sg13g2_decap_4
X_0984_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1536_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6 Tile_X0Y0_N2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1605_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10 Tile_X0Y0_WW4BEG[10]
+ VPWR VGND sg13g2_buf_1
XFILLER_59_0 VPWR VGND sg13g2_fill_2
X_0418_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q Tile_X0Y0_E2MID[1]
+ Tile_X0Y0_E2END[1] Tile_X0Y0_E6END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6
+ VPWR VGND sg13g2_mux4_1
XFILLER_86_159 VPWR VGND sg13g2_fill_2
X_1398_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1467_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0349_ _0048_ VPWR _0049_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y1_E2END[3] sg13g2_o21ai_1
XFILLER_103_58 VPWR VGND sg13g2_fill_1
XFILLER_52_7 VPWR VGND sg13g2_fill_1
XFILLER_68_115 VPWR VGND sg13g2_decap_8
X_1321_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1252_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1183_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0967_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1519_ Tile_X0Y1_FrameStrobe[13] Tile_X0Y0_FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
X_0898_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_126 VPWR VGND sg13g2_decap_4
XFILLER_48_95 VPWR VGND sg13g2_fill_2
XFILLER_73_140 VPWR VGND sg13g2_decap_4
X_0752_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q VPWR
+ _0195_ VGND _0192_ _0193_ sg13g2_o21ai_1
X_0821_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0257_ VPWR VGND sg13g2_nor2b_1
X_0683_ VGND VPWR Tile_X0Y1_E2END[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ _0164_ _0163_ sg13g2_a21oi_1
X_1304_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1235_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1166_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1097_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_173 VPWR VGND sg13g2_fill_1
XFILLER_64_195 VPWR VGND sg13g2_decap_4
XFILLER_59_50 VPWR VGND sg13g2_decap_8
X_1020_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_198 VPWR VGND sg13g2_fill_2
X_0735_ _0178_ VPWR _0179_ VGND _0019_ _0161_ sg13g2_o21ai_1
X_0804_ _0031_ _0083_ _0242_ VPWR VGND sg13g2_nor2_1
X_0597_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ _0152_ VPWR VGND sg13g2_nor2b_1
X_0666_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q DOUT_SRAM2
+ DOUT_SRAM14 _0160_ _0078_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 VPWR VGND sg13g2_mux4_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_1149_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_151 VPWR VGND sg13g2_fill_2
X_1218_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_101 VPWR VGND sg13g2_fill_2
XFILLER_20_11 VPWR VGND sg13g2_fill_2
XFILLER_20_44 VPWR VGND sg13g2_fill_1
XFILLER_20_66 VPWR VGND sg13g2_decap_4
XFILLER_43_121 VPWR VGND sg13g2_fill_1
XANTENNA_6 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
X_0520_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y0_EE4END[3]
+ Tile_X0Y0_EE4END[11] Tile_X0Y0_E6END[11] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q BM_SRAM27
+ VPWR VGND sg13g2_mux4_1
X_0451_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q DOUT_SRAM23
+ DOUT_SRAM31 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7
+ VPWR VGND sg13g2_mux4_1
X_0382_ Tile_X0Y1_N1END[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q _0075_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_86_70 VPWR VGND sg13g2_decap_8
X_1003_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_89_0 VPWR VGND sg13g2_decap_4
XFILLER_34_187 VPWR VGND sg13g2_decap_8
XFILLER_34_198 VPWR VGND sg13g2_fill_2
X_1698_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 Tile_X0Y1_W2BEGb[7]
+ VPWR VGND sg13g2_buf_1
X_0718_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y1_EE4END[1]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_E6END[1] _0160_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
+ BM_SRAM1 VPWR VGND sg13g2_mux4_1
X_0649_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0060_ Tile_X0Y0_S4END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 VPWR VGND sg13g2_mux4_1
XFILLER_15_33 VPWR VGND sg13g2_fill_2
X_1552_ Tile_X0Y1_N4END[14] Tile_X0Y0_N4BEG[6] VPWR VGND sg13g2_buf_1
X_1621_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData_O[10] VPWR VGND sg13g2_buf_1
X_0503_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[10] Tile_X0Y0_E6END[10] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q DIN_SRAM26
+ VPWR VGND sg13g2_mux4_1
X_1483_ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[9] VPWR VGND sg13g2_buf_1
X_0365_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 Tile_X0Y1_E6END[5]
+ _0063_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ VPWR VGND sg13g2_mux4_1
X_0434_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ DOUT_SRAM16 Tile_X0Y0_S1END[2] DOUT_SRAM21 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 VPWR VGND sg13g2_mux4_1
XFILLER_22_113 VPWR VGND sg13g2_decap_8
XFILLER_77_17 VPWR VGND sg13g2_fill_1
XFILLER_67_83 VPWR VGND sg13g2_fill_1
XFILLER_83_71 VPWR VGND sg13g2_fill_2
X_0983_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1535_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5 Tile_X0Y0_N2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_1604_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9 Tile_X0Y0_WW4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_0417_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6
+ Tile_X0Y0_S2MID[6] Tile_X0Y1_N2MID[6] Tile_X0Y0_S2END[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_94_171 VPWR VGND sg13g2_decap_8
X_1397_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1466_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0348_ _0048_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0002_ VPWR VGND sg13g2_nand2_1
XFILLER_12_67 VPWR VGND sg13g2_decap_8
XFILLER_12_45 VPWR VGND sg13g2_fill_1
XFILLER_12_23 VPWR VGND sg13g2_fill_1
XFILLER_77_116 VPWR VGND sg13g2_fill_2
XFILLER_37_31 VPWR VGND sg13g2_fill_1
X_1320_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1182_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1251_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_91_174 VPWR VGND sg13g2_fill_2
XFILLER_91_163 VPWR VGND sg13g2_decap_8
X_0897_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_0 VPWR VGND sg13g2_fill_2
X_0966_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1518_ Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
X_1449_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_141 VPWR VGND sg13g2_fill_1
XFILLER_82_130 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_fill_2
XFILLER_23_66 VPWR VGND sg13g2_decap_8
XFILLER_23_99 VPWR VGND sg13g2_fill_2
XFILLER_80_72 VPWR VGND sg13g2_decap_8
X_0820_ VGND VPWR _0249_ _0251_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3
+ _0256_ sg13g2_a21oi_1
X_0751_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q _0194_ VPWR
+ VGND sg13g2_mux2_1
X_1303_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0682_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q Tile_X0Y1_E2MID[0]
+ _0163_ VPWR VGND sg13g2_nor2b_1
X_1096_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1165_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1234_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_108 VPWR VGND sg13g2_fill_1
X_0949_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_166 VPWR VGND sg13g2_decap_4
XFILLER_34_54 VPWR VGND sg13g2_fill_1
XFILLER_55_141 VPWR VGND sg13g2_fill_2
X_0665_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0060_ Tile_X0Y0_S4END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
+ _0160_ VPWR VGND sg13g2_mux4_1
X_0734_ VPWR _0178_ _0177_ VGND sg13g2_inv_1
X_0803_ VGND VPWR _0032_ _0240_ _0241_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
+ sg13g2_a21oi_1
X_0596_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q _0151_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_34_0 VPWR VGND sg13g2_decap_8
X_1148_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1079_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1217_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_199 VPWR VGND sg13g2_fill_1
XFILLER_106_179 VPWR VGND sg13g2_fill_1
XFILLER_43_177 VPWR VGND sg13g2_fill_2
XFILLER_45_86 VPWR VGND sg13g2_fill_2
XANTENNA_7 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
X_0381_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E6END[11] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15
+ _0073_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q _0074_
+ VPWR VGND sg13g2_mux4_1
X_0450_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q DOUT_SRAM22
+ DOUT_SRAM30 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6
+ VPWR VGND sg13g2_mux4_1
XFILLER_86_93 VPWR VGND sg13g2_decap_8
X_1002_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_174 VPWR VGND sg13g2_fill_2
XFILLER_96_2 VPWR VGND sg13g2_fill_1
X_1697_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 Tile_X0Y1_W2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_0648_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q DOUT_SRAM5
+ DOUT_SRAM9 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 _0079_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5
+ VPWR VGND sg13g2_mux4_1
X_0717_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_EE4END[8] Tile_X0Y1_E6END[0] _0161_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
+ BM_SRAM0 VPWR VGND sg13g2_mux4_1
X_0579_ _0134_ _0136_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0
+ VPWR VGND sg13g2_nor2_1
XFILLER_25_177 VPWR VGND sg13g2_fill_2
XFILLER_40_114 VPWR VGND sg13g2_decap_4
X_1482_ Tile_X0Y0_FrameData[8] Tile_X0Y0_FrameData_O[8] VPWR VGND sg13g2_buf_1
X_1551_ Tile_X0Y1_N4END[13] Tile_X0Y0_N4BEG[5] VPWR VGND sg13g2_buf_1
X_1620_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[9] VPWR VGND sg13g2_buf_1
X_0502_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y0_EE4END[1]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_E6END[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q DIN_SRAM25
+ VPWR VGND sg13g2_mux4_1
XFILLER_97_70 VPWR VGND sg13g2_decap_8
X_0364_ VPWR VGND _0061_ _0062_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
+ _0009_ _0063_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a221oi_1
X_0433_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ DOUT_SRAM19 Tile_X0Y0_S1END[1] DOUT_SRAM22 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_22_169 VPWR VGND sg13g2_fill_2
XFILLER_89_114 VPWR VGND sg13g2_fill_2
XFILLER_13_114 VPWR VGND sg13g2_fill_2
XFILLER_95_106 VPWR VGND sg13g2_fill_2
X_0982_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1534_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4 Tile_X0Y0_N2BEG[4]
+ VPWR VGND sg13g2_buf_1
X_1603_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8 Tile_X0Y0_WW4BEG[8]
+ VPWR VGND sg13g2_buf_1
X_1465_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_2 VPWR VGND sg13g2_fill_1
XFILLER_103_38 VPWR VGND sg13g2_fill_1
X_1396_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0416_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q Tile_X0Y1_E2MID[1]
+ Tile_X0Y1_E6END[1] Tile_X0Y1_E2END[1] _0083_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 VPWR VGND sg13g2_mux4_1
X_0347_ _0044_ _0046_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0047_ VPWR VGND sg13g2_nand3_1
XFILLER_78_94 VPWR VGND sg13g2_fill_2
XFILLER_78_83 VPWR VGND sg13g2_decap_8
XFILLER_38_7 VPWR VGND sg13g2_decap_4
XFILLER_68_139 VPWR VGND sg13g2_fill_2
X_1181_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1250_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_91_197 VPWR VGND sg13g2_fill_2
X_0896_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0965_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_0 VPWR VGND sg13g2_decap_8
X_1517_ Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
X_1448_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1379_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_38 VPWR VGND sg13g2_fill_1
XFILLER_23_34 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_fill_2
XFILLER_73_197 VPWR VGND sg13g2_fill_2
XFILLER_73_175 VPWR VGND sg13g2_fill_1
XFILLER_9_25 VPWR VGND sg13g2_fill_2
X_0681_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q _0043_
+ _0162_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ sg13g2_nand3b_1
X_0750_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q VPWR
+ _0193_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
X_1302_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1233_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1095_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1164_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_39 VPWR VGND sg13g2_fill_1
X_0948_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_109_59 VPWR VGND sg13g2_fill_2
X_0879_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_55_164 VPWR VGND sg13g2_fill_2
XFILLER_55_197 VPWR VGND sg13g2_fill_2
XFILLER_109_199 VPWR VGND sg13g2_fill_1
XFILLER_75_51 VPWR VGND sg13g2_fill_1
XFILLER_46_197 VPWR VGND sg13g2_fill_2
XFILLER_98_6 VPWR VGND sg13g2_decap_4
XFILLER_91_72 VPWR VGND sg13g2_decap_4
XFILLER_91_50 VPWR VGND sg13g2_fill_1
X_0802_ Tile_X0Y1_E1END[2] Tile_X0Y1_EE4END[14] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ _0240_ VPWR VGND sg13g2_mux2_1
X_0664_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q DOUT_SRAM1
+ DOUT_SRAM13 _0159_ _0079_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 VPWR VGND sg13g2_mux4_1
X_0733_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q VPWR
+ _0177_ VGND Tile_X0Y1_E6END[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ sg13g2_o21ai_1
X_0595_ _0148_ _0150_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2
+ VPWR VGND sg13g2_nor2_1
X_1216_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_29_109 VPWR VGND sg13g2_fill_1
X_1147_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_153 VPWR VGND sg13g2_fill_1
X_1078_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_103 VPWR VGND sg13g2_fill_1
XFILLER_20_13 VPWR VGND sg13g2_fill_1
XFILLER_20_35 VPWR VGND sg13g2_decap_8
XFILLER_45_65 VPWR VGND sg13g2_decap_8
XANTENNA_8 VPWR VGND Tile_X0Y0_S2MID[4] sg13g2_antennanp
X_0380_ VPWR VGND _0071_ _0072_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ _0005_ _0073_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a221oi_1
X_1001_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0578_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q _0135_
+ _0136_ VPWR VGND sg13g2_nor2_1
X_1696_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 Tile_X0Y1_W2BEGb[5]
+ VPWR VGND sg13g2_buf_1
X_0647_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0067_ Tile_X0Y0_S4END[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 VPWR VGND sg13g2_mux4_1
X_0716_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[15] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q DIN_SRAM15
+ VPWR VGND sg13g2_mux4_1
XFILLER_15_57 VPWR VGND sg13g2_fill_1
XFILLER_15_35 VPWR VGND sg13g2_fill_1
XFILLER_31_89 VPWR VGND sg13g2_fill_2
XFILLER_16_178 VPWR VGND sg13g2_decap_4
XFILLER_56_53 VPWR VGND sg13g2_fill_1
XFILLER_31_137 VPWR VGND sg13g2_fill_2
XFILLER_98_159 VPWR VGND sg13g2_fill_1
X_0501_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[8] Tile_X0Y0_E6END[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q DIN_SRAM24
+ VPWR VGND sg13g2_mux4_1
X_0432_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ DOUT_SRAM18 Tile_X0Y0_S1END[0] DOUT_SRAM23 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
X_1481_ Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData_O[7] VPWR VGND sg13g2_buf_1
X_1550_ Tile_X0Y1_N4END[12] Tile_X0Y0_N4BEG[4] VPWR VGND sg13g2_buf_1
X_0363_ Tile_X0Y1_N1END[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q _0062_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_94_0 VPWR VGND sg13g2_decap_4
X_1679_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 Tile_X0Y1_W1BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_26_67 VPWR VGND sg13g2_decap_8
XFILLER_88_170 VPWR VGND sg13g2_fill_2
X_0981_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1602_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7 Tile_X0Y0_WW4BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1533_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3 Tile_X0Y0_N2BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1395_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0415_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q Tile_X0Y1_N2MID[6]
+ Tile_X0Y1_N2END[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6
+ Tile_X0Y0_S2MID[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
+ _0083_ VPWR VGND sg13g2_mux4_1
X_1464_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0346_ _0046_ _0045_ Tile_X0Y1_E2END[4] Tile_X0Y0_S2MID[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_37_22 VPWR VGND sg13g2_decap_8
XFILLER_5_199 VPWR VGND sg13g2_fill_1
XFILLER_5_177 VPWR VGND sg13g2_fill_1
X_1180_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_2 VPWR VGND sg13g2_fill_1
X_0964_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1516_ Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
X_0895_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_57_0 VPWR VGND sg13g2_decap_4
X_1378_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1447_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0329_ VPWR _0032_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ VGND sg13g2_inv_1
XFILLER_82_198 VPWR VGND sg13g2_fill_2
XFILLER_64_53 VPWR VGND sg13g2_decap_4
X_0680_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q DOUT_SRAM3
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 _0161_ _0084_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11
+ VPWR VGND sg13g2_mux4_1
XFILLER_50_7 VPWR VGND sg13g2_decap_8
X_1301_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1232_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1094_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1163_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0947_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0878_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_102 VPWR VGND sg13g2_fill_2
XFILLER_55_154 VPWR VGND sg13g2_fill_1
XFILLER_55_187 VPWR VGND sg13g2_fill_2
XFILLER_109_112 VPWR VGND sg13g2_fill_2
XFILLER_59_64 VPWR VGND sg13g2_decap_8
XFILLER_61_146 VPWR VGND sg13g2_fill_1
XFILLER_61_168 VPWR VGND sg13g2_decap_8
XFILLER_91_95 VPWR VGND sg13g2_decap_8
X_0801_ _0238_ VPWR _0239_ VGND _0031_ _0159_ sg13g2_o21ai_1
X_0594_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q _0149_
+ _0150_ VPWR VGND sg13g2_nor2_1
X_0663_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0067_ Tile_X0Y0_S4END[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0159_ VPWR VGND sg13g2_mux4_1
X_0732_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[15] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q BM_SRAM15
+ VPWR VGND sg13g2_mux4_1
X_1146_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1215_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_198 VPWR VGND sg13g2_fill_2
XFILLER_52_102 VPWR VGND sg13g2_decap_4
XFILLER_52_124 VPWR VGND sg13g2_fill_2
X_1077_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_9 VPWR VGND Tile_X0Y0_S2MID[4] sg13g2_antennanp
XFILLER_10_91 VPWR VGND sg13g2_decap_8
X_1000_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_198 VPWR VGND sg13g2_fill_2
XFILLER_34_124 VPWR VGND sg13g2_fill_2
X_0715_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[14] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q DIN_SRAM14
+ VPWR VGND sg13g2_mux4_1
XFILLER_106_17 VPWR VGND sg13g2_fill_2
X_0577_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_E6END[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q _0135_ VPWR
+ VGND sg13g2_mux4_1
X_0646_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q DOUT_SRAM4
+ DOUT_SRAM8 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 _0080_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4
+ VPWR VGND sg13g2_mux4_1
X_1695_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 Tile_X0Y1_W2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_1129_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_32 VPWR VGND sg13g2_decap_8
XFILLER_72_53 VPWR VGND sg13g2_fill_2
XFILLER_56_76 VPWR VGND sg13g2_decap_8
XFILLER_56_87 VPWR VGND sg13g2_decap_8
XFILLER_98_127 VPWR VGND sg13g2_fill_1
X_0500_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y0_EE4END[7]
+ Tile_X0Y0_EE4END[15] Tile_X0Y0_E6END[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q DIN_SRAM23
+ VPWR VGND sg13g2_mux4_1
X_1480_ Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData_O[6] VPWR VGND sg13g2_buf_1
X_0431_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 Tile_X0Y1_E6END[4]
+ _0091_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ VPWR VGND sg13g2_mux4_1
X_0362_ _0061_ _0060_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_87_0 VPWR VGND sg13g2_decap_8
X_1678_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3 Tile_X0Y1_S4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_0629_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q DOUT_SRAM4
+ DOUT_SRAM12 _0080_ _0081_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 VPWR VGND sg13g2_mux4_1
XFILLER_13_149 VPWR VGND sg13g2_fill_1
XFILLER_13_116 VPWR VGND sg13g2_fill_1
XFILLER_26_24 VPWR VGND sg13g2_decap_4
XFILLER_42_67 VPWR VGND sg13g2_fill_1
XFILLER_95_108 VPWR VGND sg13g2_fill_1
XFILLER_3_28 VPWR VGND sg13g2_fill_1
X_0980_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_120 VPWR VGND sg13g2_fill_1
X_1532_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2 Tile_X0Y0_N2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1601_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6 Tile_X0Y0_WW4BEG[6]
+ VPWR VGND sg13g2_buf_1
X_0414_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6
+ VPWR VGND sg13g2_mux4_1
XFILLER_79_193 VPWR VGND sg13g2_fill_2
X_1394_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0345_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0045_ VPWR VGND sg13g2_nor2_1
X_1463_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_85_196 VPWR VGND sg13g2_decap_4
XFILLER_85_163 VPWR VGND sg13g2_decap_4
XFILLER_85_130 VPWR VGND sg13g2_decap_4
XFILLER_53_66 VPWR VGND sg13g2_fill_2
XFILLER_78_41 VPWR VGND sg13g2_decap_8
XFILLER_68_108 VPWR VGND sg13g2_decap_8
XFILLER_91_199 VPWR VGND sg13g2_fill_1
X_0894_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0963_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1515_ Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
XFILLER_59_119 VPWR VGND sg13g2_decap_8
X_1377_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1446_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0328_ VPWR _0031_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ VGND sg13g2_inv_1
XFILLER_82_166 VPWR VGND sg13g2_decap_8
XFILLER_73_199 VPWR VGND sg13g2_fill_1
XFILLER_73_144 VPWR VGND sg13g2_fill_1
XFILLER_73_133 VPWR VGND sg13g2_decap_8
XFILLER_80_97 VPWR VGND sg13g2_decap_4
XFILLER_80_53 VPWR VGND sg13g2_fill_2
XFILLER_43_7 VPWR VGND sg13g2_fill_2
X_1300_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1162_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1231_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1093_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_166 VPWR VGND sg13g2_decap_8
XFILLER_64_199 VPWR VGND sg13g2_fill_1
X_0877_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0946_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1429_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_199 VPWR VGND sg13g2_fill_1
XFILLER_46_199 VPWR VGND sg13g2_fill_1
X_0800_ VPWR _0238_ _0237_ VGND sg13g2_inv_1
X_0731_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_EE4END[6] Tile_X0Y1_EE4END[14] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q BM_SRAM14
+ VPWR VGND sg13g2_mux4_1
X_0593_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E6END[6] Tile_X0Y0_EE4END[14] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q _0149_ VPWR
+ VGND sg13g2_mux4_1
X_0662_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q DOUT_SRAM0
+ DOUT_SRAM12 _0158_ _0080_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 VPWR VGND sg13g2_mux4_1
X_1145_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1214_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1076_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0929_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_24 VPWR VGND sg13g2_fill_2
XFILLER_19_100 VPWR VGND sg13g2_fill_2
XFILLER_42_191 VPWR VGND sg13g2_decap_8
X_0645_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0074_ Tile_X0Y0_S4END[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 VPWR VGND sg13g2_mux4_1
X_1694_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 Tile_X0Y1_W2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_0714_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[13] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q DIN_SRAM13
+ VPWR VGND sg13g2_mux4_1
X_0576_ VGND VPWR _0015_ _0130_ _0134_ _0133_ sg13g2_a21oi_1
X_1128_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_15_15 VPWR VGND sg13g2_fill_1
X_1059_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_40_139 VPWR VGND sg13g2_fill_1
XFILLER_72_32 VPWR VGND sg13g2_decap_4
XFILLER_31_139 VPWR VGND sg13g2_fill_1
XFILLER_97_84 VPWR VGND sg13g2_decap_4
X_0361_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13
+ _0059_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q _0060_
+ VPWR VGND sg13g2_mux4_1
X_0430_ VPWR VGND _0090_ _0089_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
+ _0010_ _0091_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_a221oi_1
XFILLER_22_106 VPWR VGND sg13g2_decap_8
X_1677_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2 Tile_X0Y1_S4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_0628_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q DOUT_SRAM3
+ DOUT_SRAM11 _0080_ _0081_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 VPWR VGND sg13g2_mux4_1
X_0559_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q VPWR
+ _0119_ VGND _0117_ _0118_ sg13g2_o21ai_1
XFILLER_42_24 VPWR VGND sg13g2_decap_8
XFILLER_21_150 VPWR VGND sg13g2_fill_1
XFILLER_88_194 VPWR VGND sg13g2_decap_4
XFILLER_88_172 VPWR VGND sg13g2_fill_1
X_1531_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1 Tile_X0Y0_N2BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_8_198 VPWR VGND sg13g2_fill_2
X_1462_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1600_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5 Tile_X0Y0_WW4BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0413_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q Tile_X0Y0_E2MID[2]
+ Tile_X0Y0_E2END[2] Tile_X0Y0_E6END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5
+ VPWR VGND sg13g2_mux4_1
X_1393_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0344_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q VPWR
+ _0044_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 sg13g2_o21ai_1
XFILLER_5_135 VPWR VGND sg13g2_fill_1
XFILLER_76_164 VPWR VGND sg13g2_fill_2
XFILLER_91_123 VPWR VGND sg13g2_fill_2
X_0893_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0962_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1514_ Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_1445_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_197 VPWR VGND sg13g2_fill_2
XFILLER_67_164 VPWR VGND sg13g2_fill_2
X_1376_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0327_ VPWR _0030_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ VGND sg13g2_inv_1
XFILLER_58_131 VPWR VGND sg13g2_decap_8
XFILLER_58_175 VPWR VGND sg13g2_fill_1
XFILLER_58_197 VPWR VGND sg13g2_fill_2
XFILLER_36_7 VPWR VGND sg13g2_decap_8
X_1092_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1161_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_186 VPWR VGND sg13g2_fill_2
XFILLER_49_197 VPWR VGND sg13g2_fill_2
X_1230_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0876_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0945_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_62_0 VPWR VGND sg13g2_fill_2
X_1428_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_159 VPWR VGND sg13g2_decap_8
X_1359_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_48 VPWR VGND sg13g2_fill_2
XFILLER_109_158 VPWR VGND sg13g2_fill_1
XFILLER_46_123 VPWR VGND sg13g2_decap_4
XFILLER_61_115 VPWR VGND sg13g2_decap_8
X_0661_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0074_ Tile_X0Y0_S4END[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
+ _0158_ VPWR VGND sg13g2_mux4_1
X_0730_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[13] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q BM_SRAM13
+ VPWR VGND sg13g2_mux4_1
X_0592_ VGND VPWR _0017_ _0144_ _0148_ _0147_ sg13g2_a21oi_1
X_1213_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1144_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1075_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0928_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0859_ Tile_X0Y1_E2END[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q _0294_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_45_35 VPWR VGND sg13g2_decap_8
XFILLER_45_79 VPWR VGND sg13g2_decap_8
XFILLER_86_86 VPWR VGND sg13g2_decap_8
XFILLER_34_148 VPWR VGND sg13g2_fill_1
X_1693_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 Tile_X0Y1_W2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_0644_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q DOUT_SRAM3
+ DOUT_SRAM15 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 _0081_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3
+ VPWR VGND sg13g2_mux4_1
X_0713_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_EE4END[4] Tile_X0Y1_EE4END[12] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q DIN_SRAM12
+ VPWR VGND sg13g2_mux4_1
X_0575_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q VPWR
+ _0133_ VGND _0131_ _0132_ sg13g2_o21ai_1
X_1127_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1058_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_40_107 VPWR VGND sg13g2_decap_8
XFILLER_40_118 VPWR VGND sg13g2_fill_1
XFILLER_16_148 VPWR VGND sg13g2_decap_4
X_0360_ VPWR VGND _0057_ _0058_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ _0003_ _0059_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a221oi_1
X_0558_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q VPWR
+ _0118_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
X_0627_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q DOUT_SRAM2
+ DOUT_SRAM10 _0079_ _0082_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 VPWR VGND sg13g2_mux4_1
X_1676_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1 Tile_X0Y1_S4BEG[13]
+ VPWR VGND sg13g2_buf_1
X_0489_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q DOUT_SRAM16
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 VPWR VGND sg13g2_mux4_1
XFILLER_88_151 VPWR VGND sg13g2_fill_2
XFILLER_12_140 VPWR VGND sg13g2_fill_1
XFILLER_8_177 VPWR VGND sg13g2_decap_4
XFILLER_8_111 VPWR VGND sg13g2_decap_8
X_0412_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5
+ Tile_X0Y0_S2MID[5] Tile_X0Y1_N2MID[5] Tile_X0Y0_S2END[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 VPWR VGND sg13g2_mux4_1
X_1530_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0 Tile_X0Y0_N2BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_79_151 VPWR VGND sg13g2_decap_4
X_1392_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1461_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_0343_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0
+ Tile_X0Y0_S2MID[0] Tile_X0Y1_N2MID[0] Tile_X0Y0_S2END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_79_195 VPWR VGND sg13g2_fill_1
X_1659_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4 Tile_X0Y1_S2BEGb[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_78_76 VPWR VGND sg13g2_decap_8
XFILLER_94_31 VPWR VGND sg13g2_fill_1
X_0961_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0892_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1513_ Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
XFILLER_67_132 VPWR VGND sg13g2_fill_2
X_1375_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1444_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0326_ VPWR _0029_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ VGND sg13g2_inv_1
XFILLER_13_71 VPWR VGND sg13g2_decap_4
XFILLER_43_9 VPWR VGND sg13g2_fill_1
X_1091_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1160_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_90 VPWR VGND sg13g2_decap_8
XFILLER_49_143 VPWR VGND sg13g2_decap_4
X_0944_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0875_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_0 VPWR VGND sg13g2_decap_8
X_1358_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1427_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0309_ VPWR _0012_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q
+ VGND sg13g2_inv_1
X_1289_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_50_14 VPWR VGND sg13g2_fill_1
XFILLER_75_44 VPWR VGND sg13g2_decap_8
XFILLER_75_22 VPWR VGND sg13g2_fill_1
XFILLER_91_76 VPWR VGND sg13g2_fill_2
XFILLER_91_43 VPWR VGND sg13g2_decap_8
XFILLER_91_21 VPWR VGND sg13g2_fill_1
X_0591_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q VPWR
+ _0147_ VGND _0145_ _0146_ sg13g2_o21ai_1
X_0660_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q DOUT_SRAM7
+ DOUT_SRAM11 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 _0081_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11
+ VPWR VGND sg13g2_mux4_1
X_1212_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1143_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1074_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0927_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0789_ VPWR _0228_ _0227_ VGND sg13g2_inv_1
X_0858_ VGND VPWR Tile_X0Y0_S2MID[2] _0037_ _0293_ _0292_ sg13g2_a21oi_1
XFILLER_28_135 VPWR VGND sg13g2_fill_2
XFILLER_61_24 VPWR VGND sg13g2_fill_2
XFILLER_105_151 VPWR VGND sg13g2_fill_1
XFILLER_86_21 VPWR VGND sg13g2_fill_1
XFILLER_10_61 VPWR VGND sg13g2_fill_2
X_0574_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q VPWR
+ _0132_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
X_0643_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q DOUT_SRAM2
+ DOUT_SRAM14 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 _0082_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2
+ VPWR VGND sg13g2_mux4_1
X_1692_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 Tile_X0Y1_W2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_0712_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q Tile_X0Y1_EE4END[3]
+ Tile_X0Y1_EE4END[11] Tile_X0Y1_E6END[11] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q DIN_SRAM11
+ VPWR VGND sg13g2_mux4_1
X_1126_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_0 VPWR VGND sg13g2_fill_2
X_1057_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_138 VPWR VGND sg13g2_decap_4
XFILLER_31_49 VPWR VGND sg13g2_fill_2
XFILLER_56_46 VPWR VGND sg13g2_decap_8
XFILLER_94_4 VPWR VGND sg13g2_fill_1
X_0557_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ _0117_ VPWR VGND sg13g2_nor2b_1
X_1675_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0 Tile_X0Y1_S4BEG[12]
+ VPWR VGND sg13g2_buf_1
X_0626_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q DOUT_SRAM1
+ DOUT_SRAM9 _0078_ _0083_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 VPWR VGND sg13g2_mux4_1
X_1109_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0488_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q DOUT_SRAM23
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 VPWR VGND sg13g2_mux4_1
XFILLER_67_89 VPWR VGND sg13g2_fill_1
XFILLER_83_44 VPWR VGND sg13g2_decap_4
XFILLER_16_82 VPWR VGND sg13g2_decap_4
XFILLER_79_174 VPWR VGND sg13g2_fill_2
X_1391_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0342_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q Tile_X0Y1_E2MID[7]
+ Tile_X0Y1_E2END[7] Tile_X0Y1_E6END[7] _0043_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 VPWR VGND sg13g2_mux4_1
X_0411_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q Tile_X0Y1_E2MID[2]
+ Tile_X0Y1_E6END[2] Tile_X0Y1_E2END[2] _0082_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 VPWR VGND sg13g2_mux4_1
X_1460_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_85_0 VPWR VGND sg13g2_decap_8
X_1658_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 Tile_X0Y1_S2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_1589_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 Tile_X0Y0_W6BEG[6]
+ VPWR VGND sg13g2_buf_1
X_0609_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_E6END[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12
+ _0091_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0
+ VPWR VGND sg13g2_mux4_1
XFILLER_76_166 VPWR VGND sg13g2_fill_1
X_0960_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1512_ Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
X_0891_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_166 VPWR VGND sg13g2_fill_1
XFILLER_67_111 VPWR VGND sg13g2_decap_4
X_1374_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0325_ VPWR _0028_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
+ VGND sg13g2_inv_1
X_1443_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_199 VPWR VGND sg13g2_fill_1
XFILLER_67_188 VPWR VGND sg13g2_fill_1
XFILLER_73_114 VPWR VGND sg13g2_fill_2
XFILLER_58_199 VPWR VGND sg13g2_fill_1
XFILLER_89_54 VPWR VGND sg13g2_fill_1
XFILLER_89_32 VPWR VGND sg13g2_decap_4
X_1090_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_188 VPWR VGND sg13g2_fill_1
XFILLER_49_199 VPWR VGND sg13g2_fill_1
X_0874_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0943_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_62_2 VPWR VGND sg13g2_fill_1
X_0308_ VPWR _0011_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
+ VGND sg13g2_inv_1
X_1357_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1426_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1288_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_103 VPWR VGND sg13g2_decap_4
XFILLER_55_147 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_1__leaf_Tile_X0Y1_UserCLK
+ VPWR VGND sg13g2_buf_8
XFILLER_59_57 VPWR VGND sg13g2_decap_8
XFILLER_61_139 VPWR VGND sg13g2_decap_8
X_0590_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q VPWR
+ _0146_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
X_1142_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1211_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1073_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_45_191 VPWR VGND sg13g2_decap_8
XFILLER_52_106 VPWR VGND sg13g2_fill_1
XFILLER_60_150 VPWR VGND sg13g2_fill_1
X_0926_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0857_ VGND VPWR _0001_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ _0292_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q sg13g2_a21oi_1
X_1409_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0788_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q VPWR
+ _0227_ VGND Tile_X0Y1_E6END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ sg13g2_o21ai_1
XFILLER_101_43 VPWR VGND sg13g2_decap_8
XFILLER_51_150 VPWR VGND sg13g2_fill_1
XFILLER_61_47 VPWR VGND sg13g2_decap_4
XFILLER_86_77 VPWR VGND sg13g2_fill_1
XFILLER_10_84 VPWR VGND sg13g2_decap_8
XFILLER_42_161 VPWR VGND sg13g2_decap_8
XFILLER_42_172 VPWR VGND sg13g2_fill_2
X_1691_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 Tile_X0Y1_W2BEGb[0]
+ VPWR VGND sg13g2_buf_1
X_0711_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y1_EE4END[2]
+ Tile_X0Y1_EE4END[10] Tile_X0Y1_E6END[10] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q DIN_SRAM10
+ VPWR VGND sg13g2_mux4_1
X_0573_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ _0131_ VPWR VGND sg13g2_nor2b_1
X_0642_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q DOUT_SRAM1
+ DOUT_SRAM13 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 _0083_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1
+ VPWR VGND sg13g2_mux4_1
X_1125_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_117 VPWR VGND sg13g2_decap_4
X_1056_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0909_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_199 VPWR VGND sg13g2_fill_1
XFILLER_30_164 VPWR VGND sg13g2_fill_2
X_1674_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3 Tile_X0Y1_S4BEG[11]
+ VPWR VGND sg13g2_buf_1
X_0625_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q DOUT_SRAM0
+ DOUT_SRAM8 _0043_ _0084_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 VPWR VGND sg13g2_mux4_1
X_0556_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q _0116_ VPWR
+ VGND sg13g2_mux2_1
X_0487_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q DOUT_SRAM22
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_30_0 VPWR VGND sg13g2_decap_8
X_1108_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1039_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_26_17 VPWR VGND sg13g2_decap_8
XFILLER_26_28 VPWR VGND sg13g2_fill_1
XFILLER_67_79 VPWR VGND sg13g2_decap_4
XFILLER_83_67 VPWR VGND sg13g2_decap_4
XFILLER_12_197 VPWR VGND sg13g2_fill_2
XFILLER_12_175 VPWR VGND sg13g2_fill_1
X_0410_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2END[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5
+ Tile_X0Y0_S2MID[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
+ _0082_ VPWR VGND sg13g2_mux4_1
X_0341_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q Tile_X0Y1_N2MID[0]
+ Tile_X0Y1_N2END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0
+ Tile_X0Y0_S2MID[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
+ _0043_ VPWR VGND sg13g2_mux4_1
X_1390_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_94_178 VPWR VGND sg13g2_fill_1
XFILLER_78_0 VPWR VGND sg13g2_fill_2
X_0608_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_E6END[4]
+ _0087_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1588_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 Tile_X0Y0_W6BEG[5]
+ VPWR VGND sg13g2_buf_1
X_1726_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 Tile_X0Y1_WW4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_1657_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 Tile_X0Y1_S2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_0539_ VPWR VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ _0100_ _0101_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ ADDR_SRAM9 _0042_ sg13g2_a221oi_1
XFILLER_85_189 VPWR VGND sg13g2_decap_8
XFILLER_85_167 VPWR VGND sg13g2_fill_1
XFILLER_85_156 VPWR VGND sg13g2_fill_2
XFILLER_85_134 VPWR VGND sg13g2_fill_1
XFILLER_85_123 VPWR VGND sg13g2_decap_8
XFILLER_37_49 VPWR VGND sg13g2_fill_1
XFILLER_94_66 VPWR VGND sg13g2_fill_2
XFILLER_94_22 VPWR VGND sg13g2_decap_8
X_0890_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1511_ Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
XFILLER_4_193 VPWR VGND sg13g2_decap_8
XFILLER_4_171 VPWR VGND sg13g2_fill_1
X_1442_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1373_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0324_ VPWR _0027_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ VGND sg13g2_inv_1
XFILLER_90_170 VPWR VGND sg13g2_decap_8
XFILLER_82_159 VPWR VGND sg13g2_decap_8
XFILLER_82_137 VPWR VGND sg13g2_decap_4
X_1709_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10 Tile_X0Y1_W6BEG[10]
+ VPWR VGND sg13g2_buf_1
XFILLER_58_145 VPWR VGND sg13g2_fill_2
XFILLER_64_14 VPWR VGND sg13g2_fill_1
XFILLER_80_79 VPWR VGND sg13g2_fill_1
XFILLER_80_46 VPWR VGND sg13g2_decap_8
XFILLER_8_0 VPWR VGND sg13g2_fill_2
XFILLER_49_101 VPWR VGND sg13g2_fill_2
XFILLER_64_159 VPWR VGND sg13g2_decap_8
X_0873_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0942_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1425_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_29 VPWR VGND sg13g2_fill_2
X_1356_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0307_ VPWR _0010_ Tile_X0Y1_E6END[0] VGND sg13g2_inv_1
X_1287_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_159 VPWR VGND sg13g2_fill_1
XFILLER_34_7 VPWR VGND sg13g2_decap_4
X_1141_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1072_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1210_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_104 VPWR VGND sg13g2_fill_1
X_0925_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0787_ VGND VPWR _0219_ _0221_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0
+ _0226_ sg13g2_a21oi_1
X_0856_ _0288_ _0289_ _0290_ _0291_ VPWR VGND sg13g2_nor3_1
X_1408_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_17 VPWR VGND sg13g2_decap_8
X_1339_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1690_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 Tile_X0Y1_W2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_0641_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q DOUT_SRAM0
+ DOUT_SRAM12 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 _0084_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0
+ VPWR VGND sg13g2_mux4_1
X_0710_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q Tile_X0Y1_EE4END[1]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_E6END[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q DIN_SRAM9
+ VPWR VGND sg13g2_mux4_1
X_0572_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q _0130_ VPWR
+ VGND sg13g2_mux2_1
X_1124_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1055_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_2 VPWR VGND sg13g2_fill_1
X_0839_ _0275_ Tile_X0Y1_E2END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
X_0908_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_72_25 VPWR VGND sg13g2_decap_8
XFILLER_21_40 VPWR VGND sg13g2_fill_1
XFILLER_108_0 VPWR VGND sg13g2_fill_1
XFILLER_97_77 VPWR VGND sg13g2_decap_8
X_0624_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q Tile_X0Y1_N1END[3]
+ DOUT_SRAM1 _0074_ DOUT_SRAM4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 VPWR VGND sg13g2_mux4_1
X_1673_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2 Tile_X0Y1_S4BEG[10]
+ VPWR VGND sg13g2_buf_1
X_0486_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q DOUT_SRAM21
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_23_0 VPWR VGND sg13g2_decap_8
X_0555_ _0113_ _0115_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1
+ VPWR VGND sg13g2_nor2_1
X_1107_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1038_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_42_17 VPWR VGND sg13g2_decap_8
XFILLER_21_143 VPWR VGND sg13g2_decap_8
XFILLER_107_21 VPWR VGND sg13g2_fill_2
XFILLER_88_198 VPWR VGND sg13g2_fill_2
X_0340_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q Tile_X0Y0_E2MID[7]
+ Tile_X0Y0_E2END[7] Tile_X0Y0_E6END[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0
+ VPWR VGND sg13g2_mux4_1
X_1725_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14 Tile_X0Y1_WW4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_0538_ _0101_ Tile_X0Y0_E2END[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_nand2b_1
X_1587_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 Tile_X0Y0_W6BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0607_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0074_ Tile_X0Y0_S4END[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_mux4_1
X_1656_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1 Tile_X0Y1_S2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_0469_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_5_117 VPWR VGND sg13g2_fill_1
XFILLER_76_124 VPWR VGND sg13g2_decap_4
XFILLER_84_190 VPWR VGND sg13g2_decap_4
XFILLER_27_61 VPWR VGND sg13g2_decap_8
X_1510_ Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
X_1441_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_7 VPWR VGND sg13g2_decap_8
X_1372_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0323_ VPWR _0026_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
+ VGND sg13g2_inv_1
X_1708_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9 Tile_X0Y1_W6BEG[9]
+ VPWR VGND sg13g2_buf_1
XFILLER_48_38 VPWR VGND sg13g2_decap_4
X_1639_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData_O[28] VPWR VGND sg13g2_buf_1
XFILLER_58_113 VPWR VGND sg13g2_fill_1
XFILLER_58_168 VPWR VGND sg13g2_decap_8
XFILLER_38_60 VPWR VGND sg13g2_decap_4
X_0941_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0872_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_91 VPWR VGND sg13g2_decap_8
X_1355_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1424_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0306_ VPWR _0009_ Tile_X0Y1_E6END[1] VGND sg13g2_inv_1
X_1286_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_50_39 VPWR VGND sg13g2_fill_2
XFILLER_59_26 VPWR VGND sg13g2_decap_8
X_1140_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1071_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0924_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0786_ VGND VPWR _0028_ _0224_ _0226_ _0225_ sg13g2_a21oi_1
X_0855_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q VPWR
+ _0290_ VGND Tile_X0Y0_S2MID[3] _0283_ sg13g2_o21ai_1
X_1338_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1407_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_45_28 VPWR VGND sg13g2_decap_8
X_1269_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_196 VPWR VGND sg13g2_decap_4
X_0571_ _0127_ _0129_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3
+ VPWR VGND sg13g2_nor2_1
X_0640_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q DOUT_SRAM7
+ DOUT_SRAM15 _0043_ _0084_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7 VPWR VGND sg13g2_mux4_1
X_1123_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1054_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0907_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_124 VPWR VGND sg13g2_fill_1
X_0769_ Tile_X0Y1_E1END[3] Tile_X0Y1_EE4END[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ _0210_ VPWR VGND sg13g2_mux2_1
X_0838_ _0271_ _0272_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ _0274_ VPWR VGND _0273_ sg13g2_nand4_1
XFILLER_15_174 VPWR VGND sg13g2_fill_2
X_1672_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1 Tile_X0Y1_S4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_0623_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q Tile_X0Y1_N1END[2]
+ DOUT_SRAM0 _0067_ DOUT_SRAM5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 VPWR VGND sg13g2_mux4_1
X_0554_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q _0114_
+ _0115_ VPWR VGND sg13g2_nor2_1
X_1106_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0485_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q DOUT_SRAM20
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4 VPWR VGND sg13g2_mux4_1
XFILLER_16_0 VPWR VGND sg13g2_fill_2
X_1037_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_100 VPWR VGND sg13g2_decap_4
XFILLER_21_122 VPWR VGND sg13g2_decap_4
XFILLER_88_144 VPWR VGND sg13g2_decap_8
XFILLER_88_100 VPWR VGND sg13g2_decap_4
XFILLER_12_199 VPWR VGND sg13g2_fill_1
XFILLER_12_122 VPWR VGND sg13g2_fill_1
XFILLER_8_159 VPWR VGND sg13g2_fill_1
XFILLER_32_95 VPWR VGND sg13g2_decap_4
XFILLER_79_155 VPWR VGND sg13g2_fill_2
XFILLER_78_2 VPWR VGND sg13g2_fill_1
X_1724_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13 Tile_X0Y1_WW4BEG[13]
+ VPWR VGND sg13g2_buf_1
X_1586_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 Tile_X0Y0_W6BEG[3]
+ VPWR VGND sg13g2_buf_1
X_0537_ Tile_X0Y0_E2MID[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q _0100_ VPWR
+ VGND sg13g2_nor3_1
X_1655_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 Tile_X0Y1_S2BEGb[0]
+ VPWR VGND sg13g2_buf_1
X_0606_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0067_ Tile_X0Y0_S4END[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_mux4_1
X_0399_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q Tile_X0Y0_E2MID[4]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E6END[11] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_85_158 VPWR VGND sg13g2_fill_1
X_0468_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q DOUT_SRAM21
+ DOUT_SRAM25 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9
+ VPWR VGND sg13g2_mux4_1
XFILLER_37_29 VPWR VGND sg13g2_fill_2
XFILLER_43_72 VPWR VGND sg13g2_fill_1
X_1371_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1440_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0322_ VPWR _0025_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ VGND sg13g2_inv_1
XFILLER_83_0 VPWR VGND sg13g2_fill_2
X_1707_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8 Tile_X0Y1_W6BEG[8]
+ VPWR VGND sg13g2_buf_1
X_1638_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData_O[27] VPWR VGND sg13g2_buf_1
X_1569_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2 Tile_X0Y0_W2BEG[2]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_67 VPWR VGND sg13g2_fill_2
XFILLER_81_172 VPWR VGND sg13g2_fill_1
XFILLER_13_75 VPWR VGND sg13g2_fill_1
XFILLER_13_64 VPWR VGND sg13g2_decap_8
XFILLER_13_42 VPWR VGND sg13g2_fill_1
XFILLER_8_2 VPWR VGND sg13g2_fill_1
XFILLER_1_176 VPWR VGND sg13g2_fill_2
XFILLER_38_83 VPWR VGND sg13g2_decap_8
XFILLER_49_136 VPWR VGND sg13g2_decap_8
XFILLER_49_147 VPWR VGND sg13g2_fill_1
XFILLER_57_180 VPWR VGND sg13g2_fill_1
X_0940_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_54_82 VPWR VGND sg13g2_fill_1
X_0871_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1354_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1285_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1423_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0305_ VPWR _0008_ Tile_X0Y1_E6END[2] VGND sg13g2_inv_1
XFILLER_39_180 VPWR VGND sg13g2_fill_2
X_1070_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0923_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0854_ Tile_X0Y1_E2END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q _0289_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_60_175 VPWR VGND sg13g2_fill_2
X_0785_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q VPWR
+ _0225_ VGND _0222_ _0223_ sg13g2_o21ai_1
X_1337_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1268_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1406_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_79 VPWR VGND sg13g2_fill_2
X_1199_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_105_199 VPWR VGND sg13g2_fill_1
XFILLER_19_96 VPWR VGND sg13g2_decap_4
X_0570_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q _0128_
+ _0129_ VPWR VGND sg13g2_nor2_1
XFILLER_51_83 VPWR VGND sg13g2_fill_1
XFILLER_51_94 VPWR VGND sg13g2_fill_1
X_1122_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_197 VPWR VGND sg13g2_fill_2
X_1053_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0906_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0837_ VGND VPWR _0273_ _0258_ Tile_X0Y0_S2MID[3] sg13g2_or2_1
X_0699_ VGND VPWR Tile_X0Y1_E2END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ _0176_ _0175_ sg13g2_a21oi_1
X_0768_ _0208_ VPWR _0209_ VGND _0025_ _0158_ sg13g2_o21ai_1
XFILLER_56_39 VPWR VGND sg13g2_decap_8
XFILLER_97_46 VPWR VGND sg13g2_fill_2
XFILLER_97_24 VPWR VGND sg13g2_decap_4
XFILLER_21_31 VPWR VGND sg13g2_decap_8
XFILLER_15_131 VPWR VGND sg13g2_fill_2
XFILLER_87_7 VPWR VGND sg13g2_decap_4
X_1671_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0 Tile_X0Y1_S4BEG[8]
+ VPWR VGND sg13g2_buf_1
XFILLER_62_71 VPWR VGND sg13g2_decap_4
X_0484_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y1_N4END[7]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3 VPWR VGND sg13g2_mux4_1
X_0622_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q Tile_X0Y1_N1END[1]
+ DOUT_SRAM3 _0060_ DOUT_SRAM6 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 VPWR VGND sg13g2_mux4_1
X_0553_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q _0114_ VPWR
+ VGND sg13g2_mux4_1
X_1105_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1036_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_83_48 VPWR VGND sg13g2_fill_2
XFILLER_83_26 VPWR VGND sg13g2_fill_1
XFILLER_16_64 VPWR VGND sg13g2_fill_1
XFILLER_16_42 VPWR VGND sg13g2_fill_1
XFILLER_57_71 VPWR VGND sg13g2_fill_1
XFILLER_57_93 VPWR VGND sg13g2_fill_1
X_1723_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12 Tile_X0Y1_WW4BEG[12]
+ VPWR VGND sg13g2_buf_1
X_1654_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 Tile_X0Y1_S2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_0536_ VPWR VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ _0098_ _0099_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ ADDR_SRAM8 _0041_ sg13g2_a221oi_1
X_0467_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 VPWR VGND sg13g2_mux4_1
X_1585_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 Tile_X0Y0_W6BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0605_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0060_ Tile_X0Y0_S4END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_mux4_1
X_0398_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2END[5] Tile_X0Y0_E6END[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2
+ VPWR VGND sg13g2_mux4_1
X_1019_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_78_48 VPWR VGND sg13g2_decap_8
X_1370_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0321_ VPWR _0024_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
+ VGND sg13g2_inv_1
XFILLER_76_0 VPWR VGND sg13g2_fill_2
X_1706_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7 Tile_X0Y1_W6BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1637_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameData_O[26] VPWR VGND sg13g2_buf_1
X_1499_ Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData_O[25] VPWR VGND sg13g2_buf_1
X_0519_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[10] Tile_X0Y0_E6END[10] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q BM_SRAM26
+ VPWR VGND sg13g2_mux4_1
X_1568_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1 Tile_X0Y0_W2BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_89_36 VPWR VGND sg13g2_fill_1
XFILLER_89_25 VPWR VGND sg13g2_decap_8
XFILLER_49_115 VPWR VGND sg13g2_decap_4
XFILLER_38_51 VPWR VGND sg13g2_fill_1
X_0870_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1422_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1353_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1284_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0304_ VPWR _0007_ Tile_X0Y1_E6END[3] VGND sg13g2_inv_1
XFILLER_48_170 VPWR VGND sg13g2_decap_8
XFILLER_63_173 VPWR VGND sg13g2_fill_1
XFILLER_63_195 VPWR VGND sg13g2_decap_4
X_0999_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_42 VPWR VGND sg13g2_fill_1
XFILLER_6_0 VPWR VGND sg13g2_fill_2
XFILLER_49_83 VPWR VGND sg13g2_fill_1
XFILLER_45_184 VPWR VGND sg13g2_decap_8
X_0922_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0853_ _0037_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0 _0288_ VPWR VGND sg13g2_nor3_1
X_0784_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q _0224_ VPWR
+ VGND sg13g2_mux2_1
X_1405_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1336_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1198_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1267_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_105_178 VPWR VGND sg13g2_fill_1
XFILLER_42_198 VPWR VGND sg13g2_fill_2
X_1121_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_76_70 VPWR VGND sg13g2_fill_1
X_1052_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_195 VPWR VGND sg13g2_decap_4
X_0905_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0767_ VPWR _0208_ _0207_ VGND sg13g2_inv_1
X_0836_ Tile_X0Y1_E2END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q _0272_ VPWR
+ VGND sg13g2_or3_1
X_0698_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q Tile_X0Y1_E2MID[4]
+ _0175_ VPWR VGND sg13g2_nor2b_1
X_1319_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_198 VPWR VGND sg13g2_fill_2
XFILLER_15_198 VPWR VGND sg13g2_fill_2
XFILLER_15_176 VPWR VGND sg13g2_fill_1
X_1670_ Tile_X0Y0_S4END[15] Tile_X0Y1_S4BEG[7] VPWR VGND sg13g2_buf_1
X_0621_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q Tile_X0Y1_N1END[0]
+ DOUT_SRAM2 _0088_ DOUT_SRAM7 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
X_0483_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q Tile_X0Y1_N4END[6]
+ Tile_X0Y0_S4END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2 VPWR VGND sg13g2_mux4_1
X_0552_ VGND VPWR _0012_ _0109_ _0113_ _0112_ sg13g2_a21oi_1
X_1104_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1035_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_0819_ VGND VPWR _0034_ _0254_ _0256_ _0255_ sg13g2_a21oi_1
XFILLER_12_102 VPWR VGND sg13g2_fill_2
X_1584_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 Tile_X0Y0_W6BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1722_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11 Tile_X0Y1_WW4BEG[11]
+ VPWR VGND sg13g2_buf_1
X_0604_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0088_ Tile_X0Y0_S4END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_mux4_1
X_1653_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 Tile_X0Y1_S2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_0535_ _0099_ Tile_X0Y0_E2END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_nand2b_1
X_0397_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2
+ Tile_X0Y1_N2MID[2] Tile_X0Y0_S2MID[2] Tile_X0Y0_S2END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 VPWR VGND sg13g2_mux4_1
X_0466_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q DOUT_SRAM20
+ DOUT_SRAM24 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8
+ VPWR VGND sg13g2_mux4_1
XFILLER_21_0 VPWR VGND sg13g2_decap_8
X_1018_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_76_116 VPWR VGND sg13g2_decap_4
XFILLER_4_164 VPWR VGND sg13g2_decap_8
X_0320_ VPWR _0023_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ VGND sg13g2_inv_1
XFILLER_90_163 VPWR VGND sg13g2_decap_8
XFILLER_69_0 VPWR VGND sg13g2_fill_1
X_1705_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6 Tile_X0Y1_W6BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1636_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData_O[25] VPWR VGND sg13g2_buf_1
X_1567_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0 Tile_X0Y0_W2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0518_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y0_EE4END[1]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_E6END[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q BM_SRAM25
+ VPWR VGND sg13g2_mux4_1
X_1498_ Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData_O[24] VPWR VGND sg13g2_buf_1
XFILLER_58_138 VPWR VGND sg13g2_decap_8
X_0449_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q DOUT_SRAM21
+ DOUT_SRAM29 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5
+ VPWR VGND sg13g2_mux4_1
XFILLER_80_39 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_fill_2
XFILLER_1_178 VPWR VGND sg13g2_fill_1
XFILLER_54_40 VPWR VGND sg13g2_fill_2
XFILLER_70_50 VPWR VGND sg13g2_fill_2
X_1421_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0303_ VPWR _0006_ Tile_X0Y0_E6END[0] VGND sg13g2_inv_1
X_1352_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1283_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_141 VPWR VGND sg13g2_decap_8
X_0998_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1619_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_39_182 VPWR VGND sg13g2_fill_1
XFILLER_24_98 VPWR VGND sg13g2_fill_2
XFILLER_40_42 VPWR VGND sg13g2_fill_2
XFILLER_49_62 VPWR VGND sg13g2_decap_8
X_0921_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_177 VPWR VGND sg13g2_fill_1
XFILLER_81_93 VPWR VGND sg13g2_decap_8
X_0783_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q VPWR
+ _0223_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
X_0852_ _0286_ VPWR _0287_ VGND _0037_ _0279_ sg13g2_o21ai_1
XFILLER_60_199 VPWR VGND sg13g2_fill_1
X_1335_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1404_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1197_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1266_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_100 VPWR VGND sg13g2_decap_4
XFILLER_10_34 VPWR VGND sg13g2_fill_2
XFILLER_19_21 VPWR VGND sg13g2_decap_4
XFILLER_35_64 VPWR VGND sg13g2_fill_1
XFILLER_42_133 VPWR VGND sg13g2_decap_8
X_1120_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_141 VPWR VGND sg13g2_fill_2
X_1051_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0904_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_122 VPWR VGND sg13g2_decap_8
XFILLER_33_199 VPWR VGND sg13g2_fill_1
X_0697_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q _0081_
+ _0174_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ sg13g2_nand3b_1
X_0766_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q VPWR
+ _0207_ VGND Tile_X0Y1_E6END[11] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ sg13g2_o21ai_1
XFILLER_51_0 VPWR VGND sg13g2_decap_8
X_0835_ _0271_ _0257_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0
+ VPWR VGND sg13g2_nand2b_1
X_1318_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1249_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_40 VPWR VGND Tile_X0Y1_N2MID[7] sg13g2_antennanp
XFILLER_97_48 VPWR VGND sg13g2_fill_1
XFILLER_15_100 VPWR VGND sg13g2_fill_2
X_0620_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_E2END[0] Tile_X0Y1_E2MID[0] _0084_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7 VPWR VGND sg13g2_mux4_1
X_0551_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q VPWR
+ _0112_ VGND _0110_ _0111_ sg13g2_o21ai_1
XFILLER_97_147 VPWR VGND sg13g2_fill_2
XFILLER_97_114 VPWR VGND sg13g2_fill_2
X_0482_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q Tile_X0Y1_N4END[5]
+ Tile_X0Y0_S4END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1 VPWR VGND sg13g2_mux4_1
X_1103_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1034_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0818_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q VPWR
+ _0255_ VGND _0252_ _0253_ sg13g2_o21ai_1
X_0749_ _0021_ _0078_ _0192_ VPWR VGND sg13g2_nor2_1
XFILLER_8_118 VPWR VGND sg13g2_fill_2
X_1721_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10 Tile_X0Y1_WW4BEG[10]
+ VPWR VGND sg13g2_buf_1
XFILLER_7_140 VPWR VGND sg13g2_fill_2
X_0603_ _0155_ _0157_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3
+ VPWR VGND sg13g2_nor2_1
X_0534_ Tile_X0Y0_E2MID[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q _0098_ VPWR
+ VGND sg13g2_nor3_1
X_1583_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 Tile_X0Y0_W6BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1652_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 Tile_X0Y1_S2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0465_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 VPWR VGND sg13g2_mux4_1
X_0396_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E6END[5] Tile_X0Y1_E2END[5] _0079_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 VPWR VGND sg13g2_mux4_1
X_1017_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_76_128 VPWR VGND sg13g2_fill_2
XFILLER_27_54 VPWR VGND sg13g2_decap_8
XFILLER_43_31 VPWR VGND sg13g2_fill_1
XFILLER_4_110 VPWR VGND sg13g2_fill_1
XFILLER_68_94 VPWR VGND sg13g2_decap_8
X_1704_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5 Tile_X0Y1_W6BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0517_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[8] Tile_X0Y0_E6END[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q BM_SRAM24
+ VPWR VGND sg13g2_mux4_1
X_1497_ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData_O[23] VPWR VGND sg13g2_buf_1
X_1635_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData_O[24] VPWR VGND sg13g2_buf_1
X_1566_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3 Tile_X0Y0_W1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_26 VPWR VGND sg13g2_fill_1
X_0379_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3 _0072_ VPWR VGND sg13g2_nor3_1
XFILLER_81_120 VPWR VGND sg13g2_fill_2
X_0448_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q DOUT_SRAM20
+ DOUT_SRAM28 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4
+ VPWR VGND sg13g2_mux4_1
XFILLER_38_64 VPWR VGND sg13g2_fill_2
XFILLER_38_97 VPWR VGND sg13g2_decap_8
XFILLER_72_197 VPWR VGND sg13g2_fill_2
XFILLER_72_186 VPWR VGND sg13g2_fill_2
XFILLER_72_131 VPWR VGND sg13g2_decap_8
X_0302_ VPWR _0005_ Tile_X0Y0_E6END[3] VGND sg13g2_inv_1
X_1351_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1420_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_7 VPWR VGND sg13g2_decap_8
X_1282_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_81_0 VPWR VGND sg13g2_fill_1
X_0997_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1618_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_59_19 VPWR VGND sg13g2_decap_8
X_1549_ Tile_X0Y1_N4END[11] Tile_X0Y0_N4BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_91_17 VPWR VGND sg13g2_decap_4
XFILLER_6_2 VPWR VGND sg13g2_fill_1
XFILLER_45_142 VPWR VGND sg13g2_decap_8
X_0920_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0782_ _0027_ _0081_ _0222_ VPWR VGND sg13g2_nor2_1
X_0851_ _0286_ _0284_ _0285_ _0282_ _0280_ VPWR VGND sg13g2_a22oi_1
X_1334_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1403_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1265_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1196_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_86_39 VPWR VGND sg13g2_fill_1
XFILLER_19_77 VPWR VGND sg13g2_fill_2
X_1050_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_7 VPWR VGND sg13g2_fill_1
X_0903_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0834_ _0266_ _0269_ _0264_ _0270_ VPWR VGND sg13g2_nand3_1
XFILLER_102_117 VPWR VGND sg13g2_decap_8
XFILLER_44_0 VPWR VGND sg13g2_decap_4
X_0765_ VGND VPWR _0199_ _0201_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A _0206_ sg13g2_a21oi_1
X_0696_ _0171_ VPWR ADDR_SRAM3 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
+ _0173_ sg13g2_o21ai_1
X_1317_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1248_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1179_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_30 VPWR VGND Tile_X0Y1_N2MID[0] sg13g2_antennanp
XANTENNA_41 VPWR VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0
+ sg13g2_antennanp
XFILLER_102_92 VPWR VGND sg13g2_decap_4
XFILLER_15_156 VPWR VGND sg13g2_fill_1
XFILLER_7_47 VPWR VGND sg13g2_fill_2
X_0550_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q VPWR
+ _0111_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
X_0481_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q Tile_X0Y1_N4END[4]
+ Tile_X0Y0_S4END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0 VPWR VGND sg13g2_mux4_1
X_1102_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1033_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_104 VPWR VGND sg13g2_fill_1
X_0817_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q _0254_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_88_104 VPWR VGND sg13g2_fill_2
X_0679_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q DOUT_SRAM2
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 _0160_ _0083_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10
+ VPWR VGND sg13g2_mux4_1
X_0748_ VGND VPWR _0022_ _0190_ _0191_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q
+ sg13g2_a21oi_1
XFILLER_12_104 VPWR VGND sg13g2_fill_1
XFILLER_32_99 VPWR VGND sg13g2_fill_1
XFILLER_94_107 VPWR VGND sg13g2_fill_1
XFILLER_85_7 VPWR VGND sg13g2_decap_8
X_1720_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9 Tile_X0Y1_WW4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_1651_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 Tile_X0Y1_S2BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0602_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q _0156_
+ _0157_ VPWR VGND sg13g2_nor2_1
X_0533_ VPWR VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ _0096_ _0097_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ ADDR_SRAM7 _0040_ sg13g2_a221oi_1
X_0464_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q DOUT_SRAM23
+ DOUT_SRAM27 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7
+ VPWR VGND sg13g2_mux4_1
X_1582_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7 Tile_X0Y0_W2BEGb[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_93_195 VPWR VGND sg13g2_decap_4
XFILLER_93_173 VPWR VGND sg13g2_decap_4
X_0395_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q Tile_X0Y1_N2MID[2]
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2 Tile_X0Y1_N2END[2]
+ Tile_X0Y0_S2MID[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
+ _0079_ VPWR VGND sg13g2_mux4_1
X_1016_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_170 VPWR VGND sg13g2_decap_8
XFILLER_27_11 VPWR VGND sg13g2_fill_2
XFILLER_84_162 VPWR VGND sg13g2_decap_8
XFILLER_4_37 VPWR VGND sg13g2_fill_2
XFILLER_90_121 VPWR VGND sg13g2_decap_4
XFILLER_90_198 VPWR VGND sg13g2_fill_2
X_1703_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4 Tile_X0Y1_W6BEG[4]
+ VPWR VGND sg13g2_buf_1
X_1634_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData_O[23] VPWR VGND sg13g2_buf_1
X_0516_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y0_EE4END[7]
+ Tile_X0Y0_EE4END[15] Tile_X0Y0_E6END[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q BM_SRAM23
+ VPWR VGND sg13g2_mux4_1
X_1496_ Tile_X0Y0_FrameData[22] Tile_X0Y0_FrameData_O[22] VPWR VGND sg13g2_buf_1
X_0447_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q DOUT_SRAM19
+ DOUT_SRAM27 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3
+ VPWR VGND sg13g2_mux4_1
X_1565_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2 Tile_X0Y0_W1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0378_ _0071_ Tile_X0Y0_S1END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_81_198 VPWR VGND sg13g2_fill_2
XFILLER_81_165 VPWR VGND sg13g2_decap_8
XFILLER_1_158 VPWR VGND sg13g2_fill_1
XFILLER_70_52 VPWR VGND sg13g2_fill_1
X_0301_ VPWR _0004_ Tile_X0Y0_E6END[2] VGND sg13g2_inv_1
X_1350_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1281_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0996_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_0 VPWR VGND sg13g2_fill_2
X_1617_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData_O[6] VPWR VGND sg13g2_buf_1
X_1479_ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData_O[5] VPWR VGND sg13g2_buf_1
X_1548_ Tile_X0Y1_N4END[10] Tile_X0Y0_N4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_108_112 VPWR VGND sg13g2_fill_2
XFILLER_45_198 VPWR VGND sg13g2_fill_2
X_0850_ VGND VPWR Tile_X0Y1_E2MID[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0285_ _0283_ sg13g2_a21oi_1
XFILLER_60_146 VPWR VGND sg13g2_decap_4
XFILLER_60_168 VPWR VGND sg13g2_decap_8
X_0781_ VGND VPWR _0028_ _0220_ _0221_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
+ sg13g2_a21oi_1
X_1402_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1333_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1264_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_17 VPWR VGND sg13g2_fill_1
X_1195_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_168 VPWR VGND sg13g2_decap_8
X_0979_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_110 VPWR VGND sg13g2_decap_4
XFILLER_42_168 VPWR VGND sg13g2_decap_4
XFILLER_92_94 VPWR VGND sg13g2_fill_1
XFILLER_18_121 VPWR VGND sg13g2_fill_2
XFILLER_18_143 VPWR VGND sg13g2_fill_1
X_0902_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0833_ _0269_ _0268_ _0257_ _0261_ _0259_ VPWR VGND sg13g2_a22oi_1
XFILLER_37_0 VPWR VGND sg13g2_decap_4
X_0764_ VGND VPWR _0024_ _0204_ _0206_ _0205_ sg13g2_a21oi_1
X_0695_ VGND VPWR Tile_X0Y1_E2END[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ _0173_ _0172_ sg13g2_a21oi_1
X_1316_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1247_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1178_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_20 VPWR VGND Tile_X0Y1_FrameStrobe[16] sg13g2_antennanp
XANTENNA_31 VPWR VGND Tile_X0Y1_N2MID[3] sg13g2_antennanp
XFILLER_97_28 VPWR VGND sg13g2_fill_1
XFILLER_21_79 VPWR VGND sg13g2_decap_4
XANTENNA_42 VPWR VGND Tile_X0Y0_S2MID[6] sg13g2_antennanp
XFILLER_99_190 VPWR VGND sg13g2_fill_2
XFILLER_15_124 VPWR VGND sg13g2_decap_8
XFILLER_15_102 VPWR VGND sg13g2_fill_1
XFILLER_62_75 VPWR VGND sg13g2_fill_2
XFILLER_97_116 VPWR VGND sg13g2_fill_1
X_0480_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q DOUT_SRAM19
+ DOUT_SRAM31 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15
+ VPWR VGND sg13g2_mux4_1
XFILLER_30_7 VPWR VGND sg13g2_fill_2
X_1101_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1032_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0816_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q VPWR
+ _0253_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
X_0747_ Tile_X0Y1_E1END[1] Tile_X0Y1_EE4END[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ _0190_ VPWR VGND sg13g2_mux2_1
X_0678_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q DOUT_SRAM1
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 _0159_ _0082_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9
+ VPWR VGND sg13g2_mux4_1
XFILLER_83_19 VPWR VGND sg13g2_decap_8
XFILLER_16_35 VPWR VGND sg13g2_decap_8
XFILLER_73_74 VPWR VGND sg13g2_fill_2
X_0601_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E6END[7] Tile_X0Y0_EE4END[15] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q _0156_ VPWR
+ VGND sg13g2_mux4_1
XFILLER_7_197 VPWR VGND sg13g2_fill_2
X_1650_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 Tile_X0Y1_S2BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1581_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6 Tile_X0Y0_W2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_0463_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8 VPWR VGND sg13g2_mux4_1
X_0394_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2END[5] Tile_X0Y0_E6END[10] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2
+ VPWR VGND sg13g2_mux4_1
X_0532_ _0097_ Tile_X0Y0_E2END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_nand2b_1
X_1015_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_91 VPWR VGND sg13g2_fill_2
XFILLER_94_29 VPWR VGND sg13g2_fill_2
XFILLER_27_34 VPWR VGND sg13g2_fill_2
XFILLER_104_0 VPWR VGND sg13g2_fill_1
XFILLER_68_41 VPWR VGND sg13g2_decap_8
X_1702_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 Tile_X0Y1_W6BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1564_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1 Tile_X0Y0_W1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1633_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameData_O[22] VPWR VGND sg13g2_buf_1
X_0377_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E6END[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14
+ _0066_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux4_1
X_1495_ Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData_O[21] VPWR VGND sg13g2_buf_1
X_0515_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q Tile_X0Y0_EE4END[6]
+ Tile_X0Y0_EE4END[14] Tile_X0Y0_E6END[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q BM_SRAM22
+ VPWR VGND sg13g2_mux4_1
X_0446_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q DOUT_SRAM18
+ DOUT_SRAM26 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_122 VPWR VGND sg13g2_fill_1
XFILLER_81_100 VPWR VGND sg13g2_fill_2
XFILLER_66_174 VPWR VGND sg13g2_decap_4
XFILLER_49_108 VPWR VGND sg13g2_decap_8
XFILLER_72_100 VPWR VGND sg13g2_decap_4
XFILLER_110_60 VPWR VGND sg13g2_fill_1
XFILLER_72_199 VPWR VGND sg13g2_fill_1
XFILLER_72_188 VPWR VGND sg13g2_fill_1
XFILLER_70_31 VPWR VGND sg13g2_fill_2
XFILLER_95_72 VPWR VGND sg13g2_fill_2
X_0300_ VPWR _0003_ Tile_X0Y0_E6END[1] VGND sg13g2_inv_1
X_1280_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_122 VPWR VGND sg13g2_fill_2
XFILLER_63_199 VPWR VGND sg13g2_fill_1
X_0995_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_0 VPWR VGND sg13g2_fill_2
X_1547_ Tile_X0Y1_N4END[9] Tile_X0Y0_N4BEG[1] VPWR VGND sg13g2_buf_1
X_1616_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData_O[5] VPWR VGND sg13g2_buf_1
X_1478_ Tile_X0Y0_FrameData[4] Tile_X0Y0_FrameData_O[4] VPWR VGND sg13g2_buf_1
X_0429_ _0090_ _0088_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_54_199 VPWR VGND sg13g2_fill_1
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_49_76 VPWR VGND sg13g2_decap_8
X_0780_ Tile_X0Y1_E1END[0] Tile_X0Y1_EE4END[12] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ _0220_ VPWR VGND sg13g2_mux2_1
X_1401_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1194_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1332_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1263_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0978_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_86_19 VPWR VGND sg13g2_fill_2
XFILLER_27_199 VPWR VGND sg13g2_fill_1
XFILLER_51_11 VPWR VGND sg13g2_fill_2
XFILLER_18_199 VPWR VGND sg13g2_fill_1
X_0901_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0763_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q VPWR
+ _0205_ VGND _0202_ _0203_ sg13g2_o21ai_1
X_0832_ VGND VPWR Tile_X0Y1_N2END[3] _0035_ _0268_ _0267_ sg13g2_a21oi_1
X_1315_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0694_ _0000_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ _0172_ VPWR VGND sg13g2_nor2_1
X_1177_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1246_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_43 VPWR VGND Tile_X0Y0_S2MID[6] sg13g2_antennanp
XANTENNA_21 VPWR VGND Tile_X0Y1_FrameStrobe[16] sg13g2_antennanp
XANTENNA_32 VPWR VGND Tile_X0Y1_N2MID[3] sg13g2_antennanp
XANTENNA_10 VPWR VGND Tile_X0Y0_S2MID[4] sg13g2_antennanp
XFILLER_7_49 VPWR VGND sg13g2_fill_1
XFILLER_62_98 VPWR VGND sg13g2_decap_4
XFILLER_87_40 VPWR VGND sg13g2_fill_1
XFILLER_11_80 VPWR VGND sg13g2_decap_8
XFILLER_23_7 VPWR VGND sg13g2_decap_4
X_1100_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1031_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_191 VPWR VGND sg13g2_decap_8
X_0815_ _0033_ _0084_ _0252_ VPWR VGND sg13g2_nor2_1
X_0746_ _0188_ VPWR _0189_ VGND _0021_ _0160_ sg13g2_o21ai_1
XFILLER_96_161 VPWR VGND sg13g2_fill_2
X_0677_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q DOUT_SRAM0
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 _0158_ _0081_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8
+ VPWR VGND sg13g2_mux4_1
X_1229_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_79_117 VPWR VGND sg13g2_decap_4
XFILLER_87_194 VPWR VGND sg13g2_decap_4
X_0600_ VGND VPWR _0018_ _0151_ _0155_ _0154_ sg13g2_a21oi_1
X_0531_ Tile_X0Y0_E2MID[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q _0096_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_7_176 VPWR VGND sg13g2_decap_4
X_1580_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5 Tile_X0Y0_W2BEGb[5]
+ VPWR VGND sg13g2_buf_1
X_0393_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q Tile_X0Y0_E2MID[6]
+ Tile_X0Y0_E2END[6] Tile_X0Y0_E6END[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1
+ VPWR VGND sg13g2_mux4_1
X_0462_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q DOUT_SRAM22
+ DOUT_SRAM26 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6
+ VPWR VGND sg13g2_mux4_1
X_1014_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_97_0 VPWR VGND sg13g2_decap_8
X_0729_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_EE4END[4] Tile_X0Y1_EE4END[12] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q BM_SRAM12
+ VPWR VGND sg13g2_mux4_1
XFILLER_76_109 VPWR VGND sg13g2_decap_8
XFILLER_27_68 VPWR VGND sg13g2_fill_1
X_1701_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 Tile_X0Y1_W6BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1494_ Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData_O[20] VPWR VGND sg13g2_buf_1
X_1563_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0 Tile_X0Y0_W1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0514_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y0_EE4END[5]
+ Tile_X0Y0_EE4END[13] Tile_X0Y0_E6END[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q BM_SRAM21
+ VPWR VGND sg13g2_mux4_1
X_1632_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData_O[21] VPWR VGND sg13g2_buf_1
X_0376_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_mux4_1
XFILLER_66_153 VPWR VGND sg13g2_decap_4
X_0445_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q DOUT_SRAM17
+ DOUT_SRAM25 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_134 VPWR VGND sg13g2_fill_2
XFILLER_72_145 VPWR VGND sg13g2_decap_8
XFILLER_70_98 VPWR VGND sg13g2_decap_4
XFILLER_48_197 VPWR VGND sg13g2_fill_2
X_0994_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_2 VPWR VGND sg13g2_fill_1
X_1477_ Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData_O[3] VPWR VGND sg13g2_buf_1
X_1546_ Tile_X0Y1_N4END[8] Tile_X0Y0_N4BEG[0] VPWR VGND sg13g2_buf_1
X_1615_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameData_O[4] VPWR VGND sg13g2_buf_1
X_0359_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1 _0058_ VPWR VGND sg13g2_nor3_1
X_0428_ Tile_X0Y1_N1END[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q _0089_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_108_125 VPWR VGND sg13g2_fill_2
XFILLER_81_53 VPWR VGND sg13g2_fill_2
XFILLER_81_42 VPWR VGND sg13g2_decap_8
XFILLER_81_20 VPWR VGND sg13g2_fill_1
XFILLER_65_98 VPWR VGND sg13g2_fill_2
XFILLER_45_112 VPWR VGND sg13g2_fill_2
X_1331_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1400_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1193_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1262_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_104 VPWR VGND sg13g2_fill_1
X_0977_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1529_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3 Tile_X0Y0_N1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_19_25 VPWR VGND sg13g2_fill_1
XFILLER_42_126 VPWR VGND sg13g2_decap_8
XFILLER_18_123 VPWR VGND sg13g2_fill_1
X_0900_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_115 VPWR VGND sg13g2_decap_8
XFILLER_41_170 VPWR VGND sg13g2_fill_1
XFILLER_41_192 VPWR VGND sg13g2_decap_8
X_0762_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q _0204_ VPWR
+ VGND sg13g2_mux2_1
X_0693_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q _0080_
+ _0171_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ sg13g2_nand3b_1
X_0831_ Tile_X0Y1_E2MID[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ _0267_ VPWR VGND sg13g2_and2_1
X_1314_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1176_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1245_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_22 VPWR VGND Tile_X0Y1_FrameStrobe[16] sg13g2_antennanp
XANTENNA_11 VPWR VGND Tile_X0Y0_S2MID[4] sg13g2_antennanp
XANTENNA_33 VPWR VGND Tile_X0Y1_N2MID[4] sg13g2_antennanp
XANTENNA_44 VPWR VGND Tile_X0Y0_S2MID[6] sg13g2_antennanp
XFILLER_102_73 VPWR VGND sg13g2_fill_2
XFILLER_15_137 VPWR VGND sg13g2_fill_2
XFILLER_7_17 VPWR VGND sg13g2_fill_1
XFILLER_30_9 VPWR VGND sg13g2_fill_1
X_1030_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0814_ VGND VPWR _0034_ _0250_ _0251_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
+ sg13g2_a21oi_1
X_0676_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q DOUT_SRAM7
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ _0080_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7
+ VPWR VGND sg13g2_mux4_1
X_0745_ VPWR _0188_ _0187_ VGND sg13g2_inv_1
X_1228_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1159_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_140 VPWR VGND sg13g2_decap_8
XFILLER_73_21 VPWR VGND sg13g2_fill_2
X_0530_ VPWR VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ _0094_ _0095_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ ADDR_SRAM6 _0039_ sg13g2_a221oi_1
XFILLER_7_199 VPWR VGND sg13g2_fill_1
XFILLER_7_133 VPWR VGND sg13g2_decap_8
X_0392_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1
+ Tile_X0Y0_S2MID[1] Tile_X0Y1_N2MID[1] Tile_X0Y0_S2END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 VPWR VGND sg13g2_mux4_1
X_0461_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9 VPWR VGND sg13g2_mux4_1
X_1013_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_93 VPWR VGND sg13g2_fill_1
X_0659_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0088_ Tile_X0Y0_S4END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 VPWR VGND sg13g2_mux4_1
X_0728_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q Tile_X0Y1_EE4END[3]
+ Tile_X0Y1_EE4END[11] Tile_X0Y1_E6END[11] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q BM_SRAM11
+ VPWR VGND sg13g2_mux4_1
XFILLER_84_198 VPWR VGND sg13g2_fill_2
XFILLER_27_36 VPWR VGND sg13g2_fill_1
XFILLER_75_132 VPWR VGND sg13g2_fill_2
XFILLER_75_110 VPWR VGND sg13g2_fill_1
XFILLER_84_97 VPWR VGND sg13g2_fill_1
XFILLER_75_198 VPWR VGND sg13g2_fill_2
X_1700_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 Tile_X0Y1_W6BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1631_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData_O[20] VPWR VGND sg13g2_buf_1
X_1562_ clknet_1_1__leaf_Tile_X0Y1_UserCLK Tile_X0Y0_UserCLKo VPWR VGND sg13g2_buf_1
X_0513_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_E6END[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q BM_SRAM20
+ VPWR VGND sg13g2_mux4_1
X_1493_ Tile_X0Y0_FrameData[19] Tile_X0Y0_FrameData_O[19] VPWR VGND sg13g2_buf_1
X_0444_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q DOUT_SRAM16
+ DOUT_SRAM24 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_102 VPWR VGND sg13g2_fill_1
X_0375_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 Tile_X0Y1_E6END[6]
+ _0070_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_157 VPWR VGND sg13g2_decap_4
XFILLER_57_132 VPWR VGND sg13g2_decap_8
XFILLER_57_198 VPWR VGND sg13g2_fill_2
XFILLER_70_11 VPWR VGND sg13g2_fill_2
XFILLER_0_172 VPWR VGND sg13g2_fill_2
X_0993_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_2 VPWR VGND sg13g2_fill_1
X_1614_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData_O[3] VPWR VGND sg13g2_buf_1
X_1545_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 Tile_X0Y0_N2BEGb[7]
+ VPWR VGND sg13g2_buf_1
X_0427_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_E6END[8]
+ _0087_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q _0088_
+ VPWR VGND sg13g2_mux4_1
X_1476_ Tile_X0Y0_FrameData[2] Tile_X0Y0_FrameData_O[2] VPWR VGND sg13g2_buf_1
X_0358_ _0057_ Tile_X0Y0_S1END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_65_66 VPWR VGND sg13g2_fill_2
XFILLER_45_135 VPWR VGND sg13g2_decap_8
X_1330_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1261_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1192_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_102 VPWR VGND sg13g2_decap_8
X_0976_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1528_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2 Tile_X0Y0_N1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1459_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_157 VPWR VGND sg13g2_decap_4
XFILLER_35_14 VPWR VGND sg13g2_fill_2
X_0830_ _0265_ VPWR _0266_ VGND _0000_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ sg13g2_o21ai_1
X_0692_ _0168_ VPWR ADDR_SRAM2 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
+ _0170_ sg13g2_o21ai_1
XFILLER_44_4 VPWR VGND sg13g2_fill_2
X_0761_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q VPWR
+ _0203_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
X_1313_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1244_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1175_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_138 VPWR VGND sg13g2_fill_2
XANTENNA_45 VPWR VGND Tile_X0Y0_S2MID[6] sg13g2_antennanp
XANTENNA_12 VPWR VGND Tile_X0Y0_S2MID[5] sg13g2_antennanp
XANTENNA_34 VPWR VGND Tile_X0Y1_N2MID[4] sg13g2_antennanp
XANTENNA_23 VPWR VGND Tile_X0Y1_FrameStrobe[17] sg13g2_antennanp
X_0959_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_38 VPWR VGND sg13g2_fill_2
XFILLER_101_198 VPWR VGND sg13g2_fill_2
XFILLER_46_24 VPWR VGND sg13g2_decap_4
XFILLER_46_46 VPWR VGND sg13g2_fill_1
XFILLER_2_0 VPWR VGND sg13g2_fill_2
X_0813_ Tile_X0Y1_E1END[3] Tile_X0Y1_EE4END[15] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ _0250_ VPWR VGND sg13g2_mux2_1
X_0675_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q DOUT_SRAM6
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ _0079_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6
+ VPWR VGND sg13g2_mux4_1
XFILLER_35_0 VPWR VGND sg13g2_decap_8
X_0744_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q VPWR
+ _0187_ VGND Tile_X0Y1_E6END[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ sg13g2_o21ai_1
X_1158_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1227_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1089_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_57_89 VPWR VGND sg13g2_decap_4
X_0460_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q DOUT_SRAM21
+ DOUT_SRAM24 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5
+ VPWR VGND sg13g2_mux4_1
XFILLER_93_177 VPWR VGND sg13g2_fill_1
X_1012_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0391_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q Tile_X0Y1_E2MID[6]
+ Tile_X0Y1_E2END[6] Tile_X0Y1_E6END[6] _0078_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 VPWR VGND sg13g2_mux4_1
XFILLER_93_199 VPWR VGND sg13g2_fill_1
X_0727_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y1_EE4END[2]
+ Tile_X0Y1_EE4END[10] Tile_X0Y1_E6END[10] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q BM_SRAM10
+ VPWR VGND sg13g2_mux4_1
X_0589_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
+ _0145_ VPWR VGND sg13g2_nor2b_1
X_0658_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q DOUT_SRAM6
+ DOUT_SRAM10 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 _0082_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10
+ VPWR VGND sg13g2_mux4_1
XFILLER_84_155 VPWR VGND sg13g2_decap_8
XFILLER_68_55 VPWR VGND sg13g2_fill_1
X_1630_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameData_O[19] VPWR VGND sg13g2_buf_1
X_1561_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3 Tile_X0Y0_N4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_0512_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y0_EE4END[3]
+ Tile_X0Y0_EE4END[11] Tile_X0Y0_E6END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q BM_SRAM19
+ VPWR VGND sg13g2_mux4_1
X_1492_ Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData_O[18] VPWR VGND sg13g2_buf_1
X_0443_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q DOUT_SRAM23
+ DOUT_SRAM31 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7
+ VPWR VGND sg13g2_mux4_1
XFILLER_3_170 VPWR VGND sg13g2_fill_2
X_0374_ VPWR VGND _0069_ _0068_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
+ _0008_ _0070_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ sg13g2_a221oi_1
XFILLER_66_199 VPWR VGND sg13g2_fill_1
XFILLER_79_76 VPWR VGND sg13g2_fill_2
XFILLER_48_177 VPWR VGND sg13g2_fill_2
XFILLER_48_199 VPWR VGND sg13g2_fill_1
XFILLER_63_169 VPWR VGND sg13g2_decap_4
X_0992_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1544_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6 Tile_X0Y0_N2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_1613_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameData_O[2] VPWR VGND sg13g2_buf_1
X_0426_ VPWR VGND _0085_ _0086_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ _0006_ _0087_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_a221oi_1
X_1475_ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData_O[1] VPWR VGND sg13g2_buf_1
X_0357_ VGND VPWR Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ _0052_ MEN_SRAM _0056_ sg13g2_a21oi_1
XFILLER_24_38 VPWR VGND sg13g2_decap_4
XFILLER_54_147 VPWR VGND sg13g2_fill_2
XFILLER_62_191 VPWR VGND sg13g2_decap_8
XFILLER_105_85 VPWR VGND sg13g2_fill_2
XFILLER_60_139 VPWR VGND sg13g2_decap_8
X_1191_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1260_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0975_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_0 VPWR VGND sg13g2_fill_2
X_1527_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1 Tile_X0Y0_N1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_0409_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_E2MID[2] Tile_X0Y0_E2END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5
+ VPWR VGND sg13g2_mux4_1
X_1389_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_103 VPWR VGND sg13g2_decap_8
XFILLER_27_114 VPWR VGND sg13g2_fill_1
X_1458_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_37 VPWR VGND sg13g2_fill_1
XFILLER_92_54 VPWR VGND sg13g2_fill_2
XFILLER_18_114 VPWR VGND sg13g2_decap_8
XFILLER_18_169 VPWR VGND sg13g2_fill_1
XFILLER_41_161 VPWR VGND sg13g2_decap_8
X_0760_ _0023_ _0079_ _0202_ VPWR VGND sg13g2_nor2_1
X_0691_ VGND VPWR Tile_X0Y1_E2END[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ _0170_ _0169_ sg13g2_a21oi_1
XFILLER_37_4 VPWR VGND sg13g2_fill_1
X_1174_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1312_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1243_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_13 VPWR VGND Tile_X0Y0_S2MID[5] sg13g2_antennanp
XANTENNA_24 VPWR VGND Tile_X0Y1_FrameStrobe[18] sg13g2_antennanp
XANTENNA_46 VPWR VGND Tile_X0Y1_FrameStrobe[15] sg13g2_antennanp
X_0889_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_35 VPWR VGND Tile_X0Y1_N2MID[5] sg13g2_antennanp
X_0958_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_80 VPWR VGND sg13g2_decap_4
X_0812_ _0248_ VPWR _0249_ VGND _0033_ _0158_ sg13g2_o21ai_1
X_0743_ VGND VPWR _0179_ _0181_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A _0186_ sg13g2_a21oi_1
XFILLER_96_153 VPWR VGND sg13g2_fill_1
X_0674_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q DOUT_SRAM5
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6
+ _0078_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5
+ VPWR VGND sg13g2_mux4_1
XFILLER_96_197 VPWR VGND sg13g2_fill_2
X_1157_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1226_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1088_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_73_67 VPWR VGND sg13g2_decap_8
XFILLER_73_45 VPWR VGND sg13g2_decap_4
XFILLER_73_23 VPWR VGND sg13g2_fill_1
XFILLER_11_197 VPWR VGND sg13g2_fill_2
X_0390_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q Tile_X0Y1_N2MID[1]
+ Tile_X0Y1_N2END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1
+ Tile_X0Y0_S2MID[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
+ _0078_ VPWR VGND sg13g2_mux4_1
XFILLER_93_112 VPWR VGND sg13g2_fill_2
XFILLER_78_197 VPWR VGND sg13g2_fill_2
X_1011_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_7 VPWR VGND sg13g2_fill_2
X_0726_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y1_EE4END[1]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_E6END[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q BM_SRAM9
+ VPWR VGND sg13g2_mux4_1
X_0588_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q _0144_ VPWR
+ VGND sg13g2_mux2_1
X_0657_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0060_ Tile_X0Y0_S4END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 VPWR VGND sg13g2_mux4_1
X_1209_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1560_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2 Tile_X0Y0_N4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_0511_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[10] Tile_X0Y0_E6END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q BM_SRAM18
+ VPWR VGND sg13g2_mux4_1
X_1491_ Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_66_112 VPWR VGND sg13g2_decap_8
X_0373_ _0069_ _0067_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_0442_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q DOUT_SRAM22
+ DOUT_SRAM30 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6
+ VPWR VGND sg13g2_mux4_1
X_1689_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 Tile_X0Y1_W2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_0709_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_EE4END[8] Tile_X0Y1_E6END[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q DIN_SRAM8
+ VPWR VGND sg13g2_mux4_1
XFILLER_72_104 VPWR VGND sg13g2_fill_2
XFILLER_70_13 VPWR VGND sg13g2_fill_1
XFILLER_0_174 VPWR VGND sg13g2_fill_1
XFILLER_0_196 VPWR VGND sg13g2_decap_4
XFILLER_63_115 VPWR VGND sg13g2_decap_8
X_0991_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1543_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5 Tile_X0Y0_N2BEGb[5]
+ VPWR VGND sg13g2_buf_1
X_1474_ Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData_O[0] VPWR VGND sg13g2_buf_1
X_1612_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData_O[1] VPWR VGND sg13g2_buf_1
X_0425_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0 _0086_ VPWR VGND sg13g2_nor3_1
X_0356_ CONFIGURED_top VPWR _0056_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ _0055_ sg13g2_o21ai_1
XFILLER_49_69 VPWR VGND sg13g2_decap_8
XFILLER_107_161 VPWR VGND sg13g2_fill_1
X_1190_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0974_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_105_109 VPWR VGND sg13g2_fill_1
X_1526_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0 Tile_X0Y0_N1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1457_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0339_ VPWR _0042_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ VGND sg13g2_inv_1
X_0408_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q Tile_X0Y0_E2MID[3]
+ Tile_X0Y0_E2END[3] Tile_X0Y0_E6END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4
+ VPWR VGND sg13g2_mux4_1
X_1388_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_104_120 VPWR VGND sg13g2_decap_8
X_0690_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q Tile_X0Y1_E2MID[2]
+ _0169_ VPWR VGND sg13g2_nor2b_1
X_1311_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_7 VPWR VGND sg13g2_decap_4
X_1173_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1242_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_25 VPWR VGND Tile_X0Y1_FrameStrobe[18] sg13g2_antennanp
XANTENNA_14 VPWR VGND Tile_X0Y0_S2MID[5] sg13g2_antennanp
XANTENNA_36 VPWR VGND Tile_X0Y1_N2MID[5] sg13g2_antennanp
XFILLER_32_195 VPWR VGND sg13g2_decap_4
X_0888_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0957_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1509_ Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
XFILLER_99_195 VPWR VGND sg13g2_fill_1
XFILLER_23_140 VPWR VGND sg13g2_decap_4
XFILLER_62_36 VPWR VGND sg13g2_fill_1
XFILLER_87_33 VPWR VGND sg13g2_decap_8
XFILLER_87_11 VPWR VGND sg13g2_fill_1
XFILLER_14_184 VPWR VGND sg13g2_decap_8
X_0673_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q DOUT_SRAM4
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7
+ _0043_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4
+ VPWR VGND sg13g2_mux4_1
X_0811_ VPWR _0248_ _0247_ VGND sg13g2_inv_1
X_0742_ VGND VPWR _0020_ _0184_ _0186_ _0185_ sg13g2_a21oi_1
X_1156_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1087_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1225_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_198 VPWR VGND sg13g2_fill_2
XFILLER_87_198 VPWR VGND sg13g2_fill_2
XFILLER_57_25 VPWR VGND sg13g2_fill_1
XFILLER_57_47 VPWR VGND sg13g2_decap_8
XFILLER_11_132 VPWR VGND sg13g2_decap_4
XFILLER_11_154 VPWR VGND sg13g2_decap_4
XFILLER_22_50 VPWR VGND sg13g2_decap_8
X_1010_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0656_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q DOUT_SRAM5
+ DOUT_SRAM9 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 _0083_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9
+ VPWR VGND sg13g2_mux4_1
X_0725_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_EE4END[8] Tile_X0Y1_E6END[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q BM_SRAM8
+ VPWR VGND sg13g2_mux4_1
XFILLER_40_0 VPWR VGND sg13g2_decap_4
X_0587_ _0141_ _0143_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1
+ VPWR VGND sg13g2_nor2_1
X_1208_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1139_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_4_128 VPWR VGND sg13g2_fill_2
XFILLER_84_67 VPWR VGND sg13g2_fill_2
XFILLER_17_72 VPWR VGND sg13g2_decap_4
XFILLER_33_60 VPWR VGND sg13g2_decap_4
X_1490_ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_3_172 VPWR VGND sg13g2_fill_1
X_0510_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q Tile_X0Y0_EE4END[1]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_E6END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q BM_SRAM17
+ VPWR VGND sg13g2_mux4_1
XFILLER_3_194 VPWR VGND sg13g2_decap_4
X_0372_ Tile_X0Y1_N1END[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q _0068_ VPWR
+ VGND sg13g2_nor3_1
X_0441_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q DOUT_SRAM21
+ DOUT_SRAM29 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_127 VPWR VGND sg13g2_decap_8
XFILLER_88_0 VPWR VGND sg13g2_decap_4
X_1688_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 Tile_X0Y1_W2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0639_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q DOUT_SRAM6
+ DOUT_SRAM14 _0078_ _0083_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6 VPWR VGND sg13g2_mux4_1
X_0708_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q Tile_X0Y1_EE4END[7]
+ Tile_X0Y1_EE4END[15] Tile_X0Y1_E6END[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q DIN_SRAM7
+ VPWR VGND sg13g2_mux4_1
XFILLER_72_138 VPWR VGND sg13g2_decap_8
XFILLER_38_49 VPWR VGND sg13g2_fill_2
XFILLER_57_168 VPWR VGND sg13g2_decap_4
XFILLER_110_65 VPWR VGND sg13g2_fill_2
XFILLER_79_78 VPWR VGND sg13g2_fill_1
XFILLER_95_99 VPWR VGND sg13g2_decap_8
XFILLER_48_135 VPWR VGND sg13g2_fill_1
XFILLER_71_171 VPWR VGND sg13g2_fill_1
XFILLER_48_179 VPWR VGND sg13g2_fill_1
X_1611_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData_O[0] VPWR VGND sg13g2_buf_1
X_0990_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1542_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 Tile_X0Y0_N2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_0424_ _0085_ Tile_X0Y0_S1END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
X_1473_ clknet_1_0__leaf_Tile_X0Y1_UserCLK CLK_SRAM VPWR VGND sg13g2_buf_1
X_0355_ _0054_ _0053_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0055_ VPWR VGND sg13g2_mux2_1
XFILLER_54_149 VPWR VGND sg13g2_fill_1
XFILLER_105_54 VPWR VGND sg13g2_fill_2
XFILLER_105_21 VPWR VGND sg13g2_fill_1
XFILLER_105_87 VPWR VGND sg13g2_fill_1
XFILLER_45_105 VPWR VGND sg13g2_decap_8
XFILLER_45_149 VPWR VGND sg13g2_fill_1
XFILLER_30_72 VPWR VGND sg13g2_fill_1
XFILLER_30_94 VPWR VGND sg13g2_fill_2
XFILLER_44_171 VPWR VGND sg13g2_fill_1
XFILLER_44_193 VPWR VGND sg13g2_decap_8
X_0973_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_2 VPWR VGND sg13g2_fill_1
X_1525_ Tile_X0Y1_FrameStrobe[19] Tile_X0Y0_FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_0407_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4
+ Tile_X0Y0_S2MID[4] Tile_X0Y1_N2MID[4] Tile_X0Y0_S2END[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4 VPWR VGND sg13g2_mux4_1
X_1387_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1456_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0338_ VPWR _0041_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3
+ VGND sg13g2_inv_1
XFILLER_42_119 VPWR VGND sg13g2_decap_8
XFILLER_50_141 VPWR VGND sg13g2_decap_8
XFILLER_50_174 VPWR VGND sg13g2_decap_4
XFILLER_104_198 VPWR VGND sg13g2_fill_2
XFILLER_110_113 VPWR VGND sg13g2_fill_2
X_1310_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1241_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1172_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_15 VPWR VGND Tile_X0Y1_FrameStrobe[10] sg13g2_antennanp
XANTENNA_26 VPWR VGND Tile_X0Y1_FrameStrobe[18] sg13g2_antennanp
X_0956_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_0 VPWR VGND sg13g2_fill_2
XANTENNA_37 VPWR VGND Tile_X0Y1_N2MID[7] sg13g2_antennanp
X_0887_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1508_ Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
X_1439_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_174 VPWR VGND sg13g2_decap_4
X_0810_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q VPWR
+ _0247_ VGND Tile_X0Y1_E6END[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ sg13g2_o21ai_1
X_0672_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q Tile_X0Y1_N4END[3]
+ Tile_X0Y0_S4END[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3 VPWR VGND sg13g2_mux4_1
X_0741_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q VPWR
+ _0185_ VGND _0182_ _0183_ sg13g2_o21ai_1
XFILLER_96_199 VPWR VGND sg13g2_fill_1
X_1224_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1155_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1086_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0939_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_11_199 VPWR VGND sg13g2_fill_1
XFILLER_78_199 VPWR VGND sg13g2_fill_1
XFILLER_0_0 VPWR VGND sg13g2_fill_1
XFILLER_21_9 VPWR VGND sg13g2_fill_1
XFILLER_47_70 VPWR VGND sg13g2_fill_2
X_0586_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q _0142_
+ _0143_ VPWR VGND sg13g2_nor2_1
X_0655_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0067_ Tile_X0Y0_S4END[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 VPWR VGND sg13g2_mux4_1
X_0724_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q Tile_X0Y1_EE4END[7]
+ Tile_X0Y1_EE4END[15] Tile_X0Y1_E6END[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q BM_SRAM7
+ VPWR VGND sg13g2_mux4_1
XFILLER_84_136 VPWR VGND sg13g2_fill_2
XFILLER_69_199 VPWR VGND sg13g2_fill_1
XFILLER_69_177 VPWR VGND sg13g2_fill_1
X_1207_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1138_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1069_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_43 VPWR VGND sg13g2_fill_1
XFILLER_83_191 VPWR VGND sg13g2_fill_2
X_0440_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q DOUT_SRAM20
+ DOUT_SRAM28 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4
+ VPWR VGND sg13g2_mux4_1
X_0371_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14
+ _0066_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q _0067_
+ VPWR VGND sg13g2_mux4_1
XFILLER_58_91 VPWR VGND sg13g2_fill_1
X_0707_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y1_EE4END[6]
+ Tile_X0Y1_EE4END[14] Tile_X0Y1_E6END[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q DIN_SRAM6
+ VPWR VGND sg13g2_mux4_1
X_0569_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E6END[11] Tile_X0Y0_EE4END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q _0128_ VPWR
+ VGND sg13g2_mux4_1
X_0638_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q DOUT_SRAM5
+ DOUT_SRAM13 _0079_ _0082_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5 VPWR VGND sg13g2_mux4_1
X_1687_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4 Tile_X0Y1_W2BEG[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_56_180 VPWR VGND sg13g2_fill_1
X_1610_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15 Tile_X0Y0_WW4BEG[15]
+ VPWR VGND sg13g2_buf_1
XFILLER_60_92 VPWR VGND sg13g2_decap_8
X_1541_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 Tile_X0Y0_N2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_0423_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2END[0] Tile_X0Y0_E6END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7
+ VPWR VGND sg13g2_mux4_1
X_1472_ VPWR VGND TIE_LOW_SRAM sg13g2_tielo
X_0354_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_N2MID[6]
+ Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3] Tile_X0Y1_E2MID[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0054_ VPWR VGND sg13g2_mux4_1
XFILLER_14_96 VPWR VGND sg13g2_fill_1
XFILLER_100_0 VPWR VGND sg13g2_fill_1
XFILLER_39_71 VPWR VGND sg13g2_fill_2
X_0972_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1524_ Tile_X0Y1_FrameStrobe[18] Tile_X0Y0_FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_0337_ VPWR _0040_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2
+ VGND sg13g2_inv_1
X_1386_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1455_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0406_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q Tile_X0Y1_E2MID[3]
+ Tile_X0Y1_E2END[3] Tile_X0Y1_E6END[3] _0081_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4 VPWR VGND sg13g2_mux4_1
XFILLER_25_95 VPWR VGND sg13g2_decap_4
X_1171_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1240_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_38 VPWR VGND Tile_X0Y1_N2MID[7] sg13g2_antennanp
XANTENNA_27 VPWR VGND Tile_X0Y1_FrameStrobe[19] sg13g2_antennanp
X_0886_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_16 VPWR VGND Tile_X0Y1_FrameStrobe[11] sg13g2_antennanp
X_0955_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1507_ Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
XFILLER_99_131 VPWR VGND sg13g2_fill_2
XFILLER_63_0 VPWR VGND sg13g2_fill_2
X_1369_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_46_17 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_fill_1
X_1438_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0740_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q _0184_ VPWR
+ VGND sg13g2_mux2_1
X_0671_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q Tile_X0Y1_N4END[2]
+ Tile_X0Y0_S4END[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2 VPWR VGND sg13g2_mux4_1
X_1154_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_134 VPWR VGND sg13g2_fill_2
X_1223_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1085_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0938_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0869_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_87_134 VPWR VGND sg13g2_fill_2
XFILLER_7_105 VPWR VGND sg13g2_decap_8
XFILLER_6_160 VPWR VGND sg13g2_fill_1
X_0723_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y1_EE4END[6]
+ Tile_X0Y1_EE4END[14] Tile_X0Y1_E6END[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q BM_SRAM6 VPWR
+ VGND sg13g2_mux4_1
X_0585_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_E6END[5] Tile_X0Y0_EE4END[13] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q _0142_ VPWR
+ VGND sg13g2_mux4_1
X_0654_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q DOUT_SRAM4
+ DOUT_SRAM8 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 _0084_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8
+ VPWR VGND sg13g2_mux4_1
X_1137_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_84_115 VPWR VGND sg13g2_decap_4
X_1206_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1068_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_77 VPWR VGND sg13g2_fill_1
XFILLER_68_48 VPWR VGND sg13g2_decap_8
X_0370_ VPWR VGND _0064_ _0065_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ _0004_ _0066_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ sg13g2_a221oi_1
XFILLER_66_137 VPWR VGND sg13g2_fill_1
X_1686_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3 Tile_X0Y1_W2BEG[3]
+ VPWR VGND sg13g2_buf_1
X_0706_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q Tile_X0Y1_EE4END[5]
+ Tile_X0Y1_EE4END[13] Tile_X0Y1_E6END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q DIN_SRAM5
+ VPWR VGND sg13g2_mux4_1
X_0568_ VGND VPWR _0014_ _0123_ _0127_ _0126_ sg13g2_a21oi_1
X_0499_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q Tile_X0Y0_EE4END[6]
+ Tile_X0Y0_EE4END[14] Tile_X0Y0_E6END[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q DIN_SRAM22
+ VPWR VGND sg13g2_mux4_1
X_0637_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q DOUT_SRAM4
+ DOUT_SRAM12 _0080_ _0081_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4 VPWR VGND sg13g2_mux4_1
XFILLER_79_58 VPWR VGND sg13g2_fill_1
XFILLER_95_46 VPWR VGND sg13g2_decap_4
XFILLER_95_24 VPWR VGND sg13g2_fill_1
XFILLER_28_95 VPWR VGND sg13g2_fill_2
X_1540_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2 Tile_X0Y0_N2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_0422_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7
+ Tile_X0Y0_S2MID[7] Tile_X0Y1_N2MID[7] Tile_X0Y0_S2END[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 VPWR VGND sg13g2_mux4_1
X_1471_ VPWR VGND TIE_HIGH_SRAM sg13g2_tiehi
X_0353_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_E2MID[3]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0053_ VPWR VGND sg13g2_mux4_1
XFILLER_47_170 VPWR VGND sg13g2_decap_8
XFILLER_93_0 VPWR VGND sg13g2_fill_2
X_1669_ Tile_X0Y0_S4END[14] Tile_X0Y1_S4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_49_17 VPWR VGND sg13g2_fill_1
XFILLER_38_192 VPWR VGND sg13g2_decap_8
XFILLER_29_181 VPWR VGND sg13g2_fill_1
X_0971_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_70 VPWR VGND sg13g2_decap_4
X_1523_ Tile_X0Y1_FrameStrobe[17] Tile_X0Y0_FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_1454_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0336_ VPWR _0039_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1
+ VGND sg13g2_inv_1
X_1385_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0405_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y1_N2MID[4]
+ Tile_X0Y1_N2END[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4
+ Tile_X0Y0_S2MID[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
+ _0081_ VPWR VGND sg13g2_mux4_1
XFILLER_41_95 VPWR VGND sg13g2_decap_4
X_1170_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_17_162 VPWR VGND sg13g2_decap_8
XANTENNA_17 VPWR VGND Tile_X0Y1_FrameStrobe[12] sg13g2_antennanp
X_0885_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0954_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_2 VPWR VGND sg13g2_fill_1
XANTENNA_39 VPWR VGND Tile_X0Y1_N2MID[7] sg13g2_antennanp
XANTENNA_28 VPWR VGND Tile_X0Y1_N2MID[0] sg13g2_antennanp
X_1506_ Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
XFILLER_101_126 VPWR VGND sg13g2_fill_1
XFILLER_99_110 VPWR VGND sg13g2_decap_4
X_1437_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_0 VPWR VGND sg13g2_decap_8
XFILLER_101_148 VPWR VGND sg13g2_fill_1
X_1368_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1299_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0319_ VPWR _0022_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
+ VGND sg13g2_inv_1
XFILLER_11_87 VPWR VGND sg13g2_fill_2
XFILLER_11_43 VPWR VGND sg13g2_fill_2
XFILLER_87_58 VPWR VGND sg13g2_fill_1
XFILLER_36_73 VPWR VGND sg13g2_decap_8
XFILLER_36_84 VPWR VGND sg13g2_fill_1
XFILLER_14_198 VPWR VGND sg13g2_fill_2
X_0670_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q Tile_X0Y1_N4END[1]
+ Tile_X0Y0_S4END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1 VPWR VGND sg13g2_mux4_1
X_1153_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_157 VPWR VGND sg13g2_decap_4
X_1222_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1084_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0937_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0868_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0799_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q VPWR
+ _0237_ VGND Tile_X0Y1_E6END[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
+ sg13g2_o21ai_1
XFILLER_87_157 VPWR VGND sg13g2_fill_2
XFILLER_73_49 VPWR VGND sg13g2_fill_1
XFILLER_22_31 VPWR VGND sg13g2_fill_2
XFILLER_78_157 VPWR VGND sg13g2_fill_2
XFILLER_47_72 VPWR VGND sg13g2_fill_1
XFILLER_47_94 VPWR VGND sg13g2_decap_4
X_0653_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0074_ Tile_X0Y0_S4END[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 VPWR VGND sg13g2_mux4_1
X_0722_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q Tile_X0Y1_EE4END[5]
+ Tile_X0Y1_EE4END[13] Tile_X0Y1_E6END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q BM_SRAM5 VPWR
+ VGND sg13g2_mux4_1
X_0584_ VGND VPWR _0016_ _0137_ _0141_ _0140_ sg13g2_a21oi_1
X_1136_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1205_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1067_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_17_97 VPWR VGND sg13g2_decap_4
X_1685_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2 Tile_X0Y1_W2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0636_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q DOUT_SRAM3
+ DOUT_SRAM11 _0080_ _0081_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3 VPWR VGND sg13g2_mux4_1
X_0705_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_E6END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q DIN_SRAM4
+ VPWR VGND sg13g2_mux4_1
X_0567_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q VPWR
+ _0126_ VGND _0124_ _0125_ sg13g2_o21ai_1
X_0498_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q Tile_X0Y0_EE4END[5]
+ Tile_X0Y0_EE4END[13] Tile_X0Y0_E6END[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q DIN_SRAM21
+ VPWR VGND sg13g2_mux4_1
X_1119_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_174 VPWR VGND sg13g2_fill_2
X_1470_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_70 VPWR VGND sg13g2_fill_2
X_0421_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2END[0] Tile_X0Y1_E6END[0] _0084_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7 VPWR VGND sg13g2_mux4_1
X_0352_ _0047_ VPWR _0052_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0051_ sg13g2_o21ai_1
XFILLER_86_0 VPWR VGND sg13g2_fill_2
X_1668_ Tile_X0Y0_S4END[13] Tile_X0Y1_S4BEG[5] VPWR VGND sg13g2_buf_1
X_1599_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4 Tile_X0Y0_WW4BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0619_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2END[1] _0083_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_81_49 VPWR VGND sg13g2_decap_4
XFILLER_53_152 VPWR VGND sg13g2_fill_1
XFILLER_107_198 VPWR VGND sg13g2_fill_2
X_0970_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1522_ Tile_X0Y1_FrameStrobe[16] Tile_X0Y0_FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
X_0404_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_E2END[3] Tile_X0Y0_E2MID[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4
+ VPWR VGND sg13g2_mux4_1
X_1453_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0335_ VPWR _0038_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0
+ VGND sg13g2_inv_1
X_1384_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_50_155 VPWR VGND sg13g2_fill_2
XFILLER_50_199 VPWR VGND sg13g2_fill_1
XFILLER_26_152 VPWR VGND sg13g2_fill_2
XFILLER_26_174 VPWR VGND sg13g2_decap_4
XFILLER_41_199 VPWR VGND sg13g2_fill_1
XFILLER_66_93 VPWR VGND sg13g2_fill_2
XANTENNA_18 VPWR VGND Tile_X0Y1_FrameStrobe[13] sg13g2_antennanp
XFILLER_82_70 VPWR VGND sg13g2_fill_1
XANTENNA_29 VPWR VGND Tile_X0Y1_N2MID[0] sg13g2_antennanp
XFILLER_32_199 VPWR VGND sg13g2_fill_1
X_0953_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0884_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_2 VPWR VGND sg13g2_fill_1
XFILLER_99_155 VPWR VGND sg13g2_fill_1
X_1505_ Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData_O[31] VPWR VGND sg13g2_buf_1
X_1367_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1436_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1298_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0318_ VPWR _0021_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
+ VGND sg13g2_inv_1
XFILLER_14_166 VPWR VGND sg13g2_fill_1
X_1221_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1152_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1083_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0936_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_114 VPWR VGND sg13g2_decap_4
XFILLER_20_147 VPWR VGND sg13g2_fill_1
X_0867_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0798_ VGND VPWR _0229_ _0231_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1
+ _0236_ sg13g2_a21oi_1
X_1419_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_11_158 VPWR VGND sg13g2_fill_1
XFILLER_11_136 VPWR VGND sg13g2_fill_1
X_0583_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q VPWR
+ _0140_ VGND _0138_ _0139_ sg13g2_o21ai_1
XFILLER_10_180 VPWR VGND sg13g2_fill_2
X_0652_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q DOUT_SRAM7
+ DOUT_SRAM11 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 _0043_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7
+ VPWR VGND sg13g2_mux4_1
X_0721_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q Tile_X0Y1_EE4END[4]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_E6END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q BM_SRAM4 VPWR
+ VGND sg13g2_mux4_1
X_1204_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1135_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1066_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0919_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_128 VPWR VGND sg13g2_decap_4
XFILLER_3_198 VPWR VGND sg13g2_fill_2
XFILLER_58_50 VPWR VGND sg13g2_fill_1
XFILLER_88_4 VPWR VGND sg13g2_fill_2
X_0566_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q VPWR
+ _0125_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
X_0635_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q DOUT_SRAM2
+ DOUT_SRAM10 _0079_ _0082_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2 VPWR VGND sg13g2_mux4_1
X_1684_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1 Tile_X0Y1_W2BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_31_0 VPWR VGND sg13g2_decap_4
X_0704_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q Tile_X0Y1_EE4END[3]
+ Tile_X0Y1_EE4END[11] Tile_X0Y1_E6END[3] _0158_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
+ DIN_SRAM3 VPWR VGND sg13g2_mux4_1
X_0497_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_E6END[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q DIN_SRAM20
+ VPWR VGND sg13g2_mux4_1
XFILLER_57_139 VPWR VGND sg13g2_decap_4
X_1118_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_197 VPWR VGND sg13g2_fill_2
X_1049_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_131 VPWR VGND sg13g2_decap_4
XFILLER_28_64 VPWR VGND sg13g2_fill_2
XFILLER_71_197 VPWR VGND sg13g2_fill_2
X_0420_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q Tile_X0Y1_N2MID[7]
+ Tile_X0Y1_N2END[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7
+ Tile_X0Y0_S2MID[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
+ _0084_ VPWR VGND sg13g2_mux4_1
X_0351_ _0050_ VPWR _0051_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0049_ sg13g2_o21ai_1
XFILLER_79_0 VPWR VGND sg13g2_fill_2
X_1667_ Tile_X0Y0_S4END[12] Tile_X0Y1_S4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_105_25 VPWR VGND sg13g2_fill_1
X_1598_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3 Tile_X0Y0_WW4BEG[3]
+ VPWR VGND sg13g2_buf_1
X_0549_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ _0110_ VPWR VGND sg13g2_nor2b_1
X_0618_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_E2MID[2] Tile_X0Y1_E2END[2] _0082_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_53_120 VPWR VGND sg13g2_decap_4
XFILLER_36_109 VPWR VGND sg13g2_decap_8
XFILLER_55_40 VPWR VGND sg13g2_fill_2
X_0403_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q Tile_X0Y0_E2MID[4]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E6END[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3
+ VPWR VGND sg13g2_mux4_1
X_1521_ Tile_X0Y1_FrameStrobe[15] Tile_X0Y0_FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_1383_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1452_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0334_ VPWR _0037_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
+ VGND sg13g2_inv_1
X_1719_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8 Tile_X0Y1_WW4BEG[8]
+ VPWR VGND sg13g2_buf_1
XFILLER_26_197 VPWR VGND sg13g2_fill_2
XFILLER_41_42 VPWR VGND sg13g2_fill_2
XFILLER_41_64 VPWR VGND sg13g2_fill_2
XFILLER_66_72 VPWR VGND sg13g2_decap_4
XANTENNA_19 VPWR VGND Tile_X0Y1_FrameStrobe[14] sg13g2_antennanp
X_0952_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0883_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1504_ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData_O[30] VPWR VGND sg13g2_buf_1
X_1366_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0317_ VPWR _0020_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q
+ VGND sg13g2_inv_1
X_1435_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_101 VPWR VGND sg13g2_fill_1
X_1297_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_178 VPWR VGND sg13g2_fill_1
XFILLER_11_89 VPWR VGND sg13g2_fill_1
XFILLER_11_45 VPWR VGND sg13g2_fill_1
X_1151_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_7 VPWR VGND sg13g2_decap_8
X_1220_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1082_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0866_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0935_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0797_ VGND VPWR _0030_ _0234_ _0236_ _0235_ sg13g2_a21oi_1
XFILLER_61_0 VPWR VGND sg13g2_fill_2
XFILLER_87_159 VPWR VGND sg13g2_fill_1
X_1349_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1418_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_22_99 VPWR VGND sg13g2_decap_8
XFILLER_78_159 VPWR VGND sg13g2_fill_1
X_0720_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q Tile_X0Y1_EE4END[3]
+ Tile_X0Y1_EE4END[11] Tile_X0Y1_E6END[3] _0158_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
+ BM_SRAM3 VPWR VGND sg13g2_mux4_1
X_0582_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q VPWR
+ _0139_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
X_0651_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0088_ Tile_X0Y0_S4END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8 VPWR VGND sg13g2_mux4_1
X_1134_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1203_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_173 VPWR VGND sg13g2_decap_8
X_1065_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0918_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0849_ _0284_ Tile_X0Y1_E2MID[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_109_0 VPWR VGND sg13g2_fill_1
XFILLER_74_50 VPWR VGND sg13g2_fill_1
X_1683_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0 Tile_X0Y1_W2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0703_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y1_EE4END[2]
+ Tile_X0Y1_EE4END[10] Tile_X0Y1_E6END[2] _0159_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
+ DIN_SRAM2 VPWR VGND sg13g2_mux4_1
X_0565_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
+ _0124_ VPWR VGND sg13g2_nor2b_1
X_0496_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q Tile_X0Y0_EE4END[3]
+ Tile_X0Y0_EE4END[11] Tile_X0Y0_E6END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q DIN_SRAM19
+ VPWR VGND sg13g2_mux4_1
X_0634_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q DOUT_SRAM1
+ DOUT_SRAM9 _0078_ _0083_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1 VPWR VGND sg13g2_mux4_1
X_1117_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1048_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_162 VPWR VGND sg13g2_decap_8
Xclkbuf_1_0__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_0__leaf_Tile_X0Y1_UserCLK
+ VPWR VGND sg13g2_buf_8
XFILLER_69_72 VPWR VGND sg13g2_fill_1
X_0350_ Tile_X0Y1_E2END[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0050_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
+ sg13g2_nand3b_1
XFILLER_47_140 VPWR VGND sg13g2_decap_8
XFILLER_62_198 VPWR VGND sg13g2_fill_2
X_1666_ Tile_X0Y0_S4END[11] Tile_X0Y1_S4BEG[3] VPWR VGND sg13g2_buf_1
X_0479_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0 VPWR VGND sg13g2_mux4_1
X_0548_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q _0109_ VPWR
+ VGND sg13g2_mux2_1
X_0617_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_E2END[3] Tile_X0Y1_E2MID[3] _0081_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4 VPWR VGND sg13g2_mux4_1
X_1597_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2 Tile_X0Y0_WW4BEG[2]
+ VPWR VGND sg13g2_buf_1
XFILLER_81_18 VPWR VGND sg13g2_fill_2
X_1520_ Tile_X0Y1_FrameStrobe[14] Tile_X0Y0_FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
X_0402_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3
+ Tile_X0Y1_N2MID[3] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 VPWR VGND sg13g2_mux4_1
X_1382_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1451_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0333_ VPWR _0036_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
+ VGND sg13g2_inv_1
X_1649_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 Tile_X0Y1_S2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1718_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7 Tile_X0Y1_WW4BEG[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_92_17 VPWR VGND sg13g2_fill_2
XFILLER_25_77 VPWR VGND sg13g2_fill_1
XFILLER_25_99 VPWR VGND sg13g2_fill_1
XFILLER_41_168 VPWR VGND sg13g2_fill_2
XFILLER_17_176 VPWR VGND sg13g2_fill_2
X_0882_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0951_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1503_ Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData_O[29] VPWR VGND sg13g2_buf_1
X_1365_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1434_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0316_ VPWR _0019_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ VGND sg13g2_inv_1
X_1296_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_173 VPWR VGND sg13g2_fill_1
X_1150_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_77_50 VPWR VGND sg13g2_fill_2
X_1081_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0865_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0934_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_194 VPWR VGND sg13g2_decap_4
XFILLER_9_172 VPWR VGND sg13g2_fill_1
XFILLER_87_127 VPWR VGND sg13g2_decap_8
X_1417_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0796_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q VPWR
+ _0235_ VGND _0232_ _0233_ sg13g2_o21ai_1
XFILLER_95_171 VPWR VGND sg13g2_decap_8
X_1348_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1279_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_6_153 VPWR VGND sg13g2_decap_8
X_0581_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
+ _0138_ VPWR VGND sg13g2_nor2b_1
X_0650_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q DOUT_SRAM6
+ DOUT_SRAM10 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9 _0078_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6
+ VPWR VGND sg13g2_mux4_1
XFILLER_77_160 VPWR VGND sg13g2_decap_4
X_1064_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1133_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1202_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0917_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0779_ _0218_ VPWR _0219_ VGND _0027_ _0161_ sg13g2_o21ai_1
X_0848_ _0283_ _0037_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_nand2_1
XFILLER_17_45 VPWR VGND sg13g2_decap_4
XFILLER_3_134 VPWR VGND sg13g2_fill_2
XFILLER_66_119 VPWR VGND sg13g2_fill_1
XFILLER_99_92 VPWR VGND sg13g2_fill_1
XFILLER_99_81 VPWR VGND sg13g2_decap_8
X_1682_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3 Tile_X0Y1_W1BEG[3]
+ VPWR VGND sg13g2_buf_1
X_0633_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q DOUT_SRAM0
+ DOUT_SRAM8 _0043_ _0084_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0 VPWR VGND sg13g2_mux4_1
X_0702_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q Tile_X0Y1_EE4END[1]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_E6END[1] _0160_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
+ DIN_SRAM1 VPWR VGND sg13g2_mux4_1
X_0564_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q _0123_ VPWR
+ VGND sg13g2_mux2_1
X_0495_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[10] Tile_X0Y0_E6END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q DIN_SRAM18
+ VPWR VGND sg13g2_mux4_1
X_1116_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1047_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_199 VPWR VGND sg13g2_fill_1
XFILLER_95_17 VPWR VGND sg13g2_decap_8
XFILLER_28_66 VPWR VGND sg13g2_fill_1
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_56_130 VPWR VGND sg13g2_fill_1
XFILLER_71_199 VPWR VGND sg13g2_fill_1
XFILLER_44_65 VPWR VGND sg13g2_fill_1
XFILLER_79_2 VPWR VGND sg13g2_fill_1
X_1665_ Tile_X0Y0_S4END[10] Tile_X0Y1_S4BEG[2] VPWR VGND sg13g2_buf_1
X_1596_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1 Tile_X0Y0_WW4BEG[1]
+ VPWR VGND sg13g2_buf_1
X_0616_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q Tile_X0Y1_E2MID[4]
+ Tile_X0Y1_E6END[11] Tile_X0Y1_E2END[4] _0080_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3 VPWR VGND sg13g2_mux4_1
X_0547_ _0106_ _0108_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0
+ VPWR VGND sg13g2_nor2_1
X_0478_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q DOUT_SRAM18
+ DOUT_SRAM30 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14
+ VPWR VGND sg13g2_mux4_1
XFILLER_14_68 VPWR VGND sg13g2_decap_8
XFILLER_107_179 VPWR VGND sg13g2_fill_2
XFILLER_44_111 VPWR VGND sg13g2_decap_4
XFILLER_71_74 VPWR VGND sg13g2_fill_1
XFILLER_71_41 VPWR VGND sg13g2_decap_8
X_1450_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1381_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0401_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q Tile_X0Y1_E2MID[4]
+ Tile_X0Y1_E6END[4] Tile_X0Y1_E2END[4] _0080_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3 VPWR VGND sg13g2_mux4_1
X_0332_ VPWR _0035_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ VGND sg13g2_inv_1
XFILLER_84_0 VPWR VGND sg13g2_decap_8
XFILLER_104_127 VPWR VGND sg13g2_fill_2
X_1579_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4 Tile_X0Y0_W2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_1717_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6 Tile_X0Y1_WW4BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1648_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 Tile_X0Y1_S2BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_26_199 VPWR VGND sg13g2_fill_1
XFILLER_41_66 VPWR VGND sg13g2_fill_1
XFILLER_17_199 VPWR VGND sg13g2_fill_1
X_0881_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0950_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_119 VPWR VGND sg13g2_decap_8
X_1502_ Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData_O[28] VPWR VGND sg13g2_buf_1
X_1433_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0315_ VPWR _0018_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
+ VGND sg13g2_inv_1
X_1364_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1295_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_136 VPWR VGND sg13g2_fill_2
XFILLER_77_73 VPWR VGND sg13g2_fill_1
X_1080_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0864_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0933_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0795_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q _0234_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_61_2 VPWR VGND sg13g2_fill_1
X_1347_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1416_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1278_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_22_24 VPWR VGND sg13g2_decap_8
XFILLER_22_57 VPWR VGND sg13g2_decap_4
XFILLER_78_117 VPWR VGND sg13g2_fill_2
XFILLER_47_98 VPWR VGND sg13g2_fill_2
XFILLER_63_97 VPWR VGND sg13g2_fill_1
X_0580_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q _0137_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_69_128 VPWR VGND sg13g2_fill_1
X_1201_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_197 VPWR VGND sg13g2_fill_2
X_1063_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1132_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0916_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0778_ VPWR _0218_ _0217_ VGND sg13g2_inv_1
X_0847_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0281_ _0282_ VPWR VGND sg13g2_nor3_1
XFILLER_83_197 VPWR VGND sg13g2_fill_2
XFILLER_83_153 VPWR VGND sg13g2_decap_4
XFILLER_74_197 VPWR VGND sg13g2_fill_2
XFILLER_90_84 VPWR VGND sg13g2_fill_2
XFILLER_90_73 VPWR VGND sg13g2_fill_2
XFILLER_90_51 VPWR VGND sg13g2_fill_1
X_0563_ _0120_ _0122_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2
+ VPWR VGND sg13g2_nor2_1
X_1681_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2 Tile_X0Y1_W1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0632_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q DOUT_SRAM7
+ DOUT_SRAM15 _0043_ _0084_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7 VPWR VGND sg13g2_mux4_1
X_0701_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_EE4END[8] Tile_X0Y1_E6END[0] _0161_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
+ DIN_SRAM0 VPWR VGND sg13g2_mux4_1
X_0494_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q Tile_X0Y0_EE4END[1]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_E6END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q DIN_SRAM17
+ VPWR VGND sg13g2_mux4_1
X_1115_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_123 VPWR VGND sg13g2_fill_2
XFILLER_80_101 VPWR VGND sg13g2_fill_1
X_1046_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_197 VPWR VGND sg13g2_fill_2
XFILLER_28_34 VPWR VGND sg13g2_fill_2
XFILLER_56_120 VPWR VGND sg13g2_decap_4
XFILLER_56_197 VPWR VGND sg13g2_fill_2
XFILLER_71_167 VPWR VGND sg13g2_decap_4
XFILLER_69_63 VPWR VGND sg13g2_decap_8
X_1664_ Tile_X0Y0_S4END[9] Tile_X0Y1_S4BEG[1] VPWR VGND sg13g2_buf_1
X_0546_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q _0107_
+ _0108_ VPWR VGND sg13g2_nor2_1
X_0615_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E2END[5] _0079_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2 VPWR VGND sg13g2_mux4_1
X_1595_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0 Tile_X0Y0_WW4BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0477_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1 VPWR VGND sg13g2_mux4_1
X_1029_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_53_134 VPWR VGND sg13g2_fill_1
XFILLER_107_136 VPWR VGND sg13g2_fill_1
XFILLER_44_167 VPWR VGND sg13g2_decap_4
X_1380_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0400_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q Tile_X0Y1_N2MID[3]
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3 Tile_X0Y1_N2END[3]
+ Tile_X0Y0_S2MID[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
+ _0080_ VPWR VGND sg13g2_mux4_1
X_0331_ VPWR _0034_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
+ VGND sg13g2_inv_1
XFILLER_35_123 VPWR VGND sg13g2_fill_2
XFILLER_50_148 VPWR VGND sg13g2_decap_8
X_1716_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5 Tile_X0Y1_WW4BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0529_ _0095_ Tile_X0Y0_E2END[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_nand2b_1
X_1578_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3 Tile_X0Y0_W2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_1647_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 Tile_X0Y1_S2BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_92_19 VPWR VGND sg13g2_fill_1
XFILLER_25_24 VPWR VGND sg13g2_fill_2
XFILLER_26_167 VPWR VGND sg13g2_decap_8
XFILLER_26_178 VPWR VGND sg13g2_fill_2
XFILLER_41_137 VPWR VGND sg13g2_decap_8
XFILLER_66_53 VPWR VGND sg13g2_fill_2
XFILLER_17_101 VPWR VGND sg13g2_fill_2
XFILLER_32_159 VPWR VGND sg13g2_fill_2
X_0880_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1501_ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData_O[27] VPWR VGND sg13g2_buf_1
X_1363_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1432_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0314_ VPWR _0017_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
+ VGND sg13g2_inv_1
X_1294_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_120 VPWR VGND sg13g2_decap_8
XFILLER_98_181 VPWR VGND sg13g2_decap_8
XFILLER_14_159 VPWR VGND sg13g2_decap_8
XFILLER_52_44 VPWR VGND sg13g2_fill_2
XFILLER_89_170 VPWR VGND sg13g2_decap_8
X_0932_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_118 VPWR VGND sg13g2_fill_1
X_0863_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0794_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q VPWR
+ _0233_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
X_1346_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1415_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1277_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_86_195 VPWR VGND sg13g2_decap_4
XFILLER_10_140 VPWR VGND sg13g2_fill_2
XFILLER_6_199 VPWR VGND sg13g2_fill_1
X_1200_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_110 VPWR VGND sg13g2_fill_2
X_1062_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1131_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_0915_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0777_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q VPWR
+ _0217_ VGND Tile_X0Y1_E6END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ sg13g2_o21ai_1
X_0846_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_N2MID[6]
+ _0281_ VPWR VGND sg13g2_nor2b_1
X_1329_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_136 VPWR VGND sg13g2_fill_1
XFILLER_59_151 VPWR VGND sg13g2_fill_1
X_0700_ _0174_ VPWR ADDR_SRAM4 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
+ _0176_ sg13g2_o21ai_1
X_0562_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q _0121_
+ _0122_ VPWR VGND sg13g2_nor2_1
X_0631_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q DOUT_SRAM6
+ DOUT_SRAM14 _0078_ _0083_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6 VPWR VGND sg13g2_mux4_1
X_1680_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1 Tile_X0Y1_W1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1114_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0493_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[8] Tile_X0Y0_E6END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q DIN_SRAM16
+ VPWR VGND sg13g2_mux4_1
XFILLER_80_146 VPWR VGND sg13g2_decap_8
X_1045_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0829_ VGND VPWR Tile_X0Y1_E2MID[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ _0265_ _0258_ sg13g2_a21oi_1
XFILLER_71_135 VPWR VGND sg13g2_fill_1
XFILLER_28_57 VPWR VGND sg13g2_decap_8
XFILLER_44_23 VPWR VGND sg13g2_decap_4
XFILLER_100_95 VPWR VGND sg13g2_decap_8
XFILLER_60_99 VPWR VGND sg13g2_fill_2
XFILLER_47_198 VPWR VGND sg13g2_fill_2
X_1663_ Tile_X0Y0_S4END[8] Tile_X0Y1_S4BEG[0] VPWR VGND sg13g2_buf_1
X_0545_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_EE4END[0] Tile_X0Y0_E6END[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q _0107_ VPWR
+ VGND sg13g2_mux4_1
X_1594_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 Tile_X0Y0_W6BEG[11]
+ VPWR VGND sg13g2_buf_1
X_0476_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q DOUT_SRAM17
+ DOUT_SRAM29 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13
+ VPWR VGND sg13g2_mux4_1
X_0614_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q Tile_X0Y1_E2MID[6]
+ Tile_X0Y1_E2END[6] Tile_X0Y1_E6END[9] _0078_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_53_113 VPWR VGND sg13g2_decap_8
XFILLER_53_124 VPWR VGND sg13g2_fill_1
X_1028_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_39_67 VPWR VGND sg13g2_decap_4
X_0330_ VPWR _0033_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
+ VGND sg13g2_inv_1
XFILLER_35_135 VPWR VGND sg13g2_fill_2
XFILLER_35_179 VPWR VGND sg13g2_decap_4
X_1715_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4 Tile_X0Y1_WW4BEG[4]
+ VPWR VGND sg13g2_buf_1
X_1646_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3 Tile_X0Y1_S1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_129 VPWR VGND sg13g2_fill_1
X_0459_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10 VPWR VGND sg13g2_mux4_1
X_0528_ Tile_X0Y0_E2MID[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q _0094_ VPWR
+ VGND sg13g2_nor3_1
X_1577_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2 Tile_X0Y0_W2BEGb[2]
+ VPWR VGND sg13g2_buf_1
XFILLER_26_124 VPWR VGND sg13g2_decap_4
XFILLER_41_35 VPWR VGND sg13g2_decap_8
XFILLER_66_21 VPWR VGND sg13g2_decap_8
XFILLER_32_138 VPWR VGND sg13g2_decap_8
X_1500_ Tile_X0Y0_FrameData[26] Tile_X0Y0_FrameData_O[26] VPWR VGND sg13g2_buf_1
X_0313_ VPWR _0016_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
+ VGND sg13g2_inv_1
X_1362_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1293_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1431_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1629_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData_O[18] VPWR VGND sg13g2_buf_1
XFILLER_52_67 VPWR VGND sg13g2_fill_2
XFILLER_93_30 VPWR VGND sg13g2_fill_1
X_0931_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_171 VPWR VGND sg13g2_decap_8
X_0862_ _0296_ VPWR REN_SRAM VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
+ _0287_ sg13g2_o21ai_1
X_0793_ _0029_ _0082_ _0232_ VPWR VGND sg13g2_nor2_1
XFILLER_95_196 VPWR VGND sg13g2_decap_4
X_1345_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1414_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1276_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_11 VPWR VGND sg13g2_fill_2
XFILLER_88_63 VPWR VGND sg13g2_fill_1
XFILLER_88_30 VPWR VGND sg13g2_decap_4
X_1130_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_199 VPWR VGND sg13g2_fill_1
XFILLER_92_155 VPWR VGND sg13g2_fill_1
X_1061_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0914_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0845_ _0280_ Tile_X0Y1_N2END[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_nand2_1
XFILLER_108_18 VPWR VGND sg13g2_fill_1
XFILLER_52_0 VPWR VGND sg13g2_decap_8
X_0776_ VGND VPWR _0209_ _0211_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A _0216_ sg13g2_a21oi_1
XFILLER_83_199 VPWR VGND sg13g2_fill_1
X_1328_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1259_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_199 VPWR VGND sg13g2_fill_1
XFILLER_90_86 VPWR VGND sg13g2_fill_1
XFILLER_23_80 VPWR VGND sg13g2_fill_2
X_0561_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_EE4END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q _0121_ VPWR
+ VGND sg13g2_mux4_1
X_0492_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q DOUT_SRAM19
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11 VPWR VGND sg13g2_mux4_1
X_0630_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q DOUT_SRAM5
+ DOUT_SRAM13 _0079_ _0082_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5 VPWR VGND sg13g2_mux4_1
X_1113_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_199 VPWR VGND sg13g2_fill_1
X_1044_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0759_ VGND VPWR _0024_ _0200_ _0201_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q
+ sg13g2_a21oi_1
X_0828_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q _0262_
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q _0264_ VPWR
+ VGND _0263_ sg13g2_nand4_1
XFILLER_44_46 VPWR VGND sg13g2_fill_1
XFILLER_56_155 VPWR VGND sg13g2_decap_8
XFILLER_56_199 VPWR VGND sg13g2_fill_1
X_1662_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7 Tile_X0Y1_S2BEGb[7]
+ VPWR VGND sg13g2_buf_1
X_0613_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q Tile_X0Y1_E2MID[7]
+ Tile_X0Y1_E2END[7] Tile_X0Y1_E6END[8] _0043_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0 VPWR VGND sg13g2_mux4_1
X_0544_ VGND VPWR _0011_ _0102_ _0106_ _0105_ sg13g2_a21oi_1
X_0475_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2 VPWR VGND sg13g2_mux4_1
X_1593_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 Tile_X0Y0_W6BEG[10]
+ VPWR VGND sg13g2_buf_1
X_1027_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_15_0 VPWR VGND sg13g2_fill_2
XFILLER_38_199 VPWR VGND sg13g2_fill_1
XFILLER_39_24 VPWR VGND sg13g2_fill_2
XFILLER_29_177 VPWR VGND sg13g2_decap_4
XFILLER_71_11 VPWR VGND sg13g2_fill_2
XFILLER_29_199 VPWR VGND sg13g2_fill_1
XFILLER_96_74 VPWR VGND sg13g2_fill_1
XFILLER_20_70 VPWR VGND sg13g2_fill_2
XFILLER_35_103 VPWR VGND sg13g2_decap_4
X_1645_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2 Tile_X0Y1_S1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1714_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3 Tile_X0Y1_WW4BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1576_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1 Tile_X0Y0_W2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_0527_ VPWR VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ _0092_ _0093_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ ADDR_SRAM5 _0038_ sg13g2_a221oi_1
X_0389_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y0_E2MID[6]
+ Tile_X0Y0_E2END[6] Tile_X0Y0_E6END[9] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1
+ VPWR VGND sg13g2_mux4_1
X_0458_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q DOUT_SRAM20
+ DOUT_SRAM24 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4
+ VPWR VGND sg13g2_mux4_1
XFILLER_103_152 VPWR VGND sg13g2_fill_1
XFILLER_2_19 VPWR VGND sg13g2_fill_2
XFILLER_17_169 VPWR VGND sg13g2_decap_8
X_1430_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_7 VPWR VGND sg13g2_fill_2
X_0312_ VPWR _0015_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ VGND sg13g2_inv_1
X_1361_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1292_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_0 VPWR VGND sg13g2_fill_2
X_1559_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1 Tile_X0Y0_N4BEG[13]
+ VPWR VGND sg13g2_buf_1
X_1628_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_100_199 VPWR VGND sg13g2_fill_1
XFILLER_36_14 VPWR VGND sg13g2_fill_1
XFILLER_52_46 VPWR VGND sg13g2_fill_1
XFILLER_52_79 VPWR VGND sg13g2_fill_1
XFILLER_89_150 VPWR VGND sg13g2_fill_2
XFILLER_77_43 VPWR VGND sg13g2_decap_8
X_0930_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_198 VPWR VGND sg13g2_fill_2
X_0792_ VGND VPWR _0030_ _0230_ _0231_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
+ sg13g2_a21oi_1
X_0861_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q VPWR
+ _0296_ VGND _0291_ _0295_ sg13g2_o21ai_1
X_1413_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_131 VPWR VGND sg13g2_fill_2
X_1344_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1275_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_103_96 VPWR VGND sg13g2_fill_1
XFILLER_77_197 VPWR VGND sg13g2_fill_2
X_1060_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0913_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0775_ VGND VPWR _0026_ _0214_ _0216_ _0215_ sg13g2_a21oi_1
X_0844_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_N2END[3]
+ Tile_X0Y1_E2MID[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0279_ VPWR VGND sg13g2_mux4_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
XFILLER_83_112 VPWR VGND sg13g2_fill_2
XFILLER_68_197 VPWR VGND sg13g2_fill_2
X_1327_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_17_38 VPWR VGND sg13g2_decap_8
XFILLER_17_49 VPWR VGND sg13g2_fill_2
X_1189_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1258_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_11 VPWR VGND sg13g2_fill_1
XFILLER_58_89 VPWR VGND sg13g2_fill_2
XFILLER_59_186 VPWR VGND sg13g2_fill_2
XFILLER_59_197 VPWR VGND sg13g2_fill_2
XFILLER_99_74 VPWR VGND sg13g2_decap_8
X_0560_ VGND VPWR _0013_ _0116_ _0120_ _0119_ sg13g2_a21oi_1
X_0491_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q DOUT_SRAM18
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10 VPWR VGND sg13g2_mux4_1
XFILLER_2_182 VPWR VGND sg13g2_fill_1
X_1112_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_41 VPWR VGND sg13g2_fill_1
X_1043_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0758_ Tile_X0Y1_E1END[2] Tile_X0Y1_EE4END[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ _0200_ VPWR VGND sg13g2_mux2_1
X_0827_ _0263_ Tile_X0Y1_E2END[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_nand2_1
X_0689_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q _0079_
+ _0168_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
+ sg13g2_nand3b_1
XFILLER_56_101 VPWR VGND sg13g2_decap_8
XFILLER_56_178 VPWR VGND sg13g2_fill_2
XFILLER_18_92 VPWR VGND sg13g2_decap_4
XFILLER_70_170 VPWR VGND sg13g2_fill_1
X_1592_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 Tile_X0Y0_W6BEG[9]
+ VPWR VGND sg13g2_buf_1
X_1661_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6 Tile_X0Y1_S2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_0612_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_E6END[11] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15
+ _0077_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3
+ VPWR VGND sg13g2_mux4_1
X_0543_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q VPWR
+ _0105_ VGND _0103_ _0104_ sg13g2_o21ai_1
X_0474_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q DOUT_SRAM16
+ DOUT_SRAM28 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12
+ VPWR VGND sg13g2_mux4_1
X_1026_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_39_47 VPWR VGND sg13g2_fill_2
XFILLER_44_104 VPWR VGND sg13g2_decap_8
XFILLER_44_115 VPWR VGND sg13g2_fill_1
XFILLER_71_34 VPWR VGND sg13g2_decap_8
X_1713_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2 Tile_X0Y1_WW4BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0526_ _0093_ Tile_X0Y0_E2END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_nand2b_1
X_1575_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0 Tile_X0Y0_W2BEGb[0]
+ VPWR VGND sg13g2_buf_1
X_1644_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1 Tile_X0Y1_S1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_0457_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11 VPWR VGND sg13g2_mux4_1
X_0388_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q Tile_X0Y0_E2MID[7]
+ Tile_X0Y0_E2END[7] Tile_X0Y0_E6END[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0
+ VPWR VGND sg13g2_mux4_1
X_1009_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1360_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0311_ VPWR _0014_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
+ VGND sg13g2_inv_1
X_1291_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_0 VPWR VGND sg13g2_fill_1
X_1558_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0 Tile_X0Y0_N4BEG[12]
+ VPWR VGND sg13g2_buf_1
XFILLER_100_134 VPWR VGND sg13g2_decap_4
XFILLER_98_195 VPWR VGND sg13g2_fill_1
X_0509_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[8] Tile_X0Y0_E6END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q BM_SRAM16
+ VPWR VGND sg13g2_mux4_1
X_1489_ Tile_X0Y0_FrameData[15] Tile_X0Y0_FrameData_O[15] VPWR VGND sg13g2_buf_1
X_1627_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_14_118 VPWR VGND sg13g2_fill_1
XFILLER_9_111 VPWR VGND sg13g2_decap_4
X_0791_ Tile_X0Y1_E1END[1] Tile_X0Y1_EE4END[13] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
+ _0230_ VPWR VGND sg13g2_mux2_1
X_0860_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q _0293_
+ _0294_ _0295_ VPWR VGND sg13g2_nor3_1
X_1343_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1412_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1274_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_22_17 VPWR VGND sg13g2_decap_8
X_0989_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_13 VPWR VGND sg13g2_fill_1
X_0912_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0774_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q VPWR
+ _0215_ VGND _0212_ _0213_ sg13g2_o21ai_1
X_0843_ WEN_SRAM _0274_ _0278_ _0270_ _0036_ VPWR VGND sg13g2_a22oi_1
X_1326_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_0 VPWR VGND sg13g2_decap_8
X_1188_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1257_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_58_46 VPWR VGND sg13g2_decap_4
X_0490_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q DOUT_SRAM17
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9 VPWR VGND sg13g2_mux4_1
X_1111_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1042_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0688_ _0165_ VPWR ADDR_SRAM1 VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
+ _0167_ sg13g2_o21ai_1
X_0757_ _0198_ VPWR _0199_ VGND _0023_ _0159_ sg13g2_o21ai_1
X_0826_ _0262_ Tile_X0Y1_E2END[1] _0035_ VPWR VGND sg13g2_nand2_1
X_1309_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_113 VPWR VGND sg13g2_decap_8
XFILLER_60_25 VPWR VGND sg13g2_decap_4
XFILLER_60_47 VPWR VGND sg13g2_decap_8
XFILLER_85_44 VPWR VGND sg13g2_fill_2
XFILLER_69_56 VPWR VGND sg13g2_decap_8
XFILLER_34_70 VPWR VGND sg13g2_decap_4
X_0542_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q VPWR
+ _0104_ VGND Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
X_1591_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8 Tile_X0Y0_W6BEG[8]
+ VPWR VGND sg13g2_buf_1
X_1660_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5 Tile_X0Y1_S2BEGb[5]
+ VPWR VGND sg13g2_buf_1
X_0611_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14
+ _0070_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2
+ VPWR VGND sg13g2_mux4_1
X_0473_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3 VPWR VGND sg13g2_mux4_1
XFILLER_15_2 VPWR VGND sg13g2_fill_1
X_1025_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_29 VPWR VGND sg13g2_fill_1
X_0809_ VGND VPWR _0239_ _0241_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2
+ _0246_ sg13g2_a21oi_1
XFILLER_39_26 VPWR VGND sg13g2_fill_1
XFILLER_55_14 VPWR VGND sg13g2_fill_2
XFILLER_52_171 VPWR VGND sg13g2_decap_4
XFILLER_29_70 VPWR VGND sg13g2_decap_4
XANTENNA_1 VPWR VGND Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A sg13g2_antennanp
X_1712_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1 Tile_X0Y1_WW4BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1643_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0 Tile_X0Y1_S1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0525_ Tile_X0Y0_E2MID[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q _0092_ VPWR
+ VGND sg13g2_nor3_1
X_0456_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q DOUT_SRAM19
+ DOUT_SRAM31 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3
+ VPWR VGND sg13g2_mux4_1
X_1574_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7 Tile_X0Y0_W2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_0387_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E6END[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15
+ _0073_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_25_17 VPWR VGND sg13g2_decap_8
X_1008_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0310_ VPWR _0013_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q
+ VGND sg13g2_inv_1
XFILLER_56_9 VPWR VGND sg13g2_fill_1
X_1290_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_2 VPWR VGND sg13g2_fill_1
XFILLER_16_182 VPWR VGND sg13g2_fill_1
XFILLER_68_0 VPWR VGND sg13g2_fill_2
X_1626_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameData_O[15] VPWR VGND sg13g2_buf_1
X_1557_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A Tile_X0Y0_N4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_100_102 VPWR VGND sg13g2_fill_1
X_0508_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[15] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q DIN_SRAM31
+ VPWR VGND sg13g2_mux4_1
X_1488_ Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData_O[14] VPWR VGND sg13g2_buf_1
X_0439_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q DOUT_SRAM19
+ DOUT_SRAM27 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_36_49 VPWR VGND sg13g2_decap_4
XFILLER_89_152 VPWR VGND sg13g2_fill_1
XFILLER_89_196 VPWR VGND sg13g2_decap_4
X_0790_ _0228_ VPWR _0229_ VGND _0029_ _0160_ sg13g2_o21ai_1
X_1342_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1411_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1273_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0988_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1609_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14 Tile_X0Y0_WW4BEG[14]
+ VPWR VGND sg13g2_buf_1
XFILLER_86_199 VPWR VGND sg13g2_fill_1
XFILLER_86_155 VPWR VGND sg13g2_decap_4
XFILLER_86_100 VPWR VGND sg13g2_decap_4
XFILLER_63_69 VPWR VGND sg13g2_fill_1
XFILLER_12_95 VPWR VGND sg13g2_decap_8
XFILLER_10_199 VPWR VGND sg13g2_fill_1
XFILLER_77_199 VPWR VGND sg13g2_fill_1
X_0911_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0842_ VGND VPWR _0035_ _0277_ _0278_ _0036_ sg13g2_a21oi_1
XFILLER_5_170 VPWR VGND sg13g2_decap_8
X_0773_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q _0214_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_83_114 VPWR VGND sg13g2_fill_1
XFILLER_68_199 VPWR VGND sg13g2_fill_1
X_1325_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1256_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1187_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_17 VPWR VGND sg13g2_fill_2
XFILLER_59_188 VPWR VGND sg13g2_fill_1
XFILLER_59_199 VPWR VGND sg13g2_fill_1
X_1110_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_91 VPWR VGND sg13g2_decap_4
X_1041_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0825_ VGND VPWR Tile_X0Y1_N2MID[6] _0035_ _0261_ _0260_ sg13g2_a21oi_1
X_0687_ VGND VPWR Tile_X0Y1_E2END[1] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ _0167_ _0166_ sg13g2_a21oi_1
X_0756_ VPWR _0198_ _0197_ VGND sg13g2_inv_1
XFILLER_50_0 VPWR VGND sg13g2_decap_8
X_1308_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1239_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_169 VPWR VGND sg13g2_fill_1
XFILLER_44_27 VPWR VGND sg13g2_fill_2
XFILLER_47_147 VPWR VGND sg13g2_fill_2
XFILLER_55_180 VPWR VGND sg13g2_fill_2
X_0541_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
+ _0103_ VPWR VGND sg13g2_nor2b_1
X_1590_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7 Tile_X0Y0_W6BEG[7]
+ VPWR VGND sg13g2_buf_1
X_0472_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q DOUT_SRAM23
+ DOUT_SRAM27 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11
+ VPWR VGND sg13g2_mux4_1
X_0610_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13
+ _0063_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1024_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_125 VPWR VGND sg13g2_fill_1
XFILLER_38_136 VPWR VGND sg13g2_fill_1
XFILLER_53_106 VPWR VGND sg13g2_decap_8
XFILLER_98_0 VPWR VGND sg13g2_fill_2
X_0808_ VGND VPWR _0032_ _0244_ _0246_ _0245_ sg13g2_a21oi_1
X_0739_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q VPWR
+ _0183_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
XFILLER_39_49 VPWR VGND sg13g2_fill_1
XFILLER_55_59 VPWR VGND sg13g2_fill_1
XANTENNA_2 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
X_1711_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0 Tile_X0Y1_WW4BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1642_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData_O[31] VPWR VGND sg13g2_buf_1
X_0455_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_mux4_1
X_0524_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[15] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q BM_SRAM31
+ VPWR VGND sg13g2_mux4_1
X_1573_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6 Tile_X0Y0_W2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_0386_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_mux4_1
X_1007_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_0 VPWR VGND sg13g2_fill_2
XFILLER_26_117 VPWR VGND sg13g2_decap_8
XFILLER_26_128 VPWR VGND sg13g2_fill_2
XFILLER_34_194 VPWR VGND sg13g2_decap_4
XFILLER_41_28 VPWR VGND sg13g2_decap_8
XFILLER_103_199 VPWR VGND sg13g2_fill_1
X_1556_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A Tile_X0Y0_N4BEG[10] VPWR VGND sg13g2_buf_1
X_1625_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData_O[14] VPWR VGND sg13g2_buf_1
X_0369_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2 _0065_ VPWR VGND sg13g2_nor3_1
X_1487_ Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData_O[13] VPWR VGND sg13g2_buf_1
X_0507_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[14] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q DIN_SRAM30
+ VPWR VGND sg13g2_mux4_1
X_0438_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q DOUT_SRAM18
+ DOUT_SRAM26 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_22_120 VPWR VGND sg13g2_decap_8
XFILLER_93_23 VPWR VGND sg13g2_decap_8
XFILLER_13_142 VPWR VGND sg13g2_decap_8
XFILLER_9_168 VPWR VGND sg13g2_decap_4
X_1410_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_178 VPWR VGND sg13g2_fill_1
X_1341_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1272_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0987_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_0 VPWR VGND sg13g2_fill_1
X_1539_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1 Tile_X0Y0_N2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_1608_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13 Tile_X0Y0_WW4BEG[13]
+ VPWR VGND sg13g2_buf_1
XFILLER_103_77 VPWR VGND sg13g2_fill_2
XFILLER_88_34 VPWR VGND sg13g2_fill_1
XFILLER_88_23 VPWR VGND sg13g2_decap_8
XFILLER_12_74 VPWR VGND sg13g2_decap_4
XFILLER_88_56 VPWR VGND sg13g2_decap_8
XFILLER_77_112 VPWR VGND sg13g2_decap_4
XFILLER_92_148 VPWR VGND sg13g2_decap_8
X_0910_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0772_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q VPWR
+ _0213_ VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
X_0841_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0276_ _0275_ _0002_ _0277_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ sg13g2_a221oi_1
XFILLER_68_101 VPWR VGND sg13g2_decap_8
X_1186_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1324_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1255_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_91_170 VPWR VGND sg13g2_decap_4
XFILLER_59_112 VPWR VGND sg13g2_decap_8
XFILLER_74_148 VPWR VGND sg13g2_fill_2
XFILLER_23_73 VPWR VGND sg13g2_decap_8
XFILLER_99_88 VPWR VGND sg13g2_decap_4
XFILLER_2_141 VPWR VGND sg13g2_fill_2
X_1040_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_22 VPWR VGND sg13g2_fill_2
X_0755_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q VPWR
+ _0197_ VGND Tile_X0Y1_E6END[10] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
+ sg13g2_o21ai_1
X_0824_ VGND VPWR _0260_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q sg13g2_or2_1
X_0686_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q Tile_X0Y1_E2MID[1]
+ _0166_ VPWR VGND sg13g2_nor2b_1
XFILLER_43_0 VPWR VGND sg13g2_decap_8
X_1169_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1307_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1238_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_148 VPWR VGND sg13g2_decap_8
XFILLER_55_170 VPWR VGND sg13g2_fill_2
X_0471_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 VPWR VGND sg13g2_mux4_1
X_0540_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q _0102_ VPWR
+ VGND sg13g2_mux2_1
X_1023_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_90 VPWR VGND sg13g2_fill_2
XFILLER_38_104 VPWR VGND sg13g2_fill_1
X_0738_ _0019_ _0043_ _0182_ VPWR VGND sg13g2_nor2_1
X_0807_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q VPWR
+ _0245_ VGND _0242_ _0243_ sg13g2_o21ai_1
X_0669_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q Tile_X0Y1_N4END[0]
+ Tile_X0Y0_S4END[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_29_115 VPWR VGND sg13g2_decap_8
XFILLER_39_17 VPWR VGND sg13g2_decap_8
XFILLER_71_48 VPWR VGND sg13g2_fill_1
XFILLER_84_7 VPWR VGND sg13g2_fill_1
X_1710_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11 Tile_X0Y1_W6BEG[11]
+ VPWR VGND sg13g2_buf_1
XANTENNA_3 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
X_1641_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData_O[30] VPWR VGND sg13g2_buf_1
X_1572_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5 Tile_X0Y0_W2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0523_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[14] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q BM_SRAM30
+ VPWR VGND sg13g2_mux4_1
X_0385_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15 Tile_X0Y1_E6END[7]
+ _0077_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
+ VPWR VGND sg13g2_mux4_1
X_0454_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q DOUT_SRAM18
+ DOUT_SRAM30 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2
+ VPWR VGND sg13g2_mux4_1
X_1006_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_110_0 VPWR VGND sg13g2_fill_1
X_1555_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A Tile_X0Y0_N4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_68_2 VPWR VGND sg13g2_fill_1
X_1624_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData_O[13] VPWR VGND sg13g2_buf_1
X_0506_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[13] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q DIN_SRAM29
+ VPWR VGND sg13g2_mux4_1
X_0368_ _0064_ Tile_X0Y0_S1END[2] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_1486_ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData_O[12] VPWR VGND sg13g2_buf_1
X_0437_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q DOUT_SRAM17
+ DOUT_SRAM25 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_22_165 VPWR VGND sg13g2_decap_4
X_0299_ VPWR _0002_ Tile_X0Y0_S2MID[2] VGND sg13g2_inv_1
XFILLER_89_110 VPWR VGND sg13g2_decap_4
X_1340_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1271_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
Xclkbuf_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VPWR VGND
+ sg13g2_buf_8
X_0986_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1538_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0 Tile_X0Y0_N2BEGb[0]
+ VPWR VGND sg13g2_buf_1
X_1607_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12 Tile_X0Y0_WW4BEG[12]
+ VPWR VGND sg13g2_buf_1
X_1469_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_103_67 VPWR VGND sg13g2_fill_1
XFILLER_103_56 VPWR VGND sg13g2_fill_2
X_0840_ Tile_X0Y1_E2END[3] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q _0276_ VPWR
+ VGND sg13g2_nor3_1
X_0771_ _0025_ _0080_ _0212_ VPWR VGND sg13g2_nor2_1
XFILLER_78_90 VPWR VGND sg13g2_decap_4
X_1323_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1185_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1254_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0969_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_90_69 VPWR VGND sg13g2_decap_4
XFILLER_23_41 VPWR VGND sg13g2_decap_4
XFILLER_80_119 VPWR VGND sg13g2_decap_4
X_0685_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q _0078_
+ _0165_ VPWR VGND Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
+ sg13g2_nand3b_1
X_0754_ VGND VPWR _0189_ _0191_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A _0196_ sg13g2_a21oi_1
X_0823_ _0259_ Tile_X0Y1_N2END[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_nand2_1
X_1306_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_0 VPWR VGND sg13g2_decap_8
X_1099_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1168_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1237_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_26 VPWR VGND sg13g2_fill_2
XFILLER_85_14 VPWR VGND sg13g2_fill_2
XFILLER_18_74 VPWR VGND sg13g2_fill_1
XFILLER_18_96 VPWR VGND sg13g2_fill_1
XFILLER_55_182 VPWR VGND sg13g2_fill_1
XFILLER_109_184 VPWR VGND sg13g2_fill_2
XFILLER_50_83 VPWR VGND sg13g2_decap_4
X_0470_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q DOUT_SRAM22
+ DOUT_SRAM26 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10
+ VPWR VGND sg13g2_mux4_1
X_1022_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0668_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q DOUT_SRAM3
+ DOUT_SRAM15 _0161_ _0043_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15 VPWR VGND sg13g2_mux4_1
X_0737_ VGND VPWR _0020_ _0180_ _0181_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q
+ sg13g2_a21oi_1
X_0806_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
+ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q _0244_ VPWR
+ VGND sg13g2_mux2_1
X_0599_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q VPWR
+ _0154_ VGND _0152_ _0153_ sg13g2_o21ai_1
XFILLER_37_171 VPWR VGND sg13g2_fill_2
XFILLER_20_42 VPWR VGND sg13g2_fill_2
XFILLER_45_72 VPWR VGND sg13g2_decap_8
XFILLER_61_93 VPWR VGND sg13g2_fill_1
XFILLER_6_11 VPWR VGND sg13g2_fill_1
XANTENNA_4 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
X_1640_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData_O[29] VPWR VGND sg13g2_buf_1
X_1571_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4 Tile_X0Y0_W2BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0522_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[13] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q BM_SRAM29
+ VPWR VGND sg13g2_mux4_1
X_0453_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q DOUT_SRAM17
+ DOUT_SRAM29 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_13_2 VPWR VGND sg13g2_fill_1
X_0384_ VPWR VGND _0076_ _0075_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
+ _0007_ _0077_ Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a221oi_1
X_1005_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_66_49 VPWR VGND sg13g2_decap_4
XFILLER_15_75 VPWR VGND sg13g2_decap_4
XFILLER_15_53 VPWR VGND sg13g2_decap_4
XFILLER_40_199 VPWR VGND sg13g2_fill_1
XFILLER_31_30 VPWR VGND sg13g2_fill_2
XFILLER_16_152 VPWR VGND sg13g2_fill_1
XFILLER_16_141 VPWR VGND sg13g2_decap_8
X_1554_ Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A Tile_X0Y0_N4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_98_199 VPWR VGND sg13g2_fill_1
XFILLER_98_188 VPWR VGND sg13g2_decap_8
X_0505_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_EE4END[4] Tile_X0Y0_EE4END[12] Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q DIN_SRAM28
+ VPWR VGND sg13g2_mux4_1
X_1485_ Tile_X0Y0_FrameData[11] Tile_X0Y0_FrameData_O[11] VPWR VGND sg13g2_buf_1
X_0436_ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q DOUT_SRAM16
+ DOUT_SRAM24 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0
+ VPWR VGND sg13g2_mux4_1
X_1623_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData_O[12] VPWR VGND sg13g2_buf_1
.ends

