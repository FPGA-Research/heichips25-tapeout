* NGSPICE file created from W_TT_IF2.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

.subckt W_TT_IF2 CLK_TT_PROJECT ENA_TT_PROJECT RST_N_TT_PROJECT Tile_X0Y0_E1BEG[0]
+ Tile_X0Y0_E1BEG[1] Tile_X0Y0_E1BEG[2] Tile_X0Y0_E1BEG[3] Tile_X0Y0_E2BEG[0] Tile_X0Y0_E2BEG[1]
+ Tile_X0Y0_E2BEG[2] Tile_X0Y0_E2BEG[3] Tile_X0Y0_E2BEG[4] Tile_X0Y0_E2BEG[5] Tile_X0Y0_E2BEG[6]
+ Tile_X0Y0_E2BEG[7] Tile_X0Y0_E2BEGb[0] Tile_X0Y0_E2BEGb[1] Tile_X0Y0_E2BEGb[2] Tile_X0Y0_E2BEGb[3]
+ Tile_X0Y0_E2BEGb[4] Tile_X0Y0_E2BEGb[5] Tile_X0Y0_E2BEGb[6] Tile_X0Y0_E2BEGb[7]
+ Tile_X0Y0_E6BEG[0] Tile_X0Y0_E6BEG[10] Tile_X0Y0_E6BEG[11] Tile_X0Y0_E6BEG[1] Tile_X0Y0_E6BEG[2]
+ Tile_X0Y0_E6BEG[3] Tile_X0Y0_E6BEG[4] Tile_X0Y0_E6BEG[5] Tile_X0Y0_E6BEG[6] Tile_X0Y0_E6BEG[7]
+ Tile_X0Y0_E6BEG[8] Tile_X0Y0_E6BEG[9] Tile_X0Y0_EE4BEG[0] Tile_X0Y0_EE4BEG[10] Tile_X0Y0_EE4BEG[11]
+ Tile_X0Y0_EE4BEG[12] Tile_X0Y0_EE4BEG[13] Tile_X0Y0_EE4BEG[14] Tile_X0Y0_EE4BEG[15]
+ Tile_X0Y0_EE4BEG[1] Tile_X0Y0_EE4BEG[2] Tile_X0Y0_EE4BEG[3] Tile_X0Y0_EE4BEG[4]
+ Tile_X0Y0_EE4BEG[5] Tile_X0Y0_EE4BEG[6] Tile_X0Y0_EE4BEG[7] Tile_X0Y0_EE4BEG[8]
+ Tile_X0Y0_EE4BEG[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2]
+ Tile_X0Y0_S1END[3] Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3]
+ Tile_X0Y0_S2END[4] Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0]
+ Tile_X0Y0_S2MID[1] Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5]
+ Tile_X0Y0_S2MID[6] Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11]
+ Tile_X0Y0_S4END[12] Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15]
+ Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2] Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5]
+ Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7] Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_UserCLKo
+ Tile_X0Y0_W1END[0] Tile_X0Y0_W1END[1] Tile_X0Y0_W1END[2] Tile_X0Y0_W1END[3] Tile_X0Y0_W2END[0]
+ Tile_X0Y0_W2END[1] Tile_X0Y0_W2END[2] Tile_X0Y0_W2END[3] Tile_X0Y0_W2END[4] Tile_X0Y0_W2END[5]
+ Tile_X0Y0_W2END[6] Tile_X0Y0_W2END[7] Tile_X0Y0_W2MID[0] Tile_X0Y0_W2MID[1] Tile_X0Y0_W2MID[2]
+ Tile_X0Y0_W2MID[3] Tile_X0Y0_W2MID[4] Tile_X0Y0_W2MID[5] Tile_X0Y0_W2MID[6] Tile_X0Y0_W2MID[7]
+ Tile_X0Y0_W6END[0] Tile_X0Y0_W6END[10] Tile_X0Y0_W6END[11] Tile_X0Y0_W6END[1] Tile_X0Y0_W6END[2]
+ Tile_X0Y0_W6END[3] Tile_X0Y0_W6END[4] Tile_X0Y0_W6END[5] Tile_X0Y0_W6END[6] Tile_X0Y0_W6END[7]
+ Tile_X0Y0_W6END[8] Tile_X0Y0_W6END[9] Tile_X0Y0_WW4END[0] Tile_X0Y0_WW4END[10] Tile_X0Y0_WW4END[11]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_WW4END[13] Tile_X0Y0_WW4END[14] Tile_X0Y0_WW4END[15]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_WW4END[2] Tile_X0Y0_WW4END[3] Tile_X0Y0_WW4END[4]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_WW4END[6] Tile_X0Y0_WW4END[7] Tile_X0Y0_WW4END[8]
+ Tile_X0Y0_WW4END[9] Tile_X0Y1_E1BEG[0] Tile_X0Y1_E1BEG[1] Tile_X0Y1_E1BEG[2] Tile_X0Y1_E1BEG[3]
+ Tile_X0Y1_E2BEG[0] Tile_X0Y1_E2BEG[1] Tile_X0Y1_E2BEG[2] Tile_X0Y1_E2BEG[3] Tile_X0Y1_E2BEG[4]
+ Tile_X0Y1_E2BEG[5] Tile_X0Y1_E2BEG[6] Tile_X0Y1_E2BEG[7] Tile_X0Y1_E2BEGb[0] Tile_X0Y1_E2BEGb[1]
+ Tile_X0Y1_E2BEGb[2] Tile_X0Y1_E2BEGb[3] Tile_X0Y1_E2BEGb[4] Tile_X0Y1_E2BEGb[5]
+ Tile_X0Y1_E2BEGb[6] Tile_X0Y1_E2BEGb[7] Tile_X0Y1_E6BEG[0] Tile_X0Y1_E6BEG[10] Tile_X0Y1_E6BEG[11]
+ Tile_X0Y1_E6BEG[1] Tile_X0Y1_E6BEG[2] Tile_X0Y1_E6BEG[3] Tile_X0Y1_E6BEG[4] Tile_X0Y1_E6BEG[5]
+ Tile_X0Y1_E6BEG[6] Tile_X0Y1_E6BEG[7] Tile_X0Y1_E6BEG[8] Tile_X0Y1_E6BEG[9] Tile_X0Y1_EE4BEG[0]
+ Tile_X0Y1_EE4BEG[10] Tile_X0Y1_EE4BEG[11] Tile_X0Y1_EE4BEG[12] Tile_X0Y1_EE4BEG[13]
+ Tile_X0Y1_EE4BEG[14] Tile_X0Y1_EE4BEG[15] Tile_X0Y1_EE4BEG[1] Tile_X0Y1_EE4BEG[2]
+ Tile_X0Y1_EE4BEG[3] Tile_X0Y1_EE4BEG[4] Tile_X0Y1_EE4BEG[5] Tile_X0Y1_EE4BEG[6]
+ Tile_X0Y1_EE4BEG[7] Tile_X0Y1_EE4BEG[8] Tile_X0Y1_EE4BEG[9] Tile_X0Y1_FrameData[0]
+ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13]
+ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17]
+ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20]
+ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24]
+ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28]
+ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31]
+ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6]
+ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0]
+ Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11] Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13]
+ Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15] Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17]
+ Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19] Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20]
+ Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22] Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24]
+ Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26] Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28]
+ Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2] Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31]
+ Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4] Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6]
+ Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8] Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0]
+ Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13]
+ Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15] Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17]
+ Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2]
+ Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6]
+ Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2] Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1]
+ Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3] Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6]
+ Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0] Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3]
+ Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5] Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0]
+ Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11] Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13]
+ Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15] Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3]
+ Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5] Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8]
+ Tile_X0Y1_N4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1] Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3]
+ Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2] Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4]
+ Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7] Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1]
+ Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3] Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5]
+ Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7] Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11]
+ Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13] Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15]
+ Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3] Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5]
+ Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8] Tile_X0Y1_S4BEG[9] Tile_X0Y1_UserCLK
+ Tile_X0Y1_W1END[0] Tile_X0Y1_W1END[1] Tile_X0Y1_W1END[2] Tile_X0Y1_W1END[3] Tile_X0Y1_W2END[0]
+ Tile_X0Y1_W2END[1] Tile_X0Y1_W2END[2] Tile_X0Y1_W2END[3] Tile_X0Y1_W2END[4] Tile_X0Y1_W2END[5]
+ Tile_X0Y1_W2END[6] Tile_X0Y1_W2END[7] Tile_X0Y1_W2MID[0] Tile_X0Y1_W2MID[1] Tile_X0Y1_W2MID[2]
+ Tile_X0Y1_W2MID[3] Tile_X0Y1_W2MID[4] Tile_X0Y1_W2MID[5] Tile_X0Y1_W2MID[6] Tile_X0Y1_W2MID[7]
+ Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[10] Tile_X0Y1_W6END[11] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[2]
+ Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[4] Tile_X0Y1_W6END[5] Tile_X0Y1_W6END[6] Tile_X0Y1_W6END[7]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W6END[9] Tile_X0Y1_WW4END[0] Tile_X0Y1_WW4END[10] Tile_X0Y1_WW4END[11]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[15]
+ Tile_X0Y1_WW4END[1] Tile_X0Y1_WW4END[2] Tile_X0Y1_WW4END[3] Tile_X0Y1_WW4END[4]
+ Tile_X0Y1_WW4END[5] Tile_X0Y1_WW4END[6] Tile_X0Y1_WW4END[7] Tile_X0Y1_WW4END[8]
+ Tile_X0Y1_WW4END[9] UIO_IN_TT_PROJECT0 UIO_IN_TT_PROJECT1 UIO_IN_TT_PROJECT2 UIO_IN_TT_PROJECT3
+ UIO_IN_TT_PROJECT4 UIO_IN_TT_PROJECT5 UIO_IN_TT_PROJECT6 UIO_IN_TT_PROJECT7 UIO_OE_TT_PROJECT0
+ UIO_OE_TT_PROJECT1 UIO_OE_TT_PROJECT2 UIO_OE_TT_PROJECT3 UIO_OE_TT_PROJECT4 UIO_OE_TT_PROJECT5
+ UIO_OE_TT_PROJECT6 UIO_OE_TT_PROJECT7 UIO_OUT_TT_PROJECT0 UIO_OUT_TT_PROJECT1 UIO_OUT_TT_PROJECT2
+ UIO_OUT_TT_PROJECT3 UIO_OUT_TT_PROJECT4 UIO_OUT_TT_PROJECT5 UIO_OUT_TT_PROJECT6
+ UIO_OUT_TT_PROJECT7 UI_IN_TT_PROJECT0 UI_IN_TT_PROJECT1 UI_IN_TT_PROJECT2 UI_IN_TT_PROJECT3
+ UI_IN_TT_PROJECT4 UI_IN_TT_PROJECT5 UI_IN_TT_PROJECT6 UI_IN_TT_PROJECT7 UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT1 UO_OUT_TT_PROJECT2 UO_OUT_TT_PROJECT3 UO_OUT_TT_PROJECT4 UO_OUT_TT_PROJECT5
+ UO_OUT_TT_PROJECT6 UO_OUT_TT_PROJECT7 VGND VPWR
X_0367_ VPWR _0297_ Tile_X0Y1_W6END[3] VGND sg13g2_inv_1
XFILLER_22_155 VPWR VGND sg13g2_fill_1
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_89_199 VPWR VGND sg13g2_fill_1
XFILLER_26_85 VPWR VGND sg13g2_fill_2
XFILLER_9_126 VPWR VGND sg13g2_fill_1
XFILLER_13_177 VPWR VGND sg13g2_fill_1
XFILLER_13_199 VPWR VGND sg13g2_fill_1
X_1270_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0985_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1606_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameData_O[4] VPWR VGND sg13g2_buf_1
X_1468_ Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData_O[3] VPWR VGND sg13g2_buf_1
X_0419_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q Tile_X0Y0_W2MID[6]
+ Tile_X0Y0_W2END[6] Tile_X0Y0_W6END[9] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG1
+ VPWR VGND sg13g2_mux4_1
X_1537_ Tile_X0Y1_N4END[8] Tile_X0Y0_N4BEG[0] VPWR VGND sg13g2_buf_1
X_1399_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_103_35 VPWR VGND sg13g2_decap_8
XFILLER_10_125 VPWR VGND sg13g2_fill_1
XFILLER_6_107 VPWR VGND sg13g2_decap_8
XFILLER_12_65 VPWR VGND sg13g2_fill_1
XFILLER_85_180 VPWR VGND sg13g2_decap_4
XFILLER_77_158 VPWR VGND sg13g2_fill_2
XFILLER_77_114 VPWR VGND sg13g2_decap_8
X_0770_ _0162_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q
+ _0163_ VPWR VGND sg13g2_nor2b_1
XFILLER_68_114 VPWR VGND sg13g2_fill_1
X_1322_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_4 VPWR VGND sg13g2_fill_1
X_1253_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_94_90 VPWR VGND sg13g2_decap_4
X_1184_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0968_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0899_ VGND VPWR Tile_X0Y1_W2MID[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0275_ _0274_ sg13g2_a21oi_1
XFILLER_59_147 VPWR VGND sg13g2_fill_1
XFILLER_82_194 VPWR VGND sg13g2_decap_4
XFILLER_99_35 VPWR VGND sg13g2_decap_8
XFILLER_23_75 VPWR VGND sg13g2_fill_2
XFILLER_2_154 VPWR VGND sg13g2_decap_8
XFILLER_2_143 VPWR VGND sg13g2_fill_1
XFILLER_2_110 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_9_33 VPWR VGND sg13g2_fill_2
X_0822_ VGND VPWR Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
+ _0207_ _0208_ _0304_ sg13g2_a21oi_1
XFILLER_89_90 VPWR VGND sg13g2_decap_8
X_0684_ _0119_ _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_nand2b_1
X_0753_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q UO_OUT_TT_PROJECT3
+ _0158_ UO_OUT_TT_PROJECT7 _0335_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG15 VPWR VGND sg13g2_mux4_1
XFILLER_56_139 VPWR VGND sg13g2_fill_1
X_1305_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_0 VPWR VGND sg13g2_decap_4
X_1236_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_14 VPWR VGND sg13g2_decap_8
X_1098_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1167_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_7 VPWR VGND sg13g2_decap_8
XFILLER_70_175 VPWR VGND sg13g2_fill_2
XFILLER_70_142 VPWR VGND sg13g2_fill_2
XFILLER_109_141 VPWR VGND sg13g2_fill_2
XFILLER_109_130 VPWR VGND sg13g2_decap_8
XFILLER_50_40 VPWR VGND sg13g2_decap_8
X_1021_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_142 VPWR VGND sg13g2_fill_1
X_0805_ _0153_ _0149_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q
+ _0193_ VPWR VGND sg13g2_mux2_1
X_0598_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q _0065_
+ _0066_ VPWR VGND sg13g2_and2_1
X_0667_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q Tile_X0Y1_W2MID[6]
+ Tile_X0Y1_W2END[6] Tile_X0Y1_W6END[9] _0342_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG1 VPWR VGND sg13g2_mux4_1
X_0736_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0007_ Tile_X0Y0_S4END[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q
+ _0150_ VPWR VGND sg13g2_mux4_1
X_1219_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_39 VPWR VGND sg13g2_decap_4
XFILLER_106_133 VPWR VGND sg13g2_decap_8
XFILLER_96_25 VPWR VGND sg13g2_fill_1
XFILLER_96_14 VPWR VGND sg13g2_decap_8
XFILLER_43_197 VPWR VGND sg13g2_fill_2
X_0521_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q
+ _0011_ VPWR VGND sg13g2_mux4_1
X_0452_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q Tile_X0Y0_W1END[0]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W2MID[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG4
+ VPWR VGND sg13g2_mux4_1
X_1570_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb4 Tile_X0Y1_E2BEGb[4]
+ VPWR VGND sg13g2_buf_1
XANTENNA_5 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0383_ Tile_X0Y1_N1END[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q _0313_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_96_0 VPWR VGND sg13g2_decap_8
X_1004_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_197 VPWR VGND sg13g2_fill_2
XFILLER_106_35 VPWR VGND sg13g2_decap_8
X_0719_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q
+ _0142_ _0141_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb5 _0348_ sg13g2_a221oi_1
XFILLER_15_32 VPWR VGND sg13g2_fill_2
XFILLER_16_120 VPWR VGND sg13g2_fill_1
XFILLER_16_142 VPWR VGND sg13g2_fill_2
X_1622_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData_O[20] VPWR VGND sg13g2_buf_1
X_1553_ clknet_1_1__leaf_Tile_X0Y1_UserCLK Tile_X0Y0_UserCLKo VPWR VGND sg13g2_buf_1
X_1484_ Tile_X0Y0_FrameData[19] Tile_X0Y0_FrameData_O[19] VPWR VGND sg13g2_buf_1
X_0504_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q UIO_OUT_TT_PROJECT3
+ UIO_OE_TT_PROJECT7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG3 VPWR VGND sg13g2_mux4_1
X_0435_ _0345_ _0346_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q
+ _0347_ VPWR VGND sg13g2_nand3_1
XFILLER_11_0 VPWR VGND sg13g2_decap_4
X_0366_ VPWR _0296_ Tile_X0Y0_S2MID[3] VGND sg13g2_inv_1
XFILLER_77_49 VPWR VGND sg13g2_fill_1
XFILLER_26_42 VPWR VGND sg13g2_fill_2
XFILLER_42_85 VPWR VGND sg13g2_decap_4
XFILLER_3_79 VPWR VGND sg13g2_decap_8
XFILLER_3_35 VPWR VGND sg13g2_decap_8
XFILLER_83_81 VPWR VGND sg13g2_fill_1
X_0984_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1536_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb7 Tile_X0Y0_N2BEGb[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_59_0 VPWR VGND sg13g2_fill_2
X_1605_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_103_14 VPWR VGND sg13g2_decap_8
X_1467_ Tile_X0Y0_FrameData[2] Tile_X0Y0_FrameData_O[2] VPWR VGND sg13g2_buf_1
X_0418_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_W2MID[7]
+ Tile_X0Y0_W2END[7] Tile_X0Y0_W6END[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG0
+ VPWR VGND sg13g2_mux4_1
X_1398_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_18 VPWR VGND sg13g2_fill_2
XFILLER_12_55 VPWR VGND sg13g2_fill_1
XFILLER_92_129 VPWR VGND sg13g2_fill_2
XFILLER_37_30 VPWR VGND sg13g2_decap_4
XFILLER_5_185 VPWR VGND sg13g2_decap_8
X_1321_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1252_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1183_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0967_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1519_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG2 Tile_X0Y0_N1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0898_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_N2END[3]
+ _0274_ VPWR VGND sg13g2_nor2b_1
XFILLER_74_107 VPWR VGND sg13g2_decap_4
XFILLER_67_181 VPWR VGND sg13g2_fill_1
XFILLER_99_14 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_fill_1
XFILLER_48_95 VPWR VGND sg13g2_fill_2
XFILLER_73_151 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_80_60 VPWR VGND sg13g2_fill_2
X_0821_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15 _0003_
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q _0207_ VPWR
+ VGND sg13g2_mux2_1
X_0752_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0007_ Tile_X0Y0_S4END[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q
+ _0158_ VPWR VGND sg13g2_mux4_1
X_0683_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q
+ _0118_ _0117_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG1 _0341_ sg13g2_a221oi_1
X_1166_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1235_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1304_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_170 VPWR VGND sg13g2_decap_8
X_1097_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_17 VPWR VGND sg13g2_fill_1
XFILLER_55_184 VPWR VGND sg13g2_fill_1
XFILLER_70_198 VPWR VGND sg13g2_fill_2
XFILLER_34_42 VPWR VGND sg13g2_fill_1
X_1020_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_60 VPWR VGND sg13g2_decap_4
XFILLER_61_198 VPWR VGND sg13g2_fill_2
XFILLER_46_162 VPWR VGND sg13g2_decap_4
X_0804_ VGND VPWR _0188_ _0190_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG0
+ _0192_ sg13g2_a21oi_1
X_0735_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT6 _0149_ _0342_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG6 VPWR VGND sg13g2_mux4_1
X_0597_ _0065_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6 VPWR VGND sg13g2_nand2b_1
X_0666_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q Tile_X0Y1_W2MID[7]
+ Tile_X0Y1_W2END[7] Tile_X0Y1_W6END[8] _0335_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG0 VPWR VGND sg13g2_mux4_1
X_1149_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1218_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_112 VPWR VGND sg13g2_decap_8
XFILLER_20_33 VPWR VGND sg13g2_fill_1
XFILLER_20_44 VPWR VGND sg13g2_fill_1
XFILLER_20_66 VPWR VGND sg13g2_fill_1
XFILLER_29_53 VPWR VGND sg13g2_fill_1
XFILLER_29_64 VPWR VGND sg13g2_fill_1
XFILLER_29_75 VPWR VGND sg13g2_fill_2
XFILLER_43_187 VPWR VGND sg13g2_fill_2
XFILLER_61_40 VPWR VGND sg13g2_decap_8
XANTENNA_6 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_6_35 VPWR VGND sg13g2_decap_8
X_0520_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q UIO_OUT_TT_PROJECT7
+ UIO_OE_TT_PROJECT3 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG11 VPWR VGND sg13g2_mux4_1
X_0451_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2END[4] Tile_X0Y0_W6END[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_6_79 VPWR VGND sg13g2_decap_8
X_0382_ _0312_ _0311_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
X_1003_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_89_0 VPWR VGND sg13g2_fill_2
XFILLER_34_187 VPWR VGND sg13g2_fill_2
X_0718_ UO_OUT_TT_PROJECT5 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q _0142_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_106_14 VPWR VGND sg13g2_decap_8
X_0649_ Tile_X0Y0_W6END[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q
+ _0105_ VPWR VGND sg13g2_nor2b_1
XFILLER_102_170 VPWR VGND sg13g2_decap_8
XFILLER_56_95 VPWR VGND sg13g2_decap_8
XFILLER_82_7 VPWR VGND sg13g2_decap_8
XFILLER_16_165 VPWR VGND sg13g2_fill_2
X_1552_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG3 Tile_X0Y0_N4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_1621_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameData_O[19] VPWR VGND sg13g2_buf_1
X_1483_ Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData_O[18] VPWR VGND sg13g2_buf_1
X_0503_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_mux4_1
X_0365_ VPWR _0295_ Tile_X0Y1_W2END[5] VGND sg13g2_inv_1
X_0434_ _0346_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y0_S2MID[2] VPWR VGND sg13g2_nand2_1
XFILLER_89_168 VPWR VGND sg13g2_fill_2
XFILLER_93_27 VPWR VGND sg13g2_decap_8
XFILLER_13_146 VPWR VGND sg13g2_fill_2
XFILLER_3_58 VPWR VGND sg13g2_decap_8
XFILLER_3_14 VPWR VGND sg13g2_decap_8
X_0983_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1535_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb6 Tile_X0Y0_N2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_1604_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameData_O[2] VPWR VGND sg13g2_buf_1
X_1466_ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData_O[1] VPWR VGND sg13g2_buf_1
X_0417_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb0
+ Tile_X0Y0_S2MID[0] Tile_X0Y1_N2MID[0] Tile_X0Y0_S2END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_94_182 VPWR VGND sg13g2_fill_2
XFILLER_94_160 VPWR VGND sg13g2_fill_1
X_1397_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_53_96 VPWR VGND sg13g2_decap_8
XFILLER_5_142 VPWR VGND sg13g2_fill_2
X_1320_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_78_82 VPWR VGND sg13g2_fill_1
XFILLER_78_71 VPWR VGND sg13g2_decap_8
XFILLER_68_138 VPWR VGND sg13g2_fill_2
X_1182_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1251_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0966_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_0 VPWR VGND sg13g2_fill_2
X_0897_ VGND VPWR Tile_X0Y1_W2MID[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0273_ _0272_ sg13g2_a21oi_1
X_1518_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG1 Tile_X0Y0_N1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1449_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG0 Tile_X0Y0_EE4BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_23_77 VPWR VGND sg13g2_fill_1
XFILLER_58_160 VPWR VGND sg13g2_fill_1
XFILLER_2_189 VPWR VGND sg13g2_decap_8
XFILLER_104_91 VPWR VGND sg13g2_decap_8
XFILLER_64_84 VPWR VGND sg13g2_fill_2
XFILLER_9_35 VPWR VGND sg13g2_fill_1
XFILLER_9_79 VPWR VGND sg13g2_fill_1
X_0820_ _0206_ _0205_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_nand2b_1
X_0751_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT6 _0157_ _0342_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG14 VPWR VGND sg13g2_mux4_1
X_0682_ UO_OUT_TT_PROJECT1 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q _0118_ VPWR
+ VGND sg13g2_nor3_1
X_1303_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_163 VPWR VGND sg13g2_fill_1
XFILLER_64_141 VPWR VGND sg13g2_fill_2
X_1096_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1234_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1165_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_160 VPWR VGND sg13g2_decap_8
XFILLER_100_49 VPWR VGND sg13g2_decap_8
XFILLER_109_47 VPWR VGND sg13g2_fill_2
X_0949_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_144 VPWR VGND sg13g2_fill_1
XFILLER_18_55 VPWR VGND sg13g2_fill_2
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_75_83 VPWR VGND sg13g2_decap_4
XFILLER_38_119 VPWR VGND sg13g2_decap_8
X_0803_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q _0191_
+ _0192_ VPWR VGND sg13g2_nor2_1
X_0665_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W6END[11] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15
+ _0328_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG3
+ VPWR VGND sg13g2_mux4_1
X_0734_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0311_ Tile_X0Y0_S4END[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q
+ _0149_ VPWR VGND sg13g2_mux4_1
X_0596_ VPWR _0064_ _0063_ VGND sg13g2_inv_1
X_1079_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1148_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1217_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_177 VPWR VGND sg13g2_decap_8
XFILLER_106_168 VPWR VGND sg13g2_decap_8
XFILLER_29_32 VPWR VGND sg13g2_fill_2
XFILLER_101_70 VPWR VGND sg13g2_decap_4
XFILLER_43_155 VPWR VGND sg13g2_decap_8
XFILLER_43_199 VPWR VGND sg13g2_fill_1
XANTENNA_7 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_6_58 VPWR VGND sg13g2_decap_8
XFILLER_6_14 VPWR VGND sg13g2_decap_8
X_0450_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb3
+ Tile_X0Y0_S2MID[3] Tile_X0Y1_N2MID[3] Tile_X0Y0_S2END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3 VPWR VGND sg13g2_mux4_1
X_0381_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q Tile_X0Y0_W1END[1]
+ Tile_X0Y0_W6END[9] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13
+ _0310_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q _0311_
+ VPWR VGND sg13g2_mux4_1
X_1002_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_199 VPWR VGND sg13g2_fill_1
X_0648_ VGND VPWR UIO_IN_TT_PROJECT5 _0104_ _0103_ sg13g2_or2_1
X_0717_ _0141_ _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_nand2b_1
X_0579_ _0048_ VPWR _0049_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ _0014_ sg13g2_o21ai_1
XFILLER_15_34 VPWR VGND sg13g2_fill_1
XFILLER_15_45 VPWR VGND sg13g2_fill_1
XFILLER_25_199 VPWR VGND sg13g2_fill_1
XFILLER_40_147 VPWR VGND sg13g2_fill_2
XFILLER_16_111 VPWR VGND sg13g2_decap_8
XFILLER_16_144 VPWR VGND sg13g2_fill_1
X_1551_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG2 Tile_X0Y0_N4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_1482_ Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData_O[17] VPWR VGND sg13g2_buf_1
X_0502_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q UIO_OUT_TT_PROJECT2
+ UIO_OE_TT_PROJECT6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG2 VPWR VGND sg13g2_mux4_1
X_1620_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData_O[18] VPWR VGND sg13g2_buf_1
X_0364_ VPWR _0294_ Tile_X0Y0_W6END[11] VGND sg13g2_inv_1
X_0433_ _0345_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG2 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_89_125 VPWR VGND sg13g2_decap_8
XFILLER_101_0 VPWR VGND sg13g2_decap_8
XFILLER_107_91 VPWR VGND sg13g2_decap_8
XFILLER_67_84 VPWR VGND sg13g2_decap_4
XFILLER_67_40 VPWR VGND sg13g2_fill_2
XFILLER_83_50 VPWR VGND sg13g2_fill_2
X_0982_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1534_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb5 Tile_X0Y0_N2BEGb[5]
+ VPWR VGND sg13g2_buf_1
X_1465_ Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData_O[0] VPWR VGND sg13g2_buf_1
X_1603_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_103_49 VPWR VGND sg13g2_decap_8
X_1396_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_0416_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q Tile_X0Y1_W2MID[7]
+ Tile_X0Y1_W2END[7] Tile_X0Y1_W6END[7] _0335_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb0 VPWR VGND sg13g2_mux4_1
XFILLER_5_7 VPWR VGND sg13g2_decap_8
XFILLER_85_150 VPWR VGND sg13g2_decap_4
XFILLER_77_128 VPWR VGND sg13g2_decap_4
XFILLER_53_53 VPWR VGND sg13g2_decap_4
XFILLER_5_121 VPWR VGND sg13g2_decap_8
XFILLER_5_154 VPWR VGND sg13g2_decap_8
XFILLER_91_120 VPWR VGND sg13g2_decap_8
X_1250_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1181_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0965_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_0 VPWR VGND sg13g2_decap_8
X_0896_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_W2MID[3]
+ _0272_ VPWR VGND sg13g2_nor2b_1
X_1517_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG0 Tile_X0Y0_N1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1448_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG11 Tile_X0Y0_E6BEG[11]
+ VPWR VGND sg13g2_buf_1
XFILLER_67_150 VPWR VGND sg13g2_fill_2
X_1379_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_49 VPWR VGND sg13g2_decap_8
XFILLER_2_168 VPWR VGND sg13g2_decap_8
XFILLER_2_135 VPWR VGND sg13g2_fill_2
XFILLER_2_124 VPWR VGND sg13g2_decap_8
XFILLER_104_70 VPWR VGND sg13g2_decap_8
XFILLER_58_150 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_4
XFILLER_48_97 VPWR VGND sg13g2_fill_1
XFILLER_64_41 VPWR VGND sg13g2_decap_4
XFILLER_9_58 VPWR VGND sg13g2_decap_4
XFILLER_9_14 VPWR VGND sg13g2_decap_4
X_0681_ _0117_ _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_nand2b_1
X_0750_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0311_ Tile_X0Y0_S4END[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q
+ _0157_ VPWR VGND sg13g2_mux4_1
X_1233_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_4 VPWR VGND sg13g2_fill_1
X_1302_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1095_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1164_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_28 VPWR VGND sg13g2_decap_8
X_0948_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_109_59 VPWR VGND sg13g2_fill_1
X_0879_ Tile_X0Y1_W2END[4] Tile_X0Y0_S2MID[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0256_ VPWR VGND sg13g2_mux2_1
XFILLER_34_88 VPWR VGND sg13g2_decap_4
XFILLER_109_155 VPWR VGND sg13g2_decap_8
XFILLER_109_122 VPWR VGND sg13g2_decap_4
XFILLER_50_98 VPWR VGND sg13g2_decap_4
XFILLER_75_40 VPWR VGND sg13g2_fill_2
X_0802_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q Tile_X0Y1_W1END[0]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_W6END[4] _0158_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
+ _0191_ VPWR VGND sg13g2_mux4_1
X_0664_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y1_W1END[2]
+ Tile_X0Y1_W6END[10] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14
+ _0321_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG2
+ VPWR VGND sg13g2_mux4_1
X_0733_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q UO_OUT_TT_PROJECT1
+ _0148_ UO_OUT_TT_PROJECT5 _0349_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG5 VPWR VGND sg13g2_mux4_1
X_0595_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q VPWR
+ _0063_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q
+ _0062_ sg13g2_o21ai_1
X_1216_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_0 VPWR VGND sg13g2_fill_2
X_1078_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1147_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_153 VPWR VGND sg13g2_decap_4
XFILLER_106_147 VPWR VGND sg13g2_decap_8
XFILLER_105_7 VPWR VGND sg13g2_decap_8
XFILLER_29_77 VPWR VGND sg13g2_fill_1
XFILLER_61_97 VPWR VGND sg13g2_decap_4
XANTENNA_8 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0380_ VPWR VGND _0308_ _0309_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q
+ _0287_ _0310_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a221oi_1
XFILLER_20_7 VPWR VGND sg13g2_decap_4
X_1001_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_89_2 VPWR VGND sg13g2_fill_1
XFILLER_106_49 VPWR VGND sg13g2_decap_8
X_0647_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q _0100_
+ _0101_ _0104_ VPWR VGND sg13g2_nor3_1
X_0578_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q _0047_
+ _0048_ VPWR VGND sg13g2_and2_1
X_0716_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q
+ _0140_ _0139_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb4 _0355_ sg13g2_a221oi_1
XFILLER_25_145 VPWR VGND sg13g2_decap_8
XFILLER_31_89 VPWR VGND sg13g2_fill_2
XFILLER_16_167 VPWR VGND sg13g2_fill_1
X_1550_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG1 Tile_X0Y0_N4BEG[13]
+ VPWR VGND sg13g2_buf_1
X_1481_ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData_O[16] VPWR VGND sg13g2_buf_1
X_0501_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q UIO_OUT_TT_PROJECT1
+ UIO_OE_TT_PROJECT5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG1 VPWR VGND sg13g2_mux4_1
X_0432_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q _0343_
+ _0344_ VPWR VGND sg13g2_nor2_1
X_0363_ VPWR _0293_ Tile_X0Y0_W6END[10] VGND sg13g2_inv_1
XFILLER_26_78 VPWR VGND sg13g2_decap_8
XFILLER_21_170 VPWR VGND sg13g2_fill_1
XFILLER_107_70 VPWR VGND sg13g2_decap_8
XFILLER_3_49 VPWR VGND sg13g2_decap_4
X_0981_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1602_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData_O[0] VPWR VGND sg13g2_buf_1
X_1533_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb4 Tile_X0Y0_N2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_1464_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG15 Tile_X0Y0_EE4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_1395_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0415_ _0330_ _0333_ _0335_ VPWR VGND sg13g2_nor2b_1
XFILLER_103_28 VPWR VGND sg13g2_decap_8
XFILLER_94_184 VPWR VGND sg13g2_fill_1
XFILLER_85_184 VPWR VGND sg13g2_fill_1
XFILLER_77_107 VPWR VGND sg13g2_decap_8
XFILLER_5_100 VPWR VGND sg13g2_decap_8
XFILLER_5_199 VPWR VGND sg13g2_fill_1
XFILLER_94_94 VPWR VGND sg13g2_fill_1
XFILLER_94_83 VPWR VGND sg13g2_decap_8
X_1180_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0964_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_57_0 VPWR VGND sg13g2_decap_8
X_1516_ Tile_X0Y1_FrameStrobe[19] Tile_X0Y0_FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_0895_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0270_ _0271_ VPWR VGND sg13g2_nor3_1
X_1447_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG10 Tile_X0Y0_E6BEG[10]
+ VPWR VGND sg13g2_buf_1
X_1378_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_198 VPWR VGND sg13g2_fill_2
XFILLER_99_28 VPWR VGND sg13g2_decap_8
XFILLER_23_57 VPWR VGND sg13g2_fill_1
XFILLER_2_147 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_80_41 VPWR VGND sg13g2_fill_2
XFILLER_9_48 VPWR VGND sg13g2_decap_4
XFILLER_89_50 VPWR VGND sg13g2_fill_2
X_0680_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q
+ _0116_ _0115_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG0 _0334_ sg13g2_a221oi_1
XFILLER_50_7 VPWR VGND sg13g2_decap_4
XFILLER_29_4 VPWR VGND sg13g2_fill_1
X_1301_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1232_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_198 VPWR VGND sg13g2_fill_2
XFILLER_64_143 VPWR VGND sg13g2_fill_1
X_1094_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1163_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0947_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0878_ _0305_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG0 _0255_ VPWR VGND sg13g2_nor3_1
XFILLER_109_101 VPWR VGND sg13g2_decap_8
XFILLER_50_11 VPWR VGND sg13g2_fill_1
XFILLER_50_33 VPWR VGND sg13g2_decap_8
XFILLER_61_135 VPWR VGND sg13g2_decap_8
XFILLER_98_7 VPWR VGND sg13g2_decap_8
XFILLER_91_73 VPWR VGND sg13g2_fill_2
XFILLER_61_179 VPWR VGND sg13g2_fill_2
X_0801_ VGND VPWR Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
+ _0189_ _0190_ _0301_ sg13g2_a21oi_1
X_0594_ _0061_ VPWR _0062_ VGND Tile_X0Y0_W6END[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ sg13g2_o21ai_1
X_0663_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q Tile_X0Y1_W1END[1]
+ Tile_X0Y1_W6END[9] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13
+ _0314_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG1
+ VPWR VGND sg13g2_mux4_1
X_0732_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0318_ Tile_X0Y0_S4END[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q
+ _0148_ VPWR VGND sg13g2_mux4_1
X_1146_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_71 VPWR VGND sg13g2_fill_1
X_1215_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1077_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_126 VPWR VGND sg13g2_decap_8
XFILLER_28_198 VPWR VGND sg13g2_fill_2
XFILLER_45_11 VPWR VGND sg13g2_fill_2
XFILLER_105_170 VPWR VGND sg13g2_decap_8
XFILLER_6_49 VPWR VGND sg13g2_decap_4
XANTENNA_9 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_105_181 VPWR VGND sg13g2_fill_1
X_1000_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0715_ UO_OUT_TT_PROJECT4 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q _0140_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_106_28 VPWR VGND sg13g2_decap_8
X_0646_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q _0102_
+ _0103_ VPWR VGND sg13g2_nor2b_1
X_0577_ _0047_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4 VPWR VGND sg13g2_nand2b_1
X_1129_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_140 VPWR VGND sg13g2_fill_2
XFILLER_56_21 VPWR VGND sg13g2_decap_4
XFILLER_56_76 VPWR VGND sg13g2_fill_2
XFILLER_24_190 VPWR VGND sg13g2_fill_2
X_1480_ Tile_X0Y0_FrameData[15] Tile_X0Y0_FrameData_O[15] VPWR VGND sg13g2_buf_1
X_0500_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q UIO_OUT_TT_PROJECT0
+ UIO_OE_TT_PROJECT4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG0 VPWR VGND sg13g2_mux4_1
X_0362_ VPWR _0292_ Tile_X0Y0_W6END[9] VGND sg13g2_inv_1
X_0431_ Tile_X0Y1_N2MID[2] Tile_X0Y1_N2END[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
+ _0343_ VPWR VGND sg13g2_mux2_1
XFILLER_7_92 VPWR VGND sg13g2_fill_1
X_0629_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q Tile_X0Y0_WW4END[2]
+ Tile_X0Y0_WW4END[10] _0012_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q _0089_ VPWR
+ VGND sg13g2_mux4_1
XFILLER_42_89 VPWR VGND sg13g2_fill_2
XFILLER_3_28 VPWR VGND sg13g2_decap_8
XFILLER_83_52 VPWR VGND sg13g2_fill_1
XFILLER_67_42 VPWR VGND sg13g2_fill_1
XFILLER_83_74 VPWR VGND sg13g2_decap_8
XFILLER_80_7 VPWR VGND sg13g2_decap_8
X_0980_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_12_171 VPWR VGND sg13g2_fill_1
X_1532_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb3 Tile_X0Y0_N2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_1601_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG15 Tile_X0Y1_EE4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_1463_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG14 Tile_X0Y0_EE4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_1394_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0414_ _0334_ _0333_ _0330_ VPWR VGND sg13g2_nand2b_1
XFILLER_12_48 VPWR VGND sg13g2_fill_2
XFILLER_12_59 VPWR VGND sg13g2_fill_1
XFILLER_37_89 VPWR VGND sg13g2_decap_4
XFILLER_5_178 VPWR VGND sg13g2_decap_8
XFILLER_91_199 VPWR VGND sg13g2_fill_1
X_0963_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0894_ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2END[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0270_ VPWR VGND sg13g2_mux2_1
X_1515_ Tile_X0Y1_FrameStrobe[18] Tile_X0Y0_FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_1446_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG9 Tile_X0Y0_E6BEG[9]
+ VPWR VGND sg13g2_buf_1
XFILLER_82_122 VPWR VGND sg13g2_decap_8
XFILLER_4_93 VPWR VGND sg13g2_decap_8
X_1377_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_11 VPWR VGND sg13g2_fill_2
XFILLER_73_199 VPWR VGND sg13g2_fill_1
X_1162_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1300_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1231_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1093_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0946_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0877_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0251_ _0253_ _0248_ _0254_ _0249_ sg13g2_a221oi_1
X_1429_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb0 Tile_X0Y0_E2BEGb[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_55_188 VPWR VGND sg13g2_decap_4
XFILLER_55_177 VPWR VGND sg13g2_decap_8
XFILLER_59_43 VPWR VGND sg13g2_decap_4
XFILLER_59_21 VPWR VGND sg13g2_fill_1
XFILLER_75_64 VPWR VGND sg13g2_fill_2
XFILLER_75_42 VPWR VGND sg13g2_fill_1
XFILLER_46_166 VPWR VGND sg13g2_fill_1
XFILLER_46_199 VPWR VGND sg13g2_fill_1
X_0800_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12 _0000_
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q _0189_ VPWR
+ VGND sg13g2_mux2_1
X_0731_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT4 _0147_ _0356_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG4 VPWR VGND sg13g2_mux4_1
X_0593_ _0061_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_nand2b_1
X_0662_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y1_W1END[0]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12
+ _0010_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG0
+ VPWR VGND sg13g2_mux4_1
XFILLER_27_2 VPWR VGND sg13g2_fill_1
X_1145_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1214_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1076_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_105 VPWR VGND sg13g2_decap_8
X_0929_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_45_34 VPWR VGND sg13g2_fill_2
XFILLER_45_78 VPWR VGND sg13g2_fill_2
XFILLER_61_11 VPWR VGND sg13g2_fill_2
XFILLER_6_28 VPWR VGND sg13g2_decap_8
X_0645_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q Tile_X0Y0_W1END[1]
+ Tile_X0Y0_WW4END[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q
+ _0102_ VPWR VGND sg13g2_mux4_1
X_0714_ _0139_ _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_nand2b_1
X_0576_ VPWR _0046_ _0045_ VGND sg13g2_inv_1
X_1059_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1128_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_31_25 VPWR VGND sg13g2_fill_1
XFILLER_31_47 VPWR VGND sg13g2_decap_4
XFILLER_110_7 VPWR VGND sg13g2_decap_8
XFILLER_102_163 VPWR VGND sg13g2_decap_8
XFILLER_98_117 VPWR VGND sg13g2_decap_4
X_0361_ VPWR _0291_ Tile_X0Y0_W6END[8] VGND sg13g2_inv_1
X_0430_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q Tile_X0Y0_W2MID[5]
+ Tile_X0Y0_W2END[5] Tile_X0Y0_W6END[10] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG2
+ VPWR VGND sg13g2_mux4_1
X_0628_ _0087_ VPWR _0088_ VGND Tile_X0Y0_W6END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q
+ sg13g2_o21ai_1
X_0559_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q VPWR
+ _0031_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q
+ _0030_ sg13g2_o21ai_1
XFILLER_8_143 VPWR VGND sg13g2_fill_1
XFILLER_12_150 VPWR VGND sg13g2_fill_1
X_1531_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb2 Tile_X0Y0_N2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_1462_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG13 Tile_X0Y0_EE4BEG[13]
+ VPWR VGND sg13g2_buf_1
X_1600_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG14 Tile_X0Y1_EE4BEG[14]
+ VPWR VGND sg13g2_buf_1
XFILLER_94_131 VPWR VGND sg13g2_fill_1
XFILLER_79_150 VPWR VGND sg13g2_decap_4
X_1393_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0413_ _0331_ _0332_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q
+ _0333_ VPWR VGND sg13g2_nand3_1
XFILLER_94_197 VPWR VGND sg13g2_fill_2
XFILLER_85_197 VPWR VGND sg13g2_fill_2
XFILLER_85_120 VPWR VGND sg13g2_decap_8
XFILLER_53_23 VPWR VGND sg13g2_fill_2
XFILLER_5_135 VPWR VGND sg13g2_decap_8
XFILLER_91_145 VPWR VGND sg13g2_decap_4
XFILLER_76_197 VPWR VGND sg13g2_fill_2
X_0962_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0893_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q _0268_
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q _0269_ VPWR
+ VGND sg13g2_nand3_1
X_1445_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG8 Tile_X0Y0_E6BEG[8]
+ VPWR VGND sg13g2_buf_1
XFILLER_4_72 VPWR VGND sg13g2_decap_8
X_1514_ Tile_X0Y1_FrameStrobe[17] Tile_X0Y0_FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_1376_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_7 VPWR VGND sg13g2_decap_8
XFILLER_2_105 VPWR VGND sg13g2_fill_1
XFILLER_104_84 VPWR VGND sg13g2_decap_8
XFILLER_64_77 VPWR VGND sg13g2_decap_8
X_1092_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1161_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1230_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0945_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0876_ VPWR _0253_ _0252_ VGND sg13g2_inv_1
X_1428_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG7 Tile_X0Y0_E2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1359_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_109_169 VPWR VGND sg13g2_decap_8
XFILLER_75_87 VPWR VGND sg13g2_fill_2
X_0661_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q Tile_X0Y0_W1END[0]
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_W6END[4]
+ _0006_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG0
+ VPWR VGND sg13g2_mux4_1
X_0730_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0325_ Tile_X0Y0_S4END[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q
+ _0147_ VPWR VGND sg13g2_mux4_1
X_0592_ VGND VPWR _0055_ _0058_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG1
+ _0060_ sg13g2_a21oi_1
X_1213_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1075_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1144_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0928_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0859_ _0238_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_nand2b_1
XFILLER_101_63 VPWR VGND sg13g2_decap_8
XFILLER_51_170 VPWR VGND sg13g2_decap_8
XFILLER_101_96 VPWR VGND sg13g2_fill_2
XFILLER_86_75 VPWR VGND sg13g2_decap_8
XFILLER_19_101 VPWR VGND sg13g2_decap_8
X_0644_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q VPWR
+ _0101_ VGND Tile_X0Y0_WW4END[13] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q
+ sg13g2_o21ai_1
X_0713_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q
+ _0138_ _0137_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb3 _0355_ sg13g2_a221oi_1
X_0575_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q VPWR
+ _0045_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q
+ _0044_ sg13g2_o21ai_1
X_1058_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1127_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_40_118 VPWR VGND sg13g2_decap_4
XFILLER_103_7 VPWR VGND sg13g2_decap_8
XFILLER_102_197 VPWR VGND sg13g2_fill_2
XFILLER_72_33 VPWR VGND sg13g2_fill_1
XFILLER_97_96 VPWR VGND sg13g2_decap_4
X_0360_ VPWR _0290_ Tile_X0Y0_W6END[0] VGND sg13g2_inv_1
XFILLER_7_72 VPWR VGND sg13g2_fill_2
XFILLER_89_118 VPWR VGND sg13g2_decap_8
X_0558_ _0029_ VPWR _0030_ VGND Tile_X0Y0_W6END[10] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ sg13g2_o21ai_1
X_0627_ VGND VPWR _0293_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q
+ _0087_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q sg13g2_a21oi_1
X_0489_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q UIO_OUT_TT_PROJECT5
+ UIO_OE_TT_PROJECT5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_21_162 VPWR VGND sg13g2_fill_2
XFILLER_107_84 VPWR VGND sg13g2_decap_8
XFILLER_67_88 VPWR VGND sg13g2_fill_2
XFILLER_67_77 VPWR VGND sg13g2_decap_8
XFILLER_83_43 VPWR VGND sg13g2_decap_8
XFILLER_8_100 VPWR VGND sg13g2_fill_1
XFILLER_32_80 VPWR VGND sg13g2_decap_8
XFILLER_32_91 VPWR VGND sg13g2_fill_2
X_1530_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb1 Tile_X0Y0_N2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_1461_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG12 Tile_X0Y0_EE4BEG[12]
+ VPWR VGND sg13g2_buf_1
X_1392_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0412_ _0332_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
+ Tile_X0Y0_S2MID[0] VPWR VGND sg13g2_nand2_1
XFILLER_92_0 VPWR VGND sg13g2_decap_8
X_1659_ Tile_X0Y0_S4END[13] Tile_X0Y1_S4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_85_154 VPWR VGND sg13g2_fill_2
XFILLER_53_46 VPWR VGND sg13g2_decap_8
XFILLER_53_57 VPWR VGND sg13g2_fill_1
XFILLER_78_43 VPWR VGND sg13g2_decap_8
XFILLER_5_147 VPWR VGND sg13g2_decap_8
XFILLER_5_114 VPWR VGND sg13g2_decap_8
XFILLER_94_31 VPWR VGND sg13g2_fill_1
XFILLER_91_113 VPWR VGND sg13g2_decap_8
X_0961_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_0892_ _0268_ Tile_X0Y1_W2END[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_nand2_1
X_1444_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG7 Tile_X0Y0_E6BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1513_ Tile_X0Y1_FrameStrobe[16] Tile_X0Y0_FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
X_1375_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_143 VPWR VGND sg13g2_decap_8
XFILLER_2_117 VPWR VGND sg13g2_decap_8
XFILLER_104_63 VPWR VGND sg13g2_decap_8
XFILLER_64_45 VPWR VGND sg13g2_fill_1
XFILLER_89_20 VPWR VGND sg13g2_fill_2
XFILLER_36_8 VPWR VGND sg13g2_decap_8
X_1091_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1160_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0944_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0875_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q Tile_X0Y1_N2END[3]
+ Tile_X0Y1_W2END[1] Tile_X0Y1_W2MID[0] Tile_X0Y1_W2END[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0252_ VPWR VGND sg13g2_mux4_1
XFILLER_55_0 VPWR VGND sg13g2_fill_2
X_1427_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG6 Tile_X0Y0_E2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1358_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1289_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_48 VPWR VGND sg13g2_fill_2
XFILLER_109_137 VPWR VGND sg13g2_decap_4
XFILLER_109_115 VPWR VGND sg13g2_decap_8
XFILLER_75_33 VPWR VGND sg13g2_decap_8
X_0660_ VGND VPWR UIO_IN_TT_PROJECT7 _0114_ _0113_ sg13g2_or2_1
X_0591_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q _0059_
+ _0060_ VPWR VGND sg13g2_nor2_1
X_1212_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1074_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1143_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_157 VPWR VGND sg13g2_fill_1
XFILLER_52_116 VPWR VGND sg13g2_fill_2
X_0927_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0858_ _0237_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q VPWR VGND
+ sg13g2_nand2b_1
X_0789_ VGND VPWR _0174_ _0177_ Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_10.A _0179_ sg13g2_a21oi_1
XFILLER_45_36 VPWR VGND sg13g2_fill_1
XFILLER_101_42 VPWR VGND sg13g2_decap_8
XFILLER_51_160 VPWR VGND sg13g2_decap_8
XFILLER_34_116 VPWR VGND sg13g2_decap_4
XFILLER_96_7 VPWR VGND sg13g2_decap_8
X_0643_ Tile_X0Y0_W6END[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q
+ _0100_ VPWR VGND sg13g2_nor2b_1
X_0574_ _0043_ VPWR _0044_ VGND Tile_X0Y0_W6END[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ sg13g2_o21ai_1
X_0712_ UO_OUT_TT_PROJECT3 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q _0138_ VPWR
+ VGND sg13g2_nor3_1
X_1126_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1057_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_127 VPWR VGND sg13g2_fill_1
XFILLER_30_174 VPWR VGND sg13g2_fill_2
X_0557_ _0029_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_nand2b_1
X_0626_ VGND VPWR Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q
+ _0084_ UIO_IN_TT_PROJECT1 _0086_ sg13g2_a21oi_1
X_0488_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q UIO_OUT_TT_PROJECT4
+ UIO_OE_TT_PROJECT4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG4 VPWR VGND sg13g2_mux4_1
X_1109_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_26_38 VPWR VGND sg13g2_decap_4
XFILLER_107_63 VPWR VGND sg13g2_decap_8
X_1460_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG11 Tile_X0Y0_EE4BEG[11]
+ VPWR VGND sg13g2_buf_1
X_1391_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0411_ _0331_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_94_199 VPWR VGND sg13g2_fill_1
XFILLER_85_0 VPWR VGND sg13g2_decap_8
X_1658_ Tile_X0Y0_S4END[12] Tile_X0Y1_S4BEG[4] VPWR VGND sg13g2_buf_1
X_0609_ _0075_ VPWR _0076_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ _0011_ sg13g2_o21ai_1
X_1589_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG3 Tile_X0Y1_EE4BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_85_199 VPWR VGND sg13g2_fill_1
XFILLER_76_199 VPWR VGND sg13g2_fill_1
XFILLER_76_188 VPWR VGND sg13g2_fill_1
X_0960_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_91 VPWR VGND sg13g2_decap_8
X_0891_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_W2END[1]
+ _0267_ VPWR VGND sg13g2_nor2b_1
X_1512_ Tile_X0Y1_FrameStrobe[15] Tile_X0Y0_FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_1443_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG6 Tile_X0Y0_E6BEG[6]
+ VPWR VGND sg13g2_buf_1
XFILLER_4_192 VPWR VGND sg13g2_decap_8
X_1374_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_199 VPWR VGND sg13g2_fill_1
XFILLER_23_17 VPWR VGND sg13g2_fill_2
XFILLER_104_42 VPWR VGND sg13g2_decap_8
XFILLER_73_158 VPWR VGND sg13g2_fill_1
XFILLER_58_199 VPWR VGND sg13g2_fill_1
XFILLER_89_43 VPWR VGND sg13g2_decap_8
X_1090_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_114 VPWR VGND sg13g2_decap_4
XFILLER_38_80 VPWR VGND sg13g2_fill_2
XFILLER_49_177 VPWR VGND sg13g2_decap_4
X_0943_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0874_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0250_ _0251_ VPWR VGND sg13g2_nor3_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_1426_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG5 Tile_X0Y0_E2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_1357_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_17 VPWR VGND sg13g2_fill_2
X_1288_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
Xclkbuf_1_1__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_1__leaf_Tile_X0Y1_UserCLK
+ VPWR VGND sg13g2_buf_8
XFILLER_59_68 VPWR VGND sg13g2_fill_2
XFILLER_108_193 VPWR VGND sg13g2_decap_8
X_0590_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q Tile_X0Y0_W1END[1]
+ Tile_X0Y0_WW4END[13] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG9 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ _0059_ VPWR VGND sg13g2_mux4_1
X_1142_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_42 VPWR VGND sg13g2_decap_4
XFILLER_37_114 VPWR VGND sg13g2_decap_4
XFILLER_37_147 VPWR VGND sg13g2_fill_2
X_1211_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1073_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_119 VPWR VGND sg13g2_decap_8
X_0926_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0857_ _0233_ VPWR UI_IN_TT_PROJECT5 VGND _0234_ _0236_ sg13g2_o21ai_1
X_1409_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0788_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q _0178_
+ _0179_ VPWR VGND sg13g2_nor2_1
XFILLER_101_21 VPWR VGND sg13g2_decap_8
XFILLER_61_47 VPWR VGND sg13g2_decap_8
XFILLER_105_163 VPWR VGND sg13g2_decap_8
XFILLER_19_125 VPWR VGND sg13g2_fill_2
XFILLER_19_147 VPWR VGND sg13g2_fill_2
X_0711_ _0137_ _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_nand2b_1
X_0573_ _0043_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_nand2b_1
X_0642_ VGND VPWR UIO_IN_TT_PROJECT4 _0099_ _0098_ sg13g2_or2_1
X_1125_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1056_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0909_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q _0282_
+ _0284_ _0285_ VPWR VGND sg13g2_nor3_1
XFILLER_102_199 VPWR VGND sg13g2_fill_1
XFILLER_102_177 VPWR VGND sg13g2_decap_4
XFILLER_102_133 VPWR VGND sg13g2_decap_8
XFILLER_56_14 VPWR VGND sg13g2_decap_8
XFILLER_24_150 VPWR VGND sg13g2_fill_2
XANTENNA_90 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XFILLER_97_21 VPWR VGND sg13g2_decap_8
XFILLER_30_142 VPWR VGND sg13g2_decap_8
X_0625_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q _0085_
+ _0086_ VPWR VGND sg13g2_nor2_1
XFILLER_7_74 VPWR VGND sg13g2_fill_1
X_0487_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q UIO_OUT_TT_PROJECT3
+ UIO_OE_TT_PROJECT3 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG3 VPWR VGND sg13g2_mux4_1
X_0556_ _0026_ _0028_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG1
+ VPWR VGND sg13g2_nor2_1
XFILLER_30_0 VPWR VGND sg13g2_fill_2
X_1039_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1108_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_42 VPWR VGND sg13g2_decap_8
XFILLER_88_197 VPWR VGND sg13g2_fill_2
X_1390_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0410_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q _0329_
+ _0330_ VPWR VGND sg13g2_nor2_1
XFILLER_94_156 VPWR VGND sg13g2_decap_4
X_0608_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q _0074_
+ _0075_ VPWR VGND sg13g2_and2_1
X_1657_ Tile_X0Y0_S4END[11] Tile_X0Y1_S4BEG[3] VPWR VGND sg13g2_buf_1
X_1588_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG2 Tile_X0Y1_EE4BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0539_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q UIO_OUT_TT_PROJECT2
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG5 _0013_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG10
+ VPWR VGND sg13g2_mux4_1
XFILLER_78_78 VPWR VGND sg13g2_decap_4
XFILLER_27_93 VPWR VGND sg13g2_decap_8
X_0890_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0266_ VPWR VGND sg13g2_nor2b_1
X_1442_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG5 Tile_X0Y0_E6BEG[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_4_171 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_decap_8
X_1511_ Tile_X0Y1_FrameStrobe[14] Tile_X0Y0_FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
XFILLER_82_115 VPWR VGND sg13g2_decap_8
XFILLER_4_86 VPWR VGND sg13g2_decap_8
XFILLER_4_53 VPWR VGND sg13g2_fill_2
X_1373_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_148 VPWR VGND sg13g2_fill_1
XFILLER_58_123 VPWR VGND sg13g2_fill_2
XFILLER_104_98 VPWR VGND sg13g2_fill_1
XFILLER_104_21 VPWR VGND sg13g2_decap_8
XFILLER_64_14 VPWR VGND sg13g2_fill_1
XFILLER_13_40 VPWR VGND sg13g2_fill_1
XFILLER_8_0 VPWR VGND sg13g2_decap_8
XFILLER_1_130 VPWR VGND sg13g2_fill_1
XFILLER_72_170 VPWR VGND sg13g2_fill_1
X_0942_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0873_ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2END[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0250_ VPWR VGND sg13g2_mux2_1
X_1425_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG4 Tile_X0Y0_E2BEG[4]
+ VPWR VGND sg13g2_buf_1
X_1356_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1287_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_137 VPWR VGND sg13g2_fill_2
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_108_183 VPWR VGND sg13g2_fill_2
XFILLER_108_172 VPWR VGND sg13g2_decap_8
X_1072_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1141_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_1_76 VPWR VGND sg13g2_fill_1
X_1210_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_80 VPWR VGND sg13g2_fill_1
XFILLER_65_90 VPWR VGND sg13g2_decap_8
XFILLER_52_118 VPWR VGND sg13g2_fill_1
X_0925_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0787_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y1_W1END[2]
+ Tile_X0Y1_W6END[10] Tile_X0Y1_WW4END[2] _0156_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ _0178_ VPWR VGND sg13g2_mux4_1
X_0856_ _0235_ VPWR _0236_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
+ _0153_ sg13g2_o21ai_1
X_1408_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1339_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_77 VPWR VGND sg13g2_fill_2
XFILLER_51_184 VPWR VGND sg13g2_fill_1
XFILLER_105_186 VPWR VGND sg13g2_fill_2
XFILLER_105_142 VPWR VGND sg13g2_decap_8
XFILLER_105_197 VPWR VGND sg13g2_fill_2
XFILLER_86_45 VPWR VGND sg13g2_fill_2
XFILLER_86_23 VPWR VGND sg13g2_fill_1
X_0641_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q _0095_
+ _0096_ _0099_ VPWR VGND sg13g2_nor3_1
X_0710_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q
+ _0136_ _0135_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb2 _0348_ sg13g2_a221oi_1
X_0572_ _0040_ _0042_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG3
+ VPWR VGND sg13g2_nor2_1
X_1055_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1124_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0908_ Tile_X0Y0_S2MID[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0284_ VPWR VGND sg13g2_nor2b_1
X_0839_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q _0219_
+ _0220_ _0222_ VPWR VGND sg13g2_nor3_1
XFILLER_16_118 VPWR VGND sg13g2_fill_2
XANTENNA_80 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_91 VPWR VGND Tile_X0Y1_N2MID[4] sg13g2_antennanp
XFILLER_108_0 VPWR VGND sg13g2_decap_8
XFILLER_15_140 VPWR VGND sg13g2_fill_2
X_0624_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q Tile_X0Y0_WW4END[1]
+ Tile_X0Y0_WW4END[9] _0013_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q _0085_ VPWR
+ VGND sg13g2_mux4_1
XFILLER_7_97 VPWR VGND sg13g2_decap_8
XFILLER_7_53 VPWR VGND sg13g2_fill_2
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_30_198 VPWR VGND sg13g2_fill_2
XFILLER_97_198 VPWR VGND sg13g2_fill_2
XFILLER_97_143 VPWR VGND sg13g2_fill_2
X_0486_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q UIO_OUT_TT_PROJECT2
+ UIO_OE_TT_PROJECT2 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG2 VPWR VGND sg13g2_mux4_1
X_0555_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q _0027_
+ _0028_ VPWR VGND sg13g2_nor2_1
X_1038_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1107_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_143 VPWR VGND sg13g2_fill_2
XFILLER_107_98 VPWR VGND sg13g2_decap_8
XFILLER_107_21 VPWR VGND sg13g2_decap_8
XFILLER_101_7 VPWR VGND sg13g2_decap_8
XFILLER_79_143 VPWR VGND sg13g2_decap_8
X_0538_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q UIO_OUT_TT_PROJECT1
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG6 _0012_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG9
+ VPWR VGND sg13g2_mux4_1
X_0607_ _0074_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7 VPWR VGND sg13g2_nand2b_1
X_1656_ Tile_X0Y0_S4END[10] Tile_X0Y1_S4BEG[2] VPWR VGND sg13g2_buf_1
X_1587_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG1 Tile_X0Y1_EE4BEG[1]
+ VPWR VGND sg13g2_buf_1
X_0469_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q Tile_X0Y1_W2MID[0]
+ Tile_X0Y1_W2END[0] Tile_X0Y1_W6END[0] _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb7 VPWR VGND sg13g2_mux4_1
XFILLER_5_128 VPWR VGND sg13g2_decap_8
XFILLER_91_127 VPWR VGND sg13g2_fill_1
X_1441_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG4 Tile_X0Y0_E6BEG[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_64_7 VPWR VGND sg13g2_decap_8
XFILLER_4_161 VPWR VGND sg13g2_decap_8
XFILLER_4_65 VPWR VGND sg13g2_decap_8
XFILLER_4_21 VPWR VGND sg13g2_decap_8
X_1510_ Tile_X0Y1_FrameStrobe[13] Tile_X0Y0_FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
XFILLER_67_124 VPWR VGND sg13g2_fill_2
X_1372_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_90_0 VPWR VGND sg13g2_decap_8
X_1639_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG1 Tile_X0Y1_S2BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_77 VPWR VGND sg13g2_decap_8
XFILLER_81_171 VPWR VGND sg13g2_decap_4
XFILLER_73_105 VPWR VGND sg13g2_decap_8
XFILLER_80_14 VPWR VGND sg13g2_fill_2
XFILLER_1_142 VPWR VGND sg13g2_fill_2
XFILLER_1_164 VPWR VGND sg13g2_fill_2
XFILLER_49_113 VPWR VGND sg13g2_fill_1
XFILLER_49_135 VPWR VGND sg13g2_decap_4
X_0941_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0872_ VGND VPWR Tile_X0Y1_W2MID[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0249_ _0247_ sg13g2_a21oi_1
X_1424_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG3 Tile_X0Y0_E2BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1355_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1286_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_116 VPWR VGND sg13g2_decap_4
XFILLER_46_116 VPWR VGND sg13g2_fill_1
XFILLER_46_138 VPWR VGND sg13g2_decap_8
XFILLER_108_151 VPWR VGND sg13g2_decap_8
X_1071_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1140_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_149 VPWR VGND sg13g2_fill_1
XFILLER_45_160 VPWR VGND sg13g2_decap_8
X_0924_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_141 VPWR VGND sg13g2_decap_4
X_0786_ _0176_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q
+ _0177_ VPWR VGND sg13g2_nor2b_1
X_0855_ _0235_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_nand2b_1
XFILLER_53_0 VPWR VGND sg13g2_decap_4
X_1407_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1338_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_56 VPWR VGND sg13g2_decap_8
XFILLER_28_149 VPWR VGND sg13g2_fill_1
X_1269_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_196 VPWR VGND sg13g2_decap_4
XFILLER_86_68 VPWR VGND sg13g2_decap_8
XFILLER_27_193 VPWR VGND sg13g2_fill_1
X_0571_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q _0041_
+ _0042_ VPWR VGND sg13g2_nor2_1
X_0640_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q _0097_
+ _0098_ VPWR VGND sg13g2_nor2b_1
X_1054_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_76_90 VPWR VGND sg13g2_fill_1
X_1123_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0907_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q VPWR
+ _0283_ VGND _0295_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ sg13g2_o21ai_1
XFILLER_102_102 VPWR VGND sg13g2_decap_8
X_0769_ VGND VPWR Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ _0334_ _0162_ _0161_ sg13g2_a21oi_1
X_0838_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y1_WW4END[2]
+ Tile_X0Y1_WW4END[10] Tile_X0Y1_W6END[2] Tile_X0Y1_W6END[10] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q
+ _0221_ VPWR VGND sg13g2_mux4_1
XFILLER_110_190 VPWR VGND sg13g2_decap_8
XANTENNA_92 VPWR VGND Tile_X0Y1_N2MID[4] sg13g2_antennanp
XANTENNA_70 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_81 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_62_70 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_97_100 VPWR VGND sg13g2_fill_1
X_0623_ _0083_ VPWR _0084_ VGND Tile_X0Y0_W6END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q
+ sg13g2_o21ai_1
X_0554_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q Tile_X0Y0_W1END[1]
+ Tile_X0Y0_WW4END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG9 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ _0027_ VPWR VGND sg13g2_mux4_1
XFILLER_7_65 VPWR VGND sg13g2_decap_8
XFILLER_97_166 VPWR VGND sg13g2_fill_2
X_0485_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q UIO_OUT_TT_PROJECT1
+ UIO_OE_TT_PROJECT1 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG1 VPWR VGND sg13g2_mux4_1
X_1106_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_16_0 VPWR VGND sg13g2_decap_4
X_1037_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_77 VPWR VGND sg13g2_decap_8
XFILLER_88_199 VPWR VGND sg13g2_fill_1
XFILLER_88_144 VPWR VGND sg13g2_decap_8
XFILLER_12_199 VPWR VGND sg13g2_fill_1
X_0537_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q UIO_OUT_TT_PROJECT0
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG7 _0011_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG8
+ VPWR VGND sg13g2_mux4_1
X_0606_ VPWR _0073_ _0072_ VGND sg13g2_inv_1
X_1655_ Tile_X0Y0_S4END[9] Tile_X0Y1_S4BEG[1] VPWR VGND sg13g2_buf_1
X_1586_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG0 Tile_X0Y1_EE4BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0399_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END3 _0323_ VPWR VGND sg13g2_nor3_1
X_0468_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q Tile_X0Y1_N2MID[7]
+ Tile_X0Y1_N2END[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG7
+ Tile_X0Y0_S2MID[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q
+ _0003_ VPWR VGND sg13g2_mux4_1
XFILLER_78_36 VPWR VGND sg13g2_decap_8
XFILLER_5_107 VPWR VGND sg13g2_decap_8
XFILLER_94_24 VPWR VGND sg13g2_decap_8
XFILLER_76_169 VPWR VGND sg13g2_fill_2
X_1440_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG3 Tile_X0Y0_E6BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_57_7 VPWR VGND sg13g2_decap_8
X_1371_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_68_91 VPWR VGND sg13g2_fill_2
XFILLER_83_0 VPWR VGND sg13g2_decap_4
X_1638_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG0 Tile_X0Y1_S2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1569_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb3 Tile_X0Y1_E2BEGb[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_56 VPWR VGND sg13g2_decap_8
XFILLER_80_37 VPWR VGND sg13g2_decap_4
XFILLER_38_61 VPWR VGND sg13g2_fill_2
X_0940_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0871_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q _0306_
+ _0248_ VPWR VGND sg13g2_nor2_1
X_1423_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG2 Tile_X0Y0_E2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1354_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1285_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_139 VPWR VGND sg13g2_fill_1
XFILLER_109_108 VPWR VGND sg13g2_decap_8
XFILLER_91_69 VPWR VGND sg13g2_decap_4
XFILLER_108_130 VPWR VGND sg13g2_decap_8
XFILLER_24_96 VPWR VGND sg13g2_fill_1
X_1070_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0923_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0854_ _0234_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q VPWR VGND
+ sg13g2_nand2b_1
X_0785_ VGND VPWR Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ _0348_ _0176_ _0175_ sg13g2_a21oi_1
X_1406_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1337_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1268_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_35 VPWR VGND sg13g2_decap_8
X_1199_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_105_199 VPWR VGND sg13g2_fill_1
XFILLER_105_188 VPWR VGND sg13g2_fill_1
XFILLER_105_177 VPWR VGND sg13g2_decap_4
XFILLER_10_98 VPWR VGND sg13g2_fill_1
XFILLER_10_76 VPWR VGND sg13g2_fill_1
XFILLER_34_109 VPWR VGND sg13g2_decap_8
XFILLER_42_153 VPWR VGND sg13g2_decap_8
X_0570_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q Tile_X0Y0_W1END[3]
+ Tile_X0Y0_WW4END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ _0041_ VPWR VGND sg13g2_mux4_1
X_1122_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_90 VPWR VGND sg13g2_decap_4
X_1053_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0906_ Tile_X0Y1_W2END[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q _0282_ VPWR
+ VGND sg13g2_nor3_1
X_0837_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q _0156_
+ _0220_ VPWR VGND sg13g2_nor2_1
X_0768_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q VPWR
+ _0161_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
X_0699_ _0129_ _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_24_197 VPWR VGND sg13g2_fill_2
XFILLER_97_35 VPWR VGND sg13g2_decap_4
XANTENNA_60 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_71 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_82 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XANTENNA_93 VPWR VGND Tile_X0Y1_N2MID[5] sg13g2_antennanp
XFILLER_15_120 VPWR VGND sg13g2_fill_2
XFILLER_30_112 VPWR VGND sg13g2_decap_8
XFILLER_46_94 VPWR VGND sg13g2_fill_1
XFILLER_30_123 VPWR VGND sg13g2_fill_2
X_0484_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q UIO_OUT_TT_PROJECT0
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG0 VPWR VGND sg13g2_mux4_1
X_0553_ VGND VPWR Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q
+ _0025_ _0026_ _0024_ sg13g2_a21oi_1
X_0622_ VGND VPWR _0292_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q
+ _0083_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q sg13g2_a21oi_1
XFILLER_87_90 VPWR VGND sg13g2_fill_2
X_1105_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1036_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_56 VPWR VGND sg13g2_decap_8
XFILLER_12_123 VPWR VGND sg13g2_fill_2
XFILLER_7_171 VPWR VGND sg13g2_decap_8
X_1654_ Tile_X0Y0_S4END[8] Tile_X0Y1_S4BEG[0] VPWR VGND sg13g2_buf_1
X_0536_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q UIO_OUT_TT_PROJECT7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG7 VPWR VGND sg13g2_mux4_1
X_0605_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q VPWR
+ _0072_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q
+ _0071_ sg13g2_o21ai_1
X_0467_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W2MID[0] Tile_X0Y0_W2END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG7
+ VPWR VGND sg13g2_mux4_1
X_1585_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG11 Tile_X0Y1_E6BEG[11]
+ VPWR VGND sg13g2_buf_1
XFILLER_93_170 VPWR VGND sg13g2_fill_2
X_1019_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0398_ _0322_ Tile_X0Y0_S1END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_4_185 VPWR VGND sg13g2_decap_8
X_1370_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_129 VPWR VGND sg13g2_fill_2
XFILLER_76_0 VPWR VGND sg13g2_fill_2
X_1637_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG3 Tile_X0Y1_S1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_35 VPWR VGND sg13g2_decap_8
X_1499_ Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
X_0519_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG4 VPWR VGND sg13g2_mux4_1
XFILLER_73_129 VPWR VGND sg13g2_fill_1
X_1568_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb2 Tile_X0Y1_E2BEGb[2]
+ VPWR VGND sg13g2_buf_1
XFILLER_1_144 VPWR VGND sg13g2_fill_1
XFILLER_1_166 VPWR VGND sg13g2_fill_1
XFILLER_1_199 VPWR VGND sg13g2_fill_1
XFILLER_64_118 VPWR VGND sg13g2_fill_2
XFILLER_64_107 VPWR VGND sg13g2_decap_8
X_0870_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_W2MID[3]
+ _0247_ VPWR VGND sg13g2_nor2b_1
X_1422_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG1 Tile_X0Y0_E2BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1353_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1284_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_170 VPWR VGND sg13g2_decap_8
X_0999_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_39_170 VPWR VGND sg13g2_fill_2
XFILLER_24_75 VPWR VGND sg13g2_decap_4
XFILLER_6_0 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_1_46 VPWR VGND sg13g2_fill_1
XFILLER_37_118 VPWR VGND sg13g2_fill_2
X_0922_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_176 VPWR VGND sg13g2_fill_2
X_0853_ _0233_ _0232_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_nand2b_1
X_1405_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0784_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q VPWR
+ _0175_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
XFILLER_39_0 VPWR VGND sg13g2_decap_4
X_1336_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1267_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1198_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_14 VPWR VGND sg13g2_decap_8
XFILLER_105_123 VPWR VGND sg13g2_fill_2
XFILLER_105_112 VPWR VGND sg13g2_decap_8
XFILLER_105_156 VPWR VGND sg13g2_decap_8
XFILLER_51_51 VPWR VGND sg13g2_fill_2
X_1052_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1121_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_33_198 VPWR VGND sg13g2_fill_2
X_0905_ _0278_ _0280_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0281_ VPWR VGND sg13g2_nand3_1
X_0767_ _0160_ _0159_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_nand2b_1
X_0836_ _0148_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q
+ _0219_ VPWR VGND sg13g2_nor2b_1
XFILLER_102_126 VPWR VGND sg13g2_decap_8
X_0698_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q
+ _0128_ _0127_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG6 _0341_ sg13g2_a221oi_1
X_1319_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_72 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_61 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_50 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_83 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XFILLER_97_14 VPWR VGND sg13g2_decap_8
XANTENNA_94 VPWR VGND Tile_X0Y1_N2MID[5] sg13g2_antennanp
XFILLER_15_176 VPWR VGND sg13g2_fill_2
X_0621_ VGND VPWR Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q
+ _0080_ UIO_IN_TT_PROJECT0 _0082_ sg13g2_a21oi_1
XFILLER_97_168 VPWR VGND sg13g2_fill_1
X_0483_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END3
+ UIO_OUT_TT_PROJECT1 Tile_X0Y0_S1END[3] UIO_OUT_TT_PROJECT4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG3 VPWR VGND sg13g2_mux4_1
X_0552_ _0013_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ _0025_ VPWR VGND sg13g2_mux2_1
X_1035_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1104_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_168 VPWR VGND sg13g2_fill_2
XFILLER_107_35 VPWR VGND sg13g2_decap_8
X_0819_ _0151_ _0147_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q
+ _0205_ VPWR VGND sg13g2_mux2_1
XFILLER_8_139 VPWR VGND sg13g2_decap_4
XFILLER_32_53 VPWR VGND sg13g2_decap_4
XFILLER_106_0 VPWR VGND sg13g2_decap_8
XFILLER_94_149 VPWR VGND sg13g2_decap_8
X_0604_ _0070_ VPWR _0071_ VGND Tile_X0Y0_W6END[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ sg13g2_o21ai_1
XFILLER_7_161 VPWR VGND sg13g2_decap_8
X_1653_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG7 Tile_X0Y1_S2BEGb[7]
+ VPWR VGND sg13g2_buf_1
X_1584_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG10 Tile_X0Y1_E6BEG[10]
+ VPWR VGND sg13g2_buf_1
X_0535_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q UIO_OUT_TT_PROJECT6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_85_127 VPWR VGND sg13g2_fill_2
X_0397_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_W1END[2]
+ Tile_X0Y0_W6END[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14
+ _0317_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux4_1
X_0466_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q Tile_X0Y0_W2MID[1]
+ Tile_X0Y0_W2END[1] Tile_X0Y0_W6END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG6
+ VPWR VGND sg13g2_mux4_1
XFILLER_93_193 VPWR VGND sg13g2_fill_2
X_1018_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_20 VPWR VGND sg13g2_fill_2
XFILLER_27_42 VPWR VGND sg13g2_fill_2
XFILLER_43_85 VPWR VGND sg13g2_fill_1
XFILLER_4_142 VPWR VGND sg13g2_fill_2
XFILLER_4_79 VPWR VGND sg13g2_decap_8
XFILLER_4_35 VPWR VGND sg13g2_decap_8
X_0518_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q UIO_OUT_TT_PROJECT6
+ UIO_OE_TT_PROJECT2 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG10 VPWR VGND sg13g2_mux4_1
XFILLER_58_105 VPWR VGND sg13g2_fill_1
X_1636_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG2 Tile_X0Y1_S1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1567_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb1 Tile_X0Y1_E2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_1498_ Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
XFILLER_104_14 VPWR VGND sg13g2_decap_8
X_0449_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2END[4] Tile_X0Y1_W6END[4] _0356_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb3 VPWR VGND sg13g2_mux4_1
XFILLER_81_152 VPWR VGND sg13g2_decap_8
XFILLER_72_196 VPWR VGND sg13g2_decap_4
XFILLER_57_171 VPWR VGND sg13g2_decap_4
XFILLER_54_51 VPWR VGND sg13g2_decap_8
XFILLER_54_62 VPWR VGND sg13g2_fill_2
XFILLER_54_84 VPWR VGND sg13g2_fill_2
X_1421_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG0 Tile_X0Y0_E2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1283_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1352_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0998_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1619_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData_O[17] VPWR VGND sg13g2_buf_1
XFILLER_39_160 VPWR VGND sg13g2_fill_2
XFILLER_54_196 VPWR VGND sg13g2_decap_4
XFILLER_24_54 VPWR VGND sg13g2_decap_4
XFILLER_108_165 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_4
X_0921_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_72 VPWR VGND sg13g2_fill_1
XFILLER_45_141 VPWR VGND sg13g2_fill_2
XFILLER_81_93 VPWR VGND sg13g2_decap_8
X_0783_ _0174_ _0173_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_nand2b_1
X_0852_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y1_W1END[1]
+ Tile_X0Y1_WW4END[13] Tile_X0Y1_WW4END[5] Tile_X0Y1_W6END[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
+ _0232_ VPWR VGND sg13g2_mux4_1
X_1335_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1404_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1266_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1197_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_177 VPWR VGND sg13g2_decap_8
XFILLER_19_21 VPWR VGND sg13g2_fill_2
XFILLER_51_74 VPWR VGND sg13g2_decap_8
X_1051_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1120_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0904_ VGND VPWR _0296_ _0266_ _0280_ _0279_ sg13g2_a21oi_1
X_0766_ _0154_ _0150_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ _0159_ VPWR VGND sg13g2_mux2_1
X_0697_ UO_OUT_TT_PROJECT6 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q _0128_ VPWR
+ VGND sg13g2_nor3_1
X_0835_ _0216_ VPWR UI_IN_TT_PROJECT1 VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q
+ _0218_ sg13g2_o21ai_1
X_1318_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_72_18 VPWR VGND sg13g2_fill_2
X_1249_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_62 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_51 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_84 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XFILLER_24_199 VPWR VGND sg13g2_fill_1
XANTENNA_95 VPWR VGND Tile_X0Y1_N2MID[7] sg13g2_antennanp
XANTENNA_40 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_73 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_101_171 VPWR VGND sg13g2_fill_1
XFILLER_102_91 VPWR VGND sg13g2_decap_8
XFILLER_15_122 VPWR VGND sg13g2_fill_1
X_0620_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q _0081_
+ _0082_ VPWR VGND sg13g2_nor2_1
X_0551_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q VPWR
+ _0024_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q
+ _0023_ sg13g2_o21ai_1
XFILLER_7_35 VPWR VGND sg13g2_decap_8
X_0482_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END2
+ UIO_OUT_TT_PROJECT0 Tile_X0Y0_S1END[2] UIO_OUT_TT_PROJECT5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG2 VPWR VGND sg13g2_mux4_1
X_1034_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1103_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_103 VPWR VGND sg13g2_fill_2
XFILLER_99_0 VPWR VGND sg13g2_decap_8
XFILLER_107_14 VPWR VGND sg13g2_decap_8
XFILLER_88_125 VPWR VGND sg13g2_fill_2
X_0818_ VGND VPWR _0200_ _0202_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG2
+ _0204_ sg13g2_a21oi_1
X_0749_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q UO_OUT_TT_PROJECT1
+ _0156_ UO_OUT_TT_PROJECT5 _0349_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG13 VPWR VGND sg13g2_mux4_1
XFILLER_12_125 VPWR VGND sg13g2_fill_1
XFILLER_16_22 VPWR VGND sg13g2_fill_2
XFILLER_32_87 VPWR VGND sg13g2_decap_4
XFILLER_87_191 VPWR VGND sg13g2_fill_1
XFILLER_92_7 VPWR VGND sg13g2_decap_4
X_0534_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q UIO_OUT_TT_PROJECT5
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG5 VPWR VGND sg13g2_mux4_1
X_0603_ _0070_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_nand2b_1
X_1652_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG6 Tile_X0Y1_S2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_1583_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG9 Tile_X0Y1_E6BEG[9]
+ VPWR VGND sg13g2_buf_1
X_0396_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_mux4_1
X_0465_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb6
+ Tile_X0Y0_S2MID[6] Tile_X0Y1_N2MID[6] Tile_X0Y0_S2END[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6 VPWR VGND sg13g2_mux4_1
X_1017_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_78_17 VPWR VGND sg13g2_fill_2
XFILLER_84_150 VPWR VGND sg13g2_fill_1
XFILLER_43_20 VPWR VGND sg13g2_fill_1
XFILLER_4_154 VPWR VGND sg13g2_decap_8
XFILLER_4_121 VPWR VGND sg13g2_decap_8
XFILLER_4_58 VPWR VGND sg13g2_decap_8
XFILLER_4_14 VPWR VGND sg13g2_decap_8
XFILLER_90_197 VPWR VGND sg13g2_fill_2
XFILLER_90_153 VPWR VGND sg13g2_fill_2
X_1497_ Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
X_0517_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG5 VPWR VGND sg13g2_mux4_1
X_1635_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG1 Tile_X0Y1_S1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1566_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb0 Tile_X0Y1_E2BEGb[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_81_164 VPWR VGND sg13g2_decap_8
X_0379_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END1 _0309_ VPWR VGND sg13g2_nor3_1
X_0448_ _0351_ _0354_ _0356_ VPWR VGND sg13g2_nor2b_1
XFILLER_13_34 VPWR VGND sg13g2_fill_1
XFILLER_49_139 VPWR VGND sg13g2_fill_1
XFILLER_72_142 VPWR VGND sg13g2_decap_8
XFILLER_70_62 VPWR VGND sg13g2_fill_1
X_1420_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG3 Tile_X0Y0_E1BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1351_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1282_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0997_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_19 VPWR VGND sg13g2_fill_2
X_1618_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData_O[16] VPWR VGND sg13g2_buf_1
X_1549_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG0 Tile_X0Y0_N4BEG[12]
+ VPWR VGND sg13g2_buf_1
XFILLER_75_18 VPWR VGND sg13g2_fill_2
XFILLER_91_17 VPWR VGND sg13g2_fill_1
XFILLER_39_172 VPWR VGND sg13g2_fill_1
XFILLER_108_144 VPWR VGND sg13g2_decap_8
XFILLER_105_91 VPWR VGND sg13g2_decap_8
X_0920_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_178 VPWR VGND sg13g2_fill_1
XFILLER_60_145 VPWR VGND sg13g2_fill_2
XANTENNA_130 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
X_0851_ _0228_ VPWR UI_IN_TT_PROJECT4 VGND _0229_ _0231_ sg13g2_o21ai_1
X_0782_ _0152_ _0148_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ _0173_ VPWR VGND sg13g2_mux2_1
XFILLER_53_4 VPWR VGND sg13g2_fill_2
X_1403_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1334_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1265_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_49 VPWR VGND sg13g2_decap_8
XFILLER_51_112 VPWR VGND sg13g2_decap_4
X_1196_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_10_24 VPWR VGND sg13g2_decap_4
XFILLER_19_55 VPWR VGND sg13g2_fill_2
X_1050_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0903_ Tile_X0Y1_W2END[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q _0279_ VPWR
+ VGND sg13g2_nor3_1
X_0834_ VPWR _0218_ _0217_ VGND sg13g2_inv_1
X_0696_ _0127_ _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_0765_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q UO_OUT_TT_PROJECT3
+ _0154_ _0158_ _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG11 VPWR VGND sg13g2_mux4_1
XFILLER_110_183 VPWR VGND sg13g2_decap_8
XFILLER_2_91 VPWR VGND sg13g2_decap_8
X_1317_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1248_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1179_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_96 VPWR VGND Tile_X0Y1_N2MID[7] sg13g2_antennanp
XANTENNA_52 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_21_45 VPWR VGND sg13g2_fill_2
XANTENNA_41 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_30 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_85 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XANTENNA_63 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_74 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_102_70 VPWR VGND sg13g2_decap_4
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_15_178 VPWR VGND sg13g2_fill_1
X_0550_ _0022_ VPWR _0023_ VGND Tile_X0Y0_W6END[9] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ sg13g2_o21ai_1
XFILLER_7_58 VPWR VGND sg13g2_decap_8
X_0481_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END1
+ UIO_OUT_TT_PROJECT3 Tile_X0Y0_S1END[1] UIO_OUT_TT_PROJECT6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG1 VPWR VGND sg13g2_mux4_1
X_1102_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_16_4 VPWR VGND sg13g2_fill_1
X_1033_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0817_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q _0203_
+ _0204_ VPWR VGND sg13g2_nor2_1
X_0679_ UO_OUT_TT_PROJECT0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q _0116_ VPWR
+ VGND sg13g2_nor3_1
X_0748_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0318_ Tile_X0Y0_S4END[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0156_ VPWR VGND sg13g2_mux4_1
XFILLER_12_148 VPWR VGND sg13g2_fill_2
XFILLER_94_129 VPWR VGND sg13g2_fill_2
XFILLER_73_84 VPWR VGND sg13g2_decap_4
XFILLER_85_7 VPWR VGND sg13g2_decap_8
X_1651_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG5 Tile_X0Y1_S2BEGb[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_98_81 VPWR VGND sg13g2_fill_2
X_0533_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q UIO_OUT_TT_PROJECT4
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG4 VPWR VGND sg13g2_mux4_1
X_0602_ VGND VPWR _0064_ _0067_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG2
+ _0069_ sg13g2_a21oi_1
X_0464_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q Tile_X0Y1_W2MID[1]
+ Tile_X0Y1_W2END[1] Tile_X0Y1_W6END[1] _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb6 VPWR VGND sg13g2_mux4_1
X_1582_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG8 Tile_X0Y1_E6BEG[8]
+ VPWR VGND sg13g2_buf_1
X_0395_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q Tile_X0Y1_W1END[2]
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14 Tile_X0Y1_W6END[6]
+ _0321_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END2
+ VPWR VGND sg13g2_mux4_1
X_1016_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_94_17 VPWR VGND sg13g2_decap_8
XFILLER_76_129 VPWR VGND sg13g2_fill_1
XFILLER_27_22 VPWR VGND sg13g2_fill_1
XFILLER_43_98 VPWR VGND sg13g2_fill_2
XFILLER_4_199 VPWR VGND sg13g2_fill_1
XFILLER_4_100 VPWR VGND sg13g2_decap_8
XFILLER_83_4 VPWR VGND sg13g2_fill_1
X_1634_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S1BEG0 Tile_X0Y1_S1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1496_ Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData_O[31] VPWR VGND sg13g2_buf_1
X_0516_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q UIO_OUT_TT_PROJECT5
+ UIO_OE_TT_PROJECT1 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG9 VPWR VGND sg13g2_mux4_1
X_0447_ _0355_ _0354_ _0351_ VPWR VGND sg13g2_nand2b_1
X_1565_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG7 Tile_X0Y1_E2BEG[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_49 VPWR VGND sg13g2_decap_8
X_0378_ _0308_ Tile_X0Y0_S1END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_13_79 VPWR VGND sg13g2_decap_4
XFILLER_72_176 VPWR VGND sg13g2_fill_2
XFILLER_54_86 VPWR VGND sg13g2_fill_1
XFILLER_110_92 VPWR VGND sg13g2_decap_8
X_1281_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1350_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_7 VPWR VGND sg13g2_decap_4
XFILLER_0_191 VPWR VGND sg13g2_decap_8
XFILLER_48_184 VPWR VGND sg13g2_fill_1
X_0996_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_0 VPWR VGND sg13g2_fill_1
X_1617_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameData_O[15] VPWR VGND sg13g2_buf_1
X_1548_ Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_11.A Tile_X0Y0_N4BEG[11] VPWR VGND sg13g2_buf_1
X_1479_ Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_108_123 VPWR VGND sg13g2_decap_8
XFILLER_105_70 VPWR VGND sg13g2_decap_8
XANTENNA_120 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XFILLER_65_52 VPWR VGND sg13g2_fill_2
XFILLER_60_113 VPWR VGND sg13g2_decap_8
XANTENNA_131 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
XFILLER_45_187 VPWR VGND sg13g2_fill_2
X_0850_ _0230_ VPWR _0231_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
+ _0154_ sg13g2_o21ai_1
XFILLER_45_198 VPWR VGND sg13g2_fill_2
X_1402_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0781_ VGND VPWR _0167_ _0170_ Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_9.A _0172_ sg13g2_a21oi_1
X_1333_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1264_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_28 VPWR VGND sg13g2_decap_8
X_1195_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0979_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_10_58 VPWR VGND sg13g2_fill_1
XFILLER_42_146 VPWR VGND sg13g2_decap_8
XFILLER_4_0 VPWR VGND sg13g2_decap_8
XFILLER_104_170 VPWR VGND sg13g2_decap_8
XFILLER_76_62 VPWR VGND sg13g2_fill_2
XFILLER_92_94 VPWR VGND sg13g2_fill_1
XFILLER_92_83 VPWR VGND sg13g2_decap_8
XFILLER_18_198 VPWR VGND sg13g2_fill_2
XFILLER_33_102 VPWR VGND sg13g2_decap_8
X_0902_ _0278_ _0265_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG0
+ VPWR VGND sg13g2_nand2b_1
X_0833_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q Tile_X0Y1_WW4END[1]
+ Tile_X0Y1_WW4END[9] Tile_X0Y1_W6END[1] Tile_X0Y1_W6END[9] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q
+ _0217_ VPWR VGND sg13g2_mux4_1
X_0695_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q
+ _0126_ _0125_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG5 _0348_ sg13g2_a221oi_1
XFILLER_37_0 VPWR VGND sg13g2_decap_4
X_0764_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q UO_OUT_TT_PROJECT2
+ _0153_ _0157_ _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG10 VPWR VGND sg13g2_mux4_1
XFILLER_110_162 VPWR VGND sg13g2_decap_8
XFILLER_2_70 VPWR VGND sg13g2_decap_8
X_1247_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1178_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1316_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_146 VPWR VGND sg13g2_decap_4
XANTENNA_20 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_31 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_97_28 VPWR VGND sg13g2_decap_8
XANTENNA_53 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_42 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_86 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XANTENNA_75 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_64 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_97 VPWR VGND Tile_X0Y1_N2MID[7] sg13g2_antennanp
XFILLER_101_140 VPWR VGND sg13g2_decap_4
XFILLER_97_39 VPWR VGND sg13g2_fill_2
XFILLER_62_42 VPWR VGND sg13g2_fill_1
XFILLER_30_149 VPWR VGND sg13g2_fill_1
X_0480_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END0
+ UIO_OUT_TT_PROJECT2 Tile_X0Y0_S1END[0] UIO_OUT_TT_PROJECT7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG0 VPWR VGND sg13g2_mux4_1
X_1032_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1101_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0816_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q Tile_X0Y1_W1END[2]
+ Tile_X0Y1_WW4END[14] Tile_X0Y1_W6END[6] _0156_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
+ _0203_ VPWR VGND sg13g2_mux4_1
X_0747_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT4 _0155_ _0356_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG12 VPWR VGND sg13g2_mux4_1
XFILLER_107_49 VPWR VGND sg13g2_decap_8
X_0678_ _0115_ _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_16_24 VPWR VGND sg13g2_fill_1
XFILLER_57_97 VPWR VGND sg13g2_decap_8
X_0601_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q _0068_
+ _0069_ VPWR VGND sg13g2_nor2_1
X_1650_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG4 Tile_X0Y1_S2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_1581_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG7 Tile_X0Y1_E6BEG[7]
+ VPWR VGND sg13g2_buf_1
X_0532_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y1_N4END[7]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG3 VPWR VGND sg13g2_mux4_1
XFILLER_78_171 VPWR VGND sg13g2_decap_4
X_0394_ VPWR VGND _0319_ _0320_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q
+ _0298_ _0321_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
+ sg13g2_a221oi_1
X_0463_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q Tile_X0Y1_N2MID[6]
+ Tile_X0Y1_N2END[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG6
+ Tile_X0Y0_S2MID[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q
+ _0002_ VPWR VGND sg13g2_mux4_1
X_1015_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_81 VPWR VGND sg13g2_decap_8
XFILLER_104_0 VPWR VGND sg13g2_decap_8
XFILLER_4_178 VPWR VGND sg13g2_decap_8
XFILLER_4_49 VPWR VGND sg13g2_decap_4
XFILLER_90_199 VPWR VGND sg13g2_fill_1
X_1633_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData_O[31] VPWR VGND sg13g2_buf_1
X_1564_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG6 Tile_X0Y1_E2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1495_ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData_O[30] VPWR VGND sg13g2_buf_1
XFILLER_104_28 VPWR VGND sg13g2_decap_8
X_0515_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG6 VPWR VGND sg13g2_mux4_1
X_0377_ VPWR _0307_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q
+ VGND sg13g2_inv_1
X_0446_ _0352_ _0353_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q
+ _0354_ VPWR VGND sg13g2_nand3_1
XFILLER_81_100 VPWR VGND sg13g2_fill_1
XFILLER_8_7 VPWR VGND sg13g2_decap_8
XFILLER_72_122 VPWR VGND sg13g2_fill_2
XFILLER_38_99 VPWR VGND sg13g2_fill_2
XFILLER_110_71 VPWR VGND sg13g2_decap_8
XFILLER_79_40 VPWR VGND sg13g2_decap_4
XFILLER_79_95 VPWR VGND sg13g2_fill_2
X_1280_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_63_199 VPWR VGND sg13g2_fill_1
X_0995_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_0 VPWR VGND sg13g2_fill_2
X_1547_ Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_10.A Tile_X0Y0_N4BEG[10] VPWR VGND sg13g2_buf_1
X_1616_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData_O[14] VPWR VGND sg13g2_buf_1
X_1478_ Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData_O[13] VPWR VGND sg13g2_buf_1
X_0429_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y0_W2MID[6]
+ Tile_X0Y0_W2END[6] Tile_X0Y0_W6END[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_108_179 VPWR VGND sg13g2_decap_4
XFILLER_108_102 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_49_76 VPWR VGND sg13g2_decap_4
XFILLER_65_97 VPWR VGND sg13g2_decap_8
XANTENNA_132 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
XANTENNA_110 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XANTENNA_121 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XFILLER_81_63 VPWR VGND sg13g2_fill_2
XFILLER_81_52 VPWR VGND sg13g2_decap_8
XFILLER_60_169 VPWR VGND sg13g2_decap_8
X_0780_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q _0171_
+ _0172_ VPWR VGND sg13g2_nor2_1
X_1401_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_39_4 VPWR VGND sg13g2_fill_1
X_1332_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1263_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1194_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_199 VPWR VGND sg13g2_fill_1
XFILLER_105_105 VPWR VGND sg13g2_decap_8
X_0978_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_105_149 VPWR VGND sg13g2_decap_8
XFILLER_86_19 VPWR VGND sg13g2_decap_4
XFILLER_19_57 VPWR VGND sg13g2_fill_1
XFILLER_19_79 VPWR VGND sg13g2_fill_1
XFILLER_27_100 VPWR VGND sg13g2_fill_2
XFILLER_27_199 VPWR VGND sg13g2_fill_1
XFILLER_18_122 VPWR VGND sg13g2_decap_4
X_0901_ _0276_ VPWR _0277_ VGND _0267_ _0269_ sg13g2_o21ai_1
X_0832_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q _0215_
+ _0216_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q
+ sg13g2_nand3b_1
X_0763_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q UO_OUT_TT_PROJECT1
+ _0152_ _0156_ _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG9 VPWR VGND sg13g2_mux4_1
XFILLER_110_141 VPWR VGND sg13g2_decap_8
X_0694_ UO_OUT_TT_PROJECT5 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q _0126_ VPWR
+ VGND sg13g2_nor3_1
X_1315_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1177_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1246_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_65 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_54 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_43 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_24_169 VPWR VGND sg13g2_fill_1
XANTENNA_21 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_32 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_10 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_108_7 VPWR VGND sg13g2_decap_8
XANTENNA_98 VPWR VGND Tile_X0Y1_N2MID[7] sg13g2_antennanp
XANTENNA_76 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_87 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XFILLER_21_47 VPWR VGND sg13g2_fill_1
XFILLER_7_49 VPWR VGND sg13g2_decap_4
XFILLER_97_139 VPWR VGND sg13g2_decap_4
XFILLER_11_80 VPWR VGND sg13g2_fill_2
X_1031_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1100_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_28 VPWR VGND sg13g2_decap_8
X_0815_ VGND VPWR Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
+ _0201_ _0202_ _0303_ sg13g2_a21oi_1
X_0746_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0325_ Tile_X0Y0_S4END[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q
+ _0155_ VPWR VGND sg13g2_mux4_1
XFILLER_96_183 VPWR VGND sg13g2_fill_2
XFILLER_96_161 VPWR VGND sg13g2_decap_4
X_0677_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y1_N1END[3]
+ UO_OUT_TT_PROJECT1 _0325_ UO_OUT_TT_PROJECT4 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG3 VPWR VGND sg13g2_mux4_1
X_1229_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_32_57 VPWR VGND sg13g2_fill_2
X_0531_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y1_N4END[6]
+ Tile_X0Y0_S4END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG2 VPWR VGND sg13g2_mux4_1
X_0600_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q Tile_X0Y0_W1END[2]
+ Tile_X0Y0_WW4END[14] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ _0068_ VPWR VGND sg13g2_mux4_1
X_1580_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG6 Tile_X0Y1_E6BEG[6]
+ VPWR VGND sg13g2_buf_1
XFILLER_78_150 VPWR VGND sg13g2_decap_4
X_0462_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q Tile_X0Y0_W1END[2]
+ Tile_X0Y0_W2MID[1] Tile_X0Y0_W2END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG6
+ VPWR VGND sg13g2_mux4_1
X_0393_ Tile_X0Y1_N1END[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q _0320_ VPWR
+ VGND sg13g2_nor3_1
X_1014_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_97_0 VPWR VGND sg13g2_decap_8
X_0729_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q UO_OUT_TT_PROJECT3
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12 UO_OUT_TT_PROJECT7
+ _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_84_197 VPWR VGND sg13g2_fill_2
XFILLER_4_135 VPWR VGND sg13g2_decap_8
XFILLER_108_60 VPWR VGND sg13g2_decap_8
XFILLER_4_28 VPWR VGND sg13g2_decap_8
XFILLER_17_90 VPWR VGND sg13g2_fill_1
XFILLER_90_7 VPWR VGND sg13g2_decap_8
X_1494_ Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData_O[29] VPWR VGND sg13g2_buf_1
X_0514_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q UIO_OUT_TT_PROJECT4
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG8 VPWR VGND sg13g2_mux4_1
X_1563_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG5 Tile_X0Y1_E2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_1632_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData_O[30] VPWR VGND sg13g2_buf_1
X_0445_ _0353_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
+ Tile_X0Y0_S2MID[3] VPWR VGND sg13g2_nand2_1
X_0376_ VPWR _0306_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ VGND sg13g2_inv_1
XFILLER_72_178 VPWR VGND sg13g2_fill_1
XFILLER_57_197 VPWR VGND sg13g2_fill_2
XFILLER_57_175 VPWR VGND sg13g2_fill_1
XFILLER_54_11 VPWR VGND sg13g2_fill_2
XFILLER_110_50 VPWR VGND sg13g2_decap_8
XFILLER_0_171 VPWR VGND sg13g2_decap_4
X_0994_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1546_ Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_9.A Tile_X0Y0_N4BEG[9] VPWR VGND sg13g2_buf_1
X_1477_ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_5_93 VPWR VGND sg13g2_decap_8
X_1615_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData_O[13] VPWR VGND sg13g2_buf_1
X_0428_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb1
+ Tile_X0Y0_S2MID[1] Tile_X0Y1_N2MID[1] Tile_X0Y0_S2END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1 VPWR VGND sg13g2_mux4_1
X_0359_ VPWR _0289_ Tile_X0Y0_W6END[3] VGND sg13g2_inv_1
XFILLER_54_112 VPWR VGND sg13g2_fill_2
XFILLER_54_178 VPWR VGND sg13g2_decap_8
XFILLER_24_36 VPWR VGND sg13g2_fill_1
XFILLER_108_158 VPWR VGND sg13g2_decap_8
XFILLER_65_32 VPWR VGND sg13g2_fill_2
XANTENNA_100 VPWR VGND UIO_OUT_TT_PROJECT0 sg13g2_antennanp
XANTENNA_133 VPWR VGND Tile_X0Y0_S4END[8] sg13g2_antennanp
XANTENNA_122 VPWR VGND Tile_X0Y0_S4END[11] sg13g2_antennanp
XANTENNA_111 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XFILLER_45_189 VPWR VGND sg13g2_fill_1
XFILLER_81_86 VPWR VGND sg13g2_decap_8
X_1400_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1331_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1262_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1193_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_137 VPWR VGND sg13g2_fill_2
X_0977_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1529_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb0 Tile_X0Y0_N2BEGb[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_76_86 VPWR VGND sg13g2_decap_4
XFILLER_76_64 VPWR VGND sg13g2_fill_1
X_0900_ VPWR VGND _0265_ _0271_ _0275_ _0266_ _0276_ _0273_ sg13g2_a221oi_1
XFILLER_33_148 VPWR VGND sg13g2_fill_2
X_0693_ _0125_ _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
X_0831_ _0157_ _0149_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q
+ _0215_ VPWR VGND sg13g2_mux2_1
X_0762_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q UO_OUT_TT_PROJECT0
+ _0151_ _0155_ _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG8 VPWR VGND sg13g2_mux4_1
XFILLER_110_120 VPWR VGND sg13g2_decap_8
X_1314_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_110_197 VPWR VGND sg13g2_fill_2
X_1176_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1245_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_99 VPWR VGND UIO_OUT_TT_PROJECT0 sg13g2_antennanp
XANTENNA_33 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_44 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_88 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XANTENNA_77 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_66 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_22 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_55 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_11 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_101_197 VPWR VGND sg13g2_fill_2
XFILLER_102_84 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_87_63 VPWR VGND sg13g2_decap_4
X_1030_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_181 VPWR VGND sg13g2_fill_1
X_0814_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14 _0002_
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q _0201_ VPWR
+ VGND sg13g2_mux2_1
X_0676_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q Tile_X0Y1_N1END[2]
+ UO_OUT_TT_PROJECT0 _0318_ UO_OUT_TT_PROJECT5 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG2 VPWR VGND sg13g2_mux4_1
X_0745_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q UO_OUT_TT_PROJECT3
+ _0154_ UO_OUT_TT_PROJECT7 _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG11 VPWR VGND sg13g2_mux4_1
X_1228_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1159_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_32_25 VPWR VGND sg13g2_fill_2
XFILLER_87_184 VPWR VGND sg13g2_decap_8
XFILLER_73_43 VPWR VGND sg13g2_decap_4
XFILLER_73_21 VPWR VGND sg13g2_fill_2
XFILLER_57_55 VPWR VGND sg13g2_decap_4
XFILLER_7_111 VPWR VGND sg13g2_decap_8
X_0530_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q Tile_X0Y1_N4END[5]
+ Tile_X0Y0_S4END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_7_199 VPWR VGND sg13g2_fill_1
XFILLER_93_110 VPWR VGND sg13g2_fill_1
X_0461_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q Tile_X0Y0_W2MID[2]
+ Tile_X0Y0_W2END[2] Tile_X0Y0_W6END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG5
+ VPWR VGND sg13g2_mux4_1
X_0392_ _0319_ _0318_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_1013_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_93 VPWR VGND sg13g2_decap_8
X_0659_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q _0110_
+ _0111_ _0114_ VPWR VGND sg13g2_nor3_1
X_0728_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT6 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13
+ _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_4_147 VPWR VGND sg13g2_decap_8
XFILLER_4_114 VPWR VGND sg13g2_decap_8
XFILLER_75_132 VPWR VGND sg13g2_fill_1
XFILLER_75_110 VPWR VGND sg13g2_fill_1
XFILLER_84_86 VPWR VGND sg13g2_fill_2
XFILLER_75_198 VPWR VGND sg13g2_fill_2
X_1631_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData_O[29] VPWR VGND sg13g2_buf_1
X_0513_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG7 VPWR VGND sg13g2_mux4_1
X_1493_ Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData_O[28] VPWR VGND sg13g2_buf_1
X_1562_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG4 Tile_X0Y1_E2BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0444_ _0352_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG3 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_nand2b_1
X_0375_ VPWR _0305_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ VGND sg13g2_inv_1
XFILLER_13_38 VPWR VGND sg13g2_fill_2
XFILLER_1_117 VPWR VGND sg13g2_fill_2
XFILLER_1_128 VPWR VGND sg13g2_fill_2
XFILLER_38_57 VPWR VGND sg13g2_decap_4
XFILLER_72_168 VPWR VGND sg13g2_fill_2
XFILLER_72_124 VPWR VGND sg13g2_fill_1
XFILLER_57_165 VPWR VGND sg13g2_fill_1
XFILLER_79_97 VPWR VGND sg13g2_fill_1
XFILLER_95_52 VPWR VGND sg13g2_decap_8
XFILLER_48_132 VPWR VGND sg13g2_decap_8
X_0993_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1614_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData_O[12] VPWR VGND sg13g2_buf_1
X_1545_ Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_8.A Tile_X0Y0_N4BEG[8] VPWR VGND sg13g2_buf_1
X_1476_ Tile_X0Y0_FrameData[11] Tile_X0Y0_FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_5_72 VPWR VGND sg13g2_decap_8
X_0427_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y1_W2MID[6]
+ Tile_X0Y1_W2END[6] Tile_X0Y1_W6END[6] _0342_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb1 VPWR VGND sg13g2_mux4_1
X_0358_ VPWR _0288_ Tile_X0Y0_W6END[2] VGND sg13g2_inv_1
XFILLER_39_198 VPWR VGND sg13g2_fill_2
XFILLER_54_135 VPWR VGND sg13g2_fill_1
XFILLER_108_137 VPWR VGND sg13g2_decap_8
XFILLER_49_45 VPWR VGND sg13g2_decap_4
XFILLER_105_84 VPWR VGND sg13g2_decap_8
XFILLER_65_11 VPWR VGND sg13g2_fill_1
XANTENNA_112 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XANTENNA_101 VPWR VGND UIO_OUT_TT_PROJECT0 sg13g2_antennanp
XANTENNA_123 VPWR VGND Tile_X0Y0_S4END[14] sg13g2_antennanp
XANTENNA_134 VPWR VGND Tile_X0Y0_S4END[12] sg13g2_antennanp
XFILLER_107_181 VPWR VGND sg13g2_decap_8
X_1330_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1261_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_105 VPWR VGND sg13g2_decap_8
X_1192_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_72_0 VPWR VGND sg13g2_fill_1
X_0976_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1528_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG7 Tile_X0Y0_N2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1459_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG10 Tile_X0Y0_EE4BEG[10]
+ VPWR VGND sg13g2_buf_1
XFILLER_19_48 VPWR VGND sg13g2_decap_8
XFILLER_27_135 VPWR VGND sg13g2_fill_2
XFILLER_50_160 VPWR VGND sg13g2_decap_8
XFILLER_51_24 VPWR VGND sg13g2_fill_2
XFILLER_104_184 VPWR VGND sg13g2_fill_1
XFILLER_33_116 VPWR VGND sg13g2_fill_1
X_0830_ _0213_ _0214_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q
+ UI_IN_TT_PROJECT0 VPWR VGND sg13g2_mux2_1
X_0692_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q
+ _0124_ _0123_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG4 _0355_ sg13g2_a221oi_1
X_0761_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q UO_OUT_TT_PROJECT7
+ _0150_ _0154_ _0356_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG7 VPWR VGND sg13g2_mux4_1
XFILLER_110_176 VPWR VGND sg13g2_decap_8
XFILLER_2_84 VPWR VGND sg13g2_decap_8
X_1313_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1244_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_105 VPWR VGND sg13g2_decap_4
X_1175_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0959_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_34 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_78 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_89 VPWR VGND Tile_X0Y1_FrameData[8] sg13g2_antennanp
XANTENNA_23 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_12 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_67 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_45 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_56 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_102_63 VPWR VGND sg13g2_decap_8
XFILLER_30_119 VPWR VGND sg13g2_decap_4
XFILLER_2_0 VPWR VGND sg13g2_decap_8
XFILLER_11_82 VPWR VGND sg13g2_fill_1
XFILLER_14_171 VPWR VGND sg13g2_fill_2
X_0813_ _0200_ _0199_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_35_0 VPWR VGND sg13g2_decap_4
X_0675_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q Tile_X0Y1_N1END[1]
+ UO_OUT_TT_PROJECT3 _0311_ UO_OUT_TT_PROJECT6 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG1 VPWR VGND sg13g2_mux4_1
X_0744_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0007_ Tile_X0Y0_S4END[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q
+ _0154_ VPWR VGND sg13g2_mux4_1
X_1158_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1227_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1089_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_16_38 VPWR VGND sg13g2_fill_2
XFILLER_79_119 VPWR VGND sg13g2_decap_8
X_0460_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb5
+ Tile_X0Y0_S2MID[5] Tile_X0Y1_N2MID[5] Tile_X0Y0_S2END[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_7_178 VPWR VGND sg13g2_decap_4
XFILLER_22_81 VPWR VGND sg13g2_fill_2
X_1012_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0391_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y0_W1END[2]
+ Tile_X0Y0_W6END[10] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14
+ _0317_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q _0318_
+ VPWR VGND sg13g2_mux4_1
XFILLER_93_199 VPWR VGND sg13g2_fill_1
XFILLER_8_50 VPWR VGND sg13g2_decap_4
X_0727_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q UO_OUT_TT_PROJECT1
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14 UO_OUT_TT_PROJECT5
+ _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG1
+ VPWR VGND sg13g2_mux4_1
X_0658_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q _0112_
+ _0113_ VPWR VGND sg13g2_nor2b_1
X_0589_ _0057_ VPWR _0058_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ _0013_ sg13g2_o21ai_1
XFILLER_84_199 VPWR VGND sg13g2_fill_1
XFILLER_108_95 VPWR VGND sg13g2_decap_8
X_1630_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData_O[28] VPWR VGND sg13g2_buf_1
X_0512_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q UIO_OUT_TT_PROJECT7
+ UIO_OE_TT_PROJECT3 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG7 VPWR VGND sg13g2_mux4_1
X_1492_ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData_O[27] VPWR VGND sg13g2_buf_1
X_1561_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG3 Tile_X0Y1_E2BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_3_192 VPWR VGND sg13g2_decap_8
X_0443_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q _0350_
+ _0351_ VPWR VGND sg13g2_nor2_1
X_0374_ VPWR _0304_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q
+ VGND sg13g2_inv_1
XFILLER_81_125 VPWR VGND sg13g2_decap_4
XFILLER_66_166 VPWR VGND sg13g2_fill_2
XFILLER_66_144 VPWR VGND sg13g2_decap_4
XFILLER_66_122 VPWR VGND sg13g2_fill_1
XFILLER_80_180 VPWR VGND sg13g2_fill_1
XFILLER_57_199 VPWR VGND sg13g2_fill_1
XFILLER_110_85 VPWR VGND sg13g2_decap_8
XFILLER_102_0 VPWR VGND sg13g2_decap_8
XFILLER_48_177 VPWR VGND sg13g2_decap_8
X_0992_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1544_ Tile_X0Y1_N4END[15] Tile_X0Y0_N4BEG[7] VPWR VGND sg13g2_buf_1
X_1613_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameData_O[11] VPWR VGND sg13g2_buf_1
X_1475_ Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData_O[10] VPWR VGND sg13g2_buf_1
X_0357_ VPWR _0287_ Tile_X0Y0_W6END[1] VGND sg13g2_inv_1
X_0426_ _0337_ _0340_ _0342_ VPWR VGND sg13g2_nor2b_1
XFILLER_108_116 VPWR VGND sg13g2_decap_8
XFILLER_6_7 VPWR VGND sg13g2_decap_8
XFILLER_105_63 VPWR VGND sg13g2_decap_8
XANTENNA_102 VPWR VGND UIO_OUT_TT_PROJECT0 sg13g2_antennanp
XFILLER_65_34 VPWR VGND sg13g2_fill_1
XANTENNA_113 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XANTENNA_124 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
XFILLER_107_160 VPWR VGND sg13g2_decap_8
X_1260_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1191_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_139 VPWR VGND sg13g2_fill_1
XFILLER_65_0 VPWR VGND sg13g2_decap_8
X_0975_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1527_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG6 Tile_X0Y0_N2BEG[6]
+ VPWR VGND sg13g2_buf_1
XFILLER_105_119 VPWR VGND sg13g2_decap_4
X_1458_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG9 Tile_X0Y0_EE4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_1389_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0409_ Tile_X0Y1_N2MID[0] Tile_X0Y1_N2END[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
+ _0329_ VPWR VGND sg13g2_mux2_1
XFILLER_27_114 VPWR VGND sg13g2_decap_4
XFILLER_51_47 VPWR VGND sg13g2_decap_4
XFILLER_104_163 VPWR VGND sg13g2_decap_8
XFILLER_76_22 VPWR VGND sg13g2_fill_2
X_0760_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q UO_OUT_TT_PROJECT6
+ _0149_ _0153_ _0349_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG6 VPWR VGND sg13g2_mux4_1
X_0691_ UO_OUT_TT_PROJECT4 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q _0124_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_37_4 VPWR VGND sg13g2_fill_1
XFILLER_110_199 VPWR VGND sg13g2_fill_1
XFILLER_110_155 VPWR VGND sg13g2_decap_8
XFILLER_2_63 VPWR VGND sg13g2_decap_8
X_1312_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1243_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1174_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_139 VPWR VGND sg13g2_decap_8
XANTENNA_13 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0958_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_35 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0889_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
+ _0265_ VPWR VGND sg13g2_nor2b_1
XANTENNA_24 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_79 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_57 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_68 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_46 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_101_122 VPWR VGND sg13g2_fill_1
XFILLER_102_42 VPWR VGND sg13g2_decap_8
XFILLER_101_199 VPWR VGND sg13g2_fill_1
XFILLER_87_21 VPWR VGND sg13g2_fill_1
X_0812_ _0152_ _0148_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q
+ _0199_ VPWR VGND sg13g2_mux2_1
X_0743_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT6 _0153_ _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG10 VPWR VGND sg13g2_mux4_1
X_0674_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q Tile_X0Y1_N1END[0]
+ UO_OUT_TT_PROJECT2 _0007_ UO_OUT_TT_PROJECT7 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_96_197 VPWR VGND sg13g2_fill_2
X_1157_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1226_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1088_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_120 VPWR VGND sg13g2_fill_1
XFILLER_106_7 VPWR VGND sg13g2_decap_8
XFILLER_11_164 VPWR VGND sg13g2_decap_4
XFILLER_98_42 VPWR VGND sg13g2_decap_8
X_0390_ VPWR VGND _0315_ _0316_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q
+ _0288_ _0317_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q
+ sg13g2_a221oi_1
X_1011_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_93_101 VPWR VGND sg13g2_decap_8
XFILLER_78_197 VPWR VGND sg13g2_fill_2
XFILLER_78_175 VPWR VGND sg13g2_fill_1
X_0726_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT4 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15
+ _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG0
+ VPWR VGND sg13g2_mux4_1
X_0657_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y0_W1END[3]
+ Tile_X0Y0_WW4END[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q
+ _0112_ VPWR VGND sg13g2_mux4_1
X_0588_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q _0056_
+ _0057_ VPWR VGND sg13g2_and2_1
XFILLER_27_38 VPWR VGND sg13g2_decap_4
X_1209_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_74 VPWR VGND sg13g2_decap_8
X_0511_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG8 VPWR VGND sg13g2_mux4_1
X_1560_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG2 Tile_X0Y1_E2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1491_ Tile_X0Y0_FrameData[26] Tile_X0Y0_FrameData_O[26] VPWR VGND sg13g2_buf_1
XFILLER_3_171 VPWR VGND sg13g2_decap_8
X_0442_ Tile_X0Y1_N2MID[3] Tile_X0Y1_N2END[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
+ _0350_ VPWR VGND sg13g2_mux2_1
X_0373_ VPWR _0303_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q
+ VGND sg13g2_inv_1
XFILLER_81_159 VPWR VGND sg13g2_fill_1
XFILLER_66_178 VPWR VGND sg13g2_fill_1
XFILLER_95_0 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_fill_1
X_0709_ UO_OUT_TT_PROJECT2 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q _0136_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_72_115 VPWR VGND sg13g2_decap_8
XFILLER_110_64 VPWR VGND sg13g2_decap_8
XFILLER_54_58 VPWR VGND sg13g2_decap_4
XFILLER_95_21 VPWR VGND sg13g2_decap_8
XFILLER_63_126 VPWR VGND sg13g2_decap_4
X_0991_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1474_ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[9] VPWR VGND sg13g2_buf_1
X_1543_ Tile_X0Y1_N4END[14] Tile_X0Y0_N4BEG[6] VPWR VGND sg13g2_buf_1
X_1612_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_10_0 VPWR VGND sg13g2_decap_8
X_0425_ _0341_ _0340_ _0337_ VPWR VGND sg13g2_nand2b_1
XFILLER_24_17 VPWR VGND sg13g2_fill_2
XFILLER_105_42 VPWR VGND sg13g2_decap_8
XANTENNA_103 VPWR VGND UIO_OUT_TT_PROJECT0 sg13g2_antennanp
XANTENNA_114 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XANTENNA_125 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
XFILLER_53_170 VPWR VGND sg13g2_decap_8
XFILLER_39_8 VPWR VGND sg13g2_decap_8
X_1190_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_90 VPWR VGND sg13g2_decap_8
X_0974_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1526_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG5 Tile_X0Y0_N2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_1457_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG8 Tile_X0Y0_EE4BEG[8]
+ VPWR VGND sg13g2_buf_1
XFILLER_58_0 VPWR VGND sg13g2_decap_8
X_0408_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q Tile_X0Y0_W2MID[7]
+ Tile_X0Y0_W2END[7] Tile_X0Y0_W6END[8] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG0
+ VPWR VGND sg13g2_mux4_1
XFILLER_27_137 VPWR VGND sg13g2_fill_1
X_1388_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_50_184 VPWR VGND sg13g2_fill_1
XFILLER_104_197 VPWR VGND sg13g2_fill_2
XFILLER_18_115 VPWR VGND sg13g2_decap_8
XFILLER_92_11 VPWR VGND sg13g2_fill_1
X_0690_ _0123_ _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_41_92 VPWR VGND sg13g2_fill_1
X_1311_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_110_134 VPWR VGND sg13g2_decap_8
XFILLER_2_42 VPWR VGND sg13g2_decap_8
X_1242_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1173_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_47 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_25 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_14 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_36 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0957_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_69 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0888_ VPWR ENA_TT_PROJECT _0264_ VGND sg13g2_inv_1
XANTENNA_58 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_1509_ Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
XFILLER_102_21 VPWR VGND sg13g2_decap_8
XFILLER_102_98 VPWR VGND sg13g2_fill_1
XFILLER_99_7 VPWR VGND sg13g2_decap_8
XFILLER_14_173 VPWR VGND sg13g2_fill_1
XFILLER_36_92 VPWR VGND sg13g2_fill_2
X_0673_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W2END[0] Tile_X0Y1_W2MID[0] _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG7 VPWR VGND sg13g2_mux4_1
X_0811_ VGND VPWR _0194_ _0196_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG1
+ _0198_ sg13g2_a21oi_1
XFILLER_52_80 VPWR VGND sg13g2_fill_1
XFILLER_52_91 VPWR VGND sg13g2_decap_8
X_0742_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0311_ Tile_X0Y0_S4END[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q
+ _0153_ VPWR VGND sg13g2_mux4_1
XFILLER_96_165 VPWR VGND sg13g2_fill_1
X_1087_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1156_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1225_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_198 VPWR VGND sg13g2_fill_2
XFILLER_57_14 VPWR VGND sg13g2_decap_4
XFILLER_98_21 VPWR VGND sg13g2_decap_8
X_1010_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_30 VPWR VGND sg13g2_fill_1
X_0656_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q VPWR
+ _0111_ VGND Tile_X0Y0_WW4END[15] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q
+ sg13g2_o21ai_1
X_0725_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q
+ _0146_ _0145_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb7 _0334_ sg13g2_a221oi_1
XFILLER_40_0 VPWR VGND sg13g2_decap_8
XFILLER_84_168 VPWR VGND sg13g2_decap_4
X_0587_ _0056_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5 VPWR VGND sg13g2_nand2b_1
X_1208_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1139_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_4_128 VPWR VGND sg13g2_decap_8
XFILLER_108_53 VPWR VGND sg13g2_decap_8
XFILLER_90_149 VPWR VGND sg13g2_decap_4
X_1490_ Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData_O[25] VPWR VGND sg13g2_buf_1
X_0510_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q UIO_OUT_TT_PROJECT6
+ UIO_OE_TT_PROJECT2 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_3_161 VPWR VGND sg13g2_decap_8
X_0441_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q Tile_X0Y0_W2MID[4]
+ Tile_X0Y0_W2END[4] Tile_X0Y0_W6END[11] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG3
+ VPWR VGND sg13g2_mux4_1
X_0372_ VPWR _0302_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q
+ VGND sg13g2_inv_1
XFILLER_88_0 VPWR VGND sg13g2_fill_1
X_0639_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y0_W1END[0]
+ Tile_X0Y0_WW4END[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q
+ _0097_ VPWR VGND sg13g2_mux4_1
X_0708_ _0135_ _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_72_149 VPWR VGND sg13g2_fill_2
XFILLER_110_43 VPWR VGND sg13g2_decap_8
XFILLER_110_21 VPWR VGND sg13g2_decap_8
XFILLER_0_164 VPWR VGND sg13g2_decap_8
X_0990_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1611_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[9] VPWR VGND sg13g2_buf_1
X_1473_ Tile_X0Y0_FrameData[8] Tile_X0Y0_FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_5_86 VPWR VGND sg13g2_decap_8
XFILLER_5_53 VPWR VGND sg13g2_fill_2
XFILLER_5_42 VPWR VGND sg13g2_decap_8
X_1542_ Tile_X0Y1_N4END[13] Tile_X0Y0_N4BEG[5] VPWR VGND sg13g2_buf_1
X_0424_ _0338_ _0339_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q
+ _0340_ VPWR VGND sg13g2_nand3_1
XFILLER_105_21 VPWR VGND sg13g2_decap_8
XFILLER_105_98 VPWR VGND sg13g2_decap_8
XANTENNA_104 VPWR VGND UIO_OUT_TT_PROJECT0 sg13g2_antennanp
XANTENNA_115 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XANTENNA_126 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
XFILLER_53_160 VPWR VGND sg13g2_decap_8
XFILLER_107_195 VPWR VGND sg13g2_decap_4
XFILLER_44_160 VPWR VGND sg13g2_fill_1
XFILLER_71_90 VPWR VGND sg13g2_fill_2
X_0973_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1525_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG4 Tile_X0Y0_N2BEG[4]
+ VPWR VGND sg13g2_buf_1
X_1456_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG7 Tile_X0Y0_EE4BEG[7]
+ VPWR VGND sg13g2_buf_1
X_0407_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W6END[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15
+ _0324_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG3
+ VPWR VGND sg13g2_mux4_1
X_1387_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_26_182 VPWR VGND sg13g2_fill_1
XFILLER_110_113 VPWR VGND sg13g2_decap_8
XFILLER_2_21 VPWR VGND sg13g2_decap_8
X_1310_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1241_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_98 VPWR VGND sg13g2_decap_8
X_1172_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_0956_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_70_0 VPWR VGND sg13g2_fill_2
XANTENNA_15 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_26 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_59 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_48 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_37 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0887_ _0263_ VPWR _0264_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q
+ _0254_ sg13g2_o21ai_1
X_1439_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG2 Tile_X0Y0_E6BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1508_ Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
XFILLER_46_38 VPWR VGND sg13g2_decap_4
XFILLER_102_77 VPWR VGND sg13g2_decap_8
XFILLER_23_163 VPWR VGND sg13g2_fill_1
XFILLER_87_67 VPWR VGND sg13g2_fill_2
XFILLER_87_56 VPWR VGND sg13g2_decap_8
X_0810_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q _0197_
+ _0198_ VPWR VGND sg13g2_nor2_1
X_0672_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q Tile_X0Y1_W1END[2]
+ Tile_X0Y1_W2END[1] Tile_X0Y1_W2MID[1] _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG6 VPWR VGND sg13g2_mux4_1
X_0741_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q UO_OUT_TT_PROJECT1
+ _0152_ UO_OUT_TT_PROJECT5 _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG9 VPWR VGND sg13g2_mux4_1
XFILLER_96_199 VPWR VGND sg13g2_fill_1
X_1224_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1086_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1155_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0939_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_144 VPWR VGND sg13g2_fill_2
XFILLER_73_47 VPWR VGND sg13g2_fill_1
XFILLER_57_37 VPWR VGND sg13g2_fill_1
XFILLER_7_104 VPWR VGND sg13g2_fill_2
XFILLER_98_77 VPWR VGND sg13g2_decap_4
XFILLER_7_137 VPWR VGND sg13g2_decap_8
XFILLER_78_199 VPWR VGND sg13g2_fill_1
XFILLER_78_100 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_69_144 VPWR VGND sg13g2_fill_2
XFILLER_69_122 VPWR VGND sg13g2_fill_1
X_0655_ Tile_X0Y0_W6END[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q
+ _0110_ VPWR VGND sg13g2_nor2b_1
X_0586_ VPWR _0055_ _0054_ VGND sg13g2_inv_1
X_0724_ UO_OUT_TT_PROJECT7 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q _0146_ VPWR
+ VGND sg13g2_nor3_1
X_1207_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1069_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1138_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_32 VPWR VGND sg13g2_fill_2
XFILLER_4_107 VPWR VGND sg13g2_decap_8
X_0440_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q Tile_X0Y0_W2MID[5]
+ Tile_X0Y0_W2END[5] Tile_X0Y0_W6END[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG2
+ VPWR VGND sg13g2_mux4_1
X_0371_ VPWR _0301_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q
+ VGND sg13g2_inv_1
X_0707_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q
+ _0134_ _0133_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb1 _0341_ sg13g2_a221oi_1
X_0569_ VGND VPWR Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q
+ _0039_ _0040_ _0038_ sg13g2_a21oi_1
X_0638_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q VPWR
+ _0096_ VGND Tile_X0Y0_WW4END[12] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q
+ sg13g2_o21ai_1
XFILLER_110_99 VPWR VGND sg13g2_decap_8
XFILLER_95_45 VPWR VGND sg13g2_decap_8
XFILLER_0_198 VPWR VGND sg13g2_fill_2
XFILLER_5_21 VPWR VGND sg13g2_decap_8
X_1610_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameData_O[8] VPWR VGND sg13g2_buf_1
X_1472_ Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_5_65 VPWR VGND sg13g2_decap_8
X_1541_ Tile_X0Y1_N4END[12] Tile_X0Y0_N4BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_39_125 VPWR VGND sg13g2_fill_1
X_0423_ _0339_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
+ Tile_X0Y0_S2MID[1] VPWR VGND sg13g2_nand2_1
XFILLER_105_77 VPWR VGND sg13g2_decap_8
XFILLER_49_38 VPWR VGND sg13g2_decap_8
XFILLER_49_49 VPWR VGND sg13g2_fill_2
XANTENNA_105 VPWR VGND UIO_OUT_TT_PROJECT0 sg13g2_antennanp
XANTENNA_116 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XFILLER_38_191 VPWR VGND sg13g2_fill_1
XANTENNA_127 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
XFILLER_14_63 VPWR VGND sg13g2_fill_2
XFILLER_107_174 VPWR VGND sg13g2_decap_8
XFILLER_100_0 VPWR VGND sg13g2_decap_8
X_0972_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1524_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG3 Tile_X0Y0_N2BEG[3]
+ VPWR VGND sg13g2_buf_1
X_0406_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_mux4_1
X_1455_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG6 Tile_X0Y0_EE4BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1386_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_17 VPWR VGND sg13g2_decap_8
XFILLER_104_177 VPWR VGND sg13g2_decap_8
XFILLER_104_144 VPWR VGND sg13g2_decap_4
XFILLER_4_7 VPWR VGND sg13g2_decap_8
XFILLER_104_199 VPWR VGND sg13g2_fill_1
XFILLER_33_109 VPWR VGND sg13g2_decap_8
XFILLER_110_169 VPWR VGND sg13g2_decap_8
XFILLER_2_77 VPWR VGND sg13g2_decap_8
X_1240_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1171_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_66_91 VPWR VGND sg13g2_decap_8
XFILLER_32_131 VPWR VGND sg13g2_fill_2
X_0955_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_16 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0886_ _0262_ VPWR _0263_ VGND _0255_ _0257_ sg13g2_o21ai_1
XFILLER_32_153 VPWR VGND sg13g2_fill_1
XANTENNA_27 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_38 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_49 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_63_0 VPWR VGND sg13g2_fill_1
X_1507_ Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
XFILLER_101_169 VPWR VGND sg13g2_fill_2
X_1438_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG1 Tile_X0Y0_E6BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1369_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_56 VPWR VGND sg13g2_decap_8
XFILLER_62_38 VPWR VGND sg13g2_decap_4
XFILLER_11_86 VPWR VGND sg13g2_fill_2
XFILLER_14_131 VPWR VGND sg13g2_fill_1
X_0740_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0318_ Tile_X0Y0_S4END[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q
+ _0152_ VPWR VGND sg13g2_mux4_1
X_0671_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q Tile_X0Y1_W1END[1]
+ Tile_X0Y1_W2END[2] Tile_X0Y1_W2MID[2] _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_35_4 VPWR VGND sg13g2_fill_1
X_1154_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1223_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1085_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0938_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0869_ _0243_ VPWR UI_IN_TT_PROJECT7 VGND _0244_ _0246_ sg13g2_o21ai_1
XFILLER_11_134 VPWR VGND sg13g2_fill_2
XFILLER_98_56 VPWR VGND sg13g2_fill_1
XFILLER_8_54 VPWR VGND sg13g2_fill_1
XFILLER_8_43 VPWR VGND sg13g2_decap_8
XFILLER_8_21 VPWR VGND sg13g2_decap_8
XFILLER_6_171 VPWR VGND sg13g2_decap_8
X_0723_ _0145_ _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_nand2b_1
X_0654_ VGND VPWR UIO_IN_TT_PROJECT6 _0109_ _0108_ sg13g2_or2_1
X_0585_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q VPWR
+ _0054_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q
+ _0053_ sg13g2_o21ai_1
X_1137_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1206_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1068_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_104_7 VPWR VGND sg13g2_decap_8
XFILLER_108_88 VPWR VGND sg13g2_decap_8
XFILLER_33_95 VPWR VGND sg13g2_decap_8
X_0370_ VPWR _0300_ Tile_X0Y1_W6END[0] VGND sg13g2_inv_1
XFILLER_3_185 VPWR VGND sg13g2_decap_8
XFILLER_81_129 VPWR VGND sg13g2_fill_2
XFILLER_81_118 VPWR VGND sg13g2_decap_8
XFILLER_66_148 VPWR VGND sg13g2_fill_1
X_0706_ UO_OUT_TT_PROJECT1 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q _0134_ VPWR
+ VGND sg13g2_nor3_1
X_0499_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q UIO_OUT_TT_PROJECT7
+ UIO_OE_TT_PROJECT7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb7 VPWR VGND sg13g2_mux4_1
X_0568_ _0011_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ _0039_ VPWR VGND sg13g2_mux2_1
X_0637_ Tile_X0Y0_W6END[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q
+ _0095_ VPWR VGND sg13g2_nor2b_1
XFILLER_57_104 VPWR VGND sg13g2_decap_4
XFILLER_80_173 VPWR VGND sg13g2_decap_8
XFILLER_110_78 VPWR VGND sg13g2_decap_8
X_1540_ Tile_X0Y1_N4END[11] Tile_X0Y0_N4BEG[3] VPWR VGND sg13g2_buf_1
X_1471_ Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData_O[6] VPWR VGND sg13g2_buf_1
X_0422_ _0338_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG1 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_62_140 VPWR VGND sg13g2_fill_1
XFILLER_47_170 VPWR VGND sg13g2_decap_8
XFILLER_108_109 VPWR VGND sg13g2_decap_8
XFILLER_93_0 VPWR VGND sg13g2_fill_2
X_1669_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG3 Tile_X0Y1_S4BEG[15]
+ VPWR VGND sg13g2_buf_1
XFILLER_105_56 VPWR VGND sg13g2_decap_8
XANTENNA_106 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XFILLER_81_59 VPWR VGND sg13g2_decap_4
XANTENNA_117 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XANTENNA_128 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
XFILLER_53_184 VPWR VGND sg13g2_fill_1
XFILLER_107_153 VPWR VGND sg13g2_decap_8
XFILLER_14_86 VPWR VGND sg13g2_decap_4
XFILLER_39_94 VPWR VGND sg13g2_fill_2
X_0971_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1523_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG2 Tile_X0Y0_N2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1454_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG5 Tile_X0Y0_EE4BEG[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_27_107 VPWR VGND sg13g2_decap_8
X_0405_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15 Tile_X0Y1_W6END[7]
+ _0328_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END3
+ VPWR VGND sg13g2_mux4_1
X_1385_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_41_110 VPWR VGND sg13g2_fill_2
XFILLER_41_73 VPWR VGND sg13g2_fill_2
XFILLER_110_148 VPWR VGND sg13g2_decap_8
XFILLER_2_56 VPWR VGND sg13g2_fill_2
X_1170_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0954_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_17 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0885_ _0261_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q
+ _0262_ VPWR VGND sg13g2_nor2b_1
XANTENNA_39 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_32_198 VPWR VGND sg13g2_fill_2
XANTENNA_28 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XFILLER_101_115 VPWR VGND sg13g2_decap_8
XFILLER_99_143 VPWR VGND sg13g2_fill_2
X_1437_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG0 Tile_X0Y0_E6BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_56_0 VPWR VGND sg13g2_decap_8
X_1506_ Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
XFILLER_102_35 VPWR VGND sg13g2_decap_8
X_1368_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1299_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_11_21 VPWR VGND sg13g2_decap_4
XFILLER_11_43 VPWR VGND sg13g2_fill_2
X_0670_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q Tile_X0Y1_W1END[0]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W2MID[3] _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG4 VPWR VGND sg13g2_mux4_1
X_1084_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1153_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1222_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_102 VPWR VGND sg13g2_decap_8
X_0937_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0799_ _0188_ _0187_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_20_179 VPWR VGND sg13g2_fill_1
X_0868_ _0245_ VPWR _0246_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0151_ sg13g2_o21ai_1
XFILLER_7_106 VPWR VGND sg13g2_fill_1
XFILLER_98_35 VPWR VGND sg13g2_decap_8
XFILLER_97_7 VPWR VGND sg13g2_decap_8
X_0653_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q _0105_
+ _0106_ _0109_ VPWR VGND sg13g2_nor3_1
XFILLER_6_161 VPWR VGND sg13g2_decap_8
X_0722_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q
+ _0144_ _0143_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb6 _0341_ sg13g2_a221oi_1
XFILLER_69_168 VPWR VGND sg13g2_fill_2
X_0584_ _0052_ VPWR _0053_ VGND Tile_X0Y0_W6END[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ sg13g2_o21ai_1
X_1067_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1136_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_0 VPWR VGND sg13g2_decap_4
X_1205_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_67 VPWR VGND sg13g2_decap_8
XFILLER_108_34 VPWR VGND sg13g2_fill_1
XFILLER_3_142 VPWR VGND sg13g2_fill_2
X_0636_ VGND VPWR Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q
+ _0092_ UIO_IN_TT_PROJECT3 _0094_ sg13g2_a21oi_1
X_0705_ _0133_ _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
X_0498_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q UIO_OUT_TT_PROJECT6
+ UIO_OE_TT_PROJECT6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb6 VPWR VGND sg13g2_mux4_1
X_0567_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q VPWR
+ _0038_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q
+ _0037_ sg13g2_o21ai_1
XFILLER_110_57 VPWR VGND sg13g2_decap_8
X_1119_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_14 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_71_141 VPWR VGND sg13g2_fill_1
XFILLER_28_41 VPWR VGND sg13g2_fill_1
X_1470_ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_60_50 VPWR VGND sg13g2_fill_1
X_0421_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q _0336_
+ _0337_ VPWR VGND sg13g2_nor2_1
XFILLER_54_108 VPWR VGND sg13g2_decap_4
XFILLER_62_163 VPWR VGND sg13g2_fill_1
XFILLER_86_0 VPWR VGND sg13g2_fill_2
X_0619_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y0_WW4END[0]
+ Tile_X0Y0_WW4END[8] _0014_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q _0081_ VPWR
+ VGND sg13g2_mux4_1
X_1668_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG2 Tile_X0Y1_S4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_1599_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG13 Tile_X0Y1_EE4BEG[13]
+ VPWR VGND sg13g2_buf_1
XFILLER_105_35 VPWR VGND sg13g2_decap_8
XANTENNA_107 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XANTENNA_118 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XANTENNA_129 VPWR VGND Tile_X0Y1_FrameData[31] sg13g2_antennanp
XFILLER_38_160 VPWR VGND sg13g2_fill_2
XFILLER_45_119 VPWR VGND sg13g2_fill_2
XFILLER_14_65 VPWR VGND sg13g2_fill_1
XFILLER_53_196 VPWR VGND sg13g2_decap_4
X_0970_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1522_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG1 Tile_X0Y0_N2BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1453_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG4 Tile_X0Y0_EE4BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0404_ VPWR VGND _0326_ _0327_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q
+ _0297_ _0328_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a221oi_1
X_1384_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_130 VPWR VGND sg13g2_fill_2
XFILLER_104_157 VPWR VGND sg13g2_fill_2
XFILLER_41_122 VPWR VGND sg13g2_fill_2
XFILLER_41_63 VPWR VGND sg13g2_decap_4
XFILLER_110_127 VPWR VGND sg13g2_decap_8
XFILLER_2_35 VPWR VGND sg13g2_decap_8
XANTENNA_29 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
XANTENNA_18 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0953_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0884_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q _0259_
+ _0260_ _0261_ VPWR VGND sg13g2_nor3_1
XFILLER_99_199 VPWR VGND sg13g2_fill_1
X_1436_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb7 Tile_X0Y0_E2BEGb[7]
+ VPWR VGND sg13g2_buf_1
X_1505_ Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_1367_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_14 VPWR VGND sg13g2_decap_8
X_1298_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_11_55 VPWR VGND sg13g2_fill_1
XFILLER_36_85 VPWR VGND sg13g2_decap_8
XFILLER_14_199 VPWR VGND sg13g2_fill_1
XFILLER_52_84 VPWR VGND sg13g2_decap_8
XFILLER_96_103 VPWR VGND sg13g2_fill_2
X_1221_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1083_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1152_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0936_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0798_ _0154_ _0150_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q
+ _0187_ VPWR VGND sg13g2_mux2_1
X_0867_ _0245_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_nand2b_1
X_1419_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG2 Tile_X0Y0_E1BEG[2]
+ VPWR VGND sg13g2_buf_1
XFILLER_57_18 VPWR VGND sg13g2_fill_2
XFILLER_98_14 VPWR VGND sg13g2_decap_8
XFILLER_7_118 VPWR VGND sg13g2_fill_2
XFILLER_22_32 VPWR VGND sg13g2_fill_1
XFILLER_47_62 VPWR VGND sg13g2_fill_2
XFILLER_47_84 VPWR VGND sg13g2_fill_2
XFILLER_47_95 VPWR VGND sg13g2_fill_2
X_0652_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q _0107_
+ _0108_ VPWR VGND sg13g2_nor2b_1
X_0583_ _0052_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_nand2b_1
XFILLER_6_195 VPWR VGND sg13g2_decap_4
X_0721_ UO_OUT_TT_PROJECT6 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q _0144_ VPWR
+ VGND sg13g2_nor3_1
X_1204_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1066_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1135_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0919_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_46 VPWR VGND sg13g2_decap_8
XFILLER_75_128 VPWR VGND sg13g2_decap_4
XFILLER_75_106 VPWR VGND sg13g2_decap_4
XFILLER_33_42 VPWR VGND sg13g2_fill_2
XFILLER_3_154 VPWR VGND sg13g2_decap_8
XFILLER_3_121 VPWR VGND sg13g2_decap_8
XFILLER_74_150 VPWR VGND sg13g2_decap_8
X_0566_ _0036_ VPWR _0037_ VGND Tile_X0Y0_W6END[11] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ sg13g2_o21ai_1
X_0635_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q _0093_
+ _0094_ VPWR VGND sg13g2_nor2_1
X_0704_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q
+ _0132_ _0131_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb0 _0334_ sg13g2_a221oi_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
X_0497_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q UIO_OUT_TT_PROJECT5
+ UIO_OE_TT_PROJECT5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb5 VPWR VGND sg13g2_mux4_1
XFILLER_57_139 VPWR VGND sg13g2_fill_1
XFILLER_110_36 VPWR VGND sg13g2_decap_8
XFILLER_110_14 VPWR VGND sg13g2_decap_8
X_1049_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_197 VPWR VGND sg13g2_fill_2
X_1118_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_59 VPWR VGND sg13g2_fill_2
XFILLER_0_157 VPWR VGND sg13g2_decap_8
XFILLER_48_139 VPWR VGND sg13g2_decap_8
XFILLER_56_183 VPWR VGND sg13g2_fill_2
XFILLER_28_97 VPWR VGND sg13g2_decap_4
XFILLER_71_197 VPWR VGND sg13g2_fill_2
XFILLER_5_79 VPWR VGND sg13g2_decap_8
XFILLER_5_35 VPWR VGND sg13g2_decap_8
X_0420_ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2END[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
+ _0336_ VPWR VGND sg13g2_mux2_1
XFILLER_93_2 VPWR VGND sg13g2_fill_1
XFILLER_79_0 VPWR VGND sg13g2_fill_2
XFILLER_105_14 VPWR VGND sg13g2_decap_8
X_0618_ _0079_ VPWR _0080_ VGND Tile_X0Y0_W6END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q
+ sg13g2_o21ai_1
X_0549_ _0022_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_nand2b_1
X_1667_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG1 Tile_X0Y1_S4BEG[13]
+ VPWR VGND sg13g2_buf_1
X_1598_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG12 Tile_X0Y1_EE4BEG[12]
+ VPWR VGND sg13g2_buf_1
XANTENNA_108 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XFILLER_81_17 VPWR VGND sg13g2_fill_1
XANTENNA_119 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XFILLER_107_199 VPWR VGND sg13g2_fill_1
XFILLER_107_188 VPWR VGND sg13g2_decap_8
XFILLER_107_133 VPWR VGND sg13g2_fill_1
XFILLER_39_96 VPWR VGND sg13g2_fill_1
XFILLER_55_40 VPWR VGND sg13g2_fill_1
XFILLER_55_84 VPWR VGND sg13g2_fill_2
X_1521_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG0 Tile_X0Y0_N2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1452_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG3 Tile_X0Y0_EE4BEG[3]
+ VPWR VGND sg13g2_buf_1
X_0403_ Tile_X0Y1_N1END[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q _0327_ VPWR
+ VGND sg13g2_nor3_1
X_1383_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_164 VPWR VGND sg13g2_fill_1
XFILLER_25_65 VPWR VGND sg13g2_decap_4
XFILLER_25_87 VPWR VGND sg13g2_fill_1
XFILLER_41_42 VPWR VGND sg13g2_decap_8
XFILLER_110_106 VPWR VGND sg13g2_decap_8
XFILLER_9_0 VPWR VGND sg13g2_decap_8
XFILLER_2_14 VPWR VGND sg13g2_decap_8
XFILLER_2_58 VPWR VGND sg13g2_fill_1
X_0952_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_19 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_1504_ Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
X_0883_ Tile_X0Y1_W2END[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q _0260_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_99_145 VPWR VGND sg13g2_fill_1
X_1435_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb6 Tile_X0Y0_E2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_1366_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_123 VPWR VGND sg13g2_fill_2
X_1297_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_7 VPWR VGND sg13g2_decap_8
XFILLER_96_126 VPWR VGND sg13g2_fill_1
X_1151_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1220_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1082_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0935_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_126 VPWR VGND sg13g2_fill_1
X_0866_ _0244_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q VPWR VGND
+ sg13g2_nand2b_1
XFILLER_61_0 VPWR VGND sg13g2_decap_8
X_0797_ VGND VPWR _0181_ _0184_ Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_11.A _0186_ sg13g2_a21oi_1
XFILLER_87_148 VPWR VGND sg13g2_fill_2
X_1418_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG1 Tile_X0Y0_E1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1349_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_11_126 VPWR VGND sg13g2_fill_2
X_0720_ _0143_ _0002_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_nand2b_1
X_0651_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q Tile_X0Y0_W1END[2]
+ Tile_X0Y0_WW4END[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q
+ _0107_ VPWR VGND sg13g2_mux4_1
X_0582_ VGND VPWR _0046_ _0049_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG0
+ _0051_ sg13g2_a21oi_1
XFILLER_6_185 VPWR VGND sg13g2_decap_4
X_1134_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1203_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1065_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_14 VPWR VGND sg13g2_fill_1
X_0918_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0849_ _0230_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_nand2b_1
XFILLER_68_29 VPWR VGND sg13g2_fill_2
XFILLER_17_22 VPWR VGND sg13g2_fill_2
XFILLER_109_0 VPWR VGND sg13g2_fill_2
XFILLER_3_100 VPWR VGND sg13g2_decap_8
XFILLER_3_199 VPWR VGND sg13g2_fill_1
X_0703_ UO_OUT_TT_PROJECT0 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q _0132_ VPWR
+ VGND sg13g2_nor3_1
X_0496_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q UIO_OUT_TT_PROJECT4
+ UIO_OE_TT_PROJECT4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb4 VPWR VGND sg13g2_mux4_1
X_0565_ _0036_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_nand2b_1
X_0634_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q Tile_X0Y0_WW4END[3]
+ Tile_X0Y0_WW4END[11] _0011_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q _0093_ VPWR
+ VGND sg13g2_mux4_1
X_1117_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1048_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_7 VPWR VGND sg13g2_decap_8
XFILLER_71_121 VPWR VGND sg13g2_fill_1
XFILLER_56_195 VPWR VGND sg13g2_decap_4
Xclkbuf_1_0__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_0__leaf_Tile_X0Y1_UserCLK
+ VPWR VGND sg13g2_buf_8
XFILLER_5_58 VPWR VGND sg13g2_decap_8
XFILLER_5_14 VPWR VGND sg13g2_decap_8
XFILLER_39_118 VPWR VGND sg13g2_decap_8
XFILLER_47_184 VPWR VGND sg13g2_fill_1
XFILLER_47_195 VPWR VGND sg13g2_decap_4
XFILLER_62_198 VPWR VGND sg13g2_fill_2
X_1666_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG0 Tile_X0Y1_S4BEG[12]
+ VPWR VGND sg13g2_buf_1
X_0617_ VGND VPWR _0291_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q
+ _0079_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q sg13g2_a21oi_1
X_0548_ _0019_ _0021_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG0
+ VPWR VGND sg13g2_nor2_1
X_0479_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q Tile_X0Y1_W1END[0]
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12 Tile_X0Y1_W6END[4]
+ _0010_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END0
+ VPWR VGND sg13g2_mux4_1
X_1597_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG11 Tile_X0Y1_EE4BEG[11]
+ VPWR VGND sg13g2_buf_1
XANTENNA_109 VPWR VGND Tile_X0Y0_S2MID[3] sg13g2_antennanp
XFILLER_107_112 VPWR VGND sg13g2_decap_8
XFILLER_107_167 VPWR VGND sg13g2_decap_8
XFILLER_107_145 VPWR VGND sg13g2_decap_4
XFILLER_71_62 VPWR VGND sg13g2_fill_2
XFILLER_44_165 VPWR VGND sg13g2_decap_4
XFILLER_44_198 VPWR VGND sg13g2_fill_2
X_1520_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG3 Tile_X0Y0_N1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_65_7 VPWR VGND sg13g2_decap_4
X_1451_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG2 Tile_X0Y0_EE4BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0402_ _0326_ _0325_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
X_1382_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_132 VPWR VGND sg13g2_fill_1
XFILLER_35_198 VPWR VGND sg13g2_fill_2
XFILLER_104_148 VPWR VGND sg13g2_fill_1
XFILLER_104_126 VPWR VGND sg13g2_fill_1
X_1649_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG3 Tile_X0Y1_S2BEGb[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_25_55 VPWR VGND sg13g2_decap_8
XFILLER_106_91 VPWR VGND sg13g2_decap_8
X_0951_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0882_ _0259_ _0258_ _0305_ _0306_ Tile_X0Y1_W2END[5] VPWR VGND sg13g2_a22oi_1
XFILLER_99_124 VPWR VGND sg13g2_fill_2
X_1503_ Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
X_1434_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb5 Tile_X0Y0_E2BEGb[5]
+ VPWR VGND sg13g2_buf_1
X_1365_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1296_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_49 VPWR VGND sg13g2_decap_8
XFILLER_23_102 VPWR VGND sg13g2_decap_4
XFILLER_87_17 VPWR VGND sg13g2_decap_4
XFILLER_14_124 VPWR VGND sg13g2_decap_8
XFILLER_14_179 VPWR VGND sg13g2_fill_2
X_1150_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1081_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0934_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_161 VPWR VGND sg13g2_decap_8
XFILLER_20_116 VPWR VGND sg13g2_decap_4
X_0865_ _0243_ _0242_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_nand2b_1
X_1417_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E1BEG0 Tile_X0Y0_E1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0796_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q _0185_
+ _0186_ VPWR VGND sg13g2_nor2_1
XFILLER_54_0 VPWR VGND sg13g2_decap_8
X_1348_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1279_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_11_105 VPWR VGND sg13g2_decap_4
XFILLER_98_49 VPWR VGND sg13g2_decap_8
XFILLER_93_108 VPWR VGND sg13g2_fill_2
XFILLER_103_81 VPWR VGND sg13g2_fill_1
XFILLER_103_70 VPWR VGND sg13g2_decap_8
XFILLER_47_86 VPWR VGND sg13g2_fill_1
XFILLER_8_36 VPWR VGND sg13g2_decap_8
XFILLER_8_14 VPWR VGND sg13g2_decap_8
X_0650_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q VPWR
+ _0106_ VGND Tile_X0Y0_WW4END[14] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q
+ sg13g2_o21ai_1
X_0581_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q _0050_
+ _0051_ VPWR VGND sg13g2_nor2_1
X_1064_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_77_160 VPWR VGND sg13g2_fill_1
X_1133_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1202_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0917_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0848_ _0229_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q VPWR VGND
+ sg13g2_nand2b_1
X_0779_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q Tile_X0Y1_W1END[1]
+ Tile_X0Y1_W6END[9] Tile_X0Y1_WW4END[1] _0157_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ _0171_ VPWR VGND sg13g2_mux4_1
XFILLER_83_152 VPWR VGND sg13g2_decap_8
XFILLER_3_178 VPWR VGND sg13g2_decap_8
XFILLER_74_51 VPWR VGND sg13g2_decap_8
XFILLER_58_41 VPWR VGND sg13g2_decap_4
XFILLER_95_7 VPWR VGND sg13g2_decap_8
X_0633_ _0091_ VPWR _0092_ VGND Tile_X0Y0_W6END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q
+ sg13g2_o21ai_1
X_0702_ _0131_ _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_nand2b_1
X_0495_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q UIO_OUT_TT_PROJECT3
+ UIO_OE_TT_PROJECT3 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb3 VPWR VGND sg13g2_mux4_1
X_0564_ _0033_ _0035_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N4BEG2
+ VPWR VGND sg13g2_nor2_1
XFILLER_57_108 VPWR VGND sg13g2_fill_1
X_1047_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1116_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_0_81 VPWR VGND sg13g2_fill_2
XFILLER_17_0 VPWR VGND sg13g2_decap_4
XFILLER_80_199 VPWR VGND sg13g2_fill_1
XFILLER_71_199 VPWR VGND sg13g2_fill_1
XFILLER_71_166 VPWR VGND sg13g2_fill_2
XFILLER_109_80 VPWR VGND sg13g2_decap_8
XFILLER_62_111 VPWR VGND sg13g2_decap_4
X_1665_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG3 Tile_X0Y1_S4BEG[11]
+ VPWR VGND sg13g2_buf_1
X_1596_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG10 Tile_X0Y1_EE4BEG[10]
+ VPWR VGND sg13g2_buf_1
X_0616_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0325_ Tile_X0Y0_S4END[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_mux4_1
XFILLER_105_49 VPWR VGND sg13g2_decap_8
X_0547_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q _0020_
+ _0021_ VPWR VGND sg13g2_nor2_1
X_0478_ VPWR VGND _0008_ _0009_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q
+ _0300_ _0010_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_a221oi_1
XFILLER_53_177 VPWR VGND sg13g2_decap_8
XFILLER_30_45 VPWR VGND sg13g2_decap_4
XFILLER_30_67 VPWR VGND sg13g2_fill_2
XFILLER_39_65 VPWR VGND sg13g2_fill_1
XFILLER_39_87 VPWR VGND sg13g2_decap_8
XFILLER_55_75 VPWR VGND sg13g2_decap_4
XFILLER_55_86 VPWR VGND sg13g2_fill_1
XFILLER_55_97 VPWR VGND sg13g2_fill_2
X_1450_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG1 Tile_X0Y0_EE4BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_58_7 VPWR VGND sg13g2_fill_1
XFILLER_96_71 VPWR VGND sg13g2_decap_4
X_0401_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q Tile_X0Y0_W1END[3]
+ Tile_X0Y0_W6END[11] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15
+ _0324_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q _0325_
+ VPWR VGND sg13g2_mux4_1
X_1381_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_84_0 VPWR VGND sg13g2_decap_8
X_1648_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG2 Tile_X0Y1_S2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_1579_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG5 Tile_X0Y1_E6BEG[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_26_144 VPWR VGND sg13g2_fill_1
XFILLER_106_70 VPWR VGND sg13g2_decap_8
XFILLER_103_171 VPWR VGND sg13g2_decap_8
XFILLER_2_49 VPWR VGND sg13g2_decap_8
XFILLER_17_177 VPWR VGND sg13g2_fill_2
X_0950_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0881_ _0258_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_S2MID[2] VPWR VGND sg13g2_nand2b_1
X_1433_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb4 Tile_X0Y0_E2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_1502_ Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
XFILLER_102_28 VPWR VGND sg13g2_decap_8
X_1364_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1295_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_98 VPWR VGND sg13g2_fill_1
X_1080_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_77_40 VPWR VGND sg13g2_decap_8
X_0933_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0864_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q Tile_X0Y1_W1END[3]
+ Tile_X0Y1_WW4END[15] Tile_X0Y1_WW4END[7] Tile_X0Y1_W6END[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0242_ VPWR VGND sg13g2_mux4_1
X_0795_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q Tile_X0Y1_W1END[3]
+ Tile_X0Y1_W6END[11] Tile_X0Y1_WW4END[3] _0155_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ _0185_ VPWR VGND sg13g2_mux4_1
X_1347_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1416_ clknet_1_0__leaf_Tile_X0Y1_UserCLK CLK_TT_PROJECT VPWR VGND sg13g2_buf_1
X_1278_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_11_128 VPWR VGND sg13g2_fill_1
XFILLER_98_28 VPWR VGND sg13g2_decap_8
XFILLER_86_150 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_fill_1
XFILLER_47_43 VPWR VGND sg13g2_fill_2
XFILLER_10_161 VPWR VGND sg13g2_fill_2
XFILLER_10_150 VPWR VGND sg13g2_decap_8
XFILLER_6_154 VPWR VGND sg13g2_decap_8
XFILLER_6_121 VPWR VGND sg13g2_decap_4
XFILLER_84_109 VPWR VGND sg13g2_decap_8
X_0580_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q Tile_X0Y0_W1END[0]
+ Tile_X0Y0_WW4END[12] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG8 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ _0050_ VPWR VGND sg13g2_mux4_1
XFILLER_40_7 VPWR VGND sg13g2_decap_4
X_1201_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_197 VPWR VGND sg13g2_fill_2
XFILLER_92_153 VPWR VGND sg13g2_fill_2
XFILLER_92_131 VPWR VGND sg13g2_fill_1
X_1063_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1132_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0916_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_27 VPWR VGND sg13g2_fill_1
X_0847_ _0228_ _0227_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_nand2b_1
X_0778_ _0169_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q
+ _0170_ VPWR VGND sg13g2_nor2b_1
XFILLER_83_120 VPWR VGND sg13g2_decap_8
XFILLER_83_197 VPWR VGND sg13g2_fill_2
XFILLER_17_46 VPWR VGND sg13g2_fill_2
XFILLER_109_2 VPWR VGND sg13g2_fill_1
XFILLER_3_135 VPWR VGND sg13g2_decap_8
XFILLER_58_75 VPWR VGND sg13g2_fill_2
X_0632_ VGND VPWR _0294_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q
+ _0091_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q sg13g2_a21oi_1
X_0563_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q _0034_
+ _0035_ VPWR VGND sg13g2_nor2_1
X_0701_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q
+ _0130_ _0129_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG7 _0334_ sg13g2_a221oi_1
X_0494_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q UIO_OUT_TT_PROJECT2
+ UIO_OE_TT_PROJECT2 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb2 VPWR VGND sg13g2_mux4_1
XFILLER_110_28 VPWR VGND sg13g2_decap_4
X_1046_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_134 VPWR VGND sg13g2_decap_4
X_1115_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_178 VPWR VGND sg13g2_fill_2
XFILLER_69_30 VPWR VGND sg13g2_fill_2
XFILLER_60_43 VPWR VGND sg13g2_decap_8
XFILLER_5_49 VPWR VGND sg13g2_decap_4
X_0546_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q Tile_X0Y0_W1END[0]
+ Tile_X0Y0_WW4END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG8 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ _0020_ VPWR VGND sg13g2_mux4_1
X_1664_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG2 Tile_X0Y1_S4BEG[10]
+ VPWR VGND sg13g2_buf_1
X_1595_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG9 Tile_X0Y1_EE4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_0615_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0318_ Tile_X0Y0_S4END[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_mux4_1
XFILLER_105_28 VPWR VGND sg13g2_decap_8
X_0477_ Tile_X0Y1_N1END[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q _0009_ VPWR
+ VGND sg13g2_nor3_1
X_1029_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0400_ VPWR VGND _0322_ _0323_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q
+ _0289_ _0324_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a221oi_1
X_1380_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_77_0 VPWR VGND sg13g2_decap_8
X_0529_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y1_N4END[4]
+ Tile_X0Y0_S4END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG0 VPWR VGND sg13g2_mux4_1
X_1647_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG1 Tile_X0Y1_S2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_1578_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG4 Tile_X0Y1_E6BEG[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_41_56 VPWR VGND sg13g2_decap_8
XFILLER_41_115 VPWR VGND sg13g2_fill_2
XFILLER_41_67 VPWR VGND sg13g2_fill_1
XFILLER_2_28 VPWR VGND sg13g2_decap_8
XFILLER_82_63 VPWR VGND sg13g2_fill_1
X_0880_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q VPWR
+ _0257_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0256_ sg13g2_o21ai_1
X_1501_ Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
X_1432_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb3 Tile_X0Y0_E2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_1363_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1294_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_120 VPWR VGND sg13g2_fill_2
XFILLER_36_78 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
X_0932_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0863_ _0241_ VPWR UI_IN_TT_PROJECT6 VGND _0237_ _0239_ sg13g2_o21ai_1
X_0794_ _0183_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q
+ _0184_ VPWR VGND sg13g2_nor2b_1
XFILLER_95_140 VPWR VGND sg13g2_fill_2
XFILLER_3_93 VPWR VGND sg13g2_decap_8
X_1415_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1346_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1277_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_6_199 VPWR VGND sg13g2_fill_1
XFILLER_6_100 VPWR VGND sg13g2_decap_8
XFILLER_12_91 VPWR VGND sg13g2_fill_1
X_1200_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1062_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1131_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0915_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_39 VPWR VGND sg13g2_decap_8
X_0846_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q Tile_X0Y1_W1END[0]
+ Tile_X0Y1_WW4END[12] Tile_X0Y1_WW4END[4] Tile_X0Y1_W6END[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
+ _0227_ VPWR VGND sg13g2_mux4_1
X_0777_ VGND VPWR Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ _0341_ _0169_ _0168_ sg13g2_a21oi_1
X_1329_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_114 VPWR VGND sg13g2_decap_8
XFILLER_58_98 VPWR VGND sg13g2_decap_8
XFILLER_3_147 VPWR VGND sg13g2_decap_8
X_0700_ UO_OUT_TT_PROJECT7 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q _0130_ VPWR
+ VGND sg13g2_nor3_1
X_0562_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q Tile_X0Y0_W1END[2]
+ Tile_X0Y0_WW4END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ _0034_ VPWR VGND sg13g2_mux4_1
X_0631_ VGND VPWR Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q
+ _0088_ UIO_IN_TT_PROJECT2 _0090_ sg13g2_a21oi_1
X_0493_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q UIO_OUT_TT_PROJECT1
+ UIO_OE_TT_PROJECT1 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb1 VPWR VGND sg13g2_mux4_1
X_1114_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1045_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_94 VPWR VGND sg13g2_fill_1
X_0829_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q _0211_
+ _0212_ _0214_ VPWR VGND sg13g2_nor3_1
XFILLER_56_165 VPWR VGND sg13g2_fill_1
XFILLER_107_0 VPWR VGND sg13g2_decap_8
XFILLER_5_28 VPWR VGND sg13g2_decap_8
X_1663_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG1 Tile_X0Y1_S4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_0545_ VGND VPWR Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q
+ _0018_ _0019_ _0017_ sg13g2_a21oi_1
X_0476_ _0008_ _0007_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_22_0 VPWR VGND sg13g2_decap_4
X_1594_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG8 Tile_X0Y1_EE4BEG[8]
+ VPWR VGND sg13g2_buf_1
X_0614_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0311_ Tile_X0Y0_S4END[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_mux4_1
X_1028_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_126 VPWR VGND sg13g2_decap_8
XFILLER_100_7 VPWR VGND sg13g2_decap_8
XFILLER_30_69 VPWR VGND sg13g2_fill_1
XFILLER_71_43 VPWR VGND sg13g2_fill_2
XFILLER_35_157 VPWR VGND sg13g2_fill_2
XFILLER_6_93 VPWR VGND sg13g2_decap_8
X_1646_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG0 Tile_X0Y1_S2BEGb[0]
+ VPWR VGND sg13g2_buf_1
X_0528_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q UIO_OUT_TT_PROJECT3
+ UIO_OE_TT_PROJECT7 _0014_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG15
+ VPWR VGND sg13g2_mux4_1
X_0459_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y1_W2MID[2]
+ Tile_X0Y1_W2END[2] Tile_X0Y1_W6END[2] _0001_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb5 VPWR VGND sg13g2_mux4_1
X_1577_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG3 Tile_X0Y1_E6BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_66_98 VPWR VGND sg13g2_decap_8
XFILLER_66_32 VPWR VGND sg13g2_decap_4
X_1500_ Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
XFILLER_99_105 VPWR VGND sg13g2_fill_2
X_1431_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb2 Tile_X0Y0_E2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_1362_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1293_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1629_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData_O[27] VPWR VGND sg13g2_buf_1
XFILLER_52_78 VPWR VGND sg13g2_fill_2
X_0931_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0862_ _0241_ _0240_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_0793_ VGND VPWR Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ _0355_ _0183_ _0182_ sg13g2_a21oi_1
XFILLER_3_72 VPWR VGND sg13g2_decap_8
X_1414_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1345_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1276_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_28 VPWR VGND sg13g2_fill_2
XFILLER_6_189 VPWR VGND sg13g2_fill_1
XFILLER_6_178 VPWR VGND sg13g2_decap_8
X_1130_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_199 VPWR VGND sg13g2_fill_1
X_1061_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0914_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0845_ _0225_ _0226_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q
+ UI_IN_TT_PROJECT3 VPWR VGND sg13g2_mux2_1
X_0776_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q VPWR
+ _0168_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
XFILLER_52_0 VPWR VGND sg13g2_decap_8
XFILLER_83_199 VPWR VGND sg13g2_fill_1
XFILLER_83_166 VPWR VGND sg13g2_fill_2
X_1328_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1259_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_111 VPWR VGND sg13g2_fill_1
XFILLER_59_196 VPWR VGND sg13g2_decap_4
XFILLER_90_97 VPWR VGND sg13g2_fill_1
X_0492_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q UIO_OUT_TT_PROJECT0
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb0 VPWR VGND sg13g2_mux4_1
X_0561_ VGND VPWR Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q
+ _0032_ _0033_ _0031_ sg13g2_a21oi_1
X_0630_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q _0089_
+ _0090_ VPWR VGND sg13g2_nor2_1
X_1044_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1113_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0828_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y1_WW4END[0]
+ Tile_X0Y1_WW4END[8] Tile_X0Y1_W6END[0] Tile_X0Y1_W6END[8] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q
+ _0213_ VPWR VGND sg13g2_mux4_1
X_0759_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q UO_OUT_TT_PROJECT5
+ _0148_ _0152_ _0342_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_56_122 VPWR VGND sg13g2_fill_2
XFILLER_0_107 VPWR VGND sg13g2_fill_1
XFILLER_71_114 VPWR VGND sg13g2_decap_8
XFILLER_56_199 VPWR VGND sg13g2_fill_1
XFILLER_56_188 VPWR VGND sg13g2_decap_8
XFILLER_109_94 VPWR VGND sg13g2_decap_8
XFILLER_69_98 VPWR VGND sg13g2_fill_2
XFILLER_69_32 VPWR VGND sg13g2_fill_1
XFILLER_47_166 VPWR VGND sg13g2_fill_1
XFILLER_47_177 VPWR VGND sg13g2_decap_8
XFILLER_47_188 VPWR VGND sg13g2_decap_8
XFILLER_47_199 VPWR VGND sg13g2_fill_1
X_1662_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG0 Tile_X0Y1_S4BEG[8]
+ VPWR VGND sg13g2_buf_1
X_0613_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0007_ Tile_X0Y0_S4END[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_mux4_1
X_0544_ _0014_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ _0018_ VPWR VGND sg13g2_mux2_1
X_0475_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q Tile_X0Y0_W1END[0]
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_W6END[8]
+ _0006_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q _0007_
+ VPWR VGND sg13g2_mux4_1
X_1593_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG7 Tile_X0Y1_EE4BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1027_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_53_103 VPWR VGND sg13g2_decap_4
XFILLER_14_38 VPWR VGND sg13g2_fill_1
XFILLER_107_138 VPWR VGND sg13g2_decap_8
XFILLER_107_105 VPWR VGND sg13g2_decap_8
XFILLER_29_144 VPWR VGND sg13g2_fill_2
XFILLER_29_199 VPWR VGND sg13g2_fill_1
XFILLER_44_158 VPWR VGND sg13g2_fill_2
XFILLER_106_193 VPWR VGND sg13g2_decap_8
XFILLER_106_182 VPWR VGND sg13g2_fill_2
XFILLER_96_96 VPWR VGND sg13g2_decap_8
XFILLER_104_119 VPWR VGND sg13g2_decap_8
XFILLER_6_72 VPWR VGND sg13g2_decap_8
X_1645_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG7 Tile_X0Y1_S2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1576_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG2 Tile_X0Y1_E6BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0527_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q
+ _0014_ VPWR VGND sg13g2_mux4_1
X_0389_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END2 _0316_ VPWR VGND sg13g2_nor3_1
X_0458_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2END[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG5
+ Tile_X0Y0_S2MID[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q
+ _0001_ VPWR VGND sg13g2_mux4_1
XFILLER_106_84 VPWR VGND sg13g2_decap_8
XFILLER_17_125 VPWR VGND sg13g2_fill_1
XFILLER_17_147 VPWR VGND sg13g2_decap_4
X_1430_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEGb1 Tile_X0Y0_E2BEGb[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_56_7 VPWR VGND sg13g2_decap_8
X_1361_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1292_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_0 VPWR VGND sg13g2_decap_8
X_1559_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG1 Tile_X0Y1_E2BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1628_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameData_O[26] VPWR VGND sg13g2_buf_1
XFILLER_100_199 VPWR VGND sg13g2_fill_1
XFILLER_14_117 VPWR VGND sg13g2_decap_8
XFILLER_93_20 VPWR VGND sg13g2_decap_8
X_0930_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_154 VPWR VGND sg13g2_decap_8
XFILLER_20_109 VPWR VGND sg13g2_decap_8
X_0861_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q Tile_X0Y1_W1END[2]
+ Tile_X0Y1_WW4END[14] Tile_X0Y1_WW4END[6] Tile_X0Y1_W6END[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
+ _0240_ VPWR VGND sg13g2_mux4_1
X_0792_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q VPWR
+ _0182_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
XFILLER_87_109 VPWR VGND sg13g2_fill_1
X_1413_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_197 VPWR VGND sg13g2_fill_2
XFILLER_95_142 VPWR VGND sg13g2_fill_1
X_1344_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1275_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_86_164 VPWR VGND sg13g2_fill_1
XFILLER_103_63 VPWR VGND sg13g2_decap_8
XFILLER_86_197 VPWR VGND sg13g2_fill_2
XFILLER_88_86 VPWR VGND sg13g2_fill_1
XFILLER_77_197 VPWR VGND sg13g2_fill_2
X_1060_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0913_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0844_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q _0223_
+ _0224_ _0226_ VPWR VGND sg13g2_nor3_1
X_0775_ _0167_ _0166_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_45_0 VPWR VGND sg13g2_decap_8
X_1327_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1258_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1189_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_90_54 VPWR VGND sg13g2_fill_2
XFILLER_74_44 VPWR VGND sg13g2_decap_8
X_0491_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q UIO_OUT_TT_PROJECT7
+ UIO_OE_TT_PROJECT7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG7 VPWR VGND sg13g2_mux4_1
X_0560_ _0012_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ _0032_ VPWR VGND sg13g2_mux2_1
XFILLER_2_182 VPWR VGND sg13g2_decap_8
X_1043_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1112_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_145 VPWR VGND sg13g2_decap_4
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_17_4 VPWR VGND sg13g2_fill_1
X_0827_ _0150_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q
+ _0212_ VPWR VGND sg13g2_nor2b_1
X_0758_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q UO_OUT_TT_PROJECT4
+ _0147_ _0151_ _0335_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG4 VPWR VGND sg13g2_mux4_1
X_0689_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q
+ _0122_ _0121_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG3 _0355_ sg13g2_a221oi_1
XFILLER_0_119 VPWR VGND sg13g2_decap_4
XFILLER_71_159 VPWR VGND sg13g2_fill_2
XFILLER_100_42 VPWR VGND sg13g2_decap_8
XFILLER_85_43 VPWR VGND sg13g2_decap_4
XFILLER_62_115 VPWR VGND sg13g2_fill_2
XFILLER_109_180 VPWR VGND sg13g2_decap_4
X_0612_ VGND VPWR _0073_ _0076_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S4BEG3
+ _0078_ sg13g2_a21oi_1
X_1661_ Tile_X0Y0_S4END[15] Tile_X0Y1_S4BEG[7] VPWR VGND sg13g2_buf_1
X_1592_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG6 Tile_X0Y1_EE4BEG[6]
+ VPWR VGND sg13g2_buf_1
X_0474_ VPWR VGND _0004_ _0005_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q
+ _0290_ _0006_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_a221oi_1
X_0543_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q VPWR
+ _0017_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q
+ _0016_ sg13g2_o21ai_1
XFILLER_38_101 VPWR VGND sg13g2_fill_1
X_1026_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_156 VPWR VGND sg13g2_decap_4
XFILLER_30_49 VPWR VGND sg13g2_fill_1
XFILLER_52_170 VPWR VGND sg13g2_fill_2
XFILLER_55_79 VPWR VGND sg13g2_fill_2
XFILLER_106_161 VPWR VGND sg13g2_decap_8
XFILLER_96_64 VPWR VGND sg13g2_decap_8
X_0526_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q UIO_OUT_TT_PROJECT2
+ UIO_OE_TT_PROJECT6 _0013_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG14
+ VPWR VGND sg13g2_mux4_1
X_1644_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG6 Tile_X0Y1_S2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1575_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG1 Tile_X0Y1_E6BEG[1]
+ VPWR VGND sg13g2_buf_1
X_0388_ _0315_ Tile_X0Y0_S1END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_0457_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q Tile_X0Y0_W1END[1]
+ Tile_X0Y0_W2MID[2] Tile_X0Y0_W2END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG5
+ VPWR VGND sg13g2_mux4_1
X_1009_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_63 VPWR VGND sg13g2_decap_8
XFILLER_103_197 VPWR VGND sg13g2_fill_2
XFILLER_103_164 VPWR VGND sg13g2_decap_8
XFILLER_103_120 VPWR VGND sg13g2_fill_2
XFILLER_82_44 VPWR VGND sg13g2_fill_2
XFILLER_15_93 VPWR VGND sg13g2_fill_1
X_1360_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1291_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_0 VPWR VGND sg13g2_fill_1
X_1489_ Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData_O[24] VPWR VGND sg13g2_buf_1
XFILLER_98_140 VPWR VGND sg13g2_decap_8
X_0509_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG9 VPWR VGND sg13g2_mux4_1
X_1558_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG0 Tile_X0Y1_E2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1627_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData_O[25] VPWR VGND sg13g2_buf_1
XFILLER_100_189 VPWR VGND sg13g2_fill_2
XFILLER_36_15 VPWR VGND sg13g2_fill_2
XFILLER_9_188 VPWR VGND sg13g2_fill_2
XFILLER_9_122 VPWR VGND sg13g2_decap_4
X_0860_ _0238_ VPWR _0239_ VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
+ _0152_ sg13g2_o21ai_1
X_0791_ _0181_ _0180_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
X_1343_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1412_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1274_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0989_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_103_42 VPWR VGND sg13g2_decap_8
XFILLER_10_143 VPWR VGND sg13g2_fill_1
XFILLER_10_121 VPWR VGND sg13g2_decap_4
XFILLER_6_147 VPWR VGND sg13g2_decap_8
XFILLER_6_125 VPWR VGND sg13g2_fill_2
XFILLER_6_114 VPWR VGND sg13g2_decap_8
XFILLER_77_121 VPWR VGND sg13g2_decap_8
XFILLER_5_0 VPWR VGND sg13g2_decap_8
XFILLER_77_132 VPWR VGND sg13g2_fill_1
X_0912_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0843_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q Tile_X0Y1_WW4END[3]
+ Tile_X0Y1_WW4END[11] Tile_X0Y1_W6END[3] Tile_X0Y1_W6END[11] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q
+ _0225_ VPWR VGND sg13g2_mux4_1
X_0774_ _0153_ _0149_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ _0166_ VPWR VGND sg13g2_mux2_1
X_1326_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_0 VPWR VGND sg13g2_decap_4
X_1188_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1257_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_128 VPWR VGND sg13g2_decap_8
XFILLER_59_143 VPWR VGND sg13g2_decap_4
XFILLER_99_42 VPWR VGND sg13g2_decap_8
X_0490_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q UIO_OUT_TT_PROJECT6
+ UIO_OE_TT_PROJECT6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E2BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_2_161 VPWR VGND sg13g2_decap_8
X_1042_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_138 VPWR VGND sg13g2_fill_1
X_1111_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_0_53 VPWR VGND sg13g2_fill_2
XFILLER_48_90 VPWR VGND sg13g2_fill_2
X_0688_ UO_OUT_TT_PROJECT3 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q _0122_ VPWR
+ VGND sg13g2_nor3_1
X_0826_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q _0158_
+ _0211_ VPWR VGND sg13g2_nor2_1
X_0757_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q Tile_X0Y1_N4END[3]
+ Tile_X0Y0_S4END[7] _0150_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_56_102 VPWR VGND sg13g2_fill_2
X_1309_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_21 VPWR VGND sg13g2_decap_8
XFILLER_69_23 VPWR VGND sg13g2_decap_8
XFILLER_62_138 VPWR VGND sg13g2_fill_2
X_0611_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q _0077_
+ _0078_ VPWR VGND sg13g2_nor2_1
X_0542_ _0015_ VPWR _0016_ VGND Tile_X0Y0_W6END[8] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ sg13g2_o21ai_1
X_1660_ Tile_X0Y0_S4END[14] Tile_X0Y1_S4BEG[6] VPWR VGND sg13g2_buf_1
X_1591_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG5 Tile_X0Y1_EE4BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0473_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END0 _0005_ VPWR VGND sg13g2_nor3_1
X_1025_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_160 VPWR VGND sg13g2_fill_2
X_0809_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q Tile_X0Y1_W1END[1]
+ Tile_X0Y1_WW4END[13] Tile_X0Y1_W6END[5] _0157_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
+ _0197_ VPWR VGND sg13g2_mux4_1
XFILLER_39_15 VPWR VGND sg13g2_decap_8
XFILLER_52_160 VPWR VGND sg13g2_decap_8
XFILLER_52_193 VPWR VGND sg13g2_decap_8
XFILLER_106_184 VPWR VGND sg13g2_fill_1
XFILLER_106_140 VPWR VGND sg13g2_decap_8
XFILLER_105_0 VPWR VGND sg13g2_decap_8
XFILLER_96_21 VPWR VGND sg13g2_decap_4
XFILLER_45_80 VPWR VGND sg13g2_fill_1
X_1643_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG5 Tile_X0Y1_S2BEG[5]
+ VPWR VGND sg13g2_buf_1
XANTENNA_1 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0525_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q
+ _0013_ VPWR VGND sg13g2_mux4_1
X_0456_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y0_W2MID[3]
+ Tile_X0Y0_W2END[3] Tile_X0Y0_W6END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG4
+ VPWR VGND sg13g2_mux4_1
X_1574_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG0 Tile_X0Y1_E6BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0387_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y0_W1END[1]
+ Tile_X0Y0_W6END[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13
+ _0310_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_20_0 VPWR VGND sg13g2_decap_8
X_1008_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_7 VPWR VGND sg13g2_decap_8
XFILLER_41_49 VPWR VGND sg13g2_decap_8
XFILLER_106_42 VPWR VGND sg13g2_decap_8
X_1290_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_31_130 VPWR VGND sg13g2_fill_1
XFILLER_68_0 VPWR VGND sg13g2_fill_2
X_1626_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData_O[24] VPWR VGND sg13g2_buf_1
X_1488_ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData_O[23] VPWR VGND sg13g2_buf_1
X_0439_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb2
+ Tile_X0Y0_S2MID[2] Tile_X0Y1_N2MID[2] Tile_X0Y0_S2END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2 VPWR VGND sg13g2_mux4_1
X_0508_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q UIO_OUT_TT_PROJECT5
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG5 VPWR VGND sg13g2_mux4_1
X_1557_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG3 Tile_X0Y1_E1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_77_67 VPWR VGND sg13g2_fill_2
XFILLER_61_7 VPWR VGND sg13g2_decap_4
X_0790_ _0151_ _0147_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ _0180_ VPWR VGND sg13g2_mux2_1
XFILLER_95_133 VPWR VGND sg13g2_decap_8
XFILLER_3_86 VPWR VGND sg13g2_decap_8
XFILLER_3_53 VPWR VGND sg13g2_fill_2
XFILLER_3_42 VPWR VGND sg13g2_decap_8
X_1342_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1411_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1273_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_199 VPWR VGND sg13g2_fill_1
X_0988_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1609_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_103_21 VPWR VGND sg13g2_decap_8
XFILLER_86_199 VPWR VGND sg13g2_fill_1
XFILLER_77_199 VPWR VGND sg13g2_fill_1
X_0911_ RST_N_TT_PROJECT _0281_ _0286_ _0277_ _0307_ VPWR VGND sg13g2_a22oi_1
X_0842_ _0147_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q
+ _0224_ VPWR VGND sg13g2_nor2b_1
XFILLER_5_192 VPWR VGND sg13g2_decap_8
X_0773_ VGND VPWR _0160_ _0163_ Tile_X0Y0_W_TT_IF2_top.N4BEG_outbuf_8.A _0165_ sg13g2_a21oi_1
XFILLER_68_199 VPWR VGND sg13g2_fill_1
XFILLER_68_133 VPWR VGND sg13g2_fill_2
X_1325_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1256_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1187_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_107 VPWR VGND sg13g2_decap_8
XFILLER_58_25 VPWR VGND sg13g2_fill_1
XFILLER_90_78 VPWR VGND sg13g2_fill_2
XFILLER_90_56 VPWR VGND sg13g2_fill_1
XFILLER_99_98 VPWR VGND sg13g2_decap_8
XFILLER_99_21 VPWR VGND sg13g2_decap_8
X_1110_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1041_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_0_87 VPWR VGND sg13g2_decap_8
XFILLER_9_41 VPWR VGND sg13g2_decap_8
X_0825_ VGND VPWR _0206_ _0208_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S4BEG3
+ _0210_ sg13g2_a21oi_1
X_0687_ _0121_ _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_nand2b_1
X_0756_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y1_N4END[2]
+ Tile_X0Y0_S4END[6] _0149_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_50_0 VPWR VGND sg13g2_decap_8
XFILLER_71_139 VPWR VGND sg13g2_fill_2
X_1308_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_17 VPWR VGND sg13g2_fill_1
X_1239_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_39 VPWR VGND sg13g2_fill_2
XFILLER_109_53 VPWR VGND sg13g2_fill_2
XFILLER_109_193 VPWR VGND sg13g2_decap_8
X_0610_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q Tile_X0Y0_W1END[3]
+ Tile_X0Y0_WW4END[15] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ _0077_ VPWR VGND sg13g2_mux4_1
X_0472_ _0004_ Tile_X0Y0_S1END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
X_0541_ _0015_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_nand2b_1
X_1590_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG4 Tile_X0Y1_EE4BEG[4]
+ VPWR VGND sg13g2_buf_1
X_1024_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_22_4 VPWR VGND sg13g2_fill_2
XFILLER_98_0 VPWR VGND sg13g2_decap_8
XFILLER_107_119 VPWR VGND sg13g2_decap_8
X_0808_ VGND VPWR Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
+ _0195_ _0196_ _0302_ sg13g2_a21oi_1
X_0739_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT4 _0151_ _0003_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG8 VPWR VGND sg13g2_mux4_1
XFILLER_29_158 VPWR VGND sg13g2_fill_1
XFILLER_71_69 VPWR VGND sg13g2_decap_4
XFILLER_52_172 VPWR VGND sg13g2_fill_1
XFILLER_20_62 VPWR VGND sg13g2_decap_4
XFILLER_20_84 VPWR VGND sg13g2_fill_1
XFILLER_43_183 VPWR VGND sg13g2_decap_4
X_1642_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG4 Tile_X0Y1_S2BEG[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_6_53 VPWR VGND sg13g2_fill_2
XFILLER_6_42 VPWR VGND sg13g2_decap_8
XANTENNA_2 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0455_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb4
+ Tile_X0Y0_S2MID[4] Tile_X0Y1_N2MID[4] Tile_X0Y0_S2END[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG4 VPWR VGND sg13g2_mux4_1
X_0524_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q UIO_OUT_TT_PROJECT1
+ UIO_OE_TT_PROJECT5 _0012_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG13
+ VPWR VGND sg13g2_mux4_1
XFILLER_6_86 VPWR VGND sg13g2_decap_8
X_1573_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb7 Tile_X0Y1_E2BEGb[7]
+ VPWR VGND sg13g2_buf_1
X_1007_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0386_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_mux4_1
XFILLER_26_117 VPWR VGND sg13g2_fill_2
XFILLER_103_122 VPWR VGND sg13g2_fill_1
XFILLER_106_98 VPWR VGND sg13g2_decap_8
XFILLER_106_21 VPWR VGND sg13g2_decap_8
XFILLER_103_199 VPWR VGND sg13g2_fill_1
XFILLER_103_144 VPWR VGND sg13g2_fill_2
XFILLER_40_197 VPWR VGND sg13g2_fill_2
X_1556_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG2 Tile_X0Y1_E1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1625_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData_O[23] VPWR VGND sg13g2_buf_1
X_1487_ Tile_X0Y0_FrameData[22] Tile_X0Y0_FrameData_O[22] VPWR VGND sg13g2_buf_1
X_0507_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG10 VPWR VGND sg13g2_mux4_1
X_0438_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y1_W2MID[5]
+ Tile_X0Y1_W2END[5] Tile_X0Y1_W6END[5] _0349_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb2 VPWR VGND sg13g2_mux4_1
XFILLER_36_17 VPWR VGND sg13g2_fill_1
X_0369_ VPWR _0299_ Tile_X0Y1_W6END[1] VGND sg13g2_inv_1
XFILLER_36_39 VPWR VGND sg13g2_fill_1
XFILLER_22_153 VPWR VGND sg13g2_fill_2
X_1410_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_54_7 VPWR VGND sg13g2_decap_4
XFILLER_3_65 VPWR VGND sg13g2_decap_8
XFILLER_3_21 VPWR VGND sg13g2_decap_8
X_1341_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1272_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_0 VPWR VGND sg13g2_decap_8
X_0987_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_190 VPWR VGND sg13g2_fill_1
X_1539_ Tile_X0Y1_N4END[10] Tile_X0Y0_N4BEG[2] VPWR VGND sg13g2_buf_1
X_1608_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData_O[6] VPWR VGND sg13g2_buf_1
XFILLER_103_77 VPWR VGND sg13g2_decap_4
XFILLER_37_82 VPWR VGND sg13g2_decap_8
X_0910_ VGND VPWR _0283_ _0285_ _0286_ _0307_ sg13g2_a21oi_1
X_0772_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q _0164_
+ _0165_ VPWR VGND sg13g2_nor2_1
X_0841_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q _0155_
+ _0223_ VPWR VGND sg13g2_nor2_1
XFILLER_68_112 VPWR VGND sg13g2_fill_2
XFILLER_5_171 VPWR VGND sg13g2_decap_8
XFILLER_83_159 VPWR VGND sg13g2_decap_8
X_1324_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1255_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1186_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_58 VPWR VGND sg13g2_fill_2
XFILLER_23_95 VPWR VGND sg13g2_fill_2
XFILLER_99_77 VPWR VGND sg13g2_fill_1
XFILLER_2_141 VPWR VGND sg13g2_fill_2
X_1040_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_196 VPWR VGND sg13g2_decap_4
XFILLER_0_77 VPWR VGND sg13g2_decap_4
XFILLER_0_99 VPWR VGND sg13g2_decap_4
XFILLER_9_97 VPWR VGND sg13g2_decap_4
X_0824_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q _0209_
+ _0210_ VPWR VGND sg13g2_nor2_1
X_0755_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q Tile_X0Y1_N4END[1]
+ Tile_X0Y0_S4END[5] _0148_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_56_104 VPWR VGND sg13g2_fill_1
X_0686_ VPWR VGND Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q
+ _0120_ _0119_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEG2 _0348_ sg13g2_a221oi_1
X_1307_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1238_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1169_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_56 VPWR VGND sg13g2_fill_1
XFILLER_109_87 VPWR VGND sg13g2_decap_8
XFILLER_18_51 VPWR VGND sg13g2_decap_4
XFILLER_55_192 VPWR VGND sg13g2_fill_1
XFILLER_55_170 VPWR VGND sg13g2_decap_8
X_0540_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q UIO_OUT_TT_PROJECT3
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG4 _0014_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.E6BEG11
+ VPWR VGND sg13g2_mux4_1
X_0471_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q Tile_X0Y0_W2MID[0]
+ Tile_X0Y0_W2END[0] Tile_X0Y0_W6END[0] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEG7
+ VPWR VGND sg13g2_mux4_1
X_1023_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_126 VPWR VGND sg13g2_decap_4
XFILLER_53_107 VPWR VGND sg13g2_fill_2
XFILLER_53_129 VPWR VGND sg13g2_decap_8
X_0807_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13 _0001_
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q _0195_ VPWR
+ VGND sg13g2_mux2_1
X_0738_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0325_ Tile_X0Y0_S4END[7] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q
+ _0151_ VPWR VGND sg13g2_mux4_1
X_0669_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q Tile_X0Y1_W2MID[4]
+ Tile_X0Y1_W2END[4] Tile_X0Y1_W6END[11] _0356_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG3 VPWR VGND sg13g2_mux4_1
XFILLER_52_184 VPWR VGND sg13g2_fill_1
XFILLER_106_175 VPWR VGND sg13g2_decap_8
XFILLER_84_7 VPWR VGND sg13g2_decap_8
XFILLER_43_162 VPWR VGND sg13g2_decap_4
XFILLER_6_65 VPWR VGND sg13g2_decap_8
XFILLER_6_21 VPWR VGND sg13g2_decap_8
X_1641_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG3 Tile_X0Y1_S2BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1572_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb6 Tile_X0Y1_E2BEGb[6]
+ VPWR VGND sg13g2_buf_1
XANTENNA_3 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0523_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q
+ _0012_ VPWR VGND sg13g2_mux4_1
X_0454_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y1_W2MID[3]
+ Tile_X0Y1_W2END[3] Tile_X0Y1_W6END[3] _0000_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb4 VPWR VGND sg13g2_mux4_1
X_0385_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q Tile_X0Y1_W1END[1]
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG13 Tile_X0Y1_W6END[5]
+ _0314_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END1
+ VPWR VGND sg13g2_mux4_1
X_1006_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_77 VPWR VGND sg13g2_decap_8
XFILLER_103_178 VPWR VGND sg13g2_decap_8
XFILLER_82_14 VPWR VGND sg13g2_fill_2
XFILLER_40_143 VPWR VGND sg13g2_decap_4
XFILLER_110_0 VPWR VGND sg13g2_decap_8
XFILLER_40_187 VPWR VGND sg13g2_fill_2
XFILLER_98_121 VPWR VGND sg13g2_fill_2
X_0506_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q UIO_OUT_TT_PROJECT4
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG4 VPWR VGND sg13g2_mux4_1
X_1555_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG1 Tile_X0Y1_E1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1624_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameData_O[22] VPWR VGND sg13g2_buf_1
X_1486_ Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData_O[21] VPWR VGND sg13g2_buf_1
XFILLER_98_198 VPWR VGND sg13g2_fill_2
X_0368_ VPWR _0298_ Tile_X0Y1_W6END[2] VGND sg13g2_inv_1
X_0437_ _0344_ _0347_ _0349_ VPWR VGND sg13g2_nor2b_1
XFILLER_22_198 VPWR VGND sg13g2_fill_2
XFILLER_89_132 VPWR VGND sg13g2_fill_2
XFILLER_77_47 VPWR VGND sg13g2_fill_2
XFILLER_77_14 VPWR VGND sg13g2_fill_2
XFILLER_9_147 VPWR VGND sg13g2_decap_8
X_1340_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1271_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
Xclkbuf_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VPWR VGND
+ sg13g2_buf_8
XFILLER_73_0 VPWR VGND sg13g2_decap_4
X_0986_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1469_ Tile_X0Y0_FrameData[4] Tile_X0Y0_FrameData_O[4] VPWR VGND sg13g2_buf_1
X_1538_ Tile_X0Y1_N4END[9] Tile_X0Y0_N4BEG[1] VPWR VGND sg13g2_buf_1
X_1607_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_47_17 VPWR VGND sg13g2_decap_4
XFILLER_103_56 VPWR VGND sg13g2_decap_8
XFILLER_86_157 VPWR VGND sg13g2_decap_8
XFILLER_47_39 VPWR VGND sg13g2_decap_4
XFILLER_10_157 VPWR VGND sg13g2_decap_4
XFILLER_92_149 VPWR VGND sg13g2_decap_4
X_0771_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q Tile_X0Y1_W1END[0]
+ Tile_X0Y1_W6END[8] Tile_X0Y1_WW4END[0] _0158_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ _0164_ VPWR VGND sg13g2_mux4_1
X_0840_ _0221_ _0222_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q
+ UI_IN_TT_PROJECT2 VPWR VGND sg13g2_mux2_1
XFILLER_5_161 VPWR VGND sg13g2_decap_8
X_1323_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_83_127 VPWR VGND sg13g2_decap_4
XFILLER_68_157 VPWR VGND sg13g2_fill_2
X_1254_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1185_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0969_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_90_14 VPWR VGND sg13g2_fill_2
XFILLER_99_56 VPWR VGND sg13g2_fill_1
XFILLER_3_0 VPWR VGND sg13g2_decap_8
XFILLER_2_175 VPWR VGND sg13g2_decap_8
XFILLER_65_138 VPWR VGND sg13g2_decap_8
X_0685_ UO_OUT_TT_PROJECT2 Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q _0120_ VPWR
+ VGND sg13g2_nor3_1
X_0823_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q Tile_X0Y1_W1END[3]
+ Tile_X0Y1_WW4END[15] Tile_X0Y1_W6END[7] _0155_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
+ _0209_ VPWR VGND sg13g2_mux4_1
X_0754_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y1_N4END[0]
+ Tile_X0Y0_S4END[4] _0147_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E6BEG0
+ VPWR VGND sg13g2_mux4_1
X_1306_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_0 VPWR VGND sg13g2_decap_4
X_1099_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1237_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1168_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_35 VPWR VGND sg13g2_decap_8
XFILLER_85_47 VPWR VGND sg13g2_fill_1
XFILLER_85_36 VPWR VGND sg13g2_decap_8
XFILLER_85_14 VPWR VGND sg13g2_fill_1
XFILLER_55_160 VPWR VGND sg13g2_decap_8
XFILLER_18_74 VPWR VGND sg13g2_fill_1
XFILLER_109_184 VPWR VGND sg13g2_fill_1
XFILLER_109_162 VPWR VGND sg13g2_decap_8
X_0470_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N2BEGb7
+ Tile_X0Y0_S2MID[7] Tile_X0Y1_N2MID[7] Tile_X0Y0_S2END[7] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG7 VPWR VGND sg13g2_mux4_1
X_1022_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0668_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y1_W2MID[5]
+ Tile_X0Y1_W2END[5] Tile_X0Y1_W6END[10] _0349_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG2 VPWR VGND sg13g2_mux4_1
X_0737_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q UO_OUT_TT_PROJECT3
+ _0150_ UO_OUT_TT_PROJECT7 _0335_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q
+ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.EE4BEG7 VPWR VGND sg13g2_mux4_1
X_0806_ _0194_ _0193_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_nand2b_1
X_0599_ _0066_ VPWR _0067_ VGND Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ _0012_ sg13g2_o21ai_1
XFILLER_29_105 VPWR VGND sg13g2_fill_1
XFILLER_44_119 VPWR VGND sg13g2_fill_1
XFILLER_106_154 VPWR VGND sg13g2_decap_8
XFILLER_29_51 VPWR VGND sg13g2_fill_2
XFILLER_77_7 VPWR VGND sg13g2_decap_8
X_0522_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q UIO_OUT_TT_PROJECT0
+ UIO_OE_TT_PROJECT4 _0011_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.EE4BEG12
+ VPWR VGND sg13g2_mux4_1
X_1640_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.S2BEG2 Tile_X0Y1_S2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1571_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E2BEGb5 Tile_X0Y1_E2BEGb[5]
+ VPWR VGND sg13g2_buf_1
XANTENNA_4 VPWR VGND Tile_X0Y1_FrameData[23] sg13g2_antennanp
X_0384_ VPWR VGND _0312_ _0313_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q
+ _0299_ _0314_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a221oi_1
X_0453_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y1_N2MID[4]
+ Tile_X0Y1_N2END[4] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.S2BEG4
+ Tile_X0Y0_S2MID[4] Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q
+ _0000_ VPWR VGND sg13g2_mux4_1
X_1005_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_56 VPWR VGND sg13g2_decap_8
XFILLER_103_146 VPWR VGND sg13g2_fill_1
XFILLER_82_37 VPWR VGND sg13g2_decap_8
XFILLER_15_86 VPWR VGND sg13g2_decap_8
XFILLER_40_122 VPWR VGND sg13g2_fill_1
XFILLER_40_199 VPWR VGND sg13g2_fill_1
XFILLER_103_0 VPWR VGND sg13g2_decap_8
XFILLER_16_185 VPWR VGND sg13g2_fill_1
XFILLER_31_144 VPWR VGND sg13g2_fill_2
X_0505_ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q
+ Tile_X0Y0_W_TT_IF2_top.Inst_W_TT_IF2_top_switch_matrix.J_NS4_BEG11 VPWR VGND sg13g2_mux4_1
XFILLER_100_116 VPWR VGND sg13g2_decap_4
X_1485_ Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData_O[20] VPWR VGND sg13g2_buf_1
X_1554_ Tile_X0Y1_W_TT_IF2_bot.Inst_W_TT_IF2_bot_switch_matrix.E1BEG0 Tile_X0Y1_E1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0436_ _0348_ _0347_ _0344_ VPWR VGND sg13g2_nand2b_1
X_1623_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData_O[21] VPWR VGND sg13g2_buf_1
.ends

