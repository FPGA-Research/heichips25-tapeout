magic
tech ihp-sg13g2
magscale 1 2
timestamp 1753873013
<< metal1 >>
rect 1152 84692 20352 84716
rect 1152 84652 3688 84692
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 4056 84652 18808 84692
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 19176 84652 20352 84692
rect 1152 84628 20352 84652
rect 5163 84524 5205 84533
rect 5163 84484 5164 84524
rect 5204 84484 5205 84524
rect 5163 84475 5205 84484
rect 13131 84524 13173 84533
rect 13131 84484 13132 84524
rect 13172 84484 13173 84524
rect 13131 84475 13173 84484
rect 18891 84524 18933 84533
rect 18891 84484 18892 84524
rect 18932 84484 18933 84524
rect 18891 84475 18933 84484
rect 1515 84440 1557 84449
rect 1515 84400 1516 84440
rect 1556 84400 1557 84440
rect 1515 84391 1557 84400
rect 1899 84440 1941 84449
rect 1899 84400 1900 84440
rect 1940 84400 1941 84440
rect 1899 84391 1941 84400
rect 7275 84440 7317 84449
rect 7275 84400 7276 84440
rect 7316 84400 7317 84440
rect 7275 84391 7317 84400
rect 7851 84440 7893 84449
rect 7851 84400 7852 84440
rect 7892 84400 7893 84440
rect 7851 84391 7893 84400
rect 8043 84440 8085 84449
rect 8043 84400 8044 84440
rect 8084 84400 8085 84440
rect 8043 84391 8085 84400
rect 19275 84440 19317 84449
rect 19275 84400 19276 84440
rect 19316 84400 19317 84440
rect 19275 84391 19317 84400
rect 20043 84440 20085 84449
rect 20043 84400 20044 84440
rect 20084 84400 20085 84440
rect 20043 84391 20085 84400
rect 1315 84356 1373 84357
rect 1315 84316 1324 84356
rect 1364 84316 1373 84356
rect 1315 84315 1373 84316
rect 1699 84356 1757 84357
rect 1699 84316 1708 84356
rect 1748 84316 1757 84356
rect 1699 84315 1757 84316
rect 7075 84356 7133 84357
rect 7075 84316 7084 84356
rect 7124 84316 7133 84356
rect 7075 84315 7133 84316
rect 7651 84356 7709 84357
rect 7651 84316 7660 84356
rect 7700 84316 7709 84356
rect 7651 84315 7709 84316
rect 8227 84356 8285 84357
rect 8227 84316 8236 84356
rect 8276 84316 8285 84356
rect 8227 84315 8285 84316
rect 11787 84356 11829 84365
rect 11787 84316 11788 84356
rect 11828 84316 11829 84356
rect 11787 84307 11829 84316
rect 12259 84356 12317 84357
rect 12259 84316 12268 84356
rect 12308 84316 12317 84356
rect 12259 84315 12317 84316
rect 12931 84356 12989 84357
rect 12931 84316 12940 84356
rect 12980 84316 12989 84356
rect 12931 84315 12989 84316
rect 13507 84356 13565 84357
rect 13507 84316 13516 84356
rect 13556 84316 13565 84356
rect 13507 84315 13565 84316
rect 19075 84356 19133 84357
rect 19075 84316 19084 84356
rect 19124 84316 19133 84356
rect 19075 84315 19133 84316
rect 19459 84356 19517 84357
rect 19459 84316 19468 84356
rect 19508 84316 19517 84356
rect 19459 84315 19517 84316
rect 19843 84356 19901 84357
rect 19843 84316 19852 84356
rect 19892 84316 19901 84356
rect 19843 84315 19901 84316
rect 20227 84356 20285 84357
rect 20227 84316 20236 84356
rect 20276 84316 20285 84356
rect 20227 84315 20285 84316
rect 2083 84272 2141 84273
rect 2083 84232 2092 84272
rect 2132 84232 2141 84272
rect 2083 84231 2141 84232
rect 3331 84272 3389 84273
rect 3331 84232 3340 84272
rect 3380 84232 3389 84272
rect 3331 84231 3389 84232
rect 3715 84272 3773 84273
rect 3715 84232 3724 84272
rect 3764 84232 3773 84272
rect 3715 84231 3773 84232
rect 4963 84272 5021 84273
rect 4963 84232 4972 84272
rect 5012 84232 5021 84272
rect 4963 84231 5021 84232
rect 5539 84272 5597 84273
rect 5539 84232 5548 84272
rect 5588 84232 5597 84272
rect 5539 84231 5597 84232
rect 6787 84272 6845 84273
rect 6787 84232 6796 84272
rect 6836 84232 6845 84272
rect 6787 84231 6845 84232
rect 8419 84272 8477 84273
rect 8419 84232 8428 84272
rect 8468 84232 8477 84272
rect 8419 84231 8477 84232
rect 9667 84272 9725 84273
rect 9667 84232 9676 84272
rect 9716 84232 9725 84272
rect 9667 84231 9725 84232
rect 10243 84272 10301 84273
rect 10243 84232 10252 84272
rect 10292 84232 10301 84272
rect 10243 84231 10301 84232
rect 11491 84272 11549 84273
rect 11491 84232 11500 84272
rect 11540 84232 11549 84272
rect 11491 84231 11549 84232
rect 11691 84272 11733 84281
rect 11691 84232 11692 84272
rect 11732 84232 11733 84272
rect 11691 84223 11733 84232
rect 11883 84272 11925 84281
rect 11883 84232 11884 84272
rect 11924 84232 11925 84272
rect 11883 84223 11925 84232
rect 13699 84272 13757 84273
rect 13699 84232 13708 84272
rect 13748 84232 13757 84272
rect 13699 84231 13757 84232
rect 14947 84272 15005 84273
rect 14947 84232 14956 84272
rect 14996 84232 15005 84272
rect 14947 84231 15005 84232
rect 15331 84272 15389 84273
rect 15331 84232 15340 84272
rect 15380 84232 15389 84272
rect 15331 84231 15389 84232
rect 16579 84272 16637 84273
rect 16579 84232 16588 84272
rect 16628 84232 16637 84272
rect 16579 84231 16637 84232
rect 17251 84272 17309 84273
rect 17251 84232 17260 84272
rect 17300 84232 17309 84272
rect 17251 84231 17309 84232
rect 18499 84272 18557 84273
rect 18499 84232 18508 84272
rect 18548 84232 18557 84272
rect 18499 84231 18557 84232
rect 3531 84104 3573 84113
rect 3531 84064 3532 84104
rect 3572 84064 3573 84104
rect 3531 84055 3573 84064
rect 5355 84104 5397 84113
rect 5355 84064 5356 84104
rect 5396 84064 5397 84104
rect 5355 84055 5397 84064
rect 9867 84104 9909 84113
rect 9867 84064 9868 84104
rect 9908 84064 9909 84104
rect 9867 84055 9909 84064
rect 10059 84104 10101 84113
rect 10059 84064 10060 84104
rect 10100 84064 10101 84104
rect 10059 84055 10101 84064
rect 12459 84104 12501 84113
rect 12459 84064 12460 84104
rect 12500 84064 12501 84104
rect 12459 84055 12501 84064
rect 12739 84104 12797 84105
rect 12739 84064 12748 84104
rect 12788 84064 12797 84104
rect 12739 84063 12797 84064
rect 13323 84104 13365 84113
rect 13323 84064 13324 84104
rect 13364 84064 13365 84104
rect 13323 84055 13365 84064
rect 15147 84104 15189 84113
rect 15147 84064 15148 84104
rect 15188 84064 15189 84104
rect 15147 84055 15189 84064
rect 16779 84104 16821 84113
rect 16779 84064 16780 84104
rect 16820 84064 16821 84104
rect 16779 84055 16821 84064
rect 17059 84104 17117 84105
rect 17059 84064 17068 84104
rect 17108 84064 17117 84104
rect 17059 84063 17117 84064
rect 18699 84104 18741 84113
rect 18699 84064 18700 84104
rect 18740 84064 18741 84104
rect 18699 84055 18741 84064
rect 19659 84104 19701 84113
rect 19659 84064 19660 84104
rect 19700 84064 19701 84104
rect 19659 84055 19701 84064
rect 1152 83936 20452 83960
rect 1152 83896 4928 83936
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 5296 83896 20048 83936
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20416 83896 20452 83936
rect 1152 83872 20452 83896
rect 1515 83768 1557 83777
rect 1515 83728 1516 83768
rect 1556 83728 1557 83768
rect 1515 83719 1557 83728
rect 6699 83768 6741 83777
rect 6699 83728 6700 83768
rect 6740 83728 6741 83768
rect 6699 83719 6741 83728
rect 7075 83768 7133 83769
rect 7075 83728 7084 83768
rect 7124 83728 7133 83768
rect 7075 83727 7133 83728
rect 9003 83768 9045 83777
rect 9003 83728 9004 83768
rect 9044 83728 9045 83768
rect 9003 83719 9045 83728
rect 18507 83768 18549 83777
rect 18507 83728 18508 83768
rect 18548 83728 18549 83768
rect 18507 83719 18549 83728
rect 19563 83768 19605 83777
rect 19563 83728 19564 83768
rect 19604 83728 19605 83768
rect 19563 83719 19605 83728
rect 19947 83768 19989 83777
rect 19947 83728 19948 83768
rect 19988 83728 19989 83768
rect 19947 83719 19989 83728
rect 11787 83684 11829 83693
rect 11787 83644 11788 83684
rect 11828 83644 11829 83684
rect 11787 83635 11829 83644
rect 19083 83642 19125 83651
rect 1699 83600 1757 83601
rect 1699 83560 1708 83600
rect 1748 83560 1757 83600
rect 1699 83559 1757 83560
rect 2947 83600 3005 83601
rect 2947 83560 2956 83600
rect 2996 83560 3005 83600
rect 2947 83559 3005 83560
rect 3331 83600 3389 83601
rect 3331 83560 3340 83600
rect 3380 83560 3389 83600
rect 3331 83559 3389 83560
rect 4579 83600 4637 83601
rect 4579 83560 4588 83600
rect 4628 83560 4637 83600
rect 4579 83559 4637 83560
rect 4963 83600 5021 83601
rect 4963 83560 4972 83600
rect 5012 83560 5021 83600
rect 4963 83559 5021 83560
rect 6211 83600 6269 83601
rect 6211 83560 6220 83600
rect 6260 83560 6269 83600
rect 6211 83559 6269 83560
rect 7363 83600 7421 83601
rect 7363 83560 7372 83600
rect 7412 83560 7421 83600
rect 7363 83559 7421 83560
rect 8611 83600 8669 83601
rect 8611 83560 8620 83600
rect 8660 83560 8669 83600
rect 8611 83559 8669 83560
rect 10059 83600 10101 83609
rect 10059 83560 10060 83600
rect 10100 83560 10101 83600
rect 10059 83551 10101 83560
rect 10155 83600 10197 83609
rect 19083 83602 19084 83642
rect 19124 83602 19125 83642
rect 10155 83560 10156 83600
rect 10196 83560 10197 83600
rect 10155 83551 10197 83560
rect 11107 83600 11165 83601
rect 11107 83560 11116 83600
rect 11156 83560 11165 83600
rect 13987 83600 14045 83601
rect 11107 83559 11165 83560
rect 11595 83586 11637 83595
rect 11595 83546 11596 83586
rect 11636 83546 11637 83586
rect 13987 83560 13996 83600
rect 14036 83560 14045 83600
rect 13987 83559 14045 83560
rect 15235 83600 15293 83601
rect 15235 83560 15244 83600
rect 15284 83560 15293 83600
rect 15235 83559 15293 83560
rect 16483 83600 16541 83601
rect 16483 83560 16492 83600
rect 16532 83560 16541 83600
rect 16483 83559 16541 83560
rect 17731 83600 17789 83601
rect 17731 83560 17740 83600
rect 17780 83560 17789 83600
rect 19083 83593 19125 83602
rect 19275 83600 19317 83609
rect 17731 83559 17789 83560
rect 19275 83560 19276 83600
rect 19316 83560 19317 83600
rect 19275 83551 19317 83560
rect 19363 83600 19421 83601
rect 19363 83560 19372 83600
rect 19412 83560 19421 83600
rect 19363 83559 19421 83560
rect 11595 83537 11637 83546
rect 1315 83516 1373 83517
rect 1315 83476 1324 83516
rect 1364 83476 1373 83516
rect 1315 83475 1373 83476
rect 9187 83516 9245 83517
rect 9187 83476 9196 83516
rect 9236 83476 9245 83516
rect 9187 83475 9245 83476
rect 10539 83516 10581 83525
rect 10539 83476 10540 83516
rect 10580 83476 10581 83516
rect 10539 83467 10581 83476
rect 10635 83516 10677 83525
rect 10635 83476 10636 83516
rect 10676 83476 10677 83516
rect 10635 83467 10677 83476
rect 12163 83516 12221 83517
rect 12163 83476 12172 83516
rect 12212 83476 12221 83516
rect 12163 83475 12221 83476
rect 12739 83516 12797 83517
rect 12739 83476 12748 83516
rect 12788 83476 12797 83516
rect 12739 83475 12797 83476
rect 13411 83516 13469 83517
rect 13411 83476 13420 83516
rect 13460 83476 13469 83516
rect 13411 83475 13469 83476
rect 13795 83516 13853 83517
rect 13795 83476 13804 83516
rect 13844 83476 13853 83516
rect 13795 83475 13853 83476
rect 15811 83516 15869 83517
rect 15811 83476 15820 83516
rect 15860 83476 15869 83516
rect 15811 83475 15869 83476
rect 16195 83516 16253 83517
rect 16195 83476 16204 83516
rect 16244 83476 16253 83516
rect 16195 83475 16253 83476
rect 18307 83516 18365 83517
rect 18307 83476 18316 83516
rect 18356 83476 18365 83516
rect 18307 83475 18365 83476
rect 18691 83516 18749 83517
rect 18691 83476 18700 83516
rect 18740 83476 18749 83516
rect 18691 83475 18749 83476
rect 19747 83516 19805 83517
rect 19747 83476 19756 83516
rect 19796 83476 19805 83516
rect 19747 83475 19805 83476
rect 20120 83513 20162 83522
rect 20120 83473 20121 83513
rect 20161 83473 20162 83513
rect 20120 83464 20162 83473
rect 6603 83432 6645 83441
rect 6603 83392 6604 83432
rect 6644 83392 6645 83432
rect 6603 83383 6645 83392
rect 7179 83432 7221 83441
rect 7179 83392 7180 83432
rect 7220 83392 7221 83432
rect 7179 83383 7221 83392
rect 9483 83432 9525 83441
rect 9483 83392 9484 83432
rect 9524 83392 9525 83432
rect 9483 83383 9525 83392
rect 9675 83432 9717 83441
rect 9675 83392 9676 83432
rect 9716 83392 9717 83432
rect 9675 83383 9717 83392
rect 12555 83432 12597 83441
rect 12555 83392 12556 83432
rect 12596 83392 12597 83432
rect 12555 83383 12597 83392
rect 12939 83432 12981 83441
rect 12939 83392 12940 83432
rect 12980 83392 12981 83432
rect 12939 83383 12981 83392
rect 19083 83432 19125 83441
rect 19083 83392 19084 83432
rect 19124 83392 19125 83432
rect 19083 83383 19125 83392
rect 3147 83348 3189 83357
rect 3147 83308 3148 83348
rect 3188 83308 3189 83348
rect 3147 83299 3189 83308
rect 4779 83348 4821 83357
rect 4779 83308 4780 83348
rect 4820 83308 4821 83348
rect 4779 83299 4821 83308
rect 6411 83348 6453 83357
rect 6411 83308 6412 83348
rect 6452 83308 6453 83348
rect 6411 83299 6453 83308
rect 8811 83348 8853 83357
rect 8811 83308 8812 83348
rect 8852 83308 8853 83348
rect 8811 83299 8853 83308
rect 12363 83348 12405 83357
rect 12363 83308 12364 83348
rect 12404 83308 12405 83348
rect 12363 83299 12405 83308
rect 13227 83348 13269 83357
rect 13227 83308 13228 83348
rect 13268 83308 13269 83348
rect 13227 83299 13269 83308
rect 13611 83348 13653 83357
rect 13611 83308 13612 83348
rect 13652 83308 13653 83348
rect 13611 83299 13653 83308
rect 15435 83348 15477 83357
rect 15435 83308 15436 83348
rect 15476 83308 15477 83348
rect 15435 83299 15477 83308
rect 15627 83348 15669 83357
rect 15627 83308 15628 83348
rect 15668 83308 15669 83348
rect 15627 83299 15669 83308
rect 16011 83348 16053 83357
rect 16011 83308 16012 83348
rect 16052 83308 16053 83348
rect 16011 83299 16053 83308
rect 17931 83348 17973 83357
rect 17931 83308 17932 83348
rect 17972 83308 17973 83348
rect 17931 83299 17973 83308
rect 18123 83348 18165 83357
rect 18123 83308 18124 83348
rect 18164 83308 18165 83348
rect 18123 83299 18165 83308
rect 1152 83180 20352 83204
rect 1152 83140 3688 83180
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 4056 83140 18808 83180
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 19176 83140 20352 83180
rect 1152 83116 20352 83140
rect 5643 83012 5685 83021
rect 5643 82972 5644 83012
rect 5684 82972 5685 83012
rect 5643 82963 5685 82972
rect 6027 83012 6069 83021
rect 6027 82972 6028 83012
rect 6068 82972 6069 83012
rect 6027 82963 6069 82972
rect 6411 83012 6453 83021
rect 6411 82972 6412 83012
rect 6452 82972 6453 83012
rect 6411 82963 6453 82972
rect 11787 83012 11829 83021
rect 11787 82972 11788 83012
rect 11828 82972 11829 83012
rect 11787 82963 11829 82972
rect 19075 83012 19133 83013
rect 19075 82972 19084 83012
rect 19124 82972 19133 83012
rect 19075 82971 19133 82972
rect 20043 83012 20085 83021
rect 20043 82972 20044 83012
rect 20084 82972 20085 83012
rect 20043 82963 20085 82972
rect 5163 82928 5205 82937
rect 5163 82888 5164 82928
rect 5204 82888 5205 82928
rect 5163 82879 5205 82888
rect 3043 82844 3101 82845
rect 3043 82804 3052 82844
rect 3092 82804 3101 82844
rect 3043 82803 3101 82804
rect 5443 82844 5501 82845
rect 5443 82804 5452 82844
rect 5492 82804 5501 82844
rect 5443 82803 5501 82804
rect 5827 82844 5885 82845
rect 5827 82804 5836 82844
rect 5876 82804 5885 82844
rect 5827 82803 5885 82804
rect 6211 82844 6269 82845
rect 6211 82804 6220 82844
rect 6260 82804 6269 82844
rect 6211 82803 6269 82804
rect 7179 82844 7221 82853
rect 7179 82804 7180 82844
rect 7220 82804 7221 82844
rect 13603 82844 13661 82845
rect 7179 82795 7221 82804
rect 8283 82802 8325 82811
rect 13603 82804 13612 82844
rect 13652 82804 13661 82844
rect 13603 82803 13661 82804
rect 14475 82844 14517 82853
rect 14475 82804 14476 82844
rect 14516 82804 14517 82844
rect 1315 82760 1373 82761
rect 1315 82720 1324 82760
rect 1364 82720 1373 82760
rect 1315 82719 1373 82720
rect 2563 82760 2621 82761
rect 2563 82720 2572 82760
rect 2612 82720 2621 82760
rect 2563 82719 2621 82720
rect 4675 82760 4733 82761
rect 4675 82720 4684 82760
rect 4724 82720 4733 82760
rect 4675 82719 4733 82720
rect 6699 82760 6741 82769
rect 6699 82720 6700 82760
rect 6740 82720 6741 82760
rect 3427 82718 3485 82719
rect 3427 82678 3436 82718
rect 3476 82678 3485 82718
rect 6699 82711 6741 82720
rect 6795 82760 6837 82769
rect 6795 82720 6796 82760
rect 6836 82720 6837 82760
rect 6795 82711 6837 82720
rect 7275 82760 7317 82769
rect 8283 82762 8284 82802
rect 8324 82762 8325 82802
rect 14475 82795 14517 82804
rect 20227 82844 20285 82845
rect 20227 82804 20236 82844
rect 20276 82804 20285 82844
rect 20227 82803 20285 82804
rect 15435 82774 15477 82783
rect 7275 82720 7276 82760
rect 7316 82720 7317 82760
rect 7275 82711 7317 82720
rect 7747 82760 7805 82761
rect 7747 82720 7756 82760
rect 7796 82720 7805 82760
rect 8283 82753 8325 82762
rect 8707 82760 8765 82761
rect 7747 82719 7805 82720
rect 8707 82720 8716 82760
rect 8756 82720 8765 82760
rect 8707 82719 8765 82720
rect 9955 82760 10013 82761
rect 9955 82720 9964 82760
rect 10004 82720 10013 82760
rect 9955 82719 10013 82720
rect 10339 82760 10397 82761
rect 10339 82720 10348 82760
rect 10388 82720 10397 82760
rect 10339 82719 10397 82720
rect 11587 82760 11645 82761
rect 11587 82720 11596 82760
rect 11636 82720 11645 82760
rect 11587 82719 11645 82720
rect 12459 82760 12501 82769
rect 12459 82720 12460 82760
rect 12500 82720 12501 82760
rect 12459 82711 12501 82720
rect 12555 82760 12597 82769
rect 12555 82720 12556 82760
rect 12596 82720 12597 82760
rect 12555 82711 12597 82720
rect 12651 82760 12693 82769
rect 12651 82720 12652 82760
rect 12692 82720 12693 82760
rect 12651 82711 12693 82720
rect 13899 82760 13941 82769
rect 13899 82720 13900 82760
rect 13940 82720 13941 82760
rect 13899 82711 13941 82720
rect 13995 82760 14037 82769
rect 13995 82720 13996 82760
rect 14036 82720 14037 82760
rect 13995 82711 14037 82720
rect 14379 82760 14421 82769
rect 14379 82720 14380 82760
rect 14420 82720 14421 82760
rect 14379 82711 14421 82720
rect 14947 82760 15005 82761
rect 14947 82720 14956 82760
rect 14996 82720 15005 82760
rect 15435 82734 15436 82774
rect 15476 82734 15477 82774
rect 15435 82725 15477 82734
rect 15811 82760 15869 82761
rect 14947 82719 15005 82720
rect 15811 82720 15820 82760
rect 15860 82720 15869 82760
rect 15811 82719 15869 82720
rect 17059 82760 17117 82761
rect 17059 82720 17068 82760
rect 17108 82720 17117 82760
rect 17059 82719 17117 82720
rect 17443 82760 17501 82761
rect 17443 82720 17452 82760
rect 17492 82720 17501 82760
rect 17443 82719 17501 82720
rect 18691 82760 18749 82761
rect 18691 82720 18700 82760
rect 18740 82720 18749 82760
rect 18691 82719 18749 82720
rect 19467 82760 19509 82769
rect 19467 82720 19468 82760
rect 19508 82720 19509 82760
rect 19467 82711 19509 82720
rect 19747 82760 19805 82761
rect 19747 82720 19756 82760
rect 19796 82720 19805 82760
rect 19747 82719 19805 82720
rect 3427 82677 3485 82678
rect 10155 82676 10197 82685
rect 10155 82636 10156 82676
rect 10196 82636 10197 82676
rect 10155 82627 10197 82636
rect 18891 82676 18933 82685
rect 18891 82636 18892 82676
rect 18932 82636 18933 82676
rect 18891 82627 18933 82636
rect 19371 82676 19413 82685
rect 19371 82636 19372 82676
rect 19412 82636 19413 82676
rect 19371 82627 19413 82636
rect 2763 82592 2805 82601
rect 2763 82552 2764 82592
rect 2804 82552 2805 82592
rect 2763 82543 2805 82552
rect 3243 82592 3285 82601
rect 3243 82552 3244 82592
rect 3284 82552 3285 82592
rect 3243 82543 3285 82552
rect 4875 82592 4917 82601
rect 4875 82552 4876 82592
rect 4916 82552 4917 82592
rect 4875 82543 4917 82552
rect 8427 82592 8469 82601
rect 8427 82552 8428 82592
rect 8468 82552 8469 82592
rect 8427 82543 8469 82552
rect 12163 82592 12221 82593
rect 12163 82552 12172 82592
rect 12212 82552 12221 82592
rect 12163 82551 12221 82552
rect 12739 82592 12797 82593
rect 12739 82552 12748 82592
rect 12788 82552 12797 82592
rect 12739 82551 12797 82552
rect 12931 82592 12989 82593
rect 12931 82552 12940 82592
rect 12980 82552 12989 82592
rect 12931 82551 12989 82552
rect 13419 82592 13461 82601
rect 13419 82552 13420 82592
rect 13460 82552 13461 82592
rect 13419 82543 13461 82552
rect 15627 82592 15669 82601
rect 15627 82552 15628 82592
rect 15668 82552 15669 82592
rect 15627 82543 15669 82552
rect 17259 82592 17301 82601
rect 17259 82552 17260 82592
rect 17300 82552 17301 82592
rect 17259 82543 17301 82552
rect 1152 82424 20452 82448
rect 1152 82384 4928 82424
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 5296 82384 20048 82424
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20416 82384 20452 82424
rect 1152 82360 20452 82384
rect 3051 82256 3093 82265
rect 3051 82216 3052 82256
rect 3092 82216 3093 82256
rect 3051 82207 3093 82216
rect 3627 82256 3669 82265
rect 3627 82216 3628 82256
rect 3668 82216 3669 82256
rect 3627 82207 3669 82216
rect 4011 82256 4053 82265
rect 4011 82216 4012 82256
rect 4052 82216 4053 82256
rect 4011 82207 4053 82216
rect 4395 82256 4437 82265
rect 4395 82216 4396 82256
rect 4436 82216 4437 82256
rect 4395 82207 4437 82216
rect 6595 82256 6653 82257
rect 6595 82216 6604 82256
rect 6644 82216 6653 82256
rect 6595 82215 6653 82216
rect 6883 82256 6941 82257
rect 6883 82216 6892 82256
rect 6932 82216 6941 82256
rect 6883 82215 6941 82216
rect 7179 82256 7221 82265
rect 7179 82216 7180 82256
rect 7220 82216 7221 82256
rect 7179 82207 7221 82216
rect 10635 82256 10677 82265
rect 10635 82216 10636 82256
rect 10676 82216 10677 82256
rect 10635 82207 10677 82216
rect 11019 82256 11061 82265
rect 11019 82216 11020 82256
rect 11060 82216 11061 82256
rect 11019 82207 11061 82216
rect 12363 82256 12405 82265
rect 12363 82216 12364 82256
rect 12404 82216 12405 82256
rect 12363 82207 12405 82216
rect 6411 82172 6453 82181
rect 6411 82132 6412 82172
rect 6452 82132 6453 82172
rect 6411 82123 6453 82132
rect 14091 82172 14133 82181
rect 14091 82132 14092 82172
rect 14132 82132 14133 82172
rect 14091 82123 14133 82132
rect 16203 82172 16245 82181
rect 16203 82132 16204 82172
rect 16244 82132 16245 82172
rect 16203 82123 16245 82132
rect 1219 82088 1277 82089
rect 1219 82048 1228 82088
rect 1268 82048 1277 82088
rect 1219 82047 1277 82048
rect 2467 82088 2525 82089
rect 2467 82048 2476 82088
rect 2516 82048 2525 82088
rect 2467 82047 2525 82048
rect 4683 82088 4725 82097
rect 4683 82048 4684 82088
rect 4724 82048 4725 82088
rect 4683 82039 4725 82048
rect 4779 82088 4821 82097
rect 4779 82048 4780 82088
rect 4820 82048 4821 82088
rect 4779 82039 4821 82048
rect 5163 82088 5205 82097
rect 5163 82048 5164 82088
rect 5204 82048 5205 82088
rect 5163 82039 5205 82048
rect 5731 82088 5789 82089
rect 5731 82048 5740 82088
rect 5780 82048 5789 82088
rect 5731 82047 5789 82048
rect 6219 82083 6261 82092
rect 6219 82043 6220 82083
rect 6260 82043 6261 82083
rect 7555 82088 7613 82089
rect 7555 82048 7564 82088
rect 7604 82048 7613 82088
rect 7555 82047 7613 82048
rect 8803 82088 8861 82089
rect 8803 82048 8812 82088
rect 8852 82048 8861 82088
rect 8803 82047 8861 82048
rect 9187 82088 9245 82089
rect 9187 82048 9196 82088
rect 9236 82048 9245 82088
rect 9187 82047 9245 82048
rect 10435 82088 10493 82089
rect 10435 82048 10444 82088
rect 10484 82048 10493 82088
rect 10435 82047 10493 82048
rect 10827 82088 10869 82097
rect 10827 82048 10828 82088
rect 10868 82048 10869 82088
rect 6219 82034 6261 82043
rect 10827 82039 10869 82048
rect 11115 82088 11157 82097
rect 11115 82048 11116 82088
rect 11156 82048 11157 82088
rect 11115 82039 11157 82048
rect 11395 82088 11453 82089
rect 11395 82048 11404 82088
rect 11444 82048 11453 82088
rect 11395 82047 11453 82048
rect 11691 82088 11733 82097
rect 11691 82048 11692 82088
rect 11732 82048 11733 82088
rect 11691 82039 11733 82048
rect 11787 82088 11829 82097
rect 11787 82048 11788 82088
rect 11828 82048 11829 82088
rect 11787 82039 11829 82048
rect 12267 82088 12309 82097
rect 12267 82048 12268 82088
rect 12308 82048 12309 82088
rect 12267 82039 12309 82048
rect 12459 82088 12501 82097
rect 12459 82048 12460 82088
rect 12500 82048 12501 82088
rect 12459 82039 12501 82048
rect 12643 82088 12701 82089
rect 12643 82048 12652 82088
rect 12692 82048 12701 82088
rect 12643 82047 12701 82048
rect 13891 82088 13949 82089
rect 13891 82048 13900 82088
rect 13940 82048 13949 82088
rect 13891 82047 13949 82048
rect 14475 82088 14517 82097
rect 14475 82048 14476 82088
rect 14516 82048 14517 82088
rect 14475 82039 14517 82048
rect 14571 82088 14613 82097
rect 14571 82048 14572 82088
rect 14612 82048 14613 82088
rect 14571 82039 14613 82048
rect 15523 82088 15581 82089
rect 15523 82048 15532 82088
rect 15572 82048 15581 82088
rect 15523 82047 15581 82048
rect 16011 82083 16053 82092
rect 16011 82043 16012 82083
rect 16052 82043 16053 82083
rect 16771 82088 16829 82089
rect 16771 82048 16780 82088
rect 16820 82048 16829 82088
rect 16771 82047 16829 82048
rect 18019 82088 18077 82089
rect 18019 82048 18028 82088
rect 18068 82048 18077 82088
rect 18019 82047 18077 82048
rect 18595 82088 18653 82089
rect 18595 82048 18604 82088
rect 18644 82048 18653 82088
rect 18595 82047 18653 82048
rect 19843 82088 19901 82089
rect 19843 82048 19852 82088
rect 19892 82048 19901 82088
rect 19843 82047 19901 82048
rect 16011 82034 16053 82043
rect 2851 82004 2909 82005
rect 2851 81964 2860 82004
rect 2900 81964 2909 82004
rect 2851 81963 2909 81964
rect 3427 82004 3485 82005
rect 3427 81964 3436 82004
rect 3476 81964 3485 82004
rect 3427 81963 3485 81964
rect 3811 82004 3869 82005
rect 3811 81964 3820 82004
rect 3860 81964 3869 82004
rect 3811 81963 3869 81964
rect 4195 82004 4253 82005
rect 4195 81964 4204 82004
rect 4244 81964 4253 82004
rect 4195 81963 4253 81964
rect 5259 82004 5301 82013
rect 5259 81964 5260 82004
rect 5300 81964 5301 82004
rect 5259 81955 5301 81964
rect 7363 82004 7421 82005
rect 7363 81964 7372 82004
rect 7412 81964 7421 82004
rect 7363 81963 7421 81964
rect 14955 82004 14997 82013
rect 14955 81964 14956 82004
rect 14996 81964 14997 82004
rect 14955 81955 14997 81964
rect 15051 82004 15093 82013
rect 15051 81964 15052 82004
rect 15092 81964 15093 82004
rect 15051 81955 15093 81964
rect 16491 81920 16533 81929
rect 16491 81880 16492 81920
rect 16532 81880 16533 81920
rect 16491 81871 16533 81880
rect 2667 81836 2709 81845
rect 2667 81796 2668 81836
rect 2708 81796 2709 81836
rect 2667 81787 2709 81796
rect 9003 81836 9045 81845
rect 9003 81796 9004 81836
rect 9044 81796 9045 81836
rect 9003 81787 9045 81796
rect 12067 81836 12125 81837
rect 12067 81796 12076 81836
rect 12116 81796 12125 81836
rect 12067 81795 12125 81796
rect 18219 81836 18261 81845
rect 18219 81796 18220 81836
rect 18260 81796 18261 81836
rect 18219 81787 18261 81796
rect 20043 81836 20085 81845
rect 20043 81796 20044 81836
rect 20084 81796 20085 81836
rect 20043 81787 20085 81796
rect 1152 81668 20352 81692
rect 1152 81628 3688 81668
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 4056 81628 18808 81668
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 19176 81628 20352 81668
rect 1152 81604 20352 81628
rect 5355 81500 5397 81509
rect 5355 81460 5356 81500
rect 5396 81460 5397 81500
rect 5355 81451 5397 81460
rect 11691 81500 11733 81509
rect 11691 81460 11692 81500
rect 11732 81460 11733 81500
rect 11691 81451 11733 81460
rect 13611 81500 13653 81509
rect 13611 81460 13612 81500
rect 13652 81460 13653 81500
rect 13611 81451 13653 81460
rect 15723 81500 15765 81509
rect 15723 81460 15724 81500
rect 15764 81460 15765 81500
rect 15723 81451 15765 81460
rect 16587 81500 16629 81509
rect 16587 81460 16588 81500
rect 16628 81460 16629 81500
rect 16587 81451 16629 81460
rect 3051 81416 3093 81425
rect 3051 81376 3052 81416
rect 3092 81376 3093 81416
rect 3051 81367 3093 81376
rect 18603 81416 18645 81425
rect 18603 81376 18604 81416
rect 18644 81376 18645 81416
rect 18603 81367 18645 81376
rect 4011 81332 4053 81341
rect 4011 81292 4012 81332
rect 4052 81292 4053 81332
rect 4011 81283 4053 81292
rect 5539 81332 5597 81333
rect 5539 81292 5548 81332
rect 5588 81292 5597 81332
rect 5539 81291 5597 81292
rect 15907 81332 15965 81333
rect 15907 81292 15916 81332
rect 15956 81292 15965 81332
rect 15907 81291 15965 81292
rect 16387 81332 16445 81333
rect 16387 81292 16396 81332
rect 16436 81292 16445 81332
rect 16387 81291 16445 81292
rect 8899 81290 8957 81291
rect 4971 81262 5013 81271
rect 1219 81248 1277 81249
rect 1219 81208 1228 81248
rect 1268 81208 1277 81248
rect 1219 81207 1277 81208
rect 2467 81248 2525 81249
rect 2467 81208 2476 81248
rect 2516 81208 2525 81248
rect 2467 81207 2525 81208
rect 3435 81248 3477 81257
rect 3435 81208 3436 81248
rect 3476 81208 3477 81248
rect 3435 81199 3477 81208
rect 3531 81248 3573 81257
rect 3531 81208 3532 81248
rect 3572 81208 3573 81248
rect 3531 81199 3573 81208
rect 3915 81248 3957 81257
rect 3915 81208 3916 81248
rect 3956 81208 3957 81248
rect 3915 81199 3957 81208
rect 4483 81248 4541 81249
rect 4483 81208 4492 81248
rect 4532 81208 4541 81248
rect 4971 81222 4972 81262
rect 5012 81222 5013 81262
rect 4971 81213 5013 81222
rect 5731 81248 5789 81249
rect 4483 81207 4541 81208
rect 5731 81208 5740 81248
rect 5780 81208 5789 81248
rect 5731 81207 5789 81208
rect 6979 81248 7037 81249
rect 6979 81208 6988 81248
rect 7028 81208 7037 81248
rect 6979 81207 7037 81208
rect 7371 81248 7413 81257
rect 8899 81250 8908 81290
rect 8948 81250 8957 81290
rect 8899 81249 8957 81250
rect 7371 81208 7372 81248
rect 7412 81208 7413 81248
rect 7371 81199 7413 81208
rect 7651 81248 7709 81249
rect 7651 81208 7660 81248
rect 7700 81208 7709 81248
rect 7651 81207 7709 81208
rect 9475 81248 9533 81249
rect 9475 81208 9484 81248
rect 9524 81208 9533 81248
rect 9475 81207 9533 81208
rect 10723 81248 10781 81249
rect 10723 81208 10732 81248
rect 10772 81208 10781 81248
rect 10723 81207 10781 81208
rect 11211 81248 11253 81257
rect 11211 81208 11212 81248
rect 11252 81208 11253 81248
rect 11211 81199 11253 81208
rect 11307 81248 11349 81257
rect 11307 81208 11308 81248
rect 11348 81208 11349 81248
rect 11307 81199 11349 81208
rect 11403 81248 11445 81257
rect 11403 81208 11404 81248
rect 11444 81208 11445 81248
rect 11403 81199 11445 81208
rect 11499 81248 11541 81257
rect 11499 81208 11500 81248
rect 11540 81208 11541 81248
rect 11499 81199 11541 81208
rect 11691 81248 11733 81257
rect 11691 81208 11692 81248
rect 11732 81208 11733 81248
rect 11691 81199 11733 81208
rect 11883 81248 11925 81257
rect 11883 81208 11884 81248
rect 11924 81208 11925 81248
rect 11883 81199 11925 81208
rect 11971 81248 12029 81249
rect 11971 81208 11980 81248
rect 12020 81208 12029 81248
rect 11971 81207 12029 81208
rect 12163 81248 12221 81249
rect 12163 81208 12172 81248
rect 12212 81208 12221 81248
rect 12163 81207 12221 81208
rect 13411 81248 13469 81249
rect 13411 81208 13420 81248
rect 13460 81208 13469 81248
rect 13411 81207 13469 81208
rect 13795 81248 13853 81249
rect 13795 81208 13804 81248
rect 13844 81208 13853 81248
rect 13795 81207 13853 81208
rect 15043 81248 15101 81249
rect 15043 81208 15052 81248
rect 15092 81208 15101 81248
rect 15043 81207 15101 81208
rect 16771 81248 16829 81249
rect 16771 81208 16780 81248
rect 16820 81208 16829 81248
rect 16771 81207 16829 81208
rect 18019 81248 18077 81249
rect 18019 81208 18028 81248
rect 18068 81208 18077 81248
rect 18019 81207 18077 81208
rect 18787 81248 18845 81249
rect 18787 81208 18796 81248
rect 18836 81208 18845 81248
rect 18787 81207 18845 81208
rect 20035 81248 20093 81249
rect 20035 81208 20044 81248
rect 20084 81208 20093 81248
rect 20035 81207 20093 81208
rect 5163 81164 5205 81173
rect 5163 81124 5164 81164
rect 5204 81124 5205 81164
rect 5163 81115 5205 81124
rect 2667 81080 2709 81089
rect 2667 81040 2668 81080
rect 2708 81040 2709 81080
rect 2667 81031 2709 81040
rect 3147 81080 3189 81089
rect 3147 81040 3148 81080
rect 3188 81040 3189 81080
rect 3147 81031 3189 81040
rect 7179 81080 7221 81089
rect 7179 81040 7180 81080
rect 7220 81040 7221 81080
rect 7179 81031 7221 81040
rect 9099 81080 9141 81089
rect 9099 81040 9100 81080
rect 9140 81040 9141 81080
rect 9099 81031 9141 81040
rect 9291 81080 9333 81089
rect 9291 81040 9292 81080
rect 9332 81040 9333 81080
rect 9291 81031 9333 81040
rect 15243 81080 15285 81089
rect 15243 81040 15244 81080
rect 15284 81040 15285 81080
rect 15243 81031 15285 81040
rect 15435 81080 15477 81089
rect 15435 81040 15436 81080
rect 15476 81040 15477 81080
rect 15435 81031 15477 81040
rect 16099 81080 16157 81081
rect 16099 81040 16108 81080
rect 16148 81040 16157 81080
rect 16099 81039 16157 81040
rect 18219 81080 18261 81089
rect 18219 81040 18220 81080
rect 18260 81040 18261 81080
rect 18219 81031 18261 81040
rect 18499 81080 18557 81081
rect 18499 81040 18508 81080
rect 18548 81040 18557 81080
rect 18499 81039 18557 81040
rect 20235 81080 20277 81089
rect 20235 81040 20236 81080
rect 20276 81040 20277 81080
rect 20235 81031 20277 81040
rect 1152 80912 20452 80936
rect 1152 80872 4928 80912
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 5296 80872 20048 80912
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20416 80872 20452 80912
rect 1152 80848 20452 80872
rect 3331 80744 3389 80745
rect 3331 80704 3340 80744
rect 3380 80704 3389 80744
rect 3331 80703 3389 80704
rect 3723 80744 3765 80753
rect 3723 80704 3724 80744
rect 3764 80704 3765 80744
rect 3723 80695 3765 80704
rect 11883 80744 11925 80753
rect 11883 80704 11884 80744
rect 11924 80704 11925 80744
rect 11883 80695 11925 80704
rect 3051 80660 3093 80669
rect 3051 80620 3052 80660
rect 3092 80620 3093 80660
rect 3051 80611 3093 80620
rect 9195 80660 9237 80669
rect 9195 80620 9196 80660
rect 9236 80620 9237 80660
rect 9195 80611 9237 80620
rect 11499 80660 11541 80669
rect 11499 80620 11500 80660
rect 11540 80620 11541 80660
rect 11499 80611 11541 80620
rect 13515 80660 13557 80669
rect 13515 80620 13516 80660
rect 13556 80620 13557 80660
rect 13515 80611 13557 80620
rect 15531 80660 15573 80669
rect 15531 80620 15532 80660
rect 15572 80620 15573 80660
rect 15531 80611 15573 80620
rect 1323 80576 1365 80585
rect 1323 80536 1324 80576
rect 1364 80536 1365 80576
rect 1323 80527 1365 80536
rect 1419 80576 1461 80585
rect 1419 80536 1420 80576
rect 1460 80536 1461 80576
rect 1419 80527 1461 80536
rect 2371 80576 2429 80577
rect 2371 80536 2380 80576
rect 2420 80536 2429 80576
rect 2371 80535 2429 80536
rect 2859 80571 2901 80580
rect 2859 80531 2860 80571
rect 2900 80531 2901 80571
rect 4387 80576 4445 80577
rect 2859 80522 2901 80531
rect 3867 80534 3909 80543
rect 4387 80536 4396 80576
rect 4436 80536 4445 80576
rect 4387 80535 4445 80536
rect 4971 80576 5013 80585
rect 4971 80536 4972 80576
rect 5012 80536 5013 80576
rect 1803 80492 1845 80501
rect 1803 80452 1804 80492
rect 1844 80452 1845 80492
rect 1803 80443 1845 80452
rect 1899 80492 1941 80501
rect 1899 80452 1900 80492
rect 1940 80452 1941 80492
rect 3867 80494 3868 80534
rect 3908 80494 3909 80534
rect 4971 80527 5013 80536
rect 5355 80576 5397 80585
rect 5355 80536 5356 80576
rect 5396 80536 5397 80576
rect 5355 80527 5397 80536
rect 5451 80576 5493 80585
rect 5451 80536 5452 80576
rect 5492 80536 5493 80576
rect 5451 80527 5493 80536
rect 6027 80576 6069 80585
rect 6027 80536 6028 80576
rect 6068 80536 6069 80576
rect 6027 80527 6069 80536
rect 6219 80576 6261 80585
rect 6219 80536 6220 80576
rect 6260 80536 6261 80576
rect 6219 80527 6261 80536
rect 6603 80576 6645 80585
rect 6603 80536 6604 80576
rect 6644 80536 6645 80576
rect 6603 80527 6645 80536
rect 6891 80576 6933 80585
rect 6891 80536 6892 80576
rect 6932 80536 6933 80576
rect 6891 80527 6933 80536
rect 7467 80576 7509 80585
rect 7467 80536 7468 80576
rect 7508 80536 7509 80576
rect 7467 80527 7509 80536
rect 7563 80576 7605 80585
rect 7563 80536 7564 80576
rect 7604 80536 7605 80576
rect 7563 80527 7605 80536
rect 8515 80576 8573 80577
rect 8515 80536 8524 80576
rect 8564 80536 8573 80576
rect 8515 80535 8573 80536
rect 9003 80571 9045 80580
rect 9003 80531 9004 80571
rect 9044 80531 9045 80571
rect 9003 80522 9045 80531
rect 9771 80576 9813 80585
rect 9771 80536 9772 80576
rect 9812 80536 9813 80576
rect 9771 80527 9813 80536
rect 9867 80576 9909 80585
rect 9867 80536 9868 80576
rect 9908 80536 9909 80576
rect 9867 80527 9909 80536
rect 10819 80576 10877 80577
rect 10819 80536 10828 80576
rect 10868 80536 10877 80576
rect 11779 80576 11837 80577
rect 10819 80535 10877 80536
rect 11355 80566 11397 80575
rect 11355 80526 11356 80566
rect 11396 80526 11397 80566
rect 11779 80536 11788 80576
rect 11828 80536 11837 80576
rect 11779 80535 11837 80536
rect 12067 80576 12125 80577
rect 12067 80536 12076 80576
rect 12116 80536 12125 80576
rect 12067 80535 12125 80536
rect 13315 80576 13373 80577
rect 13315 80536 13324 80576
rect 13364 80536 13373 80576
rect 13315 80535 13373 80536
rect 13803 80576 13845 80585
rect 13803 80536 13804 80576
rect 13844 80536 13845 80576
rect 13803 80527 13845 80536
rect 13899 80576 13941 80585
rect 13899 80536 13900 80576
rect 13940 80536 13941 80576
rect 13899 80527 13941 80536
rect 14379 80576 14421 80585
rect 14379 80536 14380 80576
rect 14420 80536 14421 80576
rect 14379 80527 14421 80536
rect 14851 80576 14909 80577
rect 14851 80536 14860 80576
rect 14900 80536 14909 80576
rect 14851 80535 14909 80536
rect 15339 80571 15381 80580
rect 15339 80531 15340 80571
rect 15380 80531 15381 80571
rect 11355 80517 11397 80526
rect 15339 80522 15381 80531
rect 15819 80576 15861 80585
rect 15819 80536 15820 80576
rect 15860 80536 15861 80576
rect 15819 80527 15861 80536
rect 16011 80576 16053 80585
rect 16011 80536 16012 80576
rect 16052 80536 16053 80576
rect 16011 80527 16053 80536
rect 16203 80576 16245 80585
rect 16203 80536 16204 80576
rect 16244 80536 16245 80576
rect 16203 80527 16245 80536
rect 16491 80576 16533 80585
rect 16491 80536 16492 80576
rect 16532 80536 16533 80576
rect 16491 80527 16533 80536
rect 16867 80576 16925 80577
rect 16867 80536 16876 80576
rect 16916 80536 16925 80576
rect 16867 80535 16925 80536
rect 18115 80576 18173 80577
rect 18115 80536 18124 80576
rect 18164 80536 18173 80576
rect 18115 80535 18173 80536
rect 18883 80576 18941 80577
rect 18883 80536 18892 80576
rect 18932 80536 18941 80576
rect 18883 80535 18941 80536
rect 20131 80534 20189 80535
rect 3867 80485 3909 80494
rect 4875 80492 4917 80501
rect 1899 80443 1941 80452
rect 4875 80452 4876 80492
rect 4916 80452 4917 80492
rect 4875 80443 4917 80452
rect 5739 80492 5781 80501
rect 5739 80452 5740 80492
rect 5780 80452 5781 80492
rect 5739 80443 5781 80452
rect 6795 80492 6837 80501
rect 6795 80452 6796 80492
rect 6836 80452 6837 80492
rect 6795 80443 6837 80452
rect 7083 80492 7125 80501
rect 7083 80452 7084 80492
rect 7124 80452 7125 80492
rect 7083 80443 7125 80452
rect 7947 80492 7989 80501
rect 7947 80452 7948 80492
rect 7988 80452 7989 80492
rect 7947 80443 7989 80452
rect 8043 80492 8085 80501
rect 8043 80452 8044 80492
rect 8084 80452 8085 80492
rect 8043 80443 8085 80452
rect 10251 80492 10293 80501
rect 10251 80452 10252 80492
rect 10292 80452 10293 80492
rect 10251 80443 10293 80452
rect 10347 80492 10389 80501
rect 10347 80452 10348 80492
rect 10388 80452 10389 80492
rect 10347 80443 10389 80452
rect 14283 80492 14325 80501
rect 20131 80494 20140 80534
rect 20180 80494 20189 80534
rect 20131 80493 20189 80494
rect 14283 80452 14284 80492
rect 14324 80452 14325 80492
rect 14283 80443 14325 80452
rect 6027 80408 6069 80417
rect 6027 80368 6028 80408
rect 6068 80368 6069 80408
rect 6027 80359 6069 80368
rect 18507 80408 18549 80417
rect 18507 80368 18508 80408
rect 18548 80368 18549 80408
rect 18507 80359 18549 80368
rect 15819 80324 15861 80333
rect 15819 80284 15820 80324
rect 15860 80284 15861 80324
rect 15819 80275 15861 80284
rect 16203 80324 16245 80333
rect 16203 80284 16204 80324
rect 16244 80284 16245 80324
rect 16203 80275 16245 80284
rect 16683 80324 16725 80333
rect 16683 80284 16684 80324
rect 16724 80284 16725 80324
rect 16683 80275 16725 80284
rect 18699 80324 18741 80333
rect 18699 80284 18700 80324
rect 18740 80284 18741 80324
rect 18699 80275 18741 80284
rect 1152 80156 20352 80180
rect 1152 80116 3688 80156
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 4056 80116 18808 80156
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 19176 80116 20352 80156
rect 1152 80092 20352 80116
rect 3531 79988 3573 79997
rect 3531 79948 3532 79988
rect 3572 79948 3573 79988
rect 3531 79939 3573 79948
rect 15531 79988 15573 79997
rect 15531 79948 15532 79988
rect 15572 79948 15573 79988
rect 15531 79939 15573 79948
rect 7467 79820 7509 79829
rect 7467 79780 7468 79820
rect 7508 79780 7509 79820
rect 7467 79771 7509 79780
rect 16299 79820 16341 79829
rect 16299 79780 16300 79820
rect 16340 79780 16341 79820
rect 16299 79771 16341 79780
rect 16395 79820 16437 79829
rect 16395 79780 16396 79820
rect 16436 79780 16437 79820
rect 16395 79771 16437 79780
rect 12355 79757 12413 79758
rect 1406 79736 1464 79737
rect 1406 79696 1415 79736
rect 1455 79696 1464 79736
rect 1406 79695 1464 79696
rect 1515 79736 1557 79745
rect 1515 79696 1516 79736
rect 1556 79696 1557 79736
rect 1515 79687 1557 79696
rect 1611 79736 1653 79745
rect 1611 79696 1612 79736
rect 1652 79696 1653 79736
rect 1611 79687 1653 79696
rect 1795 79736 1853 79737
rect 1795 79696 1804 79736
rect 1844 79696 1853 79736
rect 1795 79695 1853 79696
rect 1891 79736 1949 79737
rect 1891 79696 1900 79736
rect 1940 79696 1949 79736
rect 1891 79695 1949 79696
rect 2083 79736 2141 79737
rect 2083 79696 2092 79736
rect 2132 79696 2141 79736
rect 2083 79695 2141 79696
rect 3331 79736 3389 79737
rect 3331 79696 3340 79736
rect 3380 79696 3389 79736
rect 3331 79695 3389 79696
rect 4003 79736 4061 79737
rect 4003 79696 4012 79736
rect 4052 79696 4061 79736
rect 4003 79695 4061 79696
rect 5251 79736 5309 79737
rect 5251 79696 5260 79736
rect 5300 79696 5309 79736
rect 5251 79695 5309 79696
rect 5731 79736 5789 79737
rect 5731 79696 5740 79736
rect 5780 79696 5789 79736
rect 5731 79695 5789 79696
rect 6979 79736 7037 79737
rect 6979 79696 6988 79736
rect 7028 79696 7037 79736
rect 6979 79695 7037 79696
rect 7843 79736 7901 79737
rect 7843 79696 7852 79736
rect 7892 79696 7901 79736
rect 7843 79695 7901 79696
rect 9091 79736 9149 79737
rect 9091 79696 9100 79736
rect 9140 79696 9149 79736
rect 9091 79695 9149 79696
rect 9475 79736 9533 79737
rect 9475 79696 9484 79736
rect 9524 79696 9533 79736
rect 9475 79695 9533 79696
rect 10723 79736 10781 79737
rect 10723 79696 10732 79736
rect 10772 79696 10781 79736
rect 10723 79695 10781 79696
rect 11107 79736 11165 79737
rect 11107 79696 11116 79736
rect 11156 79696 11165 79736
rect 12355 79717 12364 79757
rect 12404 79717 12413 79757
rect 17355 79750 17397 79759
rect 12355 79716 12413 79717
rect 13699 79736 13757 79737
rect 11107 79695 11165 79696
rect 13699 79696 13708 79736
rect 13748 79696 13757 79736
rect 13699 79695 13757 79696
rect 14947 79736 15005 79737
rect 14947 79696 14956 79736
rect 14996 79696 15005 79736
rect 14947 79695 15005 79696
rect 15339 79736 15381 79745
rect 15339 79696 15340 79736
rect 15380 79696 15381 79736
rect 15339 79687 15381 79696
rect 15531 79736 15573 79745
rect 15531 79696 15532 79736
rect 15572 79696 15573 79736
rect 15531 79687 15573 79696
rect 15819 79736 15861 79745
rect 15819 79696 15820 79736
rect 15860 79696 15861 79736
rect 15819 79687 15861 79696
rect 15915 79736 15957 79745
rect 15915 79696 15916 79736
rect 15956 79696 15957 79736
rect 15915 79687 15957 79696
rect 16867 79736 16925 79737
rect 16867 79696 16876 79736
rect 16916 79696 16925 79736
rect 17355 79710 17356 79750
rect 17396 79710 17397 79750
rect 17355 79701 17397 79710
rect 17931 79750 17973 79759
rect 17931 79710 17932 79750
rect 17972 79710 17973 79750
rect 19467 79755 19509 79764
rect 17931 79701 17973 79710
rect 18403 79736 18461 79737
rect 16867 79695 16925 79696
rect 18403 79696 18412 79736
rect 18452 79696 18461 79736
rect 18403 79695 18461 79696
rect 18891 79736 18933 79745
rect 18891 79696 18892 79736
rect 18932 79696 18933 79736
rect 18891 79687 18933 79696
rect 18987 79736 19029 79745
rect 18987 79696 18988 79736
rect 19028 79696 19029 79736
rect 18987 79687 19029 79696
rect 19371 79736 19413 79745
rect 19371 79696 19372 79736
rect 19412 79696 19413 79736
rect 19467 79715 19468 79755
rect 19508 79715 19509 79755
rect 19467 79706 19509 79715
rect 19755 79736 19797 79745
rect 19371 79687 19413 79696
rect 19755 79696 19756 79736
rect 19796 79696 19797 79736
rect 19755 79687 19797 79696
rect 19851 79736 19893 79745
rect 19851 79696 19852 79736
rect 19892 79696 19893 79736
rect 19851 79687 19893 79696
rect 19947 79736 19989 79745
rect 19947 79696 19948 79736
rect 19988 79696 19989 79736
rect 19947 79687 19989 79696
rect 15147 79652 15189 79661
rect 15147 79612 15148 79652
rect 15188 79612 15189 79652
rect 15147 79603 15189 79612
rect 17739 79652 17781 79661
rect 17739 79612 17740 79652
rect 17780 79612 17781 79652
rect 17739 79603 17781 79612
rect 1411 79568 1469 79569
rect 1411 79528 1420 79568
rect 1460 79528 1469 79568
rect 1411 79527 1469 79528
rect 3819 79568 3861 79577
rect 3819 79528 3820 79568
rect 3860 79528 3861 79568
rect 3819 79519 3861 79528
rect 5451 79568 5493 79577
rect 5451 79528 5452 79568
rect 5492 79528 5493 79568
rect 5451 79519 5493 79528
rect 7179 79568 7221 79577
rect 7179 79528 7180 79568
rect 7220 79528 7221 79568
rect 7179 79519 7221 79528
rect 9291 79568 9333 79577
rect 9291 79528 9292 79568
rect 9332 79528 9333 79568
rect 9291 79519 9333 79528
rect 10923 79568 10965 79577
rect 10923 79528 10924 79568
rect 10964 79528 10965 79568
rect 10923 79519 10965 79528
rect 12555 79568 12597 79577
rect 12555 79528 12556 79568
rect 12596 79528 12597 79568
rect 12555 79519 12597 79528
rect 17547 79568 17589 79577
rect 17547 79528 17548 79568
rect 17588 79528 17589 79568
rect 17547 79519 17589 79528
rect 20035 79568 20093 79569
rect 20035 79528 20044 79568
rect 20084 79528 20093 79568
rect 20035 79527 20093 79528
rect 1152 79400 20452 79424
rect 1152 79360 4928 79400
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 5296 79360 20048 79400
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20416 79360 20452 79400
rect 1152 79336 20452 79360
rect 3051 79232 3093 79241
rect 3051 79192 3052 79232
rect 3092 79192 3093 79232
rect 3051 79183 3093 79192
rect 7467 79232 7509 79241
rect 7467 79192 7468 79232
rect 7508 79192 7509 79232
rect 7467 79183 7509 79192
rect 17547 79232 17589 79241
rect 17547 79192 17548 79232
rect 17588 79192 17589 79232
rect 17547 79183 17589 79192
rect 18115 79232 18173 79233
rect 18115 79192 18124 79232
rect 18164 79192 18173 79232
rect 18115 79191 18173 79192
rect 10251 79148 10293 79157
rect 10251 79108 10252 79148
rect 10292 79108 10293 79148
rect 10251 79099 10293 79108
rect 12363 79148 12405 79157
rect 12363 79108 12364 79148
rect 12404 79108 12405 79148
rect 12363 79099 12405 79108
rect 20139 79148 20181 79157
rect 20139 79108 20140 79148
rect 20180 79108 20181 79148
rect 20139 79099 20181 79108
rect 1219 79064 1277 79065
rect 1219 79024 1228 79064
rect 1268 79024 1277 79064
rect 1219 79023 1277 79024
rect 2467 79064 2525 79065
rect 2467 79024 2476 79064
rect 2516 79024 2525 79064
rect 2467 79023 2525 79024
rect 3235 79064 3293 79065
rect 3235 79024 3244 79064
rect 3284 79024 3293 79064
rect 3235 79023 3293 79024
rect 4483 79064 4541 79065
rect 4483 79024 4492 79064
rect 4532 79024 4541 79064
rect 4483 79023 4541 79024
rect 4963 79064 5021 79065
rect 4963 79024 4972 79064
rect 5012 79024 5021 79064
rect 4963 79023 5021 79024
rect 6211 79064 6269 79065
rect 6211 79024 6220 79064
rect 6260 79024 6269 79064
rect 6211 79023 6269 79024
rect 6891 79064 6933 79073
rect 6891 79024 6892 79064
rect 6932 79024 6933 79064
rect 6891 79015 6933 79024
rect 6987 79064 7029 79073
rect 6987 79024 6988 79064
rect 7028 79024 7029 79064
rect 6987 79015 7029 79024
rect 7083 79064 7125 79073
rect 7083 79024 7084 79064
rect 7124 79024 7125 79064
rect 7083 79015 7125 79024
rect 7179 79064 7221 79073
rect 7179 79024 7180 79064
rect 7220 79024 7221 79064
rect 7179 79015 7221 79024
rect 7755 79064 7797 79073
rect 7755 79024 7756 79064
rect 7796 79024 7797 79064
rect 7755 79015 7797 79024
rect 7947 79064 7989 79073
rect 7947 79024 7948 79064
rect 7988 79024 7989 79064
rect 7947 79015 7989 79024
rect 8035 79064 8093 79065
rect 8035 79024 8044 79064
rect 8084 79024 8093 79064
rect 8035 79023 8093 79024
rect 8235 79064 8277 79073
rect 8235 79024 8236 79064
rect 8276 79024 8277 79064
rect 8235 79015 8277 79024
rect 8427 79064 8469 79073
rect 8427 79024 8428 79064
rect 8468 79024 8469 79064
rect 8427 79015 8469 79024
rect 8803 79064 8861 79065
rect 8803 79024 8812 79064
rect 8852 79024 8861 79064
rect 8803 79023 8861 79024
rect 10051 79064 10109 79065
rect 10051 79024 10060 79064
rect 10100 79024 10109 79064
rect 10051 79023 10109 79024
rect 10635 79064 10677 79073
rect 10635 79024 10636 79064
rect 10676 79024 10677 79064
rect 10635 79015 10677 79024
rect 10731 79064 10773 79073
rect 10731 79024 10732 79064
rect 10772 79024 10773 79064
rect 10731 79015 10773 79024
rect 11211 79064 11253 79073
rect 11211 79024 11212 79064
rect 11252 79024 11253 79064
rect 11211 79015 11253 79024
rect 11683 79064 11741 79065
rect 11683 79024 11692 79064
rect 11732 79024 11741 79064
rect 12547 79064 12605 79065
rect 11683 79023 11741 79024
rect 12219 79054 12261 79063
rect 12219 79014 12220 79054
rect 12260 79014 12261 79054
rect 12547 79024 12556 79064
rect 12596 79024 12605 79064
rect 12547 79023 12605 79024
rect 13795 79064 13853 79065
rect 13795 79024 13804 79064
rect 13844 79024 13853 79064
rect 13795 79023 13853 79024
rect 14371 79064 14429 79065
rect 14371 79024 14380 79064
rect 14420 79024 14429 79064
rect 14371 79023 14429 79024
rect 15619 79064 15677 79065
rect 15619 79024 15628 79064
rect 15668 79024 15677 79064
rect 15619 79023 15677 79024
rect 15907 79064 15965 79065
rect 15907 79024 15916 79064
rect 15956 79024 15965 79064
rect 15907 79023 15965 79024
rect 17155 79064 17213 79065
rect 17155 79024 17164 79064
rect 17204 79024 17213 79064
rect 17155 79023 17213 79024
rect 17635 79064 17693 79065
rect 17635 79024 17644 79064
rect 17684 79024 17693 79064
rect 17635 79023 17693 79024
rect 17835 79064 17877 79073
rect 17835 79024 17836 79064
rect 17876 79024 17877 79064
rect 17835 79015 17877 79024
rect 17931 79064 17973 79073
rect 17931 79024 17932 79064
rect 17972 79024 17973 79064
rect 17931 79015 17973 79024
rect 18027 79064 18069 79073
rect 18027 79024 18028 79064
rect 18068 79024 18069 79064
rect 19459 79064 19517 79065
rect 18027 79015 18069 79024
rect 18411 79045 18453 79054
rect 12219 79005 12261 79014
rect 18411 79005 18412 79045
rect 18452 79005 18453 79045
rect 18411 78996 18453 79005
rect 18507 79045 18549 79054
rect 18507 79005 18508 79045
rect 18548 79005 18549 79045
rect 19459 79024 19468 79064
rect 19508 79024 19517 79064
rect 19459 79023 19517 79024
rect 19947 79059 19989 79068
rect 19947 79019 19948 79059
rect 19988 79019 19989 79059
rect 19947 79010 19989 79019
rect 18507 78996 18549 79005
rect 2851 78980 2909 78981
rect 2851 78940 2860 78980
rect 2900 78940 2909 78980
rect 2851 78939 2909 78940
rect 11115 78980 11157 78989
rect 11115 78940 11116 78980
rect 11156 78940 11157 78980
rect 11115 78931 11157 78940
rect 18891 78980 18933 78989
rect 18891 78940 18892 78980
rect 18932 78940 18933 78980
rect 18891 78931 18933 78940
rect 18987 78980 19029 78989
rect 18987 78940 18988 78980
rect 19028 78940 19029 78980
rect 18987 78931 19029 78940
rect 7371 78896 7413 78905
rect 7371 78856 7372 78896
rect 7412 78856 7413 78896
rect 7371 78847 7413 78856
rect 7755 78896 7797 78905
rect 7755 78856 7756 78896
rect 7796 78856 7797 78896
rect 7755 78847 7797 78856
rect 8235 78896 8277 78905
rect 8235 78856 8236 78896
rect 8276 78856 8277 78896
rect 8235 78847 8277 78856
rect 2667 78812 2709 78821
rect 2667 78772 2668 78812
rect 2708 78772 2709 78812
rect 2667 78763 2709 78772
rect 4683 78812 4725 78821
rect 4683 78772 4684 78812
rect 4724 78772 4725 78812
rect 4683 78763 4725 78772
rect 6411 78812 6453 78821
rect 6411 78772 6412 78812
rect 6452 78772 6453 78812
rect 6411 78763 6453 78772
rect 13995 78812 14037 78821
rect 13995 78772 13996 78812
rect 14036 78772 14037 78812
rect 13995 78763 14037 78772
rect 14187 78812 14229 78821
rect 14187 78772 14188 78812
rect 14228 78772 14229 78812
rect 14187 78763 14229 78772
rect 17355 78812 17397 78821
rect 17355 78772 17356 78812
rect 17396 78772 17397 78812
rect 17355 78763 17397 78772
rect 1152 78644 20352 78668
rect 1152 78604 3688 78644
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 4056 78604 18808 78644
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 19176 78604 20352 78644
rect 1152 78580 20352 78604
rect 5355 78476 5397 78485
rect 5355 78436 5356 78476
rect 5396 78436 5397 78476
rect 5355 78427 5397 78436
rect 7083 78476 7125 78485
rect 7083 78436 7084 78476
rect 7124 78436 7125 78476
rect 7083 78427 7125 78436
rect 8035 78476 8093 78477
rect 8035 78436 8044 78476
rect 8084 78436 8093 78476
rect 8035 78435 8093 78436
rect 17643 78476 17685 78485
rect 17643 78436 17644 78476
rect 17684 78436 17685 78476
rect 17643 78427 17685 78436
rect 18507 78476 18549 78485
rect 18507 78436 18508 78476
rect 18548 78436 18549 78476
rect 18507 78427 18549 78436
rect 3531 78308 3573 78317
rect 3531 78268 3532 78308
rect 3572 78268 3573 78308
rect 3531 78259 3573 78268
rect 11115 78308 11157 78317
rect 11115 78268 11116 78308
rect 11156 78268 11157 78308
rect 11115 78259 11157 78268
rect 13803 78308 13845 78317
rect 13803 78268 13804 78308
rect 13844 78268 13845 78308
rect 13803 78259 13845 78268
rect 15819 78308 15861 78317
rect 15819 78268 15820 78308
rect 15860 78268 15861 78308
rect 15819 78259 15861 78268
rect 17443 78308 17501 78309
rect 17443 78268 17452 78308
rect 17492 78268 17501 78308
rect 17443 78267 17501 78268
rect 17827 78308 17885 78309
rect 17827 78268 17836 78308
rect 17876 78268 17885 78308
rect 17827 78267 17885 78268
rect 18027 78308 18069 78317
rect 18027 78268 18028 78308
rect 18068 78268 18069 78308
rect 18027 78259 18069 78268
rect 18307 78308 18365 78309
rect 18307 78268 18316 78308
rect 18356 78268 18365 78308
rect 18307 78267 18365 78268
rect 4491 78238 4533 78247
rect 14859 78238 14901 78247
rect 1219 78224 1277 78225
rect 1219 78184 1228 78224
rect 1268 78184 1277 78224
rect 1219 78183 1277 78184
rect 2467 78224 2525 78225
rect 2467 78184 2476 78224
rect 2516 78184 2525 78224
rect 2467 78183 2525 78184
rect 2955 78224 2997 78233
rect 2955 78184 2956 78224
rect 2996 78184 2997 78224
rect 2955 78175 2997 78184
rect 3051 78224 3093 78233
rect 3051 78184 3052 78224
rect 3092 78184 3093 78224
rect 3051 78175 3093 78184
rect 3435 78224 3477 78233
rect 3435 78184 3436 78224
rect 3476 78184 3477 78224
rect 3435 78175 3477 78184
rect 4003 78224 4061 78225
rect 4003 78184 4012 78224
rect 4052 78184 4061 78224
rect 4491 78198 4492 78238
rect 4532 78198 4533 78238
rect 4491 78189 4533 78198
rect 4875 78224 4917 78233
rect 4003 78183 4061 78184
rect 4875 78184 4876 78224
rect 4916 78184 4917 78224
rect 4875 78175 4917 78184
rect 4971 78224 5013 78233
rect 4971 78184 4972 78224
rect 5012 78184 5013 78224
rect 4971 78175 5013 78184
rect 5443 78224 5501 78225
rect 5443 78184 5452 78224
rect 5492 78184 5501 78224
rect 5443 78183 5501 78184
rect 5635 78224 5693 78225
rect 5635 78184 5644 78224
rect 5684 78184 5693 78224
rect 5635 78183 5693 78184
rect 6883 78224 6941 78225
rect 6883 78184 6892 78224
rect 6932 78184 6941 78224
rect 6883 78183 6941 78184
rect 7363 78224 7421 78225
rect 7363 78184 7372 78224
rect 7412 78184 7421 78224
rect 7363 78183 7421 78184
rect 7659 78224 7701 78233
rect 7659 78184 7660 78224
rect 7700 78184 7701 78224
rect 7659 78175 7701 78184
rect 7755 78224 7797 78233
rect 7755 78184 7756 78224
rect 7796 78184 7797 78224
rect 7755 78175 7797 78184
rect 8419 78224 8477 78225
rect 8419 78184 8428 78224
rect 8468 78184 8477 78224
rect 8419 78183 8477 78184
rect 9667 78224 9725 78225
rect 9667 78184 9676 78224
rect 9716 78184 9725 78224
rect 9667 78183 9725 78184
rect 10539 78224 10581 78233
rect 10539 78184 10540 78224
rect 10580 78184 10581 78224
rect 10539 78175 10581 78184
rect 10635 78224 10677 78233
rect 10635 78184 10636 78224
rect 10676 78184 10677 78224
rect 10635 78175 10677 78184
rect 11019 78224 11061 78233
rect 12075 78229 12117 78238
rect 11019 78184 11020 78224
rect 11060 78184 11061 78224
rect 11019 78175 11061 78184
rect 11587 78224 11645 78225
rect 11587 78184 11596 78224
rect 11636 78184 11645 78224
rect 11587 78183 11645 78184
rect 12075 78189 12076 78229
rect 12116 78189 12117 78229
rect 12075 78180 12117 78189
rect 13323 78224 13365 78233
rect 13323 78184 13324 78224
rect 13364 78184 13365 78224
rect 13323 78175 13365 78184
rect 13419 78224 13461 78233
rect 13419 78184 13420 78224
rect 13460 78184 13461 78224
rect 13419 78175 13461 78184
rect 13899 78224 13941 78233
rect 13899 78184 13900 78224
rect 13940 78184 13941 78224
rect 13899 78175 13941 78184
rect 14371 78224 14429 78225
rect 14371 78184 14380 78224
rect 14420 78184 14429 78224
rect 14859 78198 14860 78238
rect 14900 78198 14901 78238
rect 16875 78238 16917 78247
rect 14859 78189 14901 78198
rect 15339 78224 15381 78233
rect 14371 78183 14429 78184
rect 15339 78184 15340 78224
rect 15380 78184 15381 78224
rect 15339 78175 15381 78184
rect 15435 78224 15477 78233
rect 15435 78184 15436 78224
rect 15476 78184 15477 78224
rect 15435 78175 15477 78184
rect 15915 78224 15957 78233
rect 15915 78184 15916 78224
rect 15956 78184 15957 78224
rect 15915 78175 15957 78184
rect 16387 78224 16445 78225
rect 16387 78184 16396 78224
rect 16436 78184 16445 78224
rect 16875 78198 16876 78238
rect 16916 78198 16917 78238
rect 16875 78189 16917 78198
rect 18691 78224 18749 78225
rect 16387 78183 16445 78184
rect 18691 78184 18700 78224
rect 18740 78184 18749 78224
rect 18691 78183 18749 78184
rect 19939 78224 19997 78225
rect 19939 78184 19948 78224
rect 19988 78184 19997 78224
rect 19939 78183 19997 78184
rect 2667 78140 2709 78149
rect 2667 78100 2668 78140
rect 2708 78100 2709 78140
rect 2667 78091 2709 78100
rect 4683 78140 4725 78149
rect 4683 78100 4684 78140
rect 4724 78100 4725 78140
rect 4683 78091 4725 78100
rect 12267 78140 12309 78149
rect 12267 78100 12268 78140
rect 12308 78100 12309 78140
rect 12267 78091 12309 78100
rect 15051 78140 15093 78149
rect 15051 78100 15052 78140
rect 15092 78100 15093 78140
rect 15051 78091 15093 78100
rect 5155 78056 5213 78057
rect 5155 78016 5164 78056
rect 5204 78016 5213 78056
rect 5155 78015 5213 78016
rect 7083 78056 7125 78065
rect 7083 78016 7084 78056
rect 7124 78016 7125 78056
rect 7083 78007 7125 78016
rect 9867 78056 9909 78065
rect 9867 78016 9868 78056
rect 9908 78016 9909 78056
rect 9867 78007 9909 78016
rect 17067 78056 17109 78065
rect 17067 78016 17068 78056
rect 17108 78016 17109 78056
rect 17067 78007 17109 78016
rect 17259 78056 17301 78065
rect 17259 78016 17260 78056
rect 17300 78016 17301 78056
rect 17259 78007 17301 78016
rect 20139 78056 20181 78065
rect 20139 78016 20140 78056
rect 20180 78016 20181 78056
rect 20139 78007 20181 78016
rect 1152 77888 20452 77912
rect 1152 77848 4928 77888
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 5296 77848 20048 77888
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20416 77848 20452 77888
rect 1152 77824 20452 77848
rect 4971 77720 5013 77729
rect 4971 77680 4972 77720
rect 5012 77680 5013 77720
rect 4971 77671 5013 77680
rect 7851 77720 7893 77729
rect 7851 77680 7852 77720
rect 7892 77680 7893 77720
rect 7851 77671 7893 77680
rect 8323 77720 8381 77721
rect 8323 77680 8332 77720
rect 8372 77680 8381 77720
rect 8323 77679 8381 77680
rect 8619 77720 8661 77729
rect 8619 77680 8620 77720
rect 8660 77680 8661 77720
rect 14859 77720 14901 77729
rect 8619 77671 8661 77680
rect 12459 77678 12501 77687
rect 10443 77636 10485 77645
rect 10443 77596 10444 77636
rect 10484 77596 10485 77636
rect 12459 77638 12460 77678
rect 12500 77638 12501 77678
rect 14859 77680 14860 77720
rect 14900 77680 14901 77720
rect 14859 77671 14901 77680
rect 17355 77720 17397 77729
rect 17355 77680 17356 77720
rect 17396 77680 17397 77720
rect 17355 77671 17397 77680
rect 17547 77720 17589 77729
rect 17547 77680 17548 77720
rect 17588 77680 17589 77720
rect 17547 77671 17589 77680
rect 17931 77720 17973 77729
rect 17931 77680 17932 77720
rect 17972 77680 17973 77720
rect 17931 77671 17973 77680
rect 12459 77629 12501 77638
rect 10443 77587 10485 77596
rect 1219 77552 1277 77553
rect 1219 77512 1228 77552
rect 1268 77512 1277 77552
rect 1219 77511 1277 77512
rect 2467 77552 2525 77553
rect 2467 77512 2476 77552
rect 2516 77512 2525 77552
rect 2467 77511 2525 77512
rect 2947 77552 3005 77553
rect 2947 77512 2956 77552
rect 2996 77512 3005 77552
rect 2947 77511 3005 77512
rect 4195 77552 4253 77553
rect 4195 77512 4204 77552
rect 4244 77512 4253 77552
rect 4195 77511 4253 77512
rect 6123 77552 6165 77561
rect 6123 77512 6124 77552
rect 6164 77512 6165 77552
rect 6123 77503 6165 77512
rect 6219 77552 6261 77561
rect 6219 77512 6220 77552
rect 6260 77512 6261 77552
rect 6219 77503 6261 77512
rect 7171 77552 7229 77553
rect 7171 77512 7180 77552
rect 7220 77512 7229 77552
rect 7171 77511 7229 77512
rect 7659 77547 7701 77556
rect 7659 77507 7660 77547
rect 7700 77507 7701 77547
rect 7659 77498 7701 77507
rect 8043 77552 8085 77561
rect 8043 77512 8044 77552
rect 8084 77512 8085 77552
rect 8043 77503 8085 77512
rect 8139 77552 8181 77561
rect 8139 77512 8140 77552
rect 8180 77512 8181 77552
rect 8139 77503 8181 77512
rect 8235 77552 8277 77561
rect 8235 77512 8236 77552
rect 8276 77512 8277 77552
rect 8235 77503 8277 77512
rect 8515 77552 8573 77553
rect 8515 77512 8524 77552
rect 8564 77512 8573 77552
rect 8515 77511 8573 77512
rect 8995 77552 9053 77553
rect 8995 77512 9004 77552
rect 9044 77512 9053 77552
rect 8995 77511 9053 77512
rect 10243 77552 10301 77553
rect 10243 77512 10252 77552
rect 10292 77512 10301 77552
rect 10243 77511 10301 77512
rect 10731 77552 10773 77561
rect 10731 77512 10732 77552
rect 10772 77512 10773 77552
rect 10731 77503 10773 77512
rect 10827 77552 10869 77561
rect 10827 77512 10828 77552
rect 10868 77512 10869 77552
rect 10827 77503 10869 77512
rect 11307 77552 11349 77561
rect 11307 77512 11308 77552
rect 11348 77512 11349 77552
rect 11307 77503 11349 77512
rect 11779 77552 11837 77553
rect 11779 77512 11788 77552
rect 11828 77512 11837 77552
rect 13411 77552 13469 77553
rect 11779 77511 11837 77512
rect 12315 77510 12357 77519
rect 13411 77512 13420 77552
rect 13460 77512 13469 77552
rect 13411 77511 13469 77512
rect 14659 77552 14717 77553
rect 14659 77512 14668 77552
rect 14708 77512 14717 77552
rect 14659 77511 14717 77512
rect 15523 77552 15581 77553
rect 15523 77512 15532 77552
rect 15572 77512 15581 77552
rect 15523 77511 15581 77512
rect 16771 77552 16829 77553
rect 16771 77512 16780 77552
rect 16820 77512 16829 77552
rect 16771 77511 16829 77512
rect 18595 77552 18653 77553
rect 18595 77512 18604 77552
rect 18644 77512 18653 77552
rect 18595 77511 18653 77512
rect 19843 77552 19901 77553
rect 19843 77512 19852 77552
rect 19892 77512 19901 77552
rect 19843 77511 19901 77512
rect 4771 77468 4829 77469
rect 4771 77428 4780 77468
rect 4820 77428 4829 77468
rect 4771 77427 4829 77428
rect 5155 77468 5213 77469
rect 5155 77428 5164 77468
rect 5204 77428 5213 77468
rect 5155 77427 5213 77428
rect 6603 77468 6645 77477
rect 6603 77428 6604 77468
rect 6644 77428 6645 77468
rect 6603 77419 6645 77428
rect 6699 77468 6741 77477
rect 6699 77428 6700 77468
rect 6740 77428 6741 77468
rect 6699 77419 6741 77428
rect 11211 77468 11253 77477
rect 11211 77428 11212 77468
rect 11252 77428 11253 77468
rect 12315 77470 12316 77510
rect 12356 77470 12357 77510
rect 12315 77461 12357 77470
rect 15235 77468 15293 77469
rect 11211 77419 11253 77428
rect 15235 77428 15244 77468
rect 15284 77428 15293 77468
rect 15235 77427 15293 77428
rect 17155 77468 17213 77469
rect 17155 77428 17164 77468
rect 17204 77428 17213 77468
rect 17155 77427 17213 77428
rect 17731 77468 17789 77469
rect 17731 77428 17740 77468
rect 17780 77428 17789 77468
rect 17731 77427 17789 77428
rect 18115 77468 18173 77469
rect 18115 77428 18124 77468
rect 18164 77428 18173 77468
rect 18115 77427 18173 77428
rect 18315 77384 18357 77393
rect 18315 77344 18316 77384
rect 18356 77344 18357 77384
rect 18315 77335 18357 77344
rect 2667 77300 2709 77309
rect 2667 77260 2668 77300
rect 2708 77260 2709 77300
rect 2667 77251 2709 77260
rect 4395 77300 4437 77309
rect 4395 77260 4396 77300
rect 4436 77260 4437 77300
rect 4395 77251 4437 77260
rect 4587 77300 4629 77309
rect 4587 77260 4588 77300
rect 4628 77260 4629 77300
rect 4587 77251 4629 77260
rect 15051 77300 15093 77309
rect 15051 77260 15052 77300
rect 15092 77260 15093 77300
rect 15051 77251 15093 77260
rect 16971 77300 17013 77309
rect 16971 77260 16972 77300
rect 17012 77260 17013 77300
rect 16971 77251 17013 77260
rect 20043 77300 20085 77309
rect 20043 77260 20044 77300
rect 20084 77260 20085 77300
rect 20043 77251 20085 77260
rect 1152 77132 20352 77156
rect 1152 77092 3688 77132
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 4056 77092 18808 77132
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 19176 77092 20352 77132
rect 1152 77068 20352 77092
rect 2083 76880 2141 76881
rect 2083 76840 2092 76880
rect 2132 76840 2141 76880
rect 2083 76839 2141 76840
rect 4587 76880 4629 76889
rect 4587 76840 4588 76880
rect 4628 76840 4629 76880
rect 4587 76831 4629 76840
rect 12555 76880 12597 76889
rect 12555 76840 12556 76880
rect 12596 76840 12597 76880
rect 12555 76831 12597 76840
rect 17931 76880 17973 76889
rect 17931 76840 17932 76880
rect 17972 76840 17973 76880
rect 17931 76831 17973 76840
rect 1315 76796 1373 76797
rect 1315 76756 1324 76796
rect 1364 76756 1373 76796
rect 1315 76755 1373 76756
rect 1699 76796 1757 76797
rect 1699 76756 1708 76796
rect 1748 76756 1757 76796
rect 1699 76755 1757 76756
rect 3147 76796 3189 76805
rect 3147 76756 3148 76796
rect 3188 76756 3189 76796
rect 3147 76747 3189 76756
rect 4771 76796 4829 76797
rect 4771 76756 4780 76796
rect 4820 76756 4829 76796
rect 4771 76755 4829 76756
rect 8907 76796 8949 76805
rect 8907 76756 8908 76796
rect 8948 76756 8949 76796
rect 6691 76754 6749 76755
rect 4203 76726 4245 76735
rect 2091 76712 2133 76721
rect 2091 76672 2092 76712
rect 2132 76672 2133 76712
rect 2091 76663 2133 76672
rect 2187 76712 2229 76721
rect 2187 76672 2188 76712
rect 2228 76672 2229 76712
rect 2187 76663 2229 76672
rect 2379 76712 2421 76721
rect 2379 76672 2380 76712
rect 2420 76672 2421 76712
rect 2379 76663 2421 76672
rect 2667 76712 2709 76721
rect 2667 76672 2668 76712
rect 2708 76672 2709 76712
rect 2667 76663 2709 76672
rect 2763 76712 2805 76721
rect 2763 76672 2764 76712
rect 2804 76672 2805 76712
rect 2763 76663 2805 76672
rect 3243 76712 3285 76721
rect 3243 76672 3244 76712
rect 3284 76672 3285 76712
rect 3243 76663 3285 76672
rect 3715 76712 3773 76713
rect 3715 76672 3724 76712
rect 3764 76672 3773 76712
rect 4203 76686 4204 76726
rect 4244 76686 4245 76726
rect 6691 76714 6700 76754
rect 6740 76714 6749 76754
rect 8907 76747 8949 76756
rect 18115 76796 18173 76797
rect 18115 76756 18124 76796
rect 18164 76756 18173 76796
rect 18115 76755 18173 76756
rect 18891 76796 18933 76805
rect 18891 76756 18892 76796
rect 18932 76756 18933 76796
rect 18891 76747 18933 76756
rect 18987 76796 19029 76805
rect 18987 76756 18988 76796
rect 19028 76756 19029 76796
rect 18987 76747 19029 76756
rect 9963 76726 10005 76735
rect 6691 76713 6749 76714
rect 4203 76677 4245 76686
rect 5059 76712 5117 76713
rect 3715 76671 3773 76672
rect 5059 76672 5068 76712
rect 5108 76672 5117 76712
rect 5059 76671 5117 76672
rect 6307 76712 6365 76713
rect 6307 76672 6316 76712
rect 6356 76672 6365 76712
rect 6307 76671 6365 76672
rect 7939 76712 7997 76713
rect 7939 76672 7948 76712
rect 7988 76672 7997 76712
rect 7939 76671 7997 76672
rect 8427 76712 8469 76721
rect 8427 76672 8428 76712
rect 8468 76672 8469 76712
rect 8427 76663 8469 76672
rect 8523 76712 8565 76721
rect 8523 76672 8524 76712
rect 8564 76672 8565 76712
rect 8523 76663 8565 76672
rect 9003 76712 9045 76721
rect 9003 76672 9004 76712
rect 9044 76672 9045 76712
rect 9003 76663 9045 76672
rect 9475 76712 9533 76713
rect 9475 76672 9484 76712
rect 9524 76672 9533 76712
rect 9963 76686 9964 76726
rect 10004 76686 10005 76726
rect 19947 76726 19989 76735
rect 9963 76677 10005 76686
rect 11107 76712 11165 76713
rect 9475 76671 9533 76672
rect 11107 76672 11116 76712
rect 11156 76672 11165 76712
rect 11107 76671 11165 76672
rect 12355 76712 12413 76713
rect 12355 76672 12364 76712
rect 12404 76672 12413 76712
rect 12355 76671 12413 76672
rect 14563 76712 14621 76713
rect 14563 76672 14572 76712
rect 14612 76672 14621 76712
rect 14563 76671 14621 76672
rect 15811 76712 15869 76713
rect 15811 76672 15820 76712
rect 15860 76672 15869 76712
rect 15811 76671 15869 76672
rect 16195 76712 16253 76713
rect 16195 76672 16204 76712
rect 16244 76672 16253 76712
rect 16195 76671 16253 76672
rect 17443 76712 17501 76713
rect 17443 76672 17452 76712
rect 17492 76672 17501 76712
rect 17443 76671 17501 76672
rect 18411 76712 18453 76721
rect 18411 76672 18412 76712
rect 18452 76672 18453 76712
rect 18411 76663 18453 76672
rect 18507 76712 18549 76721
rect 18507 76672 18508 76712
rect 18548 76672 18549 76712
rect 18507 76663 18549 76672
rect 19459 76712 19517 76713
rect 19459 76672 19468 76712
rect 19508 76672 19517 76712
rect 19947 76686 19948 76726
rect 19988 76686 19989 76726
rect 19947 76677 19989 76686
rect 19459 76671 19517 76672
rect 4395 76628 4437 76637
rect 4395 76588 4396 76628
rect 4436 76588 4437 76628
rect 4395 76579 4437 76588
rect 8139 76628 8181 76637
rect 8139 76588 8140 76628
rect 8180 76588 8181 76628
rect 8139 76579 8181 76588
rect 1515 76544 1557 76553
rect 1515 76504 1516 76544
rect 1556 76504 1557 76544
rect 1515 76495 1557 76504
rect 1899 76544 1941 76553
rect 1899 76504 1900 76544
rect 1940 76504 1941 76544
rect 1899 76495 1941 76504
rect 6507 76544 6549 76553
rect 6507 76504 6508 76544
rect 6548 76504 6549 76544
rect 6507 76495 6549 76504
rect 10155 76544 10197 76553
rect 10155 76504 10156 76544
rect 10196 76504 10197 76544
rect 10155 76495 10197 76504
rect 16011 76544 16053 76553
rect 16011 76504 16012 76544
rect 16052 76504 16053 76544
rect 16011 76495 16053 76504
rect 17643 76544 17685 76553
rect 17643 76504 17644 76544
rect 17684 76504 17685 76544
rect 17643 76495 17685 76504
rect 20139 76544 20181 76553
rect 20139 76504 20140 76544
rect 20180 76504 20181 76544
rect 20139 76495 20181 76504
rect 1152 76376 20452 76400
rect 1152 76336 4928 76376
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 5296 76336 20048 76376
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20416 76336 20452 76376
rect 1152 76312 20452 76336
rect 1419 76208 1461 76217
rect 1419 76168 1420 76208
rect 1460 76168 1461 76208
rect 1419 76159 1461 76168
rect 6691 76208 6749 76209
rect 6691 76168 6700 76208
rect 6740 76168 6749 76208
rect 6691 76167 6749 76168
rect 7363 76208 7421 76209
rect 7363 76168 7372 76208
rect 7412 76168 7421 76208
rect 7363 76167 7421 76168
rect 19651 76208 19709 76209
rect 19651 76168 19660 76208
rect 19700 76168 19709 76208
rect 19651 76167 19709 76168
rect 20043 76208 20085 76217
rect 20043 76168 20044 76208
rect 20084 76168 20085 76208
rect 20043 76159 20085 76168
rect 6411 76124 6453 76133
rect 6411 76084 6412 76124
rect 6452 76084 6453 76124
rect 6411 76075 6453 76084
rect 15435 76124 15477 76133
rect 15435 76084 15436 76124
rect 15476 76084 15477 76124
rect 15435 76075 15477 76084
rect 1603 76040 1661 76041
rect 1603 76000 1612 76040
rect 1652 76000 1661 76040
rect 1603 75999 1661 76000
rect 2851 76040 2909 76041
rect 2851 76000 2860 76040
rect 2900 76000 2909 76040
rect 2851 75999 2909 76000
rect 3427 76040 3485 76041
rect 3427 76000 3436 76040
rect 3476 76000 3485 76040
rect 3427 75999 3485 76000
rect 4675 76040 4733 76041
rect 4675 76000 4684 76040
rect 4724 76000 4733 76040
rect 4675 75999 4733 76000
rect 4963 76040 5021 76041
rect 4963 76000 4972 76040
rect 5012 76000 5021 76040
rect 4963 75999 5021 76000
rect 6211 76040 6269 76041
rect 6211 76000 6220 76040
rect 6260 76000 6269 76040
rect 6795 76040 6837 76049
rect 6211 75999 6269 76000
rect 6637 76025 6679 76034
rect 6637 75985 6638 76025
rect 6678 75985 6679 76025
rect 6795 76000 6796 76040
rect 6836 76000 6837 76040
rect 6795 75991 6837 76000
rect 6891 76040 6933 76049
rect 6891 76000 6892 76040
rect 6932 76000 6933 76040
rect 6891 75991 6933 76000
rect 7075 76040 7133 76041
rect 7075 76000 7084 76040
rect 7124 76000 7133 76040
rect 7075 75999 7133 76000
rect 7171 76040 7229 76041
rect 7171 76000 7180 76040
rect 7220 76000 7229 76040
rect 7171 75999 7229 76000
rect 7563 76040 7605 76049
rect 7563 76000 7564 76040
rect 7604 76000 7605 76040
rect 7563 75991 7605 76000
rect 7659 76040 7701 76049
rect 7659 76000 7660 76040
rect 7700 76000 7701 76040
rect 7659 75991 7701 76000
rect 7851 76040 7893 76049
rect 7851 76000 7852 76040
rect 7892 76000 7893 76040
rect 7851 75991 7893 76000
rect 7947 76040 7989 76049
rect 7947 76000 7948 76040
rect 7988 76000 7989 76040
rect 7947 75991 7989 76000
rect 8043 76040 8085 76049
rect 8043 76000 8044 76040
rect 8084 76000 8085 76040
rect 8043 75991 8085 76000
rect 8139 76040 8181 76049
rect 8139 76000 8140 76040
rect 8180 76000 8181 76040
rect 8139 75991 8181 76000
rect 10147 76040 10205 76041
rect 10147 76000 10156 76040
rect 10196 76000 10205 76040
rect 10147 75999 10205 76000
rect 11395 76040 11453 76041
rect 11395 76000 11404 76040
rect 11444 76000 11453 76040
rect 11395 75999 11453 76000
rect 12163 76040 12221 76041
rect 12163 76000 12172 76040
rect 12212 76000 12221 76040
rect 12163 75999 12221 76000
rect 13411 76040 13469 76041
rect 13411 76000 13420 76040
rect 13460 76000 13469 76040
rect 13411 75999 13469 76000
rect 13987 76040 14045 76041
rect 13987 76000 13996 76040
rect 14036 76000 14045 76040
rect 13987 75999 14045 76000
rect 15235 76040 15293 76041
rect 15235 76000 15244 76040
rect 15284 76000 15293 76040
rect 15235 75999 15293 76000
rect 15627 76040 15669 76049
rect 15627 76000 15628 76040
rect 15668 76000 15669 76040
rect 15627 75991 15669 76000
rect 15723 76040 15765 76049
rect 15723 76000 15724 76040
rect 15764 76000 15765 76040
rect 15723 75991 15765 76000
rect 15915 76040 15957 76049
rect 15915 76000 15916 76040
rect 15956 76000 15957 76040
rect 15915 75991 15957 76000
rect 16195 76040 16253 76041
rect 16195 76000 16204 76040
rect 16244 76000 16253 76040
rect 16195 75999 16253 76000
rect 17443 76040 17501 76041
rect 17443 76000 17452 76040
rect 17492 76000 17501 76040
rect 17443 75999 17501 76000
rect 18019 76040 18077 76041
rect 18019 76000 18028 76040
rect 18068 76000 18077 76040
rect 18019 75999 18077 76000
rect 19267 76040 19325 76041
rect 19267 76000 19276 76040
rect 19316 76000 19325 76040
rect 19267 75999 19325 76000
rect 6637 75976 6679 75985
rect 1219 75956 1277 75957
rect 1219 75916 1228 75956
rect 1268 75916 1277 75956
rect 1219 75915 1277 75916
rect 20227 75956 20285 75957
rect 20227 75916 20236 75956
rect 20276 75916 20285 75956
rect 20227 75915 20285 75916
rect 15715 75872 15773 75873
rect 15715 75832 15724 75872
rect 15764 75832 15773 75872
rect 15715 75831 15773 75832
rect 3051 75788 3093 75797
rect 3051 75748 3052 75788
rect 3092 75748 3093 75788
rect 3051 75739 3093 75748
rect 3243 75788 3285 75797
rect 3243 75748 3244 75788
rect 3284 75748 3285 75788
rect 3243 75739 3285 75748
rect 11595 75788 11637 75797
rect 11595 75748 11596 75788
rect 11636 75748 11637 75788
rect 11595 75739 11637 75748
rect 13611 75788 13653 75797
rect 13611 75748 13612 75788
rect 13652 75748 13653 75788
rect 13611 75739 13653 75748
rect 17643 75788 17685 75797
rect 17643 75748 17644 75788
rect 17684 75748 17685 75788
rect 17643 75739 17685 75748
rect 17835 75788 17877 75797
rect 17835 75748 17836 75788
rect 17876 75748 17877 75788
rect 17835 75739 17877 75748
rect 1152 75620 20352 75644
rect 1152 75580 3688 75620
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 4056 75580 18808 75620
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 19176 75580 20352 75620
rect 1152 75556 20352 75580
rect 1611 75452 1653 75461
rect 1611 75412 1612 75452
rect 1652 75412 1653 75452
rect 1611 75403 1653 75412
rect 2187 75452 2229 75461
rect 2187 75412 2188 75452
rect 2228 75412 2229 75452
rect 2187 75403 2229 75412
rect 6315 75452 6357 75461
rect 6315 75412 6316 75452
rect 6356 75412 6357 75452
rect 6315 75403 6357 75412
rect 7947 75452 7989 75461
rect 7947 75412 7948 75452
rect 7988 75412 7989 75452
rect 7947 75403 7989 75412
rect 20139 75368 20181 75377
rect 20139 75328 20140 75368
rect 20180 75328 20181 75368
rect 20139 75319 20181 75328
rect 1411 75284 1469 75285
rect 1411 75244 1420 75284
rect 1460 75244 1469 75284
rect 1411 75243 1469 75244
rect 2371 75284 2429 75285
rect 2371 75244 2380 75284
rect 2420 75244 2429 75284
rect 11979 75284 12021 75293
rect 2371 75243 2429 75244
rect 4251 75242 4293 75251
rect 2667 75200 2709 75209
rect 2667 75160 2668 75200
rect 2708 75160 2709 75200
rect 2667 75151 2709 75160
rect 2763 75200 2805 75209
rect 2763 75160 2764 75200
rect 2804 75160 2805 75200
rect 2763 75151 2805 75160
rect 3147 75200 3189 75209
rect 3147 75160 3148 75200
rect 3188 75160 3189 75200
rect 3147 75151 3189 75160
rect 3243 75200 3285 75209
rect 4251 75202 4252 75242
rect 4292 75202 4293 75242
rect 11979 75244 11980 75284
rect 12020 75244 12021 75284
rect 11979 75235 12021 75244
rect 12075 75284 12117 75293
rect 12075 75244 12076 75284
rect 12116 75244 12117 75284
rect 12075 75235 12117 75244
rect 17163 75284 17205 75293
rect 17163 75244 17164 75284
rect 17204 75244 17205 75284
rect 17163 75235 17205 75244
rect 13035 75214 13077 75223
rect 3243 75160 3244 75200
rect 3284 75160 3285 75200
rect 3243 75151 3285 75160
rect 3715 75200 3773 75201
rect 3715 75160 3724 75200
rect 3764 75160 3773 75200
rect 4251 75193 4293 75202
rect 4579 75200 4637 75201
rect 3715 75159 3773 75160
rect 4579 75160 4588 75200
rect 4628 75160 4637 75200
rect 4579 75159 4637 75160
rect 5827 75200 5885 75201
rect 5827 75160 5836 75200
rect 5876 75160 5885 75200
rect 5827 75159 5885 75160
rect 6211 75200 6269 75201
rect 6211 75160 6220 75200
rect 6260 75160 6269 75200
rect 6211 75159 6269 75160
rect 6499 75200 6557 75201
rect 6499 75160 6508 75200
rect 6548 75160 6557 75200
rect 6499 75159 6557 75160
rect 7747 75200 7805 75201
rect 7747 75160 7756 75200
rect 7796 75160 7805 75200
rect 7747 75159 7805 75160
rect 8131 75200 8189 75201
rect 8131 75160 8140 75200
rect 8180 75160 8189 75200
rect 8131 75159 8189 75160
rect 9379 75200 9437 75201
rect 9379 75160 9388 75200
rect 9428 75160 9437 75200
rect 9379 75159 9437 75160
rect 9763 75200 9821 75201
rect 9763 75160 9772 75200
rect 9812 75160 9821 75200
rect 9763 75159 9821 75160
rect 11011 75200 11069 75201
rect 11011 75160 11020 75200
rect 11060 75160 11069 75200
rect 11011 75159 11069 75160
rect 11499 75200 11541 75209
rect 11499 75160 11500 75200
rect 11540 75160 11541 75200
rect 11499 75151 11541 75160
rect 11595 75200 11637 75209
rect 11595 75160 11596 75200
rect 11636 75160 11637 75200
rect 11595 75151 11637 75160
rect 12547 75200 12605 75201
rect 12547 75160 12556 75200
rect 12596 75160 12605 75200
rect 13035 75174 13036 75214
rect 13076 75174 13077 75214
rect 18219 75214 18261 75223
rect 13035 75165 13077 75174
rect 13507 75200 13565 75201
rect 12547 75159 12605 75160
rect 13507 75160 13516 75200
rect 13556 75160 13565 75200
rect 13507 75159 13565 75160
rect 14755 75200 14813 75201
rect 14755 75160 14764 75200
rect 14804 75160 14813 75200
rect 14755 75159 14813 75160
rect 15243 75200 15285 75209
rect 15243 75160 15244 75200
rect 15284 75160 15285 75200
rect 15243 75151 15285 75160
rect 15339 75200 15381 75209
rect 15339 75160 15340 75200
rect 15380 75160 15381 75200
rect 15339 75151 15381 75160
rect 15715 75200 15773 75201
rect 15715 75160 15724 75200
rect 15764 75160 15773 75200
rect 15715 75159 15773 75160
rect 15811 75200 15869 75201
rect 15811 75160 15820 75200
rect 15860 75160 15869 75200
rect 15811 75159 15869 75160
rect 16011 75200 16053 75209
rect 16011 75160 16012 75200
rect 16052 75160 16053 75200
rect 16011 75151 16053 75160
rect 16107 75200 16149 75209
rect 16107 75160 16108 75200
rect 16148 75160 16149 75200
rect 16107 75151 16149 75160
rect 16200 75200 16258 75201
rect 16200 75160 16209 75200
rect 16249 75160 16258 75200
rect 16200 75159 16258 75160
rect 16683 75200 16725 75209
rect 16683 75160 16684 75200
rect 16724 75160 16725 75200
rect 16683 75151 16725 75160
rect 16779 75200 16821 75209
rect 16779 75160 16780 75200
rect 16820 75160 16821 75200
rect 16779 75151 16821 75160
rect 17259 75200 17301 75209
rect 17259 75160 17260 75200
rect 17300 75160 17301 75200
rect 17259 75151 17301 75160
rect 17731 75200 17789 75201
rect 17731 75160 17740 75200
rect 17780 75160 17789 75200
rect 18219 75174 18220 75214
rect 18260 75174 18261 75214
rect 18219 75165 18261 75174
rect 17731 75159 17789 75160
rect 4395 75116 4437 75125
rect 4395 75076 4396 75116
rect 4436 75076 4437 75116
rect 4395 75067 4437 75076
rect 6027 75032 6069 75041
rect 6027 74992 6028 75032
rect 6068 74992 6069 75032
rect 6027 74983 6069 74992
rect 9579 75032 9621 75041
rect 9579 74992 9580 75032
rect 9620 74992 9621 75032
rect 9579 74983 9621 74992
rect 11211 75032 11253 75041
rect 11211 74992 11212 75032
rect 11252 74992 11253 75032
rect 11211 74983 11253 74992
rect 13227 75032 13269 75041
rect 13227 74992 13228 75032
rect 13268 74992 13269 75032
rect 13227 74983 13269 74992
rect 14955 75032 14997 75041
rect 14955 74992 14956 75032
rect 14996 74992 14997 75032
rect 14955 74983 14997 74992
rect 15523 75032 15581 75033
rect 15523 74992 15532 75032
rect 15572 74992 15581 75032
rect 15523 74991 15581 74992
rect 15907 75032 15965 75033
rect 15907 74992 15916 75032
rect 15956 74992 15965 75032
rect 15907 74991 15965 74992
rect 18411 75032 18453 75041
rect 18411 74992 18412 75032
rect 18452 74992 18453 75032
rect 18411 74983 18453 74992
rect 20035 75032 20093 75033
rect 20035 74992 20044 75032
rect 20084 74992 20093 75032
rect 20035 74991 20093 74992
rect 1152 74864 20452 74888
rect 1152 74824 4928 74864
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 5296 74824 20048 74864
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20416 74824 20452 74864
rect 1152 74800 20452 74824
rect 9955 74696 10013 74697
rect 9955 74656 9964 74696
rect 10004 74656 10013 74696
rect 9955 74655 10013 74656
rect 11979 74696 12021 74705
rect 11979 74656 11980 74696
rect 12020 74656 12021 74696
rect 11979 74647 12021 74656
rect 12459 74696 12501 74705
rect 12459 74656 12460 74696
rect 12500 74656 12501 74696
rect 12459 74647 12501 74656
rect 7755 74612 7797 74621
rect 7755 74572 7756 74612
rect 7796 74572 7797 74612
rect 7755 74563 7797 74572
rect 15147 74612 15189 74621
rect 15147 74572 15148 74612
rect 15188 74572 15189 74612
rect 15147 74563 15189 74572
rect 15619 74612 15677 74613
rect 15619 74572 15628 74612
rect 15668 74572 15677 74612
rect 15619 74571 15677 74572
rect 20235 74612 20277 74621
rect 20235 74572 20236 74612
rect 20276 74572 20277 74612
rect 20235 74563 20277 74572
rect 1891 74528 1949 74529
rect 1891 74488 1900 74528
rect 1940 74488 1949 74528
rect 1891 74487 1949 74488
rect 3139 74528 3197 74529
rect 3139 74488 3148 74528
rect 3188 74488 3197 74528
rect 3139 74487 3197 74488
rect 4195 74528 4253 74529
rect 4195 74488 4204 74528
rect 4244 74488 4253 74528
rect 4195 74487 4253 74488
rect 5443 74528 5501 74529
rect 5443 74488 5452 74528
rect 5492 74488 5501 74528
rect 5443 74487 5501 74488
rect 6027 74528 6069 74537
rect 6027 74488 6028 74528
rect 6068 74488 6069 74528
rect 6027 74479 6069 74488
rect 6123 74528 6165 74537
rect 6123 74488 6124 74528
rect 6164 74488 6165 74528
rect 6123 74479 6165 74488
rect 6507 74528 6549 74537
rect 6507 74488 6508 74528
rect 6548 74488 6549 74528
rect 6507 74479 6549 74488
rect 6603 74528 6645 74537
rect 6603 74488 6604 74528
rect 6644 74488 6645 74528
rect 6603 74479 6645 74488
rect 7075 74528 7133 74529
rect 7075 74488 7084 74528
rect 7124 74488 7133 74528
rect 9675 74528 9717 74537
rect 7075 74487 7133 74488
rect 7611 74518 7653 74527
rect 7611 74478 7612 74518
rect 7652 74478 7653 74518
rect 9675 74488 9676 74528
rect 9716 74488 9717 74528
rect 9675 74479 9717 74488
rect 9771 74528 9813 74537
rect 9771 74488 9772 74528
rect 9812 74488 9813 74528
rect 9771 74479 9813 74488
rect 10251 74528 10293 74537
rect 10251 74488 10252 74528
rect 10292 74488 10293 74528
rect 10251 74479 10293 74488
rect 10347 74528 10389 74537
rect 10347 74488 10348 74528
rect 10388 74488 10389 74528
rect 10347 74479 10389 74488
rect 10827 74528 10869 74537
rect 10827 74488 10828 74528
rect 10868 74488 10869 74528
rect 10827 74479 10869 74488
rect 11299 74528 11357 74529
rect 11299 74488 11308 74528
rect 11348 74488 11357 74528
rect 11299 74487 11357 74488
rect 11787 74523 11829 74532
rect 11787 74483 11788 74523
rect 11828 74483 11829 74523
rect 7611 74469 7653 74478
rect 11787 74474 11829 74483
rect 12843 74528 12885 74537
rect 12843 74488 12844 74528
rect 12884 74488 12885 74528
rect 12843 74479 12885 74488
rect 12939 74528 12981 74537
rect 12939 74488 12940 74528
rect 12980 74488 12981 74528
rect 12939 74479 12981 74488
rect 13035 74528 13077 74537
rect 13035 74488 13036 74528
rect 13076 74488 13077 74528
rect 13035 74479 13077 74488
rect 13131 74528 13173 74537
rect 13131 74488 13132 74528
rect 13172 74488 13173 74528
rect 13131 74479 13173 74488
rect 13419 74528 13461 74537
rect 13419 74488 13420 74528
rect 13460 74488 13461 74528
rect 13419 74479 13461 74488
rect 13515 74528 13557 74537
rect 13515 74488 13516 74528
rect 13556 74488 13557 74528
rect 13515 74479 13557 74488
rect 13899 74528 13941 74537
rect 13899 74488 13900 74528
rect 13940 74488 13941 74528
rect 13899 74479 13941 74488
rect 13995 74528 14037 74537
rect 13995 74488 13996 74528
rect 14036 74488 14037 74528
rect 13995 74479 14037 74488
rect 14467 74528 14525 74529
rect 14467 74488 14476 74528
rect 14516 74488 14525 74528
rect 14467 74487 14525 74488
rect 14955 74523 14997 74532
rect 14955 74483 14956 74523
rect 14996 74483 14997 74523
rect 16483 74528 16541 74529
rect 16483 74488 16492 74528
rect 16532 74488 16541 74528
rect 16483 74487 16541 74488
rect 16771 74528 16829 74529
rect 16771 74488 16780 74528
rect 16820 74488 16829 74528
rect 16771 74487 16829 74488
rect 18019 74528 18077 74529
rect 18019 74488 18028 74528
rect 18068 74488 18077 74528
rect 18019 74487 18077 74488
rect 18507 74528 18549 74537
rect 18507 74488 18508 74528
rect 18548 74488 18549 74528
rect 14955 74474 14997 74483
rect 18507 74479 18549 74488
rect 18603 74528 18645 74537
rect 18603 74488 18604 74528
rect 18644 74488 18645 74528
rect 18603 74479 18645 74488
rect 18987 74528 19029 74537
rect 18987 74488 18988 74528
rect 19028 74488 19029 74528
rect 18987 74479 19029 74488
rect 19555 74528 19613 74529
rect 19555 74488 19564 74528
rect 19604 74488 19613 74528
rect 19555 74487 19613 74488
rect 20043 74523 20085 74532
rect 20043 74483 20044 74523
rect 20084 74483 20085 74523
rect 20043 74474 20085 74483
rect 10731 74444 10773 74453
rect 10731 74404 10732 74444
rect 10772 74404 10773 74444
rect 10731 74395 10773 74404
rect 12643 74444 12701 74445
rect 12643 74404 12652 74444
rect 12692 74404 12701 74444
rect 12643 74403 12701 74404
rect 19083 74444 19125 74453
rect 19083 74404 19084 74444
rect 19124 74404 19125 74444
rect 19083 74395 19125 74404
rect 3339 74276 3381 74285
rect 3339 74236 3340 74276
rect 3380 74236 3381 74276
rect 3339 74227 3381 74236
rect 4011 74276 4053 74285
rect 4011 74236 4012 74276
rect 4052 74236 4053 74276
rect 4011 74227 4053 74236
rect 18219 74276 18261 74285
rect 18219 74236 18220 74276
rect 18260 74236 18261 74276
rect 18219 74227 18261 74236
rect 1152 74108 20352 74132
rect 1152 74068 3688 74108
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 4056 74068 18808 74108
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 19176 74068 20352 74108
rect 1152 74044 20352 74068
rect 10059 73940 10101 73949
rect 10059 73900 10060 73940
rect 10100 73900 10101 73940
rect 10059 73891 10101 73900
rect 13899 73940 13941 73949
rect 13899 73900 13900 73940
rect 13940 73900 13941 73940
rect 13899 73891 13941 73900
rect 16107 73940 16149 73949
rect 16107 73900 16108 73940
rect 16148 73900 16149 73940
rect 16107 73891 16149 73900
rect 7075 73856 7133 73857
rect 7075 73816 7084 73856
rect 7124 73816 7133 73856
rect 7075 73815 7133 73816
rect 2091 73772 2133 73781
rect 2091 73732 2092 73772
rect 2132 73732 2133 73772
rect 2091 73723 2133 73732
rect 2187 73772 2229 73781
rect 2187 73732 2188 73772
rect 2228 73732 2229 73772
rect 2187 73723 2229 73732
rect 10435 73717 10493 73718
rect 3147 73702 3189 73711
rect 1611 73688 1653 73697
rect 1611 73648 1612 73688
rect 1652 73648 1653 73688
rect 1611 73639 1653 73648
rect 1707 73688 1749 73697
rect 1707 73648 1708 73688
rect 1748 73648 1749 73688
rect 1707 73639 1749 73648
rect 2659 73688 2717 73689
rect 2659 73648 2668 73688
rect 2708 73648 2717 73688
rect 3147 73662 3148 73702
rect 3188 73662 3189 73702
rect 10155 73703 10197 73712
rect 3147 73653 3189 73662
rect 3523 73688 3581 73689
rect 2659 73647 2717 73648
rect 3523 73648 3532 73688
rect 3572 73648 3581 73688
rect 3523 73647 3581 73648
rect 4771 73688 4829 73689
rect 4771 73648 4780 73688
rect 4820 73648 4829 73688
rect 4771 73647 4829 73648
rect 5347 73688 5405 73689
rect 5347 73648 5356 73688
rect 5396 73648 5405 73688
rect 5347 73647 5405 73648
rect 6595 73688 6653 73689
rect 6595 73648 6604 73688
rect 6644 73648 6653 73688
rect 6595 73647 6653 73648
rect 6795 73688 6837 73697
rect 6795 73648 6796 73688
rect 6836 73648 6837 73688
rect 6795 73639 6837 73648
rect 6987 73688 7029 73697
rect 6987 73648 6988 73688
rect 7028 73648 7029 73688
rect 6987 73639 7029 73648
rect 7083 73688 7125 73697
rect 7083 73648 7084 73688
rect 7124 73648 7125 73688
rect 7083 73639 7125 73648
rect 7267 73688 7325 73689
rect 7267 73648 7276 73688
rect 7316 73648 7325 73688
rect 7267 73647 7325 73648
rect 7363 73688 7421 73689
rect 7363 73648 7372 73688
rect 7412 73648 7421 73688
rect 7363 73647 7421 73648
rect 7563 73688 7605 73697
rect 7563 73648 7564 73688
rect 7604 73648 7605 73688
rect 7563 73639 7605 73648
rect 7659 73688 7701 73697
rect 7659 73648 7660 73688
rect 7700 73648 7701 73688
rect 7659 73639 7701 73648
rect 7806 73688 7864 73689
rect 7806 73648 7815 73688
rect 7855 73648 7864 73688
rect 7806 73647 7864 73648
rect 8043 73688 8085 73697
rect 8043 73648 8044 73688
rect 8084 73648 8085 73688
rect 8043 73639 8085 73648
rect 8131 73688 8189 73689
rect 8131 73648 8140 73688
rect 8180 73648 8189 73688
rect 8131 73647 8189 73648
rect 8419 73688 8477 73689
rect 8419 73648 8428 73688
rect 8468 73648 8477 73688
rect 8419 73647 8477 73648
rect 9667 73688 9725 73689
rect 9667 73648 9676 73688
rect 9716 73648 9725 73688
rect 9667 73647 9725 73648
rect 10051 73688 10109 73689
rect 10051 73648 10060 73688
rect 10100 73648 10109 73688
rect 10155 73663 10156 73703
rect 10196 73663 10197 73703
rect 10155 73654 10197 73663
rect 10347 73688 10389 73697
rect 10051 73647 10109 73648
rect 10347 73648 10348 73688
rect 10388 73648 10389 73688
rect 10435 73677 10444 73717
rect 10484 73677 10493 73717
rect 10435 73676 10493 73677
rect 10536 73688 10594 73689
rect 10347 73639 10389 73648
rect 10536 73648 10545 73688
rect 10585 73648 10594 73688
rect 10536 73647 10594 73648
rect 10819 73688 10877 73689
rect 10819 73648 10828 73688
rect 10868 73648 10877 73688
rect 10819 73647 10877 73648
rect 12067 73688 12125 73689
rect 12067 73648 12076 73688
rect 12116 73648 12125 73688
rect 12067 73647 12125 73648
rect 12451 73688 12509 73689
rect 12451 73648 12460 73688
rect 12500 73648 12509 73688
rect 12451 73647 12509 73648
rect 13699 73688 13757 73689
rect 13699 73648 13708 73688
rect 13748 73648 13757 73688
rect 13699 73647 13757 73648
rect 14275 73688 14333 73689
rect 14275 73648 14284 73688
rect 14324 73648 14333 73688
rect 14275 73647 14333 73648
rect 15523 73688 15581 73689
rect 15523 73648 15532 73688
rect 15572 73648 15581 73688
rect 15523 73647 15581 73648
rect 16003 73688 16061 73689
rect 16003 73648 16012 73688
rect 16052 73648 16061 73688
rect 16003 73647 16061 73648
rect 16867 73688 16925 73689
rect 16867 73648 16876 73688
rect 16916 73648 16925 73688
rect 16867 73647 16925 73648
rect 18115 73688 18173 73689
rect 18115 73648 18124 73688
rect 18164 73648 18173 73688
rect 18115 73647 18173 73648
rect 18499 73688 18557 73689
rect 18499 73648 18508 73688
rect 18548 73648 18557 73688
rect 18499 73647 18557 73648
rect 19747 73688 19805 73689
rect 19747 73648 19756 73688
rect 19796 73648 19805 73688
rect 19747 73647 19805 73648
rect 9867 73604 9909 73613
rect 9867 73564 9868 73604
rect 9908 73564 9909 73604
rect 9867 73555 9909 73564
rect 4971 73520 5013 73529
rect 3339 73478 3381 73487
rect 3339 73438 3340 73478
rect 3380 73438 3381 73478
rect 4971 73480 4972 73520
rect 5012 73480 5013 73520
rect 4971 73471 5013 73480
rect 5163 73520 5205 73529
rect 5163 73480 5164 73520
rect 5204 73480 5205 73520
rect 5163 73471 5205 73480
rect 7651 73520 7709 73521
rect 7651 73480 7660 73520
rect 7700 73480 7709 73520
rect 7651 73479 7709 73480
rect 12267 73520 12309 73529
rect 12267 73480 12268 73520
rect 12308 73480 12309 73520
rect 12267 73471 12309 73480
rect 15723 73520 15765 73529
rect 15723 73480 15724 73520
rect 15764 73480 15765 73520
rect 15723 73471 15765 73480
rect 18315 73520 18357 73529
rect 18315 73480 18316 73520
rect 18356 73480 18357 73520
rect 18315 73471 18357 73480
rect 19947 73520 19989 73529
rect 19947 73480 19948 73520
rect 19988 73480 19989 73520
rect 19947 73471 19989 73480
rect 3339 73429 3381 73438
rect 1152 73352 20452 73376
rect 1152 73312 4928 73352
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 5296 73312 20048 73352
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20416 73312 20452 73352
rect 1152 73288 20452 73312
rect 7467 73184 7509 73193
rect 7467 73144 7468 73184
rect 7508 73144 7509 73184
rect 7467 73135 7509 73144
rect 7939 73184 7997 73185
rect 7939 73144 7948 73184
rect 7988 73144 7997 73184
rect 7939 73143 7997 73144
rect 10059 73184 10101 73193
rect 10059 73144 10060 73184
rect 10100 73144 10101 73184
rect 10059 73135 10101 73144
rect 10443 73184 10485 73193
rect 10443 73144 10444 73184
rect 10484 73144 10485 73184
rect 10443 73135 10485 73144
rect 3627 73100 3669 73109
rect 3627 73060 3628 73100
rect 3668 73060 3669 73100
rect 3627 73051 3669 73060
rect 9771 73100 9813 73109
rect 9771 73060 9772 73100
rect 9812 73060 9813 73100
rect 9771 73051 9813 73060
rect 13323 73100 13365 73109
rect 13323 73060 13324 73100
rect 13364 73060 13365 73100
rect 13323 73051 13365 73060
rect 17451 73100 17493 73109
rect 17451 73060 17452 73100
rect 17492 73060 17493 73100
rect 17451 73051 17493 73060
rect 1219 73016 1277 73017
rect 1219 72976 1228 73016
rect 1268 72976 1277 73016
rect 1219 72975 1277 72976
rect 2467 73016 2525 73017
rect 2467 72976 2476 73016
rect 2516 72976 2525 73016
rect 2467 72975 2525 72976
rect 3819 73011 3861 73020
rect 3819 72971 3820 73011
rect 3860 72971 3861 73011
rect 4291 73016 4349 73017
rect 4291 72976 4300 73016
rect 4340 72976 4349 73016
rect 4291 72975 4349 72976
rect 5259 73016 5301 73025
rect 5259 72976 5260 73016
rect 5300 72976 5301 73016
rect 3819 72962 3861 72971
rect 5259 72967 5301 72976
rect 5355 73016 5397 73025
rect 5355 72976 5356 73016
rect 5396 72976 5397 73016
rect 5355 72967 5397 72976
rect 6019 73016 6077 73017
rect 6019 72976 6028 73016
rect 6068 72976 6077 73016
rect 6019 72975 6077 72976
rect 7267 73016 7325 73017
rect 7267 72976 7276 73016
rect 7316 72976 7325 73016
rect 7267 72975 7325 72976
rect 7659 73016 7701 73025
rect 7659 72976 7660 73016
rect 7700 72976 7701 73016
rect 7659 72967 7701 72976
rect 7755 73016 7797 73025
rect 7755 72976 7756 73016
rect 7796 72976 7797 73016
rect 7755 72967 7797 72976
rect 8323 73016 8381 73017
rect 8323 72976 8332 73016
rect 8372 72976 8381 73016
rect 8323 72975 8381 72976
rect 9571 73016 9629 73017
rect 9571 72976 9580 73016
rect 9620 72976 9629 73016
rect 9571 72975 9629 72976
rect 9963 73016 10005 73025
rect 9963 72976 9964 73016
rect 10004 72976 10005 73016
rect 9963 72967 10005 72976
rect 10155 73016 10197 73025
rect 10155 72976 10156 73016
rect 10196 72976 10197 73016
rect 10155 72967 10197 72976
rect 10251 73016 10293 73025
rect 10251 72976 10252 73016
rect 10292 72976 10293 73016
rect 10251 72967 10293 72976
rect 10531 73016 10589 73017
rect 10531 72976 10540 73016
rect 10580 72976 10589 73016
rect 10531 72975 10589 72976
rect 11683 73016 11741 73017
rect 11683 72976 11692 73016
rect 11732 72976 11741 73016
rect 11683 72975 11741 72976
rect 12931 73016 12989 73017
rect 12931 72976 12940 73016
rect 12980 72976 12989 73016
rect 12931 72975 12989 72976
rect 13419 73016 13461 73025
rect 13419 72976 13420 73016
rect 13460 72976 13461 73016
rect 13419 72967 13461 72976
rect 13515 73016 13557 73025
rect 13515 72976 13516 73016
rect 13556 72976 13557 73016
rect 13515 72967 13557 72976
rect 13611 73016 13653 73025
rect 13611 72976 13612 73016
rect 13652 72976 13653 73016
rect 13611 72967 13653 72976
rect 13987 73016 14045 73017
rect 13987 72976 13996 73016
rect 14036 72976 14045 73016
rect 13987 72975 14045 72976
rect 15235 73016 15293 73017
rect 15235 72976 15244 73016
rect 15284 72976 15293 73016
rect 15819 73016 15861 73025
rect 15235 72975 15293 72976
rect 15723 72997 15765 73006
rect 15723 72957 15724 72997
rect 15764 72957 15765 72997
rect 15819 72976 15820 73016
rect 15860 72976 15861 73016
rect 15819 72967 15861 72976
rect 16771 73016 16829 73017
rect 16771 72976 16780 73016
rect 16820 72976 16829 73016
rect 16771 72975 16829 72976
rect 17259 73011 17301 73020
rect 17259 72971 17260 73011
rect 17300 72971 17301 73011
rect 18403 73016 18461 73017
rect 18403 72976 18412 73016
rect 18452 72976 18461 73016
rect 18403 72975 18461 72976
rect 19651 73016 19709 73017
rect 19651 72976 19660 73016
rect 19700 72976 19709 73016
rect 19651 72975 19709 72976
rect 17259 72962 17301 72971
rect 15723 72948 15765 72957
rect 4779 72932 4821 72941
rect 4779 72892 4780 72932
rect 4820 72892 4821 72932
rect 4779 72883 4821 72892
rect 4875 72932 4917 72941
rect 4875 72892 4876 72932
rect 4916 72892 4917 72932
rect 4875 72883 4917 72892
rect 16203 72932 16245 72941
rect 16203 72892 16204 72932
rect 16244 72892 16245 72932
rect 16203 72883 16245 72892
rect 16299 72932 16341 72941
rect 16299 72892 16300 72932
rect 16340 72892 16341 72932
rect 16299 72883 16341 72892
rect 15435 72848 15477 72857
rect 15435 72808 15436 72848
rect 15476 72808 15477 72848
rect 15435 72799 15477 72808
rect 2667 72764 2709 72773
rect 2667 72724 2668 72764
rect 2708 72724 2709 72764
rect 2667 72715 2709 72724
rect 13131 72764 13173 72773
rect 13131 72724 13132 72764
rect 13172 72724 13173 72764
rect 13131 72715 13173 72724
rect 19851 72764 19893 72773
rect 19851 72724 19852 72764
rect 19892 72724 19893 72764
rect 19851 72715 19893 72724
rect 1152 72596 20352 72620
rect 1152 72556 3688 72596
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 4056 72556 18808 72596
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 19176 72556 20352 72596
rect 1152 72532 20352 72556
rect 7371 72428 7413 72437
rect 7371 72388 7372 72428
rect 7412 72388 7413 72428
rect 7371 72379 7413 72388
rect 13323 72428 13365 72437
rect 13323 72388 13324 72428
rect 13364 72388 13365 72428
rect 13323 72379 13365 72388
rect 13611 72260 13653 72269
rect 13611 72220 13612 72260
rect 13652 72220 13653 72260
rect 13611 72211 13653 72220
rect 16299 72260 16341 72269
rect 16299 72220 16300 72260
rect 16340 72220 16341 72260
rect 16299 72211 16341 72220
rect 19083 72260 19125 72269
rect 19083 72220 19084 72260
rect 19124 72220 19125 72260
rect 19083 72211 19125 72220
rect 17259 72190 17301 72199
rect 1699 72176 1757 72177
rect 1699 72136 1708 72176
rect 1748 72136 1757 72176
rect 1699 72135 1757 72136
rect 2947 72176 3005 72177
rect 2947 72136 2956 72176
rect 2996 72136 3005 72176
rect 2947 72135 3005 72136
rect 4291 72176 4349 72177
rect 4291 72136 4300 72176
rect 4340 72136 4349 72176
rect 4291 72135 4349 72136
rect 5539 72176 5597 72177
rect 5539 72136 5548 72176
rect 5588 72136 5597 72176
rect 5539 72135 5597 72136
rect 5923 72176 5981 72177
rect 5923 72136 5932 72176
rect 5972 72136 5981 72176
rect 5923 72135 5981 72136
rect 7171 72176 7229 72177
rect 7171 72136 7180 72176
rect 7220 72136 7229 72176
rect 7171 72135 7229 72136
rect 7747 72176 7805 72177
rect 7747 72136 7756 72176
rect 7796 72136 7805 72176
rect 7747 72135 7805 72136
rect 8995 72176 9053 72177
rect 8995 72136 9004 72176
rect 9044 72136 9053 72176
rect 8995 72135 9053 72136
rect 9379 72176 9437 72177
rect 9379 72136 9388 72176
rect 9428 72136 9437 72176
rect 9379 72135 9437 72136
rect 10627 72176 10685 72177
rect 10627 72136 10636 72176
rect 10676 72136 10685 72176
rect 10627 72135 10685 72136
rect 11211 72176 11253 72185
rect 11211 72136 11212 72176
rect 11252 72136 11253 72176
rect 11211 72127 11253 72136
rect 11307 72176 11349 72185
rect 11307 72136 11308 72176
rect 11348 72136 11349 72176
rect 11307 72127 11349 72136
rect 11683 72176 11741 72177
rect 11683 72136 11692 72176
rect 11732 72136 11741 72176
rect 11683 72135 11741 72136
rect 11875 72176 11933 72177
rect 11875 72136 11884 72176
rect 11924 72136 11933 72176
rect 11875 72135 11933 72136
rect 13123 72176 13181 72177
rect 13123 72136 13132 72176
rect 13172 72136 13181 72176
rect 13123 72135 13181 72136
rect 13515 72176 13557 72185
rect 13515 72136 13516 72176
rect 13556 72136 13557 72176
rect 13515 72127 13557 72136
rect 13803 72176 13845 72185
rect 13803 72136 13804 72176
rect 13844 72136 13845 72176
rect 13803 72127 13845 72136
rect 13987 72176 14045 72177
rect 13987 72136 13996 72176
rect 14036 72136 14045 72176
rect 13987 72135 14045 72136
rect 15235 72176 15293 72177
rect 15235 72136 15244 72176
rect 15284 72136 15293 72176
rect 15235 72135 15293 72136
rect 15723 72176 15765 72185
rect 15723 72136 15724 72176
rect 15764 72136 15765 72176
rect 15723 72127 15765 72136
rect 15819 72176 15861 72185
rect 15819 72136 15820 72176
rect 15860 72136 15861 72176
rect 15819 72127 15861 72136
rect 16203 72176 16245 72185
rect 16203 72136 16204 72176
rect 16244 72136 16245 72176
rect 16203 72127 16245 72136
rect 16771 72176 16829 72177
rect 16771 72136 16780 72176
rect 16820 72136 16829 72176
rect 17259 72150 17260 72190
rect 17300 72150 17301 72190
rect 20043 72190 20085 72199
rect 17259 72141 17301 72150
rect 18507 72176 18549 72185
rect 16771 72135 16829 72136
rect 18507 72136 18508 72176
rect 18548 72136 18549 72176
rect 18507 72127 18549 72136
rect 18603 72176 18645 72185
rect 18603 72136 18604 72176
rect 18644 72136 18645 72176
rect 18603 72127 18645 72136
rect 18987 72176 19029 72185
rect 18987 72136 18988 72176
rect 19028 72136 19029 72176
rect 18987 72127 19029 72136
rect 19555 72176 19613 72177
rect 19555 72136 19564 72176
rect 19604 72136 19613 72176
rect 20043 72150 20044 72190
rect 20084 72150 20085 72190
rect 20043 72141 20085 72150
rect 19555 72135 19613 72136
rect 3147 72008 3189 72017
rect 3147 71968 3148 72008
rect 3188 71968 3189 72008
rect 3147 71959 3189 71968
rect 5739 72008 5781 72017
rect 5739 71968 5740 72008
rect 5780 71968 5781 72008
rect 5739 71959 5781 71968
rect 9195 72008 9237 72017
rect 9195 71968 9196 72008
rect 9236 71968 9237 72008
rect 9195 71959 9237 71968
rect 10827 72008 10869 72017
rect 10827 71968 10828 72008
rect 10868 71968 10869 72008
rect 10827 71959 10869 71968
rect 11011 72008 11069 72009
rect 11011 71968 11020 72008
rect 11060 71968 11069 72008
rect 11011 71967 11069 71968
rect 11595 72008 11637 72017
rect 11595 71968 11596 72008
rect 11636 71968 11637 72008
rect 11595 71959 11637 71968
rect 13323 72008 13365 72017
rect 13323 71968 13324 72008
rect 13364 71968 13365 72008
rect 13323 71959 13365 71968
rect 15435 72008 15477 72017
rect 15435 71968 15436 72008
rect 15476 71968 15477 72008
rect 15435 71959 15477 71968
rect 17451 72008 17493 72017
rect 17451 71968 17452 72008
rect 17492 71968 17493 72008
rect 17451 71959 17493 71968
rect 20235 72008 20277 72017
rect 20235 71968 20236 72008
rect 20276 71968 20277 72008
rect 20235 71959 20277 71968
rect 1152 71840 20452 71864
rect 1152 71800 4928 71840
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 5296 71800 20048 71840
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20416 71800 20452 71840
rect 1152 71776 20452 71800
rect 3243 71672 3285 71681
rect 3243 71632 3244 71672
rect 3284 71632 3285 71672
rect 3243 71623 3285 71632
rect 7659 71672 7701 71681
rect 7659 71632 7660 71672
rect 7700 71632 7701 71672
rect 7659 71623 7701 71632
rect 6027 71588 6069 71597
rect 6027 71548 6028 71588
rect 6068 71548 6069 71588
rect 6027 71539 6069 71548
rect 9675 71588 9717 71597
rect 9675 71548 9676 71588
rect 9716 71548 9717 71588
rect 9675 71539 9717 71548
rect 13995 71588 14037 71597
rect 13995 71548 13996 71588
rect 14036 71548 14037 71588
rect 13995 71539 14037 71548
rect 1515 71504 1557 71513
rect 1515 71464 1516 71504
rect 1556 71464 1557 71504
rect 1515 71455 1557 71464
rect 1611 71504 1653 71513
rect 1611 71464 1612 71504
rect 1652 71464 1653 71504
rect 1611 71455 1653 71464
rect 2091 71504 2133 71513
rect 2091 71464 2092 71504
rect 2132 71464 2133 71504
rect 2091 71455 2133 71464
rect 2563 71504 2621 71505
rect 2563 71464 2572 71504
rect 2612 71464 2621 71504
rect 2563 71463 2621 71464
rect 3051 71499 3093 71508
rect 3051 71459 3052 71499
rect 3092 71459 3093 71499
rect 3051 71450 3093 71459
rect 4299 71504 4341 71513
rect 4299 71464 4300 71504
rect 4340 71464 4341 71504
rect 4299 71455 4341 71464
rect 4395 71504 4437 71513
rect 4395 71464 4396 71504
rect 4436 71464 4437 71504
rect 4395 71455 4437 71464
rect 5347 71504 5405 71505
rect 5347 71464 5356 71504
rect 5396 71464 5405 71504
rect 5347 71463 5405 71464
rect 5835 71499 5877 71508
rect 5835 71459 5836 71499
rect 5876 71459 5877 71499
rect 6211 71504 6269 71505
rect 6211 71464 6220 71504
rect 6260 71464 6269 71504
rect 6211 71463 6269 71464
rect 7459 71504 7517 71505
rect 7459 71464 7468 71504
rect 7508 71464 7517 71504
rect 7459 71463 7517 71464
rect 7947 71504 7989 71513
rect 7947 71464 7948 71504
rect 7988 71464 7989 71504
rect 5835 71450 5877 71459
rect 7947 71455 7989 71464
rect 8043 71504 8085 71513
rect 8043 71464 8044 71504
rect 8084 71464 8085 71504
rect 8043 71455 8085 71464
rect 8523 71504 8565 71513
rect 8523 71464 8524 71504
rect 8564 71464 8565 71504
rect 8523 71455 8565 71464
rect 8995 71504 9053 71505
rect 8995 71464 9004 71504
rect 9044 71464 9053 71504
rect 8995 71463 9053 71464
rect 9483 71499 9525 71508
rect 9483 71459 9484 71499
rect 9524 71459 9525 71499
rect 9859 71504 9917 71505
rect 9859 71464 9868 71504
rect 9908 71464 9917 71504
rect 9859 71463 9917 71464
rect 11107 71504 11165 71505
rect 11107 71464 11116 71504
rect 11156 71464 11165 71504
rect 11107 71463 11165 71464
rect 11499 71504 11541 71513
rect 11499 71464 11500 71504
rect 11540 71464 11541 71504
rect 9483 71450 9525 71459
rect 11499 71455 11541 71464
rect 11595 71504 11637 71513
rect 11595 71464 11596 71504
rect 11636 71464 11637 71504
rect 11595 71455 11637 71464
rect 11787 71504 11829 71513
rect 11787 71464 11788 71504
rect 11828 71464 11829 71504
rect 11787 71455 11829 71464
rect 12267 71504 12309 71513
rect 12267 71464 12268 71504
rect 12308 71464 12309 71504
rect 12267 71455 12309 71464
rect 12363 71504 12405 71513
rect 12363 71464 12364 71504
rect 12404 71464 12405 71504
rect 12843 71504 12885 71513
rect 12363 71455 12405 71464
rect 12747 71462 12789 71471
rect 1995 71420 2037 71429
rect 1995 71380 1996 71420
rect 2036 71380 2037 71420
rect 1995 71371 2037 71380
rect 4779 71420 4821 71429
rect 4779 71380 4780 71420
rect 4820 71380 4821 71420
rect 4779 71371 4821 71380
rect 4875 71420 4917 71429
rect 4875 71380 4876 71420
rect 4916 71380 4917 71420
rect 4875 71371 4917 71380
rect 8427 71420 8469 71429
rect 8427 71380 8428 71420
rect 8468 71380 8469 71420
rect 12747 71422 12748 71462
rect 12788 71422 12789 71462
rect 12843 71464 12844 71504
rect 12884 71464 12885 71504
rect 12843 71455 12885 71464
rect 13315 71504 13373 71505
rect 13315 71464 13324 71504
rect 13364 71464 13373 71504
rect 13315 71463 13373 71464
rect 13803 71499 13845 71508
rect 13803 71459 13804 71499
rect 13844 71459 13845 71499
rect 13803 71450 13845 71459
rect 14187 71504 14229 71513
rect 14187 71464 14188 71504
rect 14228 71464 14229 71504
rect 14187 71455 14229 71464
rect 14379 71504 14421 71513
rect 14379 71464 14380 71504
rect 14420 71464 14421 71504
rect 14379 71455 14421 71464
rect 14563 71504 14621 71505
rect 14563 71464 14572 71504
rect 14612 71464 14621 71504
rect 14563 71463 14621 71464
rect 15811 71504 15869 71505
rect 15811 71464 15820 71504
rect 15860 71464 15869 71504
rect 15811 71463 15869 71464
rect 16195 71504 16253 71505
rect 16195 71464 16204 71504
rect 16244 71464 16253 71504
rect 16195 71463 16253 71464
rect 17443 71504 17501 71505
rect 17443 71464 17452 71504
rect 17492 71464 17501 71504
rect 17443 71463 17501 71464
rect 18307 71504 18365 71505
rect 18307 71464 18316 71504
rect 18356 71464 18365 71504
rect 18307 71463 18365 71464
rect 19555 71504 19613 71505
rect 19555 71464 19564 71504
rect 19604 71464 19613 71504
rect 19555 71463 19613 71464
rect 12747 71413 12789 71422
rect 8427 71371 8469 71380
rect 11491 71336 11549 71337
rect 11491 71296 11500 71336
rect 11540 71296 11549 71336
rect 11491 71295 11549 71296
rect 11307 71252 11349 71261
rect 11307 71212 11308 71252
rect 11348 71212 11349 71252
rect 11307 71203 11349 71212
rect 14379 71252 14421 71261
rect 14379 71212 14380 71252
rect 14420 71212 14421 71252
rect 14379 71203 14421 71212
rect 16011 71252 16053 71261
rect 16011 71212 16012 71252
rect 16052 71212 16053 71252
rect 16011 71203 16053 71212
rect 17643 71252 17685 71261
rect 17643 71212 17644 71252
rect 17684 71212 17685 71252
rect 17643 71203 17685 71212
rect 19755 71252 19797 71261
rect 19755 71212 19756 71252
rect 19796 71212 19797 71252
rect 19755 71203 19797 71212
rect 1152 71084 20352 71108
rect 1152 71044 3688 71084
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 4056 71044 18808 71084
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 19176 71044 20352 71084
rect 1152 71020 20352 71044
rect 10923 70916 10965 70925
rect 10923 70876 10924 70916
rect 10964 70876 10965 70916
rect 10923 70867 10965 70876
rect 12267 70916 12309 70925
rect 12267 70876 12268 70916
rect 12308 70876 12309 70916
rect 12267 70867 12309 70876
rect 12451 70832 12509 70833
rect 12451 70792 12460 70832
rect 12500 70792 12509 70832
rect 12451 70791 12509 70792
rect 4771 70706 4829 70707
rect 4771 70666 4780 70706
rect 4820 70666 4829 70706
rect 12739 70706 12797 70707
rect 9915 70673 9957 70682
rect 4771 70665 4829 70666
rect 1219 70664 1277 70665
rect 1219 70624 1228 70664
rect 1268 70624 1277 70664
rect 1219 70623 1277 70624
rect 2467 70664 2525 70665
rect 2467 70624 2476 70664
rect 2516 70624 2525 70664
rect 2467 70623 2525 70624
rect 3139 70664 3197 70665
rect 3139 70624 3148 70664
rect 3188 70624 3197 70664
rect 3139 70623 3197 70624
rect 4387 70664 4445 70665
rect 4387 70624 4396 70664
rect 4436 70624 4445 70664
rect 4387 70623 4445 70624
rect 6019 70664 6077 70665
rect 6019 70624 6028 70664
rect 6068 70624 6077 70664
rect 6019 70623 6077 70624
rect 6595 70664 6653 70665
rect 6595 70624 6604 70664
rect 6644 70624 6653 70664
rect 6595 70623 6653 70624
rect 7843 70664 7901 70665
rect 7843 70624 7852 70664
rect 7892 70624 7901 70664
rect 7843 70623 7901 70624
rect 8331 70664 8373 70673
rect 8331 70624 8332 70664
rect 8372 70624 8373 70664
rect 8331 70615 8373 70624
rect 8427 70664 8469 70673
rect 8427 70624 8428 70664
rect 8468 70624 8469 70664
rect 8427 70615 8469 70624
rect 8811 70664 8853 70673
rect 8811 70624 8812 70664
rect 8852 70624 8853 70664
rect 8811 70615 8853 70624
rect 8907 70664 8949 70673
rect 8907 70624 8908 70664
rect 8948 70624 8949 70664
rect 8907 70615 8949 70624
rect 9379 70664 9437 70665
rect 9379 70624 9388 70664
rect 9428 70624 9437 70664
rect 9915 70633 9916 70673
rect 9956 70633 9957 70673
rect 9915 70624 9957 70633
rect 10430 70664 10488 70665
rect 10430 70624 10439 70664
rect 10479 70624 10488 70664
rect 9379 70623 9437 70624
rect 10430 70623 10488 70624
rect 10539 70664 10581 70673
rect 10539 70624 10540 70664
rect 10580 70624 10581 70664
rect 10539 70615 10581 70624
rect 10635 70664 10677 70673
rect 10635 70624 10636 70664
rect 10676 70624 10677 70664
rect 10635 70615 10677 70624
rect 10819 70664 10877 70665
rect 10819 70624 10828 70664
rect 10868 70624 10877 70664
rect 10819 70623 10877 70624
rect 10915 70664 10973 70665
rect 10915 70624 10924 70664
rect 10964 70624 10973 70664
rect 10915 70623 10973 70624
rect 11203 70664 11261 70665
rect 11203 70624 11212 70664
rect 11252 70624 11261 70664
rect 11203 70623 11261 70624
rect 11971 70664 12029 70665
rect 11971 70624 11980 70664
rect 12020 70624 12029 70664
rect 11971 70623 12029 70624
rect 12075 70664 12117 70673
rect 12075 70624 12076 70664
rect 12116 70624 12117 70664
rect 12075 70615 12117 70624
rect 12267 70664 12309 70673
rect 12739 70666 12748 70706
rect 12788 70666 12797 70706
rect 12739 70665 12797 70666
rect 12267 70624 12268 70664
rect 12308 70624 12309 70664
rect 12267 70615 12309 70624
rect 12843 70664 12885 70673
rect 12843 70624 12844 70664
rect 12884 70624 12885 70664
rect 12843 70615 12885 70624
rect 13123 70664 13181 70665
rect 13123 70624 13132 70664
rect 13172 70624 13181 70664
rect 13123 70623 13181 70624
rect 13411 70664 13469 70665
rect 13411 70624 13420 70664
rect 13460 70624 13469 70664
rect 13411 70623 13469 70624
rect 14659 70664 14717 70665
rect 14659 70624 14668 70664
rect 14708 70624 14717 70664
rect 14659 70623 14717 70624
rect 15051 70664 15093 70673
rect 15051 70624 15052 70664
rect 15092 70624 15093 70664
rect 15051 70615 15093 70624
rect 15243 70664 15285 70673
rect 15243 70624 15244 70664
rect 15284 70624 15285 70664
rect 15243 70615 15285 70624
rect 16195 70664 16253 70665
rect 16195 70624 16204 70664
rect 16244 70624 16253 70664
rect 16195 70623 16253 70624
rect 17443 70664 17501 70665
rect 17443 70624 17452 70664
rect 17492 70624 17501 70664
rect 17443 70623 17501 70624
rect 18499 70664 18557 70665
rect 18499 70624 18508 70664
rect 18548 70624 18557 70664
rect 18499 70623 18557 70624
rect 19747 70664 19805 70665
rect 19747 70624 19756 70664
rect 19796 70624 19805 70664
rect 19747 70623 19805 70624
rect 8043 70580 8085 70589
rect 8043 70540 8044 70580
rect 8084 70540 8085 70580
rect 8043 70531 8085 70540
rect 10059 70580 10101 70589
rect 10059 70540 10060 70580
rect 10100 70540 10101 70580
rect 10059 70531 10101 70540
rect 11115 70580 11157 70589
rect 11115 70540 11116 70580
rect 11156 70540 11157 70580
rect 11115 70531 11157 70540
rect 15147 70580 15189 70589
rect 15147 70540 15148 70580
rect 15188 70540 15189 70580
rect 15147 70531 15189 70540
rect 17643 70580 17685 70589
rect 17643 70540 17644 70580
rect 17684 70540 17685 70580
rect 17643 70531 17685 70540
rect 2667 70496 2709 70505
rect 2667 70456 2668 70496
rect 2708 70456 2709 70496
rect 2667 70447 2709 70456
rect 4587 70496 4629 70505
rect 4587 70456 4588 70496
rect 4628 70456 4629 70496
rect 4587 70447 4629 70456
rect 6219 70496 6261 70505
rect 6219 70456 6220 70496
rect 6260 70456 6261 70496
rect 6219 70447 6261 70456
rect 14859 70496 14901 70505
rect 14859 70456 14860 70496
rect 14900 70456 14901 70496
rect 14859 70447 14901 70456
rect 19947 70496 19989 70505
rect 19947 70456 19948 70496
rect 19988 70456 19989 70496
rect 19947 70447 19989 70456
rect 1152 70328 20452 70352
rect 1152 70288 4928 70328
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 5296 70288 20048 70328
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20416 70288 20452 70328
rect 1152 70264 20452 70288
rect 5163 70160 5205 70169
rect 5163 70120 5164 70160
rect 5204 70120 5205 70160
rect 5163 70111 5205 70120
rect 10155 70160 10197 70169
rect 10155 70120 10156 70160
rect 10196 70120 10197 70160
rect 10155 70111 10197 70120
rect 7947 70076 7989 70085
rect 7947 70036 7948 70076
rect 7988 70036 7989 70076
rect 7947 70027 7989 70036
rect 12843 70076 12885 70085
rect 12843 70036 12844 70076
rect 12884 70036 12885 70076
rect 12843 70027 12885 70036
rect 14667 70076 14709 70085
rect 14667 70036 14668 70076
rect 14708 70036 14709 70076
rect 14667 70027 14709 70036
rect 16683 70076 16725 70085
rect 16683 70036 16684 70076
rect 16724 70036 16725 70076
rect 16683 70027 16725 70036
rect 19947 70076 19989 70085
rect 19947 70036 19948 70076
rect 19988 70036 19989 70076
rect 19947 70027 19989 70036
rect 1219 69992 1277 69993
rect 1219 69952 1228 69992
rect 1268 69952 1277 69992
rect 1219 69951 1277 69952
rect 2467 69992 2525 69993
rect 2467 69952 2476 69992
rect 2516 69952 2525 69992
rect 2467 69951 2525 69952
rect 3435 69992 3477 70001
rect 3435 69952 3436 69992
rect 3476 69952 3477 69992
rect 3435 69943 3477 69952
rect 3531 69992 3573 70001
rect 3531 69952 3532 69992
rect 3572 69952 3573 69992
rect 3531 69943 3573 69952
rect 3915 69992 3957 70001
rect 3915 69952 3916 69992
rect 3956 69952 3957 69992
rect 3915 69943 3957 69952
rect 4483 69992 4541 69993
rect 4483 69952 4492 69992
rect 4532 69952 4541 69992
rect 4483 69951 4541 69952
rect 4971 69987 5013 69996
rect 4971 69947 4972 69987
rect 5012 69947 5013 69987
rect 4971 69938 5013 69947
rect 6219 69992 6261 70001
rect 6219 69952 6220 69992
rect 6260 69952 6261 69992
rect 6219 69943 6261 69952
rect 6315 69992 6357 70001
rect 6315 69952 6316 69992
rect 6356 69952 6357 69992
rect 6315 69943 6357 69952
rect 6699 69992 6741 70001
rect 6699 69952 6700 69992
rect 6740 69952 6741 69992
rect 6699 69943 6741 69952
rect 6795 69992 6837 70001
rect 6795 69952 6796 69992
rect 6836 69952 6837 69992
rect 6795 69943 6837 69952
rect 7267 69992 7325 69993
rect 7267 69952 7276 69992
rect 7316 69952 7325 69992
rect 9955 69992 10013 69993
rect 7267 69951 7325 69952
rect 7755 69978 7797 69987
rect 7755 69938 7756 69978
rect 7796 69938 7797 69978
rect 9955 69952 9964 69992
rect 10004 69952 10013 69992
rect 9955 69951 10013 69952
rect 11115 69992 11157 70001
rect 11115 69952 11116 69992
rect 11156 69952 11157 69992
rect 7755 69929 7797 69938
rect 8707 69950 8765 69951
rect 4011 69908 4053 69917
rect 8707 69910 8716 69950
rect 8756 69910 8765 69950
rect 11115 69943 11157 69952
rect 11211 69992 11253 70001
rect 11211 69952 11212 69992
rect 11252 69952 11253 69992
rect 11211 69943 11253 69952
rect 11691 69992 11733 70001
rect 11691 69952 11692 69992
rect 11732 69952 11733 69992
rect 11691 69943 11733 69952
rect 12163 69992 12221 69993
rect 12163 69952 12172 69992
rect 12212 69952 12221 69992
rect 13219 69992 13277 69993
rect 12163 69951 12221 69952
rect 12651 69978 12693 69987
rect 12651 69938 12652 69978
rect 12692 69938 12693 69978
rect 13219 69952 13228 69992
rect 13268 69952 13277 69992
rect 13219 69951 13277 69952
rect 14467 69992 14525 69993
rect 14467 69952 14476 69992
rect 14516 69952 14525 69992
rect 14467 69951 14525 69952
rect 14955 69992 14997 70001
rect 14955 69952 14956 69992
rect 14996 69952 14997 69992
rect 14955 69943 14997 69952
rect 15051 69992 15093 70001
rect 15051 69952 15052 69992
rect 15092 69952 15093 69992
rect 15051 69943 15093 69952
rect 16003 69992 16061 69993
rect 16003 69952 16012 69992
rect 16052 69952 16061 69992
rect 16003 69951 16061 69952
rect 16491 69987 16533 69996
rect 16491 69947 16492 69987
rect 16532 69947 16533 69987
rect 16491 69938 16533 69947
rect 18219 69992 18261 70001
rect 18219 69952 18220 69992
rect 18260 69952 18261 69992
rect 18219 69943 18261 69952
rect 18315 69992 18357 70001
rect 18315 69952 18316 69992
rect 18356 69952 18357 69992
rect 18315 69943 18357 69952
rect 18699 69992 18741 70001
rect 18699 69952 18700 69992
rect 18740 69952 18741 69992
rect 18699 69943 18741 69952
rect 18795 69992 18837 70001
rect 18795 69952 18796 69992
rect 18836 69952 18837 69992
rect 18795 69943 18837 69952
rect 19267 69992 19325 69993
rect 19267 69952 19276 69992
rect 19316 69952 19325 69992
rect 19267 69951 19325 69952
rect 19803 69982 19845 69991
rect 19803 69942 19804 69982
rect 19844 69942 19845 69982
rect 12651 69929 12693 69938
rect 19803 69933 19845 69942
rect 8707 69909 8765 69910
rect 4011 69868 4012 69908
rect 4052 69868 4053 69908
rect 4011 69859 4053 69868
rect 11595 69908 11637 69917
rect 11595 69868 11596 69908
rect 11636 69868 11637 69908
rect 11595 69859 11637 69868
rect 15435 69908 15477 69917
rect 15435 69868 15436 69908
rect 15476 69868 15477 69908
rect 15435 69859 15477 69868
rect 15531 69908 15573 69917
rect 15531 69868 15532 69908
rect 15572 69868 15573 69908
rect 15531 69859 15573 69868
rect 2667 69740 2709 69749
rect 2667 69700 2668 69740
rect 2708 69700 2709 69740
rect 2667 69691 2709 69700
rect 1152 69572 20352 69596
rect 1152 69532 3688 69572
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 4056 69532 18808 69572
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 19176 69532 20352 69572
rect 1152 69508 20352 69532
rect 7659 69404 7701 69413
rect 7659 69364 7660 69404
rect 7700 69364 7701 69404
rect 7659 69355 7701 69364
rect 11019 69404 11061 69413
rect 11019 69364 11020 69404
rect 11060 69364 11061 69404
rect 11019 69355 11061 69364
rect 12651 69404 12693 69413
rect 12651 69364 12652 69404
rect 12692 69364 12693 69404
rect 12651 69355 12693 69364
rect 8523 69236 8565 69245
rect 8523 69196 8524 69236
rect 8564 69196 8565 69236
rect 8523 69187 8565 69196
rect 15531 69236 15573 69245
rect 15531 69196 15532 69236
rect 15572 69196 15573 69236
rect 15531 69187 15573 69196
rect 18891 69236 18933 69245
rect 18891 69196 18892 69236
rect 18932 69196 18933 69236
rect 18891 69187 18933 69196
rect 16491 69166 16533 69175
rect 1219 69152 1277 69153
rect 1219 69112 1228 69152
rect 1268 69112 1277 69152
rect 1219 69111 1277 69112
rect 2467 69152 2525 69153
rect 2467 69112 2476 69152
rect 2516 69112 2525 69152
rect 2467 69111 2525 69112
rect 2851 69152 2909 69153
rect 2851 69112 2860 69152
rect 2900 69112 2909 69152
rect 2851 69111 2909 69112
rect 4099 69152 4157 69153
rect 4099 69112 4108 69152
rect 4148 69112 4157 69152
rect 4099 69111 4157 69112
rect 4675 69152 4733 69153
rect 4675 69112 4684 69152
rect 4724 69112 4733 69152
rect 4675 69111 4733 69112
rect 5923 69152 5981 69153
rect 5923 69112 5932 69152
rect 5972 69112 5981 69152
rect 5923 69111 5981 69112
rect 6211 69152 6269 69153
rect 6211 69112 6220 69152
rect 6260 69112 6269 69152
rect 6211 69111 6269 69112
rect 7459 69152 7517 69153
rect 7459 69112 7468 69152
rect 7508 69112 7517 69152
rect 7459 69111 7517 69112
rect 8427 69152 8469 69161
rect 8427 69112 8428 69152
rect 8468 69112 8469 69152
rect 8427 69103 8469 69112
rect 8619 69152 8661 69161
rect 8619 69112 8620 69152
rect 8660 69112 8661 69152
rect 8619 69103 8661 69112
rect 8811 69152 8853 69161
rect 8811 69112 8812 69152
rect 8852 69112 8853 69152
rect 8811 69103 8853 69112
rect 8907 69152 8949 69161
rect 8907 69112 8908 69152
rect 8948 69112 8949 69152
rect 8907 69103 8949 69112
rect 9003 69152 9045 69161
rect 9003 69112 9004 69152
rect 9044 69112 9045 69152
rect 9003 69103 9045 69112
rect 9571 69152 9629 69153
rect 9571 69112 9580 69152
rect 9620 69112 9629 69152
rect 9571 69111 9629 69112
rect 10819 69152 10877 69153
rect 10819 69112 10828 69152
rect 10868 69112 10877 69152
rect 10819 69111 10877 69112
rect 11203 69152 11261 69153
rect 11203 69112 11212 69152
rect 11252 69112 11261 69152
rect 11203 69111 11261 69112
rect 12451 69152 12509 69153
rect 12451 69112 12460 69152
rect 12500 69112 12509 69152
rect 12451 69111 12509 69112
rect 13219 69152 13277 69153
rect 13219 69112 13228 69152
rect 13268 69112 13277 69152
rect 13219 69111 13277 69112
rect 14467 69152 14525 69153
rect 14467 69112 14476 69152
rect 14516 69112 14525 69152
rect 14467 69111 14525 69112
rect 14955 69152 14997 69161
rect 14955 69112 14956 69152
rect 14996 69112 14997 69152
rect 14955 69103 14997 69112
rect 15051 69152 15093 69161
rect 15051 69112 15052 69152
rect 15092 69112 15093 69152
rect 15051 69103 15093 69112
rect 15435 69152 15477 69161
rect 15435 69112 15436 69152
rect 15476 69112 15477 69152
rect 15435 69103 15477 69112
rect 16003 69152 16061 69153
rect 16003 69112 16012 69152
rect 16052 69112 16061 69152
rect 16491 69126 16492 69166
rect 16532 69126 16533 69166
rect 19851 69166 19893 69175
rect 16491 69117 16533 69126
rect 18315 69152 18357 69161
rect 16003 69111 16061 69112
rect 18315 69112 18316 69152
rect 18356 69112 18357 69152
rect 18315 69103 18357 69112
rect 18411 69152 18453 69161
rect 18411 69112 18412 69152
rect 18452 69112 18453 69152
rect 18411 69103 18453 69112
rect 18795 69152 18837 69161
rect 18795 69112 18796 69152
rect 18836 69112 18837 69152
rect 18795 69103 18837 69112
rect 19363 69152 19421 69153
rect 19363 69112 19372 69152
rect 19412 69112 19421 69152
rect 19851 69126 19852 69166
rect 19892 69126 19893 69166
rect 19851 69117 19893 69126
rect 19363 69111 19421 69112
rect 2667 68984 2709 68993
rect 2667 68944 2668 68984
rect 2708 68944 2709 68984
rect 2667 68935 2709 68944
rect 4299 68984 4341 68993
rect 4299 68944 4300 68984
rect 4340 68944 4341 68984
rect 4299 68935 4341 68944
rect 4491 68984 4533 68993
rect 4491 68944 4492 68984
rect 4532 68944 4533 68984
rect 4491 68935 4533 68944
rect 9091 68984 9149 68985
rect 9091 68944 9100 68984
rect 9140 68944 9149 68984
rect 9091 68943 9149 68944
rect 14667 68984 14709 68993
rect 14667 68944 14668 68984
rect 14708 68944 14709 68984
rect 14667 68935 14709 68944
rect 16683 68984 16725 68993
rect 16683 68944 16684 68984
rect 16724 68944 16725 68984
rect 16683 68935 16725 68944
rect 20043 68984 20085 68993
rect 20043 68944 20044 68984
rect 20084 68944 20085 68984
rect 20043 68935 20085 68944
rect 1152 68816 20452 68840
rect 1152 68776 4928 68816
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 5296 68776 20048 68816
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20416 68776 20452 68816
rect 1152 68752 20452 68776
rect 9579 68648 9621 68657
rect 9579 68608 9580 68648
rect 9620 68608 9621 68648
rect 9579 68599 9621 68608
rect 3435 68564 3477 68573
rect 3435 68524 3436 68564
rect 3476 68524 3477 68564
rect 3435 68515 3477 68524
rect 1707 68480 1749 68489
rect 1707 68440 1708 68480
rect 1748 68440 1749 68480
rect 1707 68431 1749 68440
rect 1803 68480 1845 68489
rect 1803 68440 1804 68480
rect 1844 68440 1845 68480
rect 1803 68431 1845 68440
rect 2283 68480 2325 68489
rect 2283 68440 2284 68480
rect 2324 68440 2325 68480
rect 2283 68431 2325 68440
rect 2755 68480 2813 68481
rect 2755 68440 2764 68480
rect 2804 68440 2813 68480
rect 2755 68439 2813 68440
rect 3243 68475 3285 68484
rect 3243 68435 3244 68475
rect 3284 68435 3285 68475
rect 4771 68480 4829 68481
rect 4771 68440 4780 68480
rect 4820 68440 4829 68480
rect 4771 68439 4829 68440
rect 6019 68480 6077 68481
rect 6019 68440 6028 68480
rect 6068 68440 6077 68480
rect 6019 68439 6077 68440
rect 6499 68480 6557 68481
rect 6499 68440 6508 68480
rect 6548 68440 6557 68480
rect 6499 68439 6557 68440
rect 7747 68480 7805 68481
rect 7747 68440 7756 68480
rect 7796 68440 7805 68480
rect 7747 68439 7805 68440
rect 8131 68480 8189 68481
rect 8131 68440 8140 68480
rect 8180 68440 8189 68480
rect 8131 68439 8189 68440
rect 9379 68480 9437 68481
rect 9379 68440 9388 68480
rect 9428 68440 9437 68480
rect 9379 68439 9437 68440
rect 9771 68480 9813 68489
rect 9771 68440 9772 68480
rect 9812 68440 9813 68480
rect 3243 68426 3285 68435
rect 9771 68431 9813 68440
rect 9963 68480 10005 68489
rect 9963 68440 9964 68480
rect 10004 68440 10005 68480
rect 9963 68431 10005 68440
rect 10147 68480 10205 68481
rect 10147 68440 10156 68480
rect 10196 68440 10205 68480
rect 12547 68480 12605 68481
rect 10147 68439 10205 68440
rect 11395 68459 11453 68460
rect 11395 68419 11404 68459
rect 11444 68419 11453 68459
rect 12547 68440 12556 68480
rect 12596 68440 12605 68480
rect 12547 68439 12605 68440
rect 13795 68480 13853 68481
rect 13795 68440 13804 68480
rect 13844 68440 13853 68480
rect 13795 68439 13853 68440
rect 14179 68480 14237 68481
rect 14179 68440 14188 68480
rect 14228 68440 14237 68480
rect 14179 68439 14237 68440
rect 15427 68480 15485 68481
rect 15427 68440 15436 68480
rect 15476 68440 15485 68480
rect 15427 68439 15485 68440
rect 15907 68480 15965 68481
rect 15907 68440 15916 68480
rect 15956 68440 15965 68480
rect 15907 68439 15965 68440
rect 17155 68480 17213 68481
rect 17155 68440 17164 68480
rect 17204 68440 17213 68480
rect 17155 68439 17213 68440
rect 18403 68480 18461 68481
rect 18403 68440 18412 68480
rect 18452 68440 18461 68480
rect 18403 68439 18461 68440
rect 19651 68480 19709 68481
rect 19651 68440 19660 68480
rect 19700 68440 19709 68480
rect 19651 68439 19709 68440
rect 11395 68418 11453 68419
rect 2187 68396 2229 68405
rect 2187 68356 2188 68396
rect 2228 68356 2229 68396
rect 2187 68347 2229 68356
rect 9867 68396 9909 68405
rect 9867 68356 9868 68396
rect 9908 68356 9909 68396
rect 9867 68347 9909 68356
rect 6219 68228 6261 68237
rect 6219 68188 6220 68228
rect 6260 68188 6261 68228
rect 6219 68179 6261 68188
rect 7947 68228 7989 68237
rect 7947 68188 7948 68228
rect 7988 68188 7989 68228
rect 7947 68179 7989 68188
rect 11595 68228 11637 68237
rect 11595 68188 11596 68228
rect 11636 68188 11637 68228
rect 11595 68179 11637 68188
rect 12363 68228 12405 68237
rect 12363 68188 12364 68228
rect 12404 68188 12405 68228
rect 12363 68179 12405 68188
rect 13995 68228 14037 68237
rect 13995 68188 13996 68228
rect 14036 68188 14037 68228
rect 13995 68179 14037 68188
rect 17355 68228 17397 68237
rect 17355 68188 17356 68228
rect 17396 68188 17397 68228
rect 17355 68179 17397 68188
rect 19851 68228 19893 68237
rect 19851 68188 19852 68228
rect 19892 68188 19893 68228
rect 19851 68179 19893 68188
rect 1152 68060 20352 68084
rect 1152 68020 3688 68060
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 4056 68020 18808 68060
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 19176 68020 20352 68060
rect 1152 67996 20352 68020
rect 10347 67892 10389 67901
rect 10347 67852 10348 67892
rect 10388 67852 10389 67892
rect 10347 67843 10389 67852
rect 5163 67724 5205 67733
rect 5163 67684 5164 67724
rect 5204 67684 5205 67724
rect 5163 67675 5205 67684
rect 8427 67724 8469 67733
rect 8427 67684 8428 67724
rect 8468 67684 8469 67724
rect 8427 67675 8469 67684
rect 11979 67724 12021 67733
rect 11979 67684 11980 67724
rect 12020 67684 12021 67724
rect 11979 67675 12021 67684
rect 18411 67724 18453 67733
rect 18411 67684 18412 67724
rect 18452 67684 18453 67724
rect 18411 67675 18453 67684
rect 6219 67654 6261 67663
rect 1795 67640 1853 67641
rect 1795 67600 1804 67640
rect 1844 67600 1853 67640
rect 1795 67599 1853 67600
rect 3043 67640 3101 67641
rect 3043 67600 3052 67640
rect 3092 67600 3101 67640
rect 3043 67599 3101 67600
rect 4683 67640 4725 67649
rect 4683 67600 4684 67640
rect 4724 67600 4725 67640
rect 4683 67591 4725 67600
rect 4779 67640 4821 67649
rect 4779 67600 4780 67640
rect 4820 67600 4821 67640
rect 4779 67591 4821 67600
rect 5259 67640 5301 67649
rect 5259 67600 5260 67640
rect 5300 67600 5301 67640
rect 5259 67591 5301 67600
rect 5731 67640 5789 67641
rect 5731 67600 5740 67640
rect 5780 67600 5789 67640
rect 6219 67614 6220 67654
rect 6260 67614 6261 67654
rect 9483 67654 9525 67663
rect 6219 67605 6261 67614
rect 7371 67640 7413 67649
rect 5731 67599 5789 67600
rect 7371 67600 7372 67640
rect 7412 67600 7413 67640
rect 7371 67591 7413 67600
rect 7467 67640 7509 67649
rect 7467 67600 7468 67640
rect 7508 67600 7509 67640
rect 7467 67591 7509 67600
rect 7659 67640 7701 67649
rect 7659 67600 7660 67640
rect 7700 67600 7701 67640
rect 7659 67591 7701 67600
rect 7947 67640 7989 67649
rect 7947 67600 7948 67640
rect 7988 67600 7989 67640
rect 7947 67591 7989 67600
rect 8043 67640 8085 67649
rect 8043 67600 8044 67640
rect 8084 67600 8085 67640
rect 8043 67591 8085 67600
rect 8523 67640 8565 67649
rect 8523 67600 8524 67640
rect 8564 67600 8565 67640
rect 8523 67591 8565 67600
rect 8995 67640 9053 67641
rect 8995 67600 9004 67640
rect 9044 67600 9053 67640
rect 9483 67614 9484 67654
rect 9524 67614 9525 67654
rect 13035 67654 13077 67663
rect 9483 67605 9525 67614
rect 9867 67640 9909 67649
rect 8995 67599 9053 67600
rect 9867 67600 9868 67640
rect 9908 67600 9909 67640
rect 9867 67591 9909 67600
rect 9963 67640 10005 67649
rect 9963 67600 9964 67640
rect 10004 67600 10005 67640
rect 9963 67591 10005 67600
rect 10059 67640 10101 67649
rect 10059 67600 10060 67640
rect 10100 67600 10101 67640
rect 10059 67591 10101 67600
rect 10155 67640 10197 67649
rect 10155 67600 10156 67640
rect 10196 67600 10197 67640
rect 10155 67591 10197 67600
rect 10347 67640 10389 67649
rect 10347 67600 10348 67640
rect 10388 67600 10389 67640
rect 10347 67591 10389 67600
rect 10539 67640 10581 67649
rect 10539 67600 10540 67640
rect 10580 67600 10581 67640
rect 10539 67591 10581 67600
rect 10627 67640 10685 67641
rect 10627 67600 10636 67640
rect 10676 67600 10685 67640
rect 10627 67599 10685 67600
rect 11499 67640 11541 67649
rect 11499 67600 11500 67640
rect 11540 67600 11541 67640
rect 11499 67591 11541 67600
rect 11595 67640 11637 67649
rect 11595 67600 11596 67640
rect 11636 67600 11637 67640
rect 11595 67591 11637 67600
rect 12075 67640 12117 67649
rect 12075 67600 12076 67640
rect 12116 67600 12117 67640
rect 12075 67591 12117 67600
rect 12547 67640 12605 67641
rect 12547 67600 12556 67640
rect 12596 67600 12605 67640
rect 13035 67614 13036 67654
rect 13076 67614 13077 67654
rect 19467 67654 19509 67663
rect 13035 67605 13077 67614
rect 13603 67640 13661 67641
rect 12547 67599 12605 67600
rect 13603 67600 13612 67640
rect 13652 67600 13661 67640
rect 13603 67599 13661 67600
rect 14851 67640 14909 67641
rect 14851 67600 14860 67640
rect 14900 67600 14909 67640
rect 14851 67599 14909 67600
rect 15907 67640 15965 67641
rect 15907 67600 15916 67640
rect 15956 67600 15965 67640
rect 15907 67599 15965 67600
rect 17155 67640 17213 67641
rect 17155 67600 17164 67640
rect 17204 67600 17213 67640
rect 17155 67599 17213 67600
rect 17931 67640 17973 67649
rect 17931 67600 17932 67640
rect 17972 67600 17973 67640
rect 17931 67591 17973 67600
rect 18027 67640 18069 67649
rect 18027 67600 18028 67640
rect 18068 67600 18069 67640
rect 18027 67591 18069 67600
rect 18507 67640 18549 67649
rect 18507 67600 18508 67640
rect 18548 67600 18549 67640
rect 18507 67591 18549 67600
rect 18979 67640 19037 67641
rect 18979 67600 18988 67640
rect 19028 67600 19037 67640
rect 19467 67614 19468 67654
rect 19508 67614 19509 67654
rect 19467 67605 19509 67614
rect 18979 67599 19037 67600
rect 9675 67556 9717 67565
rect 9675 67516 9676 67556
rect 9716 67516 9717 67556
rect 9675 67507 9717 67516
rect 3243 67472 3285 67481
rect 3243 67432 3244 67472
rect 3284 67432 3285 67472
rect 3243 67423 3285 67432
rect 6411 67472 6453 67481
rect 6411 67432 6412 67472
rect 6452 67432 6453 67472
rect 6411 67423 6453 67432
rect 13227 67472 13269 67481
rect 13227 67432 13228 67472
rect 13268 67432 13269 67472
rect 13227 67423 13269 67432
rect 13419 67472 13461 67481
rect 13419 67432 13420 67472
rect 13460 67432 13461 67472
rect 13419 67423 13461 67432
rect 17355 67472 17397 67481
rect 17355 67432 17356 67472
rect 17396 67432 17397 67472
rect 17355 67423 17397 67432
rect 19659 67430 19701 67439
rect 19659 67390 19660 67430
rect 19700 67390 19701 67430
rect 19659 67381 19701 67390
rect 1152 67304 20452 67328
rect 1152 67264 4928 67304
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 5296 67264 20048 67304
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20416 67264 20452 67304
rect 1152 67240 20452 67264
rect 4203 67136 4245 67145
rect 4203 67096 4204 67136
rect 4244 67096 4245 67136
rect 4203 67087 4245 67096
rect 8619 67136 8661 67145
rect 8619 67096 8620 67136
rect 8660 67096 8661 67136
rect 8619 67087 8661 67096
rect 9291 67052 9333 67061
rect 9291 67012 9292 67052
rect 9332 67012 9333 67052
rect 9291 67003 9333 67012
rect 11211 67052 11253 67061
rect 11211 67012 11212 67052
rect 11252 67012 11253 67052
rect 11211 67003 11253 67012
rect 13227 67052 13269 67061
rect 13227 67012 13228 67052
rect 13268 67012 13269 67052
rect 13227 67003 13269 67012
rect 16107 67052 16149 67061
rect 16107 67012 16108 67052
rect 16148 67012 16149 67052
rect 16107 67003 16149 67012
rect 19659 67052 19701 67061
rect 19659 67012 19660 67052
rect 19700 67012 19701 67052
rect 19659 67003 19701 67012
rect 2475 66968 2517 66977
rect 2475 66928 2476 66968
rect 2516 66928 2517 66968
rect 2475 66919 2517 66928
rect 2571 66968 2613 66977
rect 2571 66928 2572 66968
rect 2612 66928 2613 66968
rect 2571 66919 2613 66928
rect 3051 66968 3093 66977
rect 6878 66971 6920 66980
rect 3051 66928 3052 66968
rect 3092 66928 3093 66968
rect 3051 66919 3093 66928
rect 3523 66968 3581 66969
rect 3523 66928 3532 66968
rect 3572 66928 3581 66968
rect 5155 66968 5213 66969
rect 3523 66927 3581 66928
rect 4059 66958 4101 66967
rect 4059 66918 4060 66958
rect 4100 66918 4101 66958
rect 5155 66928 5164 66968
rect 5204 66928 5213 66968
rect 5155 66927 5213 66928
rect 6403 66968 6461 66969
rect 6403 66928 6412 66968
rect 6452 66928 6461 66968
rect 6403 66927 6461 66928
rect 6878 66931 6879 66971
rect 6919 66931 6920 66971
rect 6878 66922 6920 66931
rect 7171 66968 7229 66969
rect 7171 66928 7180 66968
rect 7220 66928 7229 66968
rect 7171 66927 7229 66928
rect 8419 66968 8477 66969
rect 8419 66928 8428 66968
rect 8468 66928 8477 66968
rect 8419 66927 8477 66928
rect 8899 66968 8957 66969
rect 8899 66928 8908 66968
rect 8948 66928 8957 66968
rect 8899 66927 8957 66928
rect 9195 66968 9237 66977
rect 9195 66928 9196 66968
rect 9236 66928 9237 66968
rect 9195 66919 9237 66928
rect 9763 66968 9821 66969
rect 9763 66928 9772 66968
rect 9812 66928 9821 66968
rect 9763 66927 9821 66928
rect 11011 66968 11069 66969
rect 11011 66928 11020 66968
rect 11060 66928 11069 66968
rect 11011 66927 11069 66928
rect 11499 66968 11541 66977
rect 11499 66928 11500 66968
rect 11540 66928 11541 66968
rect 11499 66919 11541 66928
rect 11595 66968 11637 66977
rect 11595 66928 11596 66968
rect 11636 66928 11637 66968
rect 11595 66919 11637 66928
rect 11979 66968 12021 66977
rect 11979 66928 11980 66968
rect 12020 66928 12021 66968
rect 11979 66919 12021 66928
rect 12547 66968 12605 66969
rect 12547 66928 12556 66968
rect 12596 66928 12605 66968
rect 14379 66968 14421 66977
rect 12547 66927 12605 66928
rect 13083 66958 13125 66967
rect 4059 66909 4101 66918
rect 13083 66918 13084 66958
rect 13124 66918 13125 66958
rect 14379 66928 14380 66968
rect 14420 66928 14421 66968
rect 14379 66919 14421 66928
rect 14475 66968 14517 66977
rect 14475 66928 14476 66968
rect 14516 66928 14517 66968
rect 14475 66919 14517 66928
rect 14859 66968 14901 66977
rect 14859 66928 14860 66968
rect 14900 66928 14901 66968
rect 14859 66919 14901 66928
rect 14955 66968 14997 66977
rect 14955 66928 14956 66968
rect 14996 66928 14997 66968
rect 14955 66919 14997 66928
rect 15427 66968 15485 66969
rect 15427 66928 15436 66968
rect 15476 66928 15485 66968
rect 15427 66927 15485 66928
rect 15915 66963 15957 66972
rect 15915 66923 15916 66963
rect 15956 66923 15957 66963
rect 16675 66968 16733 66969
rect 16675 66928 16684 66968
rect 16724 66928 16733 66968
rect 16675 66927 16733 66928
rect 17931 66968 17973 66977
rect 17931 66928 17932 66968
rect 17972 66928 17973 66968
rect 13083 66909 13125 66918
rect 15915 66914 15957 66923
rect 17931 66919 17973 66928
rect 18027 66968 18069 66977
rect 18027 66928 18028 66968
rect 18068 66928 18069 66968
rect 18027 66919 18069 66928
rect 18411 66968 18453 66977
rect 18411 66928 18412 66968
rect 18452 66928 18453 66968
rect 18411 66919 18453 66928
rect 18507 66968 18549 66977
rect 18507 66928 18508 66968
rect 18548 66928 18549 66968
rect 18507 66919 18549 66928
rect 18979 66968 19037 66969
rect 18979 66928 18988 66968
rect 19028 66928 19037 66968
rect 18979 66927 19037 66928
rect 19467 66963 19509 66972
rect 19467 66923 19468 66963
rect 19508 66923 19509 66963
rect 19467 66914 19509 66923
rect 2955 66884 2997 66893
rect 2955 66844 2956 66884
rect 2996 66844 2997 66884
rect 2955 66835 2997 66844
rect 12075 66884 12117 66893
rect 12075 66844 12076 66884
rect 12116 66844 12117 66884
rect 12075 66835 12117 66844
rect 9571 66800 9629 66801
rect 9571 66760 9580 66800
rect 9620 66760 9629 66800
rect 9571 66759 9629 66760
rect 16971 66800 17013 66809
rect 16971 66760 16972 66800
rect 17012 66760 17013 66800
rect 16971 66751 17013 66760
rect 6603 66716 6645 66725
rect 6603 66676 6604 66716
rect 6644 66676 6645 66716
rect 6603 66667 6645 66676
rect 6987 66716 7029 66725
rect 6987 66676 6988 66716
rect 7028 66676 7029 66716
rect 6987 66667 7029 66676
rect 1152 66548 20352 66572
rect 1152 66508 3688 66548
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 4056 66508 18808 66548
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 19176 66508 20352 66548
rect 1152 66484 20352 66508
rect 8995 66296 9053 66297
rect 8995 66256 9004 66296
rect 9044 66256 9053 66296
rect 8995 66255 9053 66256
rect 7075 66157 7133 66158
rect 6681 66137 6739 66138
rect 1411 66128 1469 66129
rect 1411 66088 1420 66128
rect 1460 66088 1469 66128
rect 1411 66087 1469 66088
rect 2659 66128 2717 66129
rect 2659 66088 2668 66128
rect 2708 66088 2717 66128
rect 2659 66087 2717 66088
rect 3331 66128 3389 66129
rect 3331 66088 3340 66128
rect 3380 66088 3389 66128
rect 3331 66087 3389 66088
rect 4579 66128 4637 66129
rect 4579 66088 4588 66128
rect 4628 66088 4637 66128
rect 4579 66087 4637 66088
rect 5059 66128 5117 66129
rect 5059 66088 5068 66128
rect 5108 66088 5117 66128
rect 5059 66087 5117 66088
rect 6307 66128 6365 66129
rect 6307 66088 6316 66128
rect 6356 66088 6365 66128
rect 6681 66097 6690 66137
rect 6730 66097 6739 66137
rect 6681 66096 6739 66097
rect 6787 66128 6845 66129
rect 6307 66087 6365 66088
rect 6787 66088 6796 66128
rect 6836 66088 6845 66128
rect 6787 66087 6845 66088
rect 6987 66128 7029 66137
rect 6987 66088 6988 66128
rect 7028 66088 7029 66128
rect 7075 66117 7084 66157
rect 7124 66117 7133 66157
rect 7075 66116 7133 66117
rect 7176 66128 7234 66129
rect 6987 66079 7029 66088
rect 7176 66088 7185 66128
rect 7225 66088 7234 66128
rect 7176 66087 7234 66088
rect 7467 66128 7509 66137
rect 7467 66088 7468 66128
rect 7508 66088 7509 66128
rect 7467 66079 7509 66088
rect 7563 66128 7605 66137
rect 7563 66088 7564 66128
rect 7604 66088 7605 66128
rect 7563 66079 7605 66088
rect 8715 66128 8757 66137
rect 8715 66088 8716 66128
rect 8756 66088 8757 66128
rect 8715 66079 8757 66088
rect 8907 66128 8949 66137
rect 8907 66088 8908 66128
rect 8948 66088 8949 66128
rect 8907 66079 8949 66088
rect 9003 66128 9045 66137
rect 9003 66088 9004 66128
rect 9044 66088 9045 66128
rect 9003 66079 9045 66088
rect 9187 66128 9245 66129
rect 9187 66088 9196 66128
rect 9236 66088 9245 66128
rect 9187 66087 9245 66088
rect 9291 66128 9333 66137
rect 9291 66088 9292 66128
rect 9332 66088 9333 66128
rect 9291 66079 9333 66088
rect 11203 66128 11261 66129
rect 11203 66088 11212 66128
rect 11252 66088 11261 66128
rect 11203 66087 11261 66088
rect 12451 66128 12509 66129
rect 12451 66088 12460 66128
rect 12500 66088 12509 66128
rect 12451 66087 12509 66088
rect 12835 66128 12893 66129
rect 12835 66088 12844 66128
rect 12884 66088 12893 66128
rect 12835 66087 12893 66088
rect 14083 66128 14141 66129
rect 14083 66088 14092 66128
rect 14132 66088 14141 66128
rect 14083 66087 14141 66088
rect 14467 66128 14525 66129
rect 14467 66088 14476 66128
rect 14516 66088 14525 66128
rect 14467 66087 14525 66088
rect 15715 66128 15773 66129
rect 15715 66088 15724 66128
rect 15764 66088 15773 66128
rect 15715 66087 15773 66088
rect 16675 66128 16733 66129
rect 16675 66088 16684 66128
rect 16724 66088 16733 66128
rect 16675 66087 16733 66088
rect 17923 66128 17981 66129
rect 17923 66088 17932 66128
rect 17972 66088 17981 66128
rect 17923 66087 17981 66088
rect 18307 66128 18365 66129
rect 18307 66088 18316 66128
rect 18356 66088 18365 66128
rect 18307 66087 18365 66088
rect 19555 66128 19613 66129
rect 19555 66088 19564 66128
rect 19604 66088 19613 66128
rect 19555 66087 19613 66088
rect 2859 65960 2901 65969
rect 2859 65920 2860 65960
rect 2900 65920 2901 65960
rect 2859 65911 2901 65920
rect 4779 65960 4821 65969
rect 4779 65920 4780 65960
rect 4820 65920 4821 65960
rect 4779 65911 4821 65920
rect 6507 65960 6549 65969
rect 6507 65920 6508 65960
rect 6548 65920 6549 65960
rect 6507 65911 6549 65920
rect 7075 65960 7133 65961
rect 7075 65920 7084 65960
rect 7124 65920 7133 65960
rect 7075 65919 7133 65920
rect 7747 65960 7805 65961
rect 7747 65920 7756 65960
rect 7796 65920 7805 65960
rect 7747 65919 7805 65920
rect 12651 65960 12693 65969
rect 12651 65920 12652 65960
rect 12692 65920 12693 65960
rect 12651 65911 12693 65920
rect 14283 65960 14325 65969
rect 14283 65920 14284 65960
rect 14324 65920 14325 65960
rect 14283 65911 14325 65920
rect 15915 65960 15957 65969
rect 15915 65920 15916 65960
rect 15956 65920 15957 65960
rect 15915 65911 15957 65920
rect 18123 65960 18165 65969
rect 18123 65920 18124 65960
rect 18164 65920 18165 65960
rect 18123 65911 18165 65920
rect 19755 65960 19797 65969
rect 19755 65920 19756 65960
rect 19796 65920 19797 65960
rect 19755 65911 19797 65920
rect 1152 65792 20452 65816
rect 1152 65752 4928 65792
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 5296 65752 20048 65792
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20416 65752 20452 65792
rect 1152 65728 20452 65752
rect 5739 65624 5781 65633
rect 5739 65584 5740 65624
rect 5780 65584 5781 65624
rect 5739 65575 5781 65584
rect 9195 65624 9237 65633
rect 9195 65584 9196 65624
rect 9236 65584 9237 65624
rect 9195 65575 9237 65584
rect 4587 65540 4629 65549
rect 4587 65500 4588 65540
rect 4628 65500 4629 65540
rect 4587 65491 4629 65500
rect 10827 65540 10869 65549
rect 10827 65500 10828 65540
rect 10868 65500 10869 65540
rect 10827 65491 10869 65500
rect 12843 65540 12885 65549
rect 12843 65500 12844 65540
rect 12884 65500 12885 65540
rect 12843 65491 12885 65500
rect 16011 65540 16053 65549
rect 16011 65500 16012 65540
rect 16052 65500 16053 65540
rect 16011 65491 16053 65500
rect 19179 65540 19221 65549
rect 19179 65500 19180 65540
rect 19220 65500 19221 65540
rect 19179 65491 19221 65500
rect 2859 65456 2901 65465
rect 2859 65416 2860 65456
rect 2900 65416 2901 65456
rect 2859 65407 2901 65416
rect 2955 65456 2997 65465
rect 2955 65416 2956 65456
rect 2996 65416 2997 65456
rect 2955 65407 2997 65416
rect 3435 65456 3477 65465
rect 3435 65416 3436 65456
rect 3476 65416 3477 65456
rect 3435 65407 3477 65416
rect 3907 65456 3965 65457
rect 3907 65416 3916 65456
rect 3956 65416 3965 65456
rect 5643 65456 5685 65465
rect 3907 65415 3965 65416
rect 4443 65446 4485 65455
rect 4443 65406 4444 65446
rect 4484 65406 4485 65446
rect 5643 65416 5644 65456
rect 5684 65416 5685 65456
rect 5643 65407 5685 65416
rect 5835 65456 5877 65465
rect 5835 65416 5836 65456
rect 5876 65416 5877 65456
rect 5835 65407 5877 65416
rect 5931 65456 5973 65465
rect 5931 65416 5932 65456
rect 5972 65416 5973 65456
rect 5931 65407 5973 65416
rect 6115 65456 6173 65457
rect 6115 65416 6124 65456
rect 6164 65416 6173 65456
rect 6115 65415 6173 65416
rect 7363 65456 7421 65457
rect 7363 65416 7372 65456
rect 7412 65416 7421 65456
rect 7363 65415 7421 65416
rect 7747 65456 7805 65457
rect 7747 65416 7756 65456
rect 7796 65416 7805 65456
rect 7747 65415 7805 65416
rect 9379 65456 9437 65457
rect 9379 65416 9388 65456
rect 9428 65416 9437 65456
rect 9379 65415 9437 65416
rect 10627 65456 10685 65457
rect 10627 65416 10636 65456
rect 10676 65416 10685 65456
rect 10627 65415 10685 65416
rect 11115 65456 11157 65465
rect 11115 65416 11116 65456
rect 11156 65416 11157 65456
rect 8995 65414 9053 65415
rect 4443 65397 4485 65406
rect 3339 65372 3381 65381
rect 8995 65374 9004 65414
rect 9044 65374 9053 65414
rect 11115 65407 11157 65416
rect 11211 65456 11253 65465
rect 11211 65416 11212 65456
rect 11252 65416 11253 65456
rect 11211 65407 11253 65416
rect 11595 65456 11637 65465
rect 11595 65416 11596 65456
rect 11636 65416 11637 65456
rect 11595 65407 11637 65416
rect 11691 65456 11733 65465
rect 11691 65416 11692 65456
rect 11732 65416 11733 65456
rect 11691 65407 11733 65416
rect 12163 65456 12221 65457
rect 12163 65416 12172 65456
rect 12212 65416 12221 65456
rect 12163 65415 12221 65416
rect 12651 65451 12693 65460
rect 12651 65411 12652 65451
rect 12692 65411 12693 65451
rect 12651 65402 12693 65411
rect 14283 65456 14325 65465
rect 14283 65416 14284 65456
rect 14324 65416 14325 65456
rect 14283 65407 14325 65416
rect 14379 65456 14421 65465
rect 14379 65416 14380 65456
rect 14420 65416 14421 65456
rect 14379 65407 14421 65416
rect 14763 65456 14805 65465
rect 14763 65416 14764 65456
rect 14804 65416 14805 65456
rect 14763 65407 14805 65416
rect 14859 65456 14901 65465
rect 14859 65416 14860 65456
rect 14900 65416 14901 65456
rect 14859 65407 14901 65416
rect 15331 65456 15389 65457
rect 15331 65416 15340 65456
rect 15380 65416 15389 65456
rect 17451 65456 17493 65465
rect 15331 65415 15389 65416
rect 15867 65446 15909 65455
rect 15867 65406 15868 65446
rect 15908 65406 15909 65446
rect 17451 65416 17452 65456
rect 17492 65416 17493 65456
rect 17451 65407 17493 65416
rect 17547 65456 17589 65465
rect 17547 65416 17548 65456
rect 17588 65416 17589 65456
rect 17547 65407 17589 65416
rect 18027 65456 18069 65465
rect 18027 65416 18028 65456
rect 18068 65416 18069 65456
rect 18027 65407 18069 65416
rect 18499 65456 18557 65457
rect 18499 65416 18508 65456
rect 18548 65416 18557 65456
rect 18499 65415 18557 65416
rect 18987 65451 19029 65460
rect 18987 65411 18988 65451
rect 19028 65411 19029 65451
rect 15867 65397 15909 65406
rect 18987 65402 19029 65411
rect 8995 65373 9053 65374
rect 3339 65332 3340 65372
rect 3380 65332 3381 65372
rect 3339 65323 3381 65332
rect 16483 65372 16541 65373
rect 16483 65332 16492 65372
rect 16532 65332 16541 65372
rect 16483 65331 16541 65332
rect 17931 65372 17973 65381
rect 17931 65332 17932 65372
rect 17972 65332 17973 65372
rect 17931 65323 17973 65332
rect 16683 65288 16725 65297
rect 16683 65248 16684 65288
rect 16724 65248 16725 65288
rect 16683 65239 16725 65248
rect 7563 65204 7605 65213
rect 7563 65164 7564 65204
rect 7604 65164 7605 65204
rect 7563 65155 7605 65164
rect 1152 65036 20352 65060
rect 1152 64996 3688 65036
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 4056 64996 18808 65036
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 19176 64996 20352 65036
rect 1152 64972 20352 64996
rect 9291 64868 9333 64877
rect 9291 64828 9292 64868
rect 9332 64828 9333 64868
rect 9291 64819 9333 64828
rect 2667 64700 2709 64709
rect 2667 64660 2668 64700
rect 2708 64660 2709 64700
rect 2667 64651 2709 64660
rect 6219 64700 6261 64709
rect 6219 64660 6220 64700
rect 6260 64660 6261 64700
rect 6219 64651 6261 64660
rect 18027 64700 18069 64709
rect 18027 64660 18028 64700
rect 18068 64660 18069 64700
rect 18027 64651 18069 64660
rect 18123 64700 18165 64709
rect 18123 64660 18124 64700
rect 18164 64660 18165 64700
rect 18123 64651 18165 64660
rect 19843 64700 19901 64701
rect 19843 64660 19852 64700
rect 19892 64660 19901 64700
rect 19843 64659 19901 64660
rect 9483 64639 9525 64648
rect 3627 64630 3669 64639
rect 2091 64616 2133 64625
rect 2091 64576 2092 64616
rect 2132 64576 2133 64616
rect 2091 64567 2133 64576
rect 2187 64616 2229 64625
rect 2187 64576 2188 64616
rect 2228 64576 2229 64616
rect 2187 64567 2229 64576
rect 2571 64616 2613 64625
rect 2571 64576 2572 64616
rect 2612 64576 2613 64616
rect 2571 64567 2613 64576
rect 3139 64616 3197 64617
rect 3139 64576 3148 64616
rect 3188 64576 3197 64616
rect 3627 64590 3628 64630
rect 3668 64590 3669 64630
rect 3627 64581 3669 64590
rect 4003 64616 4061 64617
rect 3139 64575 3197 64576
rect 4003 64576 4012 64616
rect 4052 64576 4061 64616
rect 4003 64575 4061 64576
rect 5251 64616 5309 64617
rect 5251 64576 5260 64616
rect 5300 64576 5309 64616
rect 5251 64575 5309 64576
rect 5739 64616 5781 64625
rect 5739 64576 5740 64616
rect 5780 64576 5781 64616
rect 5739 64567 5781 64576
rect 5835 64616 5877 64625
rect 5835 64576 5836 64616
rect 5876 64576 5877 64616
rect 5835 64567 5877 64576
rect 6315 64616 6357 64625
rect 7275 64621 7317 64630
rect 6315 64576 6316 64616
rect 6356 64576 6357 64616
rect 6315 64567 6357 64576
rect 6787 64616 6845 64617
rect 6787 64576 6796 64616
rect 6836 64576 6845 64616
rect 6787 64575 6845 64576
rect 7275 64581 7276 64621
rect 7316 64581 7317 64621
rect 7275 64572 7317 64581
rect 7843 64616 7901 64617
rect 7843 64576 7852 64616
rect 7892 64576 7901 64616
rect 7843 64575 7901 64576
rect 9091 64616 9149 64617
rect 9091 64576 9100 64616
rect 9140 64576 9149 64616
rect 9483 64599 9484 64639
rect 9524 64599 9525 64639
rect 19131 64625 19173 64634
rect 9483 64590 9525 64599
rect 9571 64616 9629 64617
rect 9091 64575 9149 64576
rect 9571 64576 9580 64616
rect 9620 64576 9629 64616
rect 9571 64575 9629 64576
rect 9771 64616 9813 64625
rect 9771 64576 9772 64616
rect 9812 64576 9813 64616
rect 9771 64567 9813 64576
rect 9867 64616 9909 64625
rect 9867 64576 9868 64616
rect 9908 64576 9909 64616
rect 9867 64567 9909 64576
rect 10014 64616 10072 64617
rect 10014 64576 10023 64616
rect 10063 64576 10072 64616
rect 10014 64575 10072 64576
rect 10243 64616 10301 64617
rect 10243 64576 10252 64616
rect 10292 64576 10301 64616
rect 10243 64575 10301 64576
rect 10347 64616 10389 64625
rect 10347 64576 10348 64616
rect 10388 64576 10389 64616
rect 10347 64567 10389 64576
rect 10819 64616 10877 64617
rect 10819 64576 10828 64616
rect 10868 64576 10877 64616
rect 10819 64575 10877 64576
rect 12067 64616 12125 64617
rect 12067 64576 12076 64616
rect 12116 64576 12125 64616
rect 12067 64575 12125 64576
rect 12643 64616 12701 64617
rect 12643 64576 12652 64616
rect 12692 64576 12701 64616
rect 12643 64575 12701 64576
rect 13891 64616 13949 64617
rect 13891 64576 13900 64616
rect 13940 64576 13949 64616
rect 13891 64575 13949 64576
rect 14467 64616 14525 64617
rect 14467 64576 14476 64616
rect 14516 64576 14525 64616
rect 14467 64575 14525 64576
rect 15715 64616 15773 64617
rect 15715 64576 15724 64616
rect 15764 64576 15773 64616
rect 15715 64575 15773 64576
rect 17547 64616 17589 64625
rect 17547 64576 17548 64616
rect 17588 64576 17589 64616
rect 17547 64567 17589 64576
rect 17643 64616 17685 64625
rect 17643 64576 17644 64616
rect 17684 64576 17685 64616
rect 17643 64567 17685 64576
rect 18595 64616 18653 64617
rect 18595 64576 18604 64616
rect 18644 64576 18653 64616
rect 19131 64585 19132 64625
rect 19172 64585 19173 64625
rect 19131 64576 19173 64585
rect 18595 64575 18653 64576
rect 3819 64532 3861 64541
rect 3819 64492 3820 64532
rect 3860 64492 3861 64532
rect 3819 64483 3861 64492
rect 9475 64532 9533 64533
rect 9475 64492 9484 64532
rect 9524 64492 9533 64532
rect 9475 64491 9533 64492
rect 5451 64448 5493 64457
rect 5451 64408 5452 64448
rect 5492 64408 5493 64448
rect 10635 64448 10677 64457
rect 5451 64399 5493 64408
rect 7467 64406 7509 64415
rect 7467 64366 7468 64406
rect 7508 64366 7509 64406
rect 10635 64408 10636 64448
rect 10676 64408 10677 64448
rect 10635 64399 10677 64408
rect 14091 64448 14133 64457
rect 14091 64408 14092 64448
rect 14132 64408 14133 64448
rect 14091 64399 14133 64408
rect 15915 64448 15957 64457
rect 15915 64408 15916 64448
rect 15956 64408 15957 64448
rect 15915 64399 15957 64408
rect 19275 64448 19317 64457
rect 19275 64408 19276 64448
rect 19316 64408 19317 64448
rect 19275 64399 19317 64408
rect 20043 64448 20085 64457
rect 20043 64408 20044 64448
rect 20084 64408 20085 64448
rect 20043 64399 20085 64408
rect 7467 64357 7509 64366
rect 1152 64280 20452 64304
rect 1152 64240 4928 64280
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 5296 64240 20048 64280
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20416 64240 20452 64280
rect 1152 64216 20452 64240
rect 8227 64112 8285 64113
rect 8227 64072 8236 64112
rect 8276 64072 8285 64112
rect 8227 64071 8285 64072
rect 15723 64028 15765 64037
rect 15723 63988 15724 64028
rect 15764 63988 15765 64028
rect 15723 63979 15765 63988
rect 1411 63944 1469 63945
rect 1411 63904 1420 63944
rect 1460 63904 1469 63944
rect 1411 63903 1469 63904
rect 2659 63944 2717 63945
rect 2659 63904 2668 63944
rect 2708 63904 2717 63944
rect 2659 63903 2717 63904
rect 3811 63944 3869 63945
rect 3811 63904 3820 63944
rect 3860 63904 3869 63944
rect 3811 63903 3869 63904
rect 5059 63944 5117 63945
rect 5059 63904 5068 63944
rect 5108 63904 5117 63944
rect 5059 63903 5117 63904
rect 6019 63944 6077 63945
rect 6019 63904 6028 63944
rect 6068 63904 6077 63944
rect 6019 63903 6077 63904
rect 7267 63944 7325 63945
rect 7267 63904 7276 63944
rect 7316 63904 7325 63944
rect 7267 63903 7325 63904
rect 8427 63944 8469 63953
rect 8427 63904 8428 63944
rect 8468 63904 8469 63944
rect 8427 63895 8469 63904
rect 8523 63944 8565 63953
rect 8523 63904 8524 63944
rect 8564 63904 8565 63944
rect 8523 63895 8565 63904
rect 8707 63944 8765 63945
rect 8707 63904 8716 63944
rect 8756 63904 8765 63944
rect 8707 63903 8765 63904
rect 9955 63944 10013 63945
rect 9955 63904 9964 63944
rect 10004 63904 10013 63944
rect 9955 63903 10013 63904
rect 10339 63944 10397 63945
rect 10339 63904 10348 63944
rect 10388 63904 10397 63944
rect 10339 63903 10397 63904
rect 11587 63944 11645 63945
rect 11587 63904 11596 63944
rect 11636 63904 11645 63944
rect 11587 63903 11645 63904
rect 12259 63944 12317 63945
rect 12259 63904 12268 63944
rect 12308 63904 12317 63944
rect 12259 63903 12317 63904
rect 13507 63944 13565 63945
rect 13507 63904 13516 63944
rect 13556 63904 13565 63944
rect 13507 63903 13565 63904
rect 13995 63944 14037 63953
rect 13995 63904 13996 63944
rect 14036 63904 14037 63944
rect 13995 63895 14037 63904
rect 14091 63944 14133 63953
rect 14091 63904 14092 63944
rect 14132 63904 14133 63944
rect 14091 63895 14133 63904
rect 14571 63944 14613 63953
rect 14571 63904 14572 63944
rect 14612 63904 14613 63944
rect 14571 63895 14613 63904
rect 15043 63944 15101 63945
rect 15043 63904 15052 63944
rect 15092 63904 15101 63944
rect 15043 63903 15101 63904
rect 15531 63939 15573 63948
rect 15531 63899 15532 63939
rect 15572 63899 15573 63939
rect 16291 63944 16349 63945
rect 16291 63904 16300 63944
rect 16340 63904 16349 63944
rect 16291 63903 16349 63904
rect 17539 63944 17597 63945
rect 17539 63904 17548 63944
rect 17588 63904 17597 63944
rect 17539 63903 17597 63904
rect 18115 63944 18173 63945
rect 18115 63904 18124 63944
rect 18164 63904 18173 63944
rect 18115 63903 18173 63904
rect 19363 63944 19421 63945
rect 19363 63904 19372 63944
rect 19412 63904 19421 63944
rect 19363 63903 19421 63904
rect 15531 63890 15573 63899
rect 14475 63860 14517 63869
rect 14475 63820 14476 63860
rect 14516 63820 14517 63860
rect 14475 63811 14517 63820
rect 19747 63860 19805 63861
rect 19747 63820 19756 63860
rect 19796 63820 19805 63860
rect 19747 63819 19805 63820
rect 2859 63692 2901 63701
rect 2859 63652 2860 63692
rect 2900 63652 2901 63692
rect 2859 63643 2901 63652
rect 5259 63692 5301 63701
rect 5259 63652 5260 63692
rect 5300 63652 5301 63692
rect 5259 63643 5301 63652
rect 7467 63692 7509 63701
rect 7467 63652 7468 63692
rect 7508 63652 7509 63692
rect 7467 63643 7509 63652
rect 10155 63692 10197 63701
rect 10155 63652 10156 63692
rect 10196 63652 10197 63692
rect 10155 63643 10197 63652
rect 11787 63692 11829 63701
rect 11787 63652 11788 63692
rect 11828 63652 11829 63692
rect 11787 63643 11829 63652
rect 13707 63692 13749 63701
rect 13707 63652 13708 63692
rect 13748 63652 13749 63692
rect 13707 63643 13749 63652
rect 17739 63692 17781 63701
rect 17739 63652 17740 63692
rect 17780 63652 17781 63692
rect 17739 63643 17781 63652
rect 17931 63692 17973 63701
rect 17931 63652 17932 63692
rect 17972 63652 17973 63692
rect 17931 63643 17973 63652
rect 19947 63692 19989 63701
rect 19947 63652 19948 63692
rect 19988 63652 19989 63692
rect 19947 63643 19989 63652
rect 1152 63524 20352 63548
rect 1152 63484 3688 63524
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 4056 63484 18808 63524
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 19176 63484 20352 63524
rect 1152 63460 20352 63484
rect 1515 63272 1557 63281
rect 1515 63232 1516 63272
rect 1556 63232 1557 63272
rect 1515 63223 1557 63232
rect 1899 63272 1941 63281
rect 1899 63232 1900 63272
rect 1940 63232 1941 63272
rect 1899 63223 1941 63232
rect 2283 63272 2325 63281
rect 2283 63232 2284 63272
rect 2324 63232 2325 63272
rect 2283 63223 2325 63232
rect 1699 63188 1757 63189
rect 1699 63148 1708 63188
rect 1748 63148 1757 63188
rect 1699 63147 1757 63148
rect 2083 63188 2141 63189
rect 2083 63148 2092 63188
rect 2132 63148 2141 63188
rect 2083 63147 2141 63148
rect 2467 63188 2525 63189
rect 2467 63148 2476 63188
rect 2516 63148 2525 63188
rect 2467 63147 2525 63148
rect 6507 63188 6549 63197
rect 6507 63148 6508 63188
rect 6548 63148 6549 63188
rect 5539 63146 5597 63147
rect 5539 63106 5548 63146
rect 5588 63106 5597 63146
rect 6507 63139 6549 63148
rect 6603 63188 6645 63197
rect 6603 63148 6604 63188
rect 6644 63148 6645 63188
rect 6603 63139 6645 63148
rect 10251 63188 10293 63197
rect 10251 63148 10252 63188
rect 10292 63148 10293 63188
rect 10251 63139 10293 63148
rect 10347 63188 10389 63197
rect 10347 63148 10348 63188
rect 10388 63148 10389 63188
rect 10347 63139 10389 63148
rect 12267 63188 12309 63197
rect 12267 63148 12268 63188
rect 12308 63148 12309 63188
rect 12267 63139 12309 63148
rect 12363 63188 12405 63197
rect 12363 63148 12364 63188
rect 12404 63148 12405 63188
rect 12363 63139 12405 63148
rect 18411 63188 18453 63197
rect 18411 63148 18412 63188
rect 18452 63148 18453 63188
rect 18411 63139 18453 63148
rect 18507 63188 18549 63197
rect 18507 63148 18508 63188
rect 18548 63148 18549 63188
rect 19843 63188 19901 63189
rect 18507 63139 18549 63148
rect 19515 63146 19557 63155
rect 19843 63148 19852 63188
rect 19892 63148 19901 63188
rect 19843 63147 19901 63148
rect 7563 63118 7605 63127
rect 11787 63123 11829 63132
rect 5539 63105 5597 63106
rect 2851 63104 2909 63105
rect 2851 63064 2860 63104
rect 2900 63064 2909 63104
rect 2851 63063 2909 63064
rect 4099 63104 4157 63105
rect 4099 63064 4108 63104
rect 4148 63064 4157 63104
rect 4099 63063 4157 63064
rect 4291 63104 4349 63105
rect 4291 63064 4300 63104
rect 4340 63064 4349 63104
rect 4291 63063 4349 63064
rect 6027 63104 6069 63113
rect 6027 63064 6028 63104
rect 6068 63064 6069 63104
rect 6027 63055 6069 63064
rect 6123 63104 6165 63113
rect 6123 63064 6124 63104
rect 6164 63064 6165 63104
rect 6123 63055 6165 63064
rect 7075 63104 7133 63105
rect 7075 63064 7084 63104
rect 7124 63064 7133 63104
rect 7563 63078 7564 63118
rect 7604 63078 7605 63118
rect 7563 63069 7605 63078
rect 8035 63104 8093 63105
rect 7075 63063 7133 63064
rect 8035 63064 8044 63104
rect 8084 63064 8093 63104
rect 8035 63063 8093 63064
rect 9283 63104 9341 63105
rect 9283 63064 9292 63104
rect 9332 63064 9341 63104
rect 9283 63063 9341 63064
rect 9771 63104 9813 63113
rect 9771 63064 9772 63104
rect 9812 63064 9813 63104
rect 9771 63055 9813 63064
rect 9867 63104 9909 63113
rect 11307 63109 11349 63118
rect 9867 63064 9868 63104
rect 9908 63064 9909 63104
rect 9867 63055 9909 63064
rect 10819 63104 10877 63105
rect 10819 63064 10828 63104
rect 10868 63064 10877 63104
rect 10819 63063 10877 63064
rect 11307 63069 11308 63109
rect 11348 63069 11349 63109
rect 11787 63083 11788 63123
rect 11828 63083 11829 63123
rect 13323 63118 13365 63127
rect 11787 63074 11829 63083
rect 11883 63104 11925 63113
rect 11307 63060 11349 63069
rect 11883 63064 11884 63104
rect 11924 63064 11925 63104
rect 11883 63055 11925 63064
rect 12835 63104 12893 63105
rect 12835 63064 12844 63104
rect 12884 63064 12893 63104
rect 13323 63078 13324 63118
rect 13364 63078 13365 63118
rect 13323 63069 13365 63078
rect 14851 63104 14909 63105
rect 12835 63063 12893 63064
rect 14851 63064 14860 63104
rect 14900 63064 14909 63104
rect 14851 63063 14909 63064
rect 16099 63104 16157 63105
rect 16099 63064 16108 63104
rect 16148 63064 16157 63104
rect 16099 63063 16157 63064
rect 17931 63104 17973 63113
rect 17931 63064 17932 63104
rect 17972 63064 17973 63104
rect 17931 63055 17973 63064
rect 18027 63104 18069 63113
rect 19515 63106 19516 63146
rect 19556 63106 19557 63146
rect 18027 63064 18028 63104
rect 18068 63064 18069 63104
rect 18027 63055 18069 63064
rect 18979 63104 19037 63105
rect 18979 63064 18988 63104
rect 19028 63064 19037 63104
rect 19515 63097 19557 63106
rect 18979 63063 19037 63064
rect 2667 63020 2709 63029
rect 2667 62980 2668 63020
rect 2708 62980 2709 63020
rect 2667 62971 2709 62980
rect 5739 63020 5781 63029
rect 5739 62980 5740 63020
rect 5780 62980 5781 63020
rect 5739 62971 5781 62980
rect 7755 62936 7797 62945
rect 7755 62896 7756 62936
rect 7796 62896 7797 62936
rect 7755 62887 7797 62896
rect 9483 62936 9525 62945
rect 9483 62896 9484 62936
rect 9524 62896 9525 62936
rect 9483 62887 9525 62896
rect 11499 62936 11541 62945
rect 11499 62896 11500 62936
rect 11540 62896 11541 62936
rect 11499 62887 11541 62896
rect 13515 62936 13557 62945
rect 13515 62896 13516 62936
rect 13556 62896 13557 62936
rect 13515 62887 13557 62896
rect 16299 62936 16341 62945
rect 16299 62896 16300 62936
rect 16340 62896 16341 62936
rect 16299 62887 16341 62896
rect 19659 62936 19701 62945
rect 19659 62896 19660 62936
rect 19700 62896 19701 62936
rect 19659 62887 19701 62896
rect 20043 62936 20085 62945
rect 20043 62896 20044 62936
rect 20084 62896 20085 62936
rect 20043 62887 20085 62896
rect 1152 62768 20452 62792
rect 1152 62728 4928 62768
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 5296 62728 20048 62768
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20416 62728 20452 62768
rect 1152 62704 20452 62728
rect 5067 62600 5109 62609
rect 5067 62560 5068 62600
rect 5108 62560 5109 62600
rect 5067 62551 5109 62560
rect 16107 62600 16149 62609
rect 16107 62560 16108 62600
rect 16148 62560 16149 62600
rect 16107 62551 16149 62560
rect 16875 62600 16917 62609
rect 16875 62560 16876 62600
rect 16916 62560 16917 62600
rect 16875 62551 16917 62560
rect 19659 62600 19701 62609
rect 19659 62560 19660 62600
rect 19700 62560 19701 62600
rect 19659 62551 19701 62560
rect 9963 62516 10005 62525
rect 9963 62476 9964 62516
rect 10004 62476 10005 62516
rect 9963 62467 10005 62476
rect 3339 62452 3381 62461
rect 1315 62432 1373 62433
rect 1315 62392 1324 62432
rect 1364 62392 1373 62432
rect 1315 62391 1373 62392
rect 2563 62432 2621 62433
rect 2563 62392 2572 62432
rect 2612 62392 2621 62432
rect 3339 62412 3340 62452
rect 3380 62412 3381 62452
rect 3339 62403 3381 62412
rect 3435 62432 3477 62441
rect 2563 62391 2621 62392
rect 3435 62392 3436 62432
rect 3476 62392 3477 62432
rect 3435 62383 3477 62392
rect 4387 62432 4445 62433
rect 4387 62392 4396 62432
rect 4436 62392 4445 62432
rect 4387 62391 4445 62392
rect 4875 62427 4917 62436
rect 4875 62387 4876 62427
rect 4916 62387 4917 62427
rect 6499 62432 6557 62433
rect 6499 62392 6508 62432
rect 6548 62392 6557 62432
rect 6499 62391 6557 62392
rect 7747 62432 7805 62433
rect 7747 62392 7756 62432
rect 7796 62392 7805 62432
rect 7747 62391 7805 62392
rect 8235 62432 8277 62441
rect 8235 62392 8236 62432
rect 8276 62392 8277 62432
rect 4875 62378 4917 62387
rect 8235 62383 8277 62392
rect 8331 62432 8373 62441
rect 8331 62392 8332 62432
rect 8372 62392 8373 62432
rect 8331 62383 8373 62392
rect 8715 62432 8757 62441
rect 8715 62392 8716 62432
rect 8756 62392 8757 62432
rect 8715 62383 8757 62392
rect 8811 62432 8853 62441
rect 8811 62392 8812 62432
rect 8852 62392 8853 62432
rect 8811 62383 8853 62392
rect 9283 62432 9341 62433
rect 9283 62392 9292 62432
rect 9332 62392 9341 62432
rect 9283 62391 9341 62392
rect 9771 62427 9813 62436
rect 9771 62387 9772 62427
rect 9812 62387 9813 62427
rect 11107 62432 11165 62433
rect 11107 62392 11116 62432
rect 11156 62392 11165 62432
rect 11107 62391 11165 62392
rect 12355 62432 12413 62433
rect 12355 62392 12364 62432
rect 12404 62392 12413 62432
rect 12355 62391 12413 62392
rect 14379 62432 14421 62441
rect 14379 62392 14380 62432
rect 14420 62392 14421 62432
rect 9771 62378 9813 62387
rect 14379 62383 14421 62392
rect 14475 62432 14517 62441
rect 14475 62392 14476 62432
rect 14516 62392 14517 62432
rect 14475 62383 14517 62392
rect 14859 62432 14901 62441
rect 14859 62392 14860 62432
rect 14900 62392 14901 62432
rect 14859 62383 14901 62392
rect 15427 62432 15485 62433
rect 15427 62392 15436 62432
rect 15476 62392 15485 62432
rect 17931 62432 17973 62441
rect 15427 62391 15485 62392
rect 15963 62422 16005 62431
rect 15963 62382 15964 62422
rect 16004 62382 16005 62422
rect 17931 62392 17932 62432
rect 17972 62392 17973 62432
rect 17931 62383 17973 62392
rect 18027 62432 18069 62441
rect 18027 62392 18028 62432
rect 18068 62392 18069 62432
rect 18027 62383 18069 62392
rect 18411 62432 18453 62441
rect 18411 62392 18412 62432
rect 18452 62392 18453 62432
rect 18411 62383 18453 62392
rect 18507 62432 18549 62441
rect 18507 62392 18508 62432
rect 18548 62392 18549 62432
rect 18507 62383 18549 62392
rect 18979 62432 19037 62433
rect 18979 62392 18988 62432
rect 19028 62392 19037 62432
rect 18979 62391 19037 62392
rect 19467 62427 19509 62436
rect 19467 62387 19468 62427
rect 19508 62387 19509 62427
rect 15963 62373 16005 62382
rect 19467 62378 19509 62387
rect 3819 62348 3861 62357
rect 3819 62308 3820 62348
rect 3860 62308 3861 62348
rect 3819 62299 3861 62308
rect 3915 62348 3957 62357
rect 3915 62308 3916 62348
rect 3956 62308 3957 62348
rect 3915 62299 3957 62308
rect 13219 62348 13277 62349
rect 13219 62308 13228 62348
rect 13268 62308 13277 62348
rect 13219 62307 13277 62308
rect 14955 62348 14997 62357
rect 14955 62308 14956 62348
rect 14996 62308 14997 62348
rect 14955 62299 14997 62308
rect 16675 62348 16733 62349
rect 16675 62308 16684 62348
rect 16724 62308 16733 62348
rect 16675 62307 16733 62308
rect 19843 62348 19901 62349
rect 19843 62308 19852 62348
rect 19892 62308 19901 62348
rect 19843 62307 19901 62308
rect 2763 62180 2805 62189
rect 2763 62140 2764 62180
rect 2804 62140 2805 62180
rect 2763 62131 2805 62140
rect 7947 62180 7989 62189
rect 7947 62140 7948 62180
rect 7988 62140 7989 62180
rect 7947 62131 7989 62140
rect 12555 62180 12597 62189
rect 12555 62140 12556 62180
rect 12596 62140 12597 62180
rect 12555 62131 12597 62140
rect 13035 62180 13077 62189
rect 13035 62140 13036 62180
rect 13076 62140 13077 62180
rect 13035 62131 13077 62140
rect 20043 62180 20085 62189
rect 20043 62140 20044 62180
rect 20084 62140 20085 62180
rect 20043 62131 20085 62140
rect 1152 62012 20352 62036
rect 1152 61972 3688 62012
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 4056 61972 18808 62012
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 19176 61972 20352 62012
rect 1152 61948 20352 61972
rect 14667 61844 14709 61853
rect 14667 61804 14668 61844
rect 14708 61804 14709 61844
rect 14667 61795 14709 61804
rect 16107 61760 16149 61769
rect 16107 61720 16108 61760
rect 16148 61720 16149 61760
rect 16107 61711 16149 61720
rect 4107 61676 4149 61685
rect 4107 61636 4108 61676
rect 4148 61636 4149 61676
rect 4107 61627 4149 61636
rect 4203 61676 4245 61685
rect 4203 61636 4204 61676
rect 4244 61636 4245 61676
rect 4203 61627 4245 61636
rect 14851 61676 14909 61677
rect 14851 61636 14860 61676
rect 14900 61636 14909 61676
rect 14851 61635 14909 61636
rect 15907 61676 15965 61677
rect 15907 61636 15916 61676
rect 15956 61636 15965 61676
rect 15907 61635 15965 61636
rect 19747 61676 19805 61677
rect 19747 61636 19756 61676
rect 19796 61636 19805 61676
rect 19747 61635 19805 61636
rect 3147 61606 3189 61615
rect 1315 61592 1373 61593
rect 1315 61552 1324 61592
rect 1364 61552 1373 61592
rect 1315 61551 1373 61552
rect 2563 61592 2621 61593
rect 2563 61552 2572 61592
rect 2612 61552 2621 61592
rect 3147 61566 3148 61606
rect 3188 61566 3189 61606
rect 3147 61557 3189 61566
rect 3619 61592 3677 61593
rect 2563 61551 2621 61552
rect 3619 61552 3628 61592
rect 3668 61552 3677 61592
rect 3619 61551 3677 61552
rect 4587 61592 4629 61601
rect 4587 61552 4588 61592
rect 4628 61552 4629 61592
rect 4587 61543 4629 61552
rect 4683 61592 4725 61601
rect 4683 61552 4684 61592
rect 4724 61552 4725 61592
rect 4683 61543 4725 61552
rect 6499 61592 6557 61593
rect 6499 61552 6508 61592
rect 6548 61552 6557 61592
rect 6499 61551 6557 61552
rect 7747 61592 7805 61593
rect 7747 61552 7756 61592
rect 7796 61552 7805 61592
rect 7747 61551 7805 61552
rect 8899 61592 8957 61593
rect 8899 61552 8908 61592
rect 8948 61552 8957 61592
rect 8899 61551 8957 61552
rect 10147 61592 10205 61593
rect 10147 61552 10156 61592
rect 10196 61552 10205 61592
rect 10147 61551 10205 61552
rect 11011 61592 11069 61593
rect 11011 61552 11020 61592
rect 11060 61552 11069 61592
rect 11011 61551 11069 61552
rect 12259 61592 12317 61593
rect 12259 61552 12268 61592
rect 12308 61552 12317 61592
rect 12259 61551 12317 61552
rect 13219 61592 13277 61593
rect 13219 61552 13228 61592
rect 13268 61552 13277 61592
rect 13219 61551 13277 61552
rect 14467 61592 14525 61593
rect 14467 61552 14476 61592
rect 14516 61552 14525 61592
rect 14467 61551 14525 61552
rect 16291 61592 16349 61593
rect 16291 61552 16300 61592
rect 16340 61552 16349 61592
rect 16291 61551 16349 61552
rect 17539 61592 17597 61593
rect 17539 61552 17548 61592
rect 17588 61552 17597 61592
rect 17539 61551 17597 61552
rect 18115 61592 18173 61593
rect 18115 61552 18124 61592
rect 18164 61552 18173 61592
rect 18115 61551 18173 61552
rect 19363 61592 19421 61593
rect 19363 61552 19372 61592
rect 19412 61552 19421 61592
rect 19363 61551 19421 61552
rect 2955 61508 2997 61517
rect 2955 61468 2956 61508
rect 2996 61468 2997 61508
rect 2955 61459 2997 61468
rect 2763 61424 2805 61433
rect 2763 61384 2764 61424
rect 2804 61384 2805 61424
rect 2763 61375 2805 61384
rect 7947 61424 7989 61433
rect 7947 61384 7948 61424
rect 7988 61384 7989 61424
rect 7947 61375 7989 61384
rect 10347 61424 10389 61433
rect 10347 61384 10348 61424
rect 10388 61384 10389 61424
rect 10347 61375 10389 61384
rect 12459 61424 12501 61433
rect 12459 61384 12460 61424
rect 12500 61384 12501 61424
rect 12459 61375 12501 61384
rect 15051 61424 15093 61433
rect 15051 61384 15052 61424
rect 15092 61384 15093 61424
rect 15051 61375 15093 61384
rect 17739 61424 17781 61433
rect 17739 61384 17740 61424
rect 17780 61384 17781 61424
rect 17739 61375 17781 61384
rect 19563 61424 19605 61433
rect 19563 61384 19564 61424
rect 19604 61384 19605 61424
rect 19563 61375 19605 61384
rect 19947 61424 19989 61433
rect 19947 61384 19948 61424
rect 19988 61384 19989 61424
rect 19947 61375 19989 61384
rect 1152 61256 20452 61280
rect 1152 61216 4928 61256
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 5296 61216 20048 61256
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20416 61216 20452 61256
rect 1152 61192 20452 61216
rect 14947 61088 15005 61089
rect 14947 61048 14956 61088
rect 14996 61048 15005 61088
rect 14947 61047 15005 61048
rect 15523 61088 15581 61089
rect 15523 61048 15532 61088
rect 15572 61048 15581 61088
rect 15523 61047 15581 61048
rect 10251 61004 10293 61013
rect 10251 60964 10252 61004
rect 10292 60964 10293 61004
rect 10251 60955 10293 60964
rect 12267 61004 12309 61013
rect 12267 60964 12268 61004
rect 12308 60964 12309 61004
rect 12267 60955 12309 60964
rect 16291 60962 16349 60963
rect 1891 60920 1949 60921
rect 1891 60880 1900 60920
rect 1940 60880 1949 60920
rect 1891 60879 1949 60880
rect 3139 60920 3197 60921
rect 3139 60880 3148 60920
rect 3188 60880 3197 60920
rect 3139 60879 3197 60880
rect 3523 60920 3581 60921
rect 3523 60880 3532 60920
rect 3572 60880 3581 60920
rect 3523 60879 3581 60880
rect 4771 60920 4829 60921
rect 4771 60880 4780 60920
rect 4820 60880 4829 60920
rect 4771 60879 4829 60880
rect 5155 60920 5213 60921
rect 5155 60880 5164 60920
rect 5204 60880 5213 60920
rect 5155 60879 5213 60880
rect 6403 60920 6461 60921
rect 6403 60880 6412 60920
rect 6452 60880 6461 60920
rect 6403 60879 6461 60880
rect 6883 60920 6941 60921
rect 6883 60880 6892 60920
rect 6932 60880 6941 60920
rect 6883 60879 6941 60880
rect 8131 60920 8189 60921
rect 8131 60880 8140 60920
rect 8180 60880 8189 60920
rect 8131 60879 8189 60880
rect 8803 60920 8861 60921
rect 8803 60880 8812 60920
rect 8852 60880 8861 60920
rect 8803 60879 8861 60880
rect 10051 60920 10109 60921
rect 10051 60880 10060 60920
rect 10100 60880 10109 60920
rect 10051 60879 10109 60880
rect 10539 60920 10581 60929
rect 10539 60880 10540 60920
rect 10580 60880 10581 60920
rect 10539 60871 10581 60880
rect 10635 60920 10677 60929
rect 10635 60880 10636 60920
rect 10676 60880 10677 60920
rect 10635 60871 10677 60880
rect 11115 60920 11157 60929
rect 11115 60880 11116 60920
rect 11156 60880 11157 60920
rect 11115 60871 11157 60880
rect 11587 60920 11645 60921
rect 11587 60880 11596 60920
rect 11636 60880 11645 60920
rect 11587 60879 11645 60880
rect 12075 60915 12117 60924
rect 12075 60875 12076 60915
rect 12116 60875 12117 60915
rect 12835 60920 12893 60921
rect 12835 60880 12844 60920
rect 12884 60880 12893 60920
rect 12835 60879 12893 60880
rect 14083 60920 14141 60921
rect 14083 60880 14092 60920
rect 14132 60880 14141 60920
rect 14083 60879 14141 60880
rect 14467 60920 14525 60921
rect 14467 60880 14476 60920
rect 14516 60880 14525 60920
rect 14467 60879 14525 60880
rect 14563 60920 14621 60921
rect 14563 60880 14572 60920
rect 14612 60880 14621 60920
rect 14563 60879 14621 60880
rect 14763 60920 14805 60929
rect 14763 60880 14764 60920
rect 14804 60880 14805 60920
rect 12075 60866 12117 60875
rect 14763 60871 14805 60880
rect 14859 60920 14901 60929
rect 14859 60880 14860 60920
rect 14900 60880 14901 60920
rect 15243 60920 15285 60929
rect 14859 60871 14901 60880
rect 15016 60905 15058 60914
rect 15016 60865 15017 60905
rect 15057 60865 15058 60905
rect 15243 60880 15244 60920
rect 15284 60880 15285 60920
rect 15243 60871 15285 60880
rect 15339 60920 15381 60929
rect 16291 60922 16300 60962
rect 16340 60922 16349 60962
rect 16291 60921 16349 60922
rect 15339 60880 15340 60920
rect 15380 60880 15381 60920
rect 15339 60871 15381 60880
rect 17539 60920 17597 60921
rect 17539 60880 17548 60920
rect 17588 60880 17597 60920
rect 17539 60879 17597 60880
rect 18115 60920 18173 60921
rect 18115 60880 18124 60920
rect 18164 60880 18173 60920
rect 18115 60879 18173 60880
rect 19363 60920 19421 60921
rect 19363 60880 19372 60920
rect 19412 60880 19421 60920
rect 19363 60879 19421 60880
rect 15016 60856 15058 60865
rect 1699 60836 1757 60837
rect 1699 60796 1708 60836
rect 1748 60796 1757 60836
rect 1699 60795 1757 60796
rect 11019 60836 11061 60845
rect 11019 60796 11020 60836
rect 11060 60796 11061 60836
rect 11019 60787 11061 60796
rect 20035 60836 20093 60837
rect 20035 60796 20044 60836
rect 20084 60796 20093 60836
rect 20035 60795 20093 60796
rect 1515 60668 1557 60677
rect 1515 60628 1516 60668
rect 1556 60628 1557 60668
rect 1515 60619 1557 60628
rect 3339 60668 3381 60677
rect 3339 60628 3340 60668
rect 3380 60628 3381 60668
rect 3339 60619 3381 60628
rect 4971 60668 5013 60677
rect 4971 60628 4972 60668
rect 5012 60628 5013 60668
rect 4971 60619 5013 60628
rect 6603 60668 6645 60677
rect 6603 60628 6604 60668
rect 6644 60628 6645 60668
rect 6603 60619 6645 60628
rect 8331 60668 8373 60677
rect 8331 60628 8332 60668
rect 8372 60628 8373 60668
rect 8331 60619 8373 60628
rect 14283 60668 14325 60677
rect 14283 60628 14284 60668
rect 14324 60628 14325 60668
rect 14283 60619 14325 60628
rect 17739 60668 17781 60677
rect 17739 60628 17740 60668
rect 17780 60628 17781 60668
rect 17739 60619 17781 60628
rect 19563 60668 19605 60677
rect 19563 60628 19564 60668
rect 19604 60628 19605 60668
rect 19563 60619 19605 60628
rect 20235 60668 20277 60677
rect 20235 60628 20236 60668
rect 20276 60628 20277 60668
rect 20235 60619 20277 60628
rect 1152 60500 20352 60524
rect 1152 60460 3688 60500
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 4056 60460 18808 60500
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 19176 60460 20352 60500
rect 1152 60436 20352 60460
rect 2955 60332 2997 60341
rect 2955 60292 2956 60332
rect 2996 60292 2997 60332
rect 2955 60283 2997 60292
rect 14091 60332 14133 60341
rect 14091 60292 14092 60332
rect 14132 60292 14133 60332
rect 14091 60283 14133 60292
rect 17163 60332 17205 60341
rect 17163 60292 17164 60332
rect 17204 60292 17205 60332
rect 17163 60283 17205 60292
rect 17547 60332 17589 60341
rect 17547 60292 17548 60332
rect 17588 60292 17589 60332
rect 17547 60283 17589 60292
rect 7083 60164 7125 60173
rect 7083 60124 7084 60164
rect 7124 60124 7125 60164
rect 7083 60115 7125 60124
rect 7179 60164 7221 60173
rect 7179 60124 7180 60164
rect 7220 60124 7221 60164
rect 11019 60164 11061 60173
rect 7179 60115 7221 60124
rect 8187 60122 8229 60131
rect 4779 60094 4821 60103
rect 1507 60080 1565 60081
rect 1507 60040 1516 60080
rect 1556 60040 1565 60080
rect 1507 60039 1565 60040
rect 2755 60080 2813 60081
rect 2755 60040 2764 60080
rect 2804 60040 2813 60080
rect 2755 60039 2813 60040
rect 3243 60080 3285 60089
rect 3243 60040 3244 60080
rect 3284 60040 3285 60080
rect 3243 60031 3285 60040
rect 3339 60080 3381 60089
rect 3339 60040 3340 60080
rect 3380 60040 3381 60080
rect 3339 60031 3381 60040
rect 3723 60080 3765 60089
rect 3723 60040 3724 60080
rect 3764 60040 3765 60080
rect 3723 60031 3765 60040
rect 3819 60080 3861 60089
rect 3819 60040 3820 60080
rect 3860 60040 3861 60080
rect 3819 60031 3861 60040
rect 4291 60080 4349 60081
rect 4291 60040 4300 60080
rect 4340 60040 4349 60080
rect 4779 60054 4780 60094
rect 4820 60054 4821 60094
rect 4779 60045 4821 60054
rect 6603 60080 6645 60089
rect 4291 60039 4349 60040
rect 6603 60040 6604 60080
rect 6644 60040 6645 60080
rect 6603 60031 6645 60040
rect 6699 60080 6741 60089
rect 8187 60082 8188 60122
rect 8228 60082 8229 60122
rect 11019 60124 11020 60164
rect 11060 60124 11061 60164
rect 11019 60115 11061 60124
rect 11115 60164 11157 60173
rect 11115 60124 11116 60164
rect 11156 60124 11157 60164
rect 16579 60164 16637 60165
rect 11115 60115 11157 60124
rect 12123 60122 12165 60131
rect 16579 60124 16588 60164
rect 16628 60124 16637 60164
rect 16579 60123 16637 60124
rect 16963 60164 17021 60165
rect 16963 60124 16972 60164
rect 17012 60124 17021 60164
rect 16963 60123 17021 60124
rect 17347 60164 17405 60165
rect 17347 60124 17356 60164
rect 17396 60124 17405 60164
rect 17347 60123 17405 60124
rect 18315 60164 18357 60173
rect 18315 60124 18316 60164
rect 18356 60124 18357 60164
rect 6699 60040 6700 60080
rect 6740 60040 6741 60080
rect 6699 60031 6741 60040
rect 7651 60080 7709 60081
rect 7651 60040 7660 60080
rect 7700 60040 7709 60080
rect 8187 60073 8229 60082
rect 10539 60080 10581 60089
rect 7651 60039 7709 60040
rect 10539 60040 10540 60080
rect 10580 60040 10581 60080
rect 10539 60031 10581 60040
rect 10635 60080 10677 60089
rect 12123 60082 12124 60122
rect 12164 60082 12165 60122
rect 18315 60115 18357 60124
rect 18411 60164 18453 60173
rect 18411 60124 18412 60164
rect 18452 60124 18453 60164
rect 19747 60164 19805 60165
rect 18411 60115 18453 60124
rect 19419 60122 19461 60131
rect 19747 60124 19756 60164
rect 19796 60124 19805 60164
rect 19747 60123 19805 60124
rect 10635 60040 10636 60080
rect 10676 60040 10677 60080
rect 10635 60031 10677 60040
rect 11587 60080 11645 60081
rect 11587 60040 11596 60080
rect 11636 60040 11645 60080
rect 12123 60073 12165 60082
rect 12643 60080 12701 60081
rect 11587 60039 11645 60040
rect 12643 60040 12652 60080
rect 12692 60040 12701 60080
rect 12643 60039 12701 60040
rect 13891 60080 13949 60081
rect 13891 60040 13900 60080
rect 13940 60040 13949 60080
rect 13891 60039 13949 60040
rect 14379 60080 14421 60089
rect 14379 60040 14380 60080
rect 14420 60040 14421 60080
rect 14379 60031 14421 60040
rect 14475 60080 14517 60089
rect 14475 60040 14476 60080
rect 14516 60040 14517 60080
rect 14475 60031 14517 60040
rect 14859 60080 14901 60089
rect 14859 60040 14860 60080
rect 14900 60040 14901 60080
rect 14859 60031 14901 60040
rect 14955 60080 14997 60089
rect 15915 60085 15957 60094
rect 14955 60040 14956 60080
rect 14996 60040 14997 60080
rect 14955 60031 14997 60040
rect 15427 60080 15485 60081
rect 15427 60040 15436 60080
rect 15476 60040 15485 60080
rect 15427 60039 15485 60040
rect 15915 60045 15916 60085
rect 15956 60045 15957 60085
rect 15915 60036 15957 60045
rect 17835 60080 17877 60089
rect 17835 60040 17836 60080
rect 17876 60040 17877 60080
rect 17835 60031 17877 60040
rect 17931 60080 17973 60089
rect 19419 60082 19420 60122
rect 19460 60082 19461 60122
rect 17931 60040 17932 60080
rect 17972 60040 17973 60080
rect 17931 60031 17973 60040
rect 18883 60080 18941 60081
rect 18883 60040 18892 60080
rect 18932 60040 18941 60080
rect 19419 60073 19461 60082
rect 18883 60039 18941 60040
rect 8331 59996 8373 60005
rect 8331 59956 8332 59996
rect 8372 59956 8373 59996
rect 8331 59947 8373 59956
rect 12267 59996 12309 60005
rect 12267 59956 12268 59996
rect 12308 59956 12309 59996
rect 12267 59947 12309 59956
rect 4971 59912 5013 59921
rect 4971 59872 4972 59912
rect 5012 59872 5013 59912
rect 4971 59863 5013 59872
rect 14091 59912 14133 59921
rect 14091 59872 14092 59912
rect 14132 59872 14133 59912
rect 14091 59863 14133 59872
rect 16107 59912 16149 59921
rect 16107 59872 16108 59912
rect 16148 59872 16149 59912
rect 16107 59863 16149 59872
rect 16779 59912 16821 59921
rect 16779 59872 16780 59912
rect 16820 59872 16821 59912
rect 16779 59863 16821 59872
rect 19563 59912 19605 59921
rect 19563 59872 19564 59912
rect 19604 59872 19605 59912
rect 19563 59863 19605 59872
rect 19947 59912 19989 59921
rect 19947 59872 19948 59912
rect 19988 59872 19989 59912
rect 19947 59863 19989 59872
rect 1152 59744 20452 59768
rect 1152 59704 4928 59744
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 5296 59704 20048 59744
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20416 59704 20452 59744
rect 1152 59680 20452 59704
rect 12747 59576 12789 59585
rect 12747 59536 12748 59576
rect 12788 59536 12789 59576
rect 12747 59527 12789 59536
rect 13035 59576 13077 59585
rect 13035 59536 13036 59576
rect 13076 59536 13077 59576
rect 13035 59527 13077 59536
rect 14763 59576 14805 59585
rect 14763 59536 14764 59576
rect 14804 59536 14805 59576
rect 14763 59527 14805 59536
rect 16395 59576 16437 59585
rect 16395 59536 16396 59576
rect 16436 59536 16437 59576
rect 16395 59527 16437 59536
rect 2955 59492 2997 59501
rect 2955 59452 2956 59492
rect 2996 59452 2997 59492
rect 2955 59443 2997 59452
rect 8043 59492 8085 59501
rect 8043 59452 8044 59492
rect 8084 59452 8085 59492
rect 8043 59443 8085 59452
rect 9771 59492 9813 59501
rect 9771 59452 9772 59492
rect 9812 59452 9813 59492
rect 9771 59443 9813 59452
rect 11787 59492 11829 59501
rect 11787 59452 11788 59492
rect 11828 59452 11829 59492
rect 11787 59443 11829 59452
rect 19563 59492 19605 59501
rect 19563 59452 19564 59492
rect 19604 59452 19605 59492
rect 19563 59443 19605 59452
rect 1219 59408 1277 59409
rect 1219 59368 1228 59408
rect 1268 59368 1277 59408
rect 1219 59367 1277 59368
rect 2467 59408 2525 59409
rect 2467 59368 2476 59408
rect 2516 59368 2525 59408
rect 2467 59367 2525 59368
rect 3147 59403 3189 59412
rect 3147 59363 3148 59403
rect 3188 59363 3189 59403
rect 3619 59408 3677 59409
rect 3619 59368 3628 59408
rect 3668 59368 3677 59408
rect 3619 59367 3677 59368
rect 4107 59408 4149 59417
rect 4107 59368 4108 59408
rect 4148 59368 4149 59408
rect 3147 59354 3189 59363
rect 4107 59359 4149 59368
rect 4587 59408 4629 59417
rect 4587 59368 4588 59408
rect 4628 59368 4629 59408
rect 4587 59359 4629 59368
rect 4683 59408 4725 59417
rect 4683 59368 4684 59408
rect 4724 59368 4725 59408
rect 4683 59359 4725 59368
rect 6315 59408 6357 59417
rect 6315 59368 6316 59408
rect 6356 59368 6357 59408
rect 6315 59359 6357 59368
rect 6411 59408 6453 59417
rect 6411 59368 6412 59408
rect 6452 59368 6453 59408
rect 6411 59359 6453 59368
rect 6891 59408 6933 59417
rect 6891 59368 6892 59408
rect 6932 59368 6933 59408
rect 6891 59359 6933 59368
rect 7363 59408 7421 59409
rect 7363 59368 7372 59408
rect 7412 59368 7421 59408
rect 7363 59367 7421 59368
rect 7851 59403 7893 59412
rect 7851 59363 7852 59403
rect 7892 59363 7893 59403
rect 8323 59408 8381 59409
rect 8323 59368 8332 59408
rect 8372 59368 8381 59408
rect 8323 59367 8381 59368
rect 9571 59408 9629 59409
rect 9571 59368 9580 59408
rect 9620 59368 9629 59408
rect 9571 59367 9629 59368
rect 10059 59408 10101 59417
rect 10059 59368 10060 59408
rect 10100 59368 10101 59408
rect 7851 59354 7893 59363
rect 10059 59359 10101 59368
rect 10155 59408 10197 59417
rect 10155 59368 10156 59408
rect 10196 59368 10197 59408
rect 10155 59359 10197 59368
rect 10539 59408 10581 59417
rect 10539 59368 10540 59408
rect 10580 59368 10581 59408
rect 10539 59359 10581 59368
rect 10635 59408 10677 59417
rect 10635 59368 10636 59408
rect 10676 59368 10677 59408
rect 10635 59359 10677 59368
rect 11107 59408 11165 59409
rect 11107 59368 11116 59408
rect 11156 59368 11165 59408
rect 12555 59408 12597 59417
rect 11107 59367 11165 59368
rect 11595 59394 11637 59403
rect 11595 59354 11596 59394
rect 11636 59354 11637 59394
rect 12555 59368 12556 59408
rect 12596 59368 12597 59408
rect 12555 59359 12597 59368
rect 12651 59408 12693 59417
rect 12651 59368 12652 59408
rect 12692 59368 12693 59408
rect 12651 59359 12693 59368
rect 12843 59408 12885 59417
rect 12843 59368 12844 59408
rect 12884 59368 12885 59408
rect 12843 59359 12885 59368
rect 13219 59408 13277 59409
rect 13219 59368 13228 59408
rect 13268 59368 13277 59408
rect 13219 59367 13277 59368
rect 14467 59408 14525 59409
rect 14467 59368 14476 59408
rect 14516 59368 14525 59408
rect 14467 59367 14525 59368
rect 14659 59408 14717 59409
rect 14659 59368 14668 59408
rect 14708 59368 14717 59408
rect 14659 59367 14717 59368
rect 14947 59408 15005 59409
rect 14947 59368 14956 59408
rect 14996 59368 15005 59408
rect 14947 59367 15005 59368
rect 16195 59408 16253 59409
rect 16195 59368 16204 59408
rect 16244 59368 16253 59408
rect 16195 59367 16253 59368
rect 17835 59408 17877 59417
rect 17835 59368 17836 59408
rect 17876 59368 17877 59408
rect 17835 59359 17877 59368
rect 17931 59408 17973 59417
rect 17931 59368 17932 59408
rect 17972 59368 17973 59408
rect 17931 59359 17973 59368
rect 18315 59408 18357 59417
rect 18315 59368 18316 59408
rect 18356 59368 18357 59408
rect 18315 59359 18357 59368
rect 18411 59408 18453 59417
rect 18411 59368 18412 59408
rect 18452 59368 18453 59408
rect 18411 59359 18453 59368
rect 18883 59408 18941 59409
rect 18883 59368 18892 59408
rect 18932 59368 18941 59408
rect 18883 59367 18941 59368
rect 19419 59398 19461 59407
rect 11595 59345 11637 59354
rect 19419 59358 19420 59398
rect 19460 59358 19461 59398
rect 19419 59349 19461 59358
rect 4203 59324 4245 59333
rect 4203 59284 4204 59324
rect 4244 59284 4245 59324
rect 4203 59275 4245 59284
rect 5155 59324 5213 59325
rect 5155 59284 5164 59324
rect 5204 59284 5213 59324
rect 5155 59283 5213 59284
rect 6795 59324 6837 59333
rect 6795 59284 6796 59324
rect 6836 59284 6837 59324
rect 6795 59275 6837 59284
rect 16963 59324 17021 59325
rect 16963 59284 16972 59324
rect 17012 59284 17021 59324
rect 16963 59283 17021 59284
rect 17347 59324 17405 59325
rect 17347 59284 17356 59324
rect 17396 59284 17405 59324
rect 17347 59283 17405 59284
rect 19747 59324 19805 59325
rect 19747 59284 19756 59324
rect 19796 59284 19805 59324
rect 19747 59283 19805 59284
rect 4971 59240 5013 59249
rect 4971 59200 4972 59240
rect 5012 59200 5013 59240
rect 4971 59191 5013 59200
rect 17163 59240 17205 59249
rect 17163 59200 17164 59240
rect 17204 59200 17205 59240
rect 17163 59191 17205 59200
rect 2667 59156 2709 59165
rect 2667 59116 2668 59156
rect 2708 59116 2709 59156
rect 2667 59107 2709 59116
rect 17547 59156 17589 59165
rect 17547 59116 17548 59156
rect 17588 59116 17589 59156
rect 17547 59107 17589 59116
rect 19947 59156 19989 59165
rect 19947 59116 19948 59156
rect 19988 59116 19989 59156
rect 19947 59107 19989 59116
rect 1152 58988 20352 59012
rect 1152 58948 3688 58988
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 4056 58948 18808 58988
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 19176 58948 20352 58988
rect 1152 58924 20352 58948
rect 11499 58820 11541 58829
rect 11499 58780 11500 58820
rect 11540 58780 11541 58820
rect 11499 58771 11541 58780
rect 9859 58652 9917 58653
rect 9859 58612 9868 58652
rect 9908 58612 9917 58652
rect 9859 58611 9917 58612
rect 12931 58652 12989 58653
rect 12931 58612 12940 58652
rect 12980 58612 12989 58652
rect 12931 58611 12989 58612
rect 17251 58652 17309 58653
rect 17251 58612 17260 58652
rect 17300 58612 17309 58652
rect 17251 58611 17309 58612
rect 17635 58652 17693 58653
rect 17635 58612 17644 58652
rect 17684 58612 17693 58652
rect 17635 58611 17693 58612
rect 19651 58652 19709 58653
rect 19651 58612 19660 58652
rect 19700 58612 19709 58652
rect 19651 58611 19709 58612
rect 20035 58652 20093 58653
rect 20035 58612 20044 58652
rect 20084 58612 20093 58652
rect 20035 58611 20093 58612
rect 1411 58568 1469 58569
rect 1411 58528 1420 58568
rect 1460 58528 1469 58568
rect 1411 58527 1469 58528
rect 2659 58568 2717 58569
rect 2659 58528 2668 58568
rect 2708 58528 2717 58568
rect 2659 58527 2717 58528
rect 3043 58568 3101 58569
rect 3043 58528 3052 58568
rect 3092 58528 3101 58568
rect 3043 58527 3101 58528
rect 4291 58568 4349 58569
rect 4291 58528 4300 58568
rect 4340 58528 4349 58568
rect 4291 58527 4349 58528
rect 4675 58568 4733 58569
rect 4675 58528 4684 58568
rect 4724 58528 4733 58568
rect 4675 58527 4733 58528
rect 5923 58568 5981 58569
rect 5923 58528 5932 58568
rect 5972 58528 5981 58568
rect 5923 58527 5981 58528
rect 6307 58568 6365 58569
rect 6307 58528 6316 58568
rect 6356 58528 6365 58568
rect 6307 58527 6365 58528
rect 7555 58568 7613 58569
rect 7555 58528 7564 58568
rect 7604 58528 7613 58568
rect 7555 58527 7613 58528
rect 8035 58568 8093 58569
rect 8035 58528 8044 58568
rect 8084 58528 8093 58568
rect 8035 58527 8093 58528
rect 9283 58568 9341 58569
rect 9283 58528 9292 58568
rect 9332 58528 9341 58568
rect 9283 58527 9341 58528
rect 10051 58568 10109 58569
rect 10051 58528 10060 58568
rect 10100 58528 10109 58568
rect 10051 58527 10109 58528
rect 11299 58568 11357 58569
rect 11299 58528 11308 58568
rect 11348 58528 11357 58568
rect 11299 58527 11357 58528
rect 13699 58568 13757 58569
rect 13699 58528 13708 58568
rect 13748 58528 13757 58568
rect 13699 58527 13757 58528
rect 14947 58568 15005 58569
rect 14947 58528 14956 58568
rect 14996 58528 15005 58568
rect 14947 58527 15005 58528
rect 15331 58568 15389 58569
rect 15331 58528 15340 58568
rect 15380 58528 15389 58568
rect 15331 58527 15389 58528
rect 16579 58568 16637 58569
rect 16579 58528 16588 58568
rect 16628 58528 16637 58568
rect 16579 58527 16637 58528
rect 18019 58568 18077 58569
rect 18019 58528 18028 58568
rect 18068 58528 18077 58568
rect 18019 58527 18077 58528
rect 19267 58568 19325 58569
rect 19267 58528 19276 58568
rect 19316 58528 19325 58568
rect 19267 58527 19325 58528
rect 2859 58400 2901 58409
rect 2859 58360 2860 58400
rect 2900 58360 2901 58400
rect 2859 58351 2901 58360
rect 4491 58400 4533 58409
rect 4491 58360 4492 58400
rect 4532 58360 4533 58400
rect 4491 58351 4533 58360
rect 6123 58400 6165 58409
rect 6123 58360 6124 58400
rect 6164 58360 6165 58400
rect 6123 58351 6165 58360
rect 7755 58400 7797 58409
rect 7755 58360 7756 58400
rect 7796 58360 7797 58400
rect 7755 58351 7797 58360
rect 9483 58400 9525 58409
rect 9483 58360 9484 58400
rect 9524 58360 9525 58400
rect 9483 58351 9525 58360
rect 9675 58400 9717 58409
rect 9675 58360 9676 58400
rect 9716 58360 9717 58400
rect 9675 58351 9717 58360
rect 12747 58400 12789 58409
rect 12747 58360 12748 58400
rect 12788 58360 12789 58400
rect 12747 58351 12789 58360
rect 15147 58400 15189 58409
rect 15147 58360 15148 58400
rect 15188 58360 15189 58400
rect 15147 58351 15189 58360
rect 16779 58400 16821 58409
rect 16779 58360 16780 58400
rect 16820 58360 16821 58400
rect 16779 58351 16821 58360
rect 17451 58400 17493 58409
rect 17451 58360 17452 58400
rect 17492 58360 17493 58400
rect 17451 58351 17493 58360
rect 17835 58400 17877 58409
rect 17835 58360 17836 58400
rect 17876 58360 17877 58400
rect 17835 58351 17877 58360
rect 19467 58400 19509 58409
rect 19467 58360 19468 58400
rect 19508 58360 19509 58400
rect 19467 58351 19509 58360
rect 19851 58400 19893 58409
rect 19851 58360 19852 58400
rect 19892 58360 19893 58400
rect 19851 58351 19893 58360
rect 20235 58400 20277 58409
rect 20235 58360 20236 58400
rect 20276 58360 20277 58400
rect 20235 58351 20277 58360
rect 1152 58232 20452 58256
rect 1152 58192 4928 58232
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 5296 58192 20048 58232
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20416 58192 20452 58232
rect 1152 58168 20452 58192
rect 9675 58064 9717 58073
rect 9675 58024 9676 58064
rect 9716 58024 9717 58064
rect 9675 58015 9717 58024
rect 3147 57980 3189 57989
rect 3147 57940 3148 57980
rect 3188 57940 3189 57980
rect 3147 57931 3189 57940
rect 5259 57980 5301 57989
rect 5259 57940 5260 57980
rect 5300 57940 5301 57980
rect 5259 57931 5301 57940
rect 1699 57896 1757 57897
rect 1699 57856 1708 57896
rect 1748 57856 1757 57896
rect 1699 57855 1757 57856
rect 2947 57896 3005 57897
rect 2947 57856 2956 57896
rect 2996 57856 3005 57896
rect 2947 57855 3005 57856
rect 3531 57896 3573 57905
rect 3531 57856 3532 57896
rect 3572 57856 3573 57896
rect 3531 57847 3573 57856
rect 3627 57896 3669 57905
rect 3627 57856 3628 57896
rect 3668 57856 3669 57896
rect 3627 57847 3669 57856
rect 4011 57896 4053 57905
rect 4011 57856 4012 57896
rect 4052 57856 4053 57896
rect 4011 57847 4053 57856
rect 4107 57896 4149 57905
rect 4107 57856 4108 57896
rect 4148 57856 4149 57896
rect 4107 57847 4149 57856
rect 4579 57896 4637 57897
rect 4579 57856 4588 57896
rect 4628 57856 4637 57896
rect 4579 57855 4637 57856
rect 5067 57891 5109 57900
rect 5067 57851 5068 57891
rect 5108 57851 5109 57891
rect 6211 57896 6269 57897
rect 6211 57856 6220 57896
rect 6260 57856 6269 57896
rect 6211 57855 6269 57856
rect 7459 57896 7517 57897
rect 7459 57856 7468 57896
rect 7508 57856 7517 57896
rect 7459 57855 7517 57856
rect 7947 57896 7989 57905
rect 7947 57856 7948 57896
rect 7988 57856 7989 57896
rect 5067 57842 5109 57851
rect 7947 57847 7989 57856
rect 8043 57896 8085 57905
rect 8043 57856 8044 57896
rect 8084 57856 8085 57896
rect 8043 57847 8085 57856
rect 8427 57896 8469 57905
rect 8427 57856 8428 57896
rect 8468 57856 8469 57896
rect 8427 57847 8469 57856
rect 8523 57896 8565 57905
rect 8523 57856 8524 57896
rect 8564 57856 8565 57896
rect 8523 57847 8565 57856
rect 8995 57896 9053 57897
rect 8995 57856 9004 57896
rect 9044 57856 9053 57896
rect 8995 57855 9053 57856
rect 9483 57891 9525 57900
rect 9483 57851 9484 57891
rect 9524 57851 9525 57891
rect 10147 57896 10205 57897
rect 10147 57856 10156 57896
rect 10196 57856 10205 57896
rect 10147 57855 10205 57856
rect 11395 57896 11453 57897
rect 11395 57856 11404 57896
rect 11444 57856 11453 57896
rect 11395 57855 11453 57856
rect 11875 57896 11933 57897
rect 11875 57856 11884 57896
rect 11924 57856 11933 57896
rect 11875 57855 11933 57856
rect 13123 57896 13181 57897
rect 13123 57856 13132 57896
rect 13172 57856 13181 57896
rect 13123 57855 13181 57856
rect 14083 57896 14141 57897
rect 14083 57856 14092 57896
rect 14132 57856 14141 57896
rect 14083 57855 14141 57856
rect 15331 57896 15389 57897
rect 15331 57856 15340 57896
rect 15380 57856 15389 57896
rect 15331 57855 15389 57856
rect 15715 57896 15773 57897
rect 15715 57856 15724 57896
rect 15764 57856 15773 57896
rect 15715 57855 15773 57856
rect 16963 57896 17021 57897
rect 16963 57856 16972 57896
rect 17012 57856 17021 57896
rect 16963 57855 17021 57856
rect 17539 57896 17597 57897
rect 17539 57856 17548 57896
rect 17588 57856 17597 57896
rect 17539 57855 17597 57856
rect 18787 57896 18845 57897
rect 18787 57856 18796 57896
rect 18836 57856 18845 57896
rect 18787 57855 18845 57856
rect 19075 57896 19133 57897
rect 19075 57856 19084 57896
rect 19124 57856 19133 57896
rect 19075 57855 19133 57856
rect 9483 57842 9525 57851
rect 1507 57812 1565 57813
rect 1507 57772 1516 57812
rect 1556 57772 1565 57812
rect 1507 57771 1565 57772
rect 1323 57728 1365 57737
rect 1323 57688 1324 57728
rect 1364 57688 1365 57728
rect 1323 57679 1365 57688
rect 7659 57644 7701 57653
rect 7659 57604 7660 57644
rect 7700 57604 7701 57644
rect 7659 57595 7701 57604
rect 11595 57644 11637 57653
rect 11595 57604 11596 57644
rect 11636 57604 11637 57644
rect 11595 57595 11637 57604
rect 13323 57644 13365 57653
rect 13323 57604 13324 57644
rect 13364 57604 13365 57644
rect 13323 57595 13365 57604
rect 15531 57644 15573 57653
rect 15531 57604 15532 57644
rect 15572 57604 15573 57644
rect 15531 57595 15573 57604
rect 17163 57644 17205 57653
rect 17163 57604 17164 57644
rect 17204 57604 17205 57644
rect 17163 57595 17205 57604
rect 17355 57644 17397 57653
rect 17355 57604 17356 57644
rect 17396 57604 17397 57644
rect 17355 57595 17397 57604
rect 19563 57644 19605 57653
rect 19563 57604 19564 57644
rect 19604 57604 19605 57644
rect 19563 57595 19605 57604
rect 1152 57476 20352 57500
rect 1152 57436 3688 57476
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 4056 57436 18808 57476
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 19176 57436 20352 57476
rect 1152 57412 20352 57436
rect 1699 57140 1757 57141
rect 1699 57100 1708 57140
rect 1748 57100 1757 57140
rect 1699 57099 1757 57100
rect 2083 57140 2141 57141
rect 2083 57100 2092 57140
rect 2132 57100 2141 57140
rect 2083 57099 2141 57100
rect 3531 57140 3573 57149
rect 3531 57100 3532 57140
rect 3572 57100 3573 57140
rect 3531 57091 3573 57100
rect 3627 57140 3669 57149
rect 3627 57100 3628 57140
rect 3668 57100 3669 57140
rect 3627 57091 3669 57100
rect 11979 57140 12021 57149
rect 11979 57100 11980 57140
rect 12020 57100 12021 57140
rect 14091 57140 14133 57149
rect 11979 57091 12021 57100
rect 13083 57098 13125 57107
rect 2571 57070 2613 57079
rect 2571 57030 2572 57070
rect 2612 57030 2613 57070
rect 7755 57070 7797 57079
rect 2571 57021 2613 57030
rect 3043 57056 3101 57057
rect 3043 57016 3052 57056
rect 3092 57016 3101 57056
rect 3043 57015 3101 57016
rect 4011 57056 4053 57065
rect 4011 57016 4012 57056
rect 4052 57016 4053 57056
rect 4011 57007 4053 57016
rect 4107 57056 4149 57065
rect 4107 57016 4108 57056
rect 4148 57016 4149 57056
rect 4107 57007 4149 57016
rect 4387 57056 4445 57057
rect 4387 57016 4396 57056
rect 4436 57016 4445 57056
rect 4387 57015 4445 57016
rect 5635 57056 5693 57057
rect 5635 57016 5644 57056
rect 5684 57016 5693 57056
rect 5635 57015 5693 57016
rect 6219 57056 6261 57065
rect 6219 57016 6220 57056
rect 6260 57016 6261 57056
rect 6219 57007 6261 57016
rect 6315 57056 6357 57065
rect 6315 57016 6316 57056
rect 6356 57016 6357 57056
rect 6315 57007 6357 57016
rect 6699 57056 6741 57065
rect 6699 57016 6700 57056
rect 6740 57016 6741 57056
rect 6699 57007 6741 57016
rect 6795 57056 6837 57065
rect 6795 57016 6796 57056
rect 6836 57016 6837 57056
rect 6795 57007 6837 57016
rect 7267 57056 7325 57057
rect 7267 57016 7276 57056
rect 7316 57016 7325 57056
rect 7755 57030 7756 57070
rect 7796 57030 7797 57070
rect 11499 57075 11541 57084
rect 7755 57021 7797 57030
rect 8131 57056 8189 57057
rect 7267 57015 7325 57016
rect 8131 57016 8140 57056
rect 8180 57016 8189 57056
rect 8131 57015 8189 57016
rect 9379 57056 9437 57057
rect 9379 57016 9388 57056
rect 9428 57016 9437 57056
rect 9379 57015 9437 57016
rect 9763 57056 9821 57057
rect 9763 57016 9772 57056
rect 9812 57016 9821 57056
rect 9763 57015 9821 57016
rect 11011 57056 11069 57057
rect 11011 57016 11020 57056
rect 11060 57016 11069 57056
rect 11499 57035 11500 57075
rect 11540 57035 11541 57075
rect 11499 57026 11541 57035
rect 11595 57056 11637 57065
rect 11011 57015 11069 57016
rect 11595 57016 11596 57056
rect 11636 57016 11637 57056
rect 11595 57007 11637 57016
rect 12075 57056 12117 57065
rect 13083 57058 13084 57098
rect 13124 57058 13125 57098
rect 14091 57100 14092 57140
rect 14132 57100 14133 57140
rect 14091 57091 14133 57100
rect 16011 57140 16053 57149
rect 16011 57100 16012 57140
rect 16052 57100 16053 57140
rect 16011 57091 16053 57100
rect 19747 57140 19805 57141
rect 19747 57100 19756 57140
rect 19796 57100 19805 57140
rect 19747 57099 19805 57100
rect 15051 57065 15093 57074
rect 19371 57070 19413 57079
rect 12075 57016 12076 57056
rect 12116 57016 12117 57056
rect 12075 57007 12117 57016
rect 12547 57056 12605 57057
rect 12547 57016 12556 57056
rect 12596 57016 12605 57056
rect 13083 57049 13125 57058
rect 13515 57056 13557 57065
rect 12547 57015 12605 57016
rect 13515 57016 13516 57056
rect 13556 57016 13557 57056
rect 13515 57007 13557 57016
rect 13611 57056 13653 57065
rect 13611 57016 13612 57056
rect 13652 57016 13653 57056
rect 13611 57007 13653 57016
rect 13995 57056 14037 57065
rect 13995 57016 13996 57056
rect 14036 57016 14037 57056
rect 13995 57007 14037 57016
rect 14563 57056 14621 57057
rect 14563 57016 14572 57056
rect 14612 57016 14621 57056
rect 15051 57025 15052 57065
rect 15092 57025 15093 57065
rect 15051 57016 15093 57025
rect 15619 57056 15677 57057
rect 15619 57016 15628 57056
rect 15668 57016 15677 57056
rect 14563 57015 14621 57016
rect 15619 57015 15677 57016
rect 15723 57056 15765 57065
rect 15723 57016 15724 57056
rect 15764 57016 15765 57056
rect 15723 57007 15765 57016
rect 15915 57056 15957 57065
rect 15915 57016 15916 57056
rect 15956 57016 15957 57056
rect 15915 57007 15957 57016
rect 16203 57056 16245 57065
rect 16203 57016 16204 57056
rect 16244 57016 16245 57056
rect 16203 57007 16245 57016
rect 16387 57056 16445 57057
rect 16387 57016 16396 57056
rect 16436 57016 16445 57056
rect 16387 57015 16445 57016
rect 16491 57056 16533 57065
rect 16491 57016 16492 57056
rect 16532 57016 16533 57056
rect 16491 57007 16533 57016
rect 16683 57056 16725 57065
rect 16683 57016 16684 57056
rect 16724 57016 16725 57056
rect 16683 57007 16725 57016
rect 16875 57056 16917 57065
rect 16875 57016 16876 57056
rect 16916 57016 16917 57056
rect 16875 57007 16917 57016
rect 16971 57056 17013 57065
rect 16971 57016 16972 57056
rect 17012 57016 17013 57056
rect 16971 57007 17013 57016
rect 17067 57056 17109 57065
rect 17067 57016 17068 57056
rect 17108 57016 17109 57056
rect 17067 57007 17109 57016
rect 17355 57056 17397 57065
rect 17355 57016 17356 57056
rect 17396 57016 17397 57056
rect 17355 57007 17397 57016
rect 17547 57056 17589 57065
rect 17547 57016 17548 57056
rect 17588 57016 17589 57056
rect 17547 57007 17589 57016
rect 17835 57056 17877 57065
rect 17835 57016 17836 57056
rect 17876 57016 17877 57056
rect 17835 57007 17877 57016
rect 17931 57056 17973 57065
rect 17931 57016 17932 57056
rect 17972 57016 17973 57056
rect 17931 57007 17973 57016
rect 18315 57056 18357 57065
rect 18315 57016 18316 57056
rect 18356 57016 18357 57056
rect 18315 57007 18357 57016
rect 18411 57056 18453 57065
rect 18411 57016 18412 57056
rect 18452 57016 18453 57056
rect 18411 57007 18453 57016
rect 18883 57056 18941 57057
rect 18883 57016 18892 57056
rect 18932 57016 18941 57056
rect 19371 57030 19372 57070
rect 19412 57030 19413 57070
rect 19371 57021 19413 57030
rect 18883 57015 18941 57016
rect 7947 56972 7989 56981
rect 7947 56932 7948 56972
rect 7988 56932 7989 56972
rect 7947 56923 7989 56932
rect 13227 56972 13269 56981
rect 13227 56932 13228 56972
rect 13268 56932 13269 56972
rect 13227 56923 13269 56932
rect 1515 56888 1557 56897
rect 1515 56848 1516 56888
rect 1556 56848 1557 56888
rect 1515 56839 1557 56848
rect 1899 56888 1941 56897
rect 1899 56848 1900 56888
rect 1940 56848 1941 56888
rect 1899 56839 1941 56848
rect 2379 56888 2421 56897
rect 2379 56848 2380 56888
rect 2420 56848 2421 56888
rect 2379 56839 2421 56848
rect 5835 56888 5877 56897
rect 5835 56848 5836 56888
rect 5876 56848 5877 56888
rect 5835 56839 5877 56848
rect 9579 56888 9621 56897
rect 9579 56848 9580 56888
rect 9620 56848 9621 56888
rect 9579 56839 9621 56848
rect 11211 56888 11253 56897
rect 11211 56848 11212 56888
rect 11252 56848 11253 56888
rect 11211 56839 11253 56848
rect 15243 56888 15285 56897
rect 15243 56848 15244 56888
rect 15284 56848 15285 56888
rect 15243 56839 15285 56848
rect 16579 56888 16637 56889
rect 16579 56848 16588 56888
rect 16628 56848 16637 56888
rect 16579 56847 16637 56848
rect 17155 56888 17213 56889
rect 17155 56848 17164 56888
rect 17204 56848 17213 56888
rect 17155 56847 17213 56848
rect 17451 56888 17493 56897
rect 17451 56848 17452 56888
rect 17492 56848 17493 56888
rect 17451 56839 17493 56848
rect 19563 56888 19605 56897
rect 19563 56848 19564 56888
rect 19604 56848 19605 56888
rect 19563 56839 19605 56848
rect 19947 56888 19989 56897
rect 19947 56848 19948 56888
rect 19988 56848 19989 56888
rect 19947 56839 19989 56848
rect 1152 56720 20452 56744
rect 1152 56680 4928 56720
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 5296 56680 20048 56720
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20416 56680 20452 56720
rect 1152 56656 20452 56680
rect 1227 56552 1269 56561
rect 1227 56512 1228 56552
rect 1268 56512 1269 56552
rect 1227 56503 1269 56512
rect 5355 56552 5397 56561
rect 5355 56512 5356 56552
rect 5396 56512 5397 56552
rect 5355 56503 5397 56512
rect 16971 56552 17013 56561
rect 16971 56512 16972 56552
rect 17012 56512 17013 56552
rect 16971 56503 17013 56512
rect 17443 56552 17501 56553
rect 17443 56512 17452 56552
rect 17492 56512 17501 56552
rect 17443 56511 17501 56512
rect 3051 56468 3093 56477
rect 3051 56428 3052 56468
rect 3092 56428 3093 56468
rect 3051 56419 3093 56428
rect 10155 56468 10197 56477
rect 10155 56428 10156 56468
rect 10196 56428 10197 56468
rect 10155 56419 10197 56428
rect 13803 56468 13845 56477
rect 13803 56428 13804 56468
rect 13844 56428 13845 56468
rect 13803 56419 13845 56428
rect 1603 56384 1661 56385
rect 1603 56344 1612 56384
rect 1652 56344 1661 56384
rect 1603 56343 1661 56344
rect 2851 56384 2909 56385
rect 2851 56344 2860 56384
rect 2900 56344 2909 56384
rect 2851 56343 2909 56344
rect 3627 56384 3669 56393
rect 3627 56344 3628 56384
rect 3668 56344 3669 56384
rect 3627 56335 3669 56344
rect 3723 56384 3765 56393
rect 3723 56344 3724 56384
rect 3764 56344 3765 56384
rect 3723 56335 3765 56344
rect 4675 56384 4733 56385
rect 4675 56344 4684 56384
rect 4724 56344 4733 56384
rect 4675 56343 4733 56344
rect 5163 56379 5205 56388
rect 5163 56339 5164 56379
rect 5204 56339 5205 56379
rect 6019 56384 6077 56385
rect 6019 56344 6028 56384
rect 6068 56344 6077 56384
rect 6019 56343 6077 56344
rect 7267 56384 7325 56385
rect 7267 56344 7276 56384
rect 7316 56344 7325 56384
rect 7267 56343 7325 56344
rect 8515 56384 8573 56385
rect 8515 56344 8524 56384
rect 8564 56344 8573 56384
rect 8515 56343 8573 56344
rect 9763 56384 9821 56385
rect 9763 56344 9772 56384
rect 9812 56344 9821 56384
rect 9763 56343 9821 56344
rect 10347 56379 10389 56388
rect 5163 56330 5205 56339
rect 10347 56339 10348 56379
rect 10388 56339 10389 56379
rect 10819 56384 10877 56385
rect 10819 56344 10828 56384
rect 10868 56344 10877 56384
rect 10819 56343 10877 56344
rect 11307 56384 11349 56393
rect 11307 56344 11308 56384
rect 11348 56344 11349 56384
rect 10347 56330 10389 56339
rect 11307 56335 11349 56344
rect 11403 56384 11445 56393
rect 11403 56344 11404 56384
rect 11444 56344 11445 56384
rect 11403 56335 11445 56344
rect 11787 56384 11829 56393
rect 11787 56344 11788 56384
rect 11828 56344 11829 56384
rect 11787 56335 11829 56344
rect 11883 56384 11925 56393
rect 11883 56344 11884 56384
rect 11924 56344 11925 56384
rect 11883 56335 11925 56344
rect 12355 56384 12413 56385
rect 12355 56344 12364 56384
rect 12404 56344 12413 56384
rect 12355 56343 12413 56344
rect 13603 56384 13661 56385
rect 13603 56344 13612 56384
rect 13652 56344 13661 56384
rect 13603 56343 13661 56344
rect 15243 56384 15285 56393
rect 15243 56344 15244 56384
rect 15284 56344 15285 56384
rect 15243 56335 15285 56344
rect 15339 56384 15381 56393
rect 15339 56344 15340 56384
rect 15380 56344 15381 56384
rect 15339 56335 15381 56344
rect 15723 56384 15765 56393
rect 15723 56344 15724 56384
rect 15764 56344 15765 56384
rect 15723 56335 15765 56344
rect 16291 56384 16349 56385
rect 16291 56344 16300 56384
rect 16340 56344 16349 56384
rect 16291 56343 16349 56344
rect 16779 56379 16821 56388
rect 16779 56339 16780 56379
rect 16820 56339 16821 56379
rect 16779 56330 16821 56339
rect 17163 56384 17205 56393
rect 17163 56344 17164 56384
rect 17204 56344 17205 56384
rect 17163 56335 17205 56344
rect 17643 56384 17685 56393
rect 17643 56344 17644 56384
rect 17684 56344 17685 56384
rect 17251 56342 17309 56343
rect 1411 56300 1469 56301
rect 1411 56260 1420 56300
rect 1460 56260 1469 56300
rect 1411 56259 1469 56260
rect 4107 56300 4149 56309
rect 4107 56260 4108 56300
rect 4148 56260 4149 56300
rect 4107 56251 4149 56260
rect 4203 56300 4245 56309
rect 4203 56260 4204 56300
rect 4244 56260 4245 56300
rect 4203 56251 4245 56260
rect 15819 56300 15861 56309
rect 17251 56302 17260 56342
rect 17300 56302 17309 56342
rect 17251 56301 17309 56302
rect 17347 56342 17405 56343
rect 17347 56302 17356 56342
rect 17396 56302 17405 56342
rect 17643 56335 17685 56344
rect 17835 56384 17877 56393
rect 17835 56344 17836 56384
rect 17876 56344 17877 56384
rect 17835 56335 17877 56344
rect 18115 56384 18173 56385
rect 18115 56344 18124 56384
rect 18164 56344 18173 56384
rect 18115 56343 18173 56344
rect 19363 56384 19421 56385
rect 19363 56344 19372 56384
rect 19412 56344 19421 56384
rect 19363 56343 19421 56344
rect 17347 56301 17405 56302
rect 15819 56260 15820 56300
rect 15860 56260 15861 56300
rect 15819 56251 15861 56260
rect 19747 56300 19805 56301
rect 19747 56260 19756 56300
rect 19796 56260 19805 56300
rect 19747 56259 19805 56260
rect 7467 56132 7509 56141
rect 7467 56092 7468 56132
rect 7508 56092 7509 56132
rect 7467 56083 7509 56092
rect 9963 56132 10005 56141
rect 9963 56092 9964 56132
rect 10004 56092 10005 56132
rect 9963 56083 10005 56092
rect 17643 56132 17685 56141
rect 17643 56092 17644 56132
rect 17684 56092 17685 56132
rect 17643 56083 17685 56092
rect 19563 56132 19605 56141
rect 19563 56092 19564 56132
rect 19604 56092 19605 56132
rect 19563 56083 19605 56092
rect 19947 56132 19989 56141
rect 19947 56092 19948 56132
rect 19988 56092 19989 56132
rect 19947 56083 19989 56092
rect 1152 55964 20352 55988
rect 1152 55924 3688 55964
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 4056 55924 18808 55964
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 19176 55924 20352 55964
rect 1152 55900 20352 55924
rect 3243 55712 3285 55721
rect 3243 55672 3244 55712
rect 3284 55672 3285 55712
rect 3243 55663 3285 55672
rect 3043 55628 3101 55629
rect 3043 55588 3052 55628
rect 3092 55588 3101 55628
rect 3043 55587 3101 55588
rect 3427 55628 3485 55629
rect 3427 55588 3436 55628
rect 3476 55588 3485 55628
rect 3427 55587 3485 55588
rect 8811 55628 8853 55637
rect 8811 55588 8812 55628
rect 8852 55588 8853 55628
rect 8811 55579 8853 55588
rect 13603 55628 13661 55629
rect 13603 55588 13612 55628
rect 13652 55588 13661 55628
rect 13603 55587 13661 55588
rect 19363 55628 19421 55629
rect 19363 55588 19372 55628
rect 19412 55588 19421 55628
rect 19363 55587 19421 55588
rect 19747 55628 19805 55629
rect 19747 55588 19756 55628
rect 19796 55588 19805 55628
rect 19747 55587 19805 55588
rect 9819 55553 9861 55562
rect 13083 55553 13125 55562
rect 1219 55544 1277 55545
rect 1219 55504 1228 55544
rect 1268 55504 1277 55544
rect 1219 55503 1277 55504
rect 2467 55544 2525 55545
rect 2467 55504 2476 55544
rect 2516 55504 2525 55544
rect 2467 55503 2525 55504
rect 4675 55544 4733 55545
rect 4675 55504 4684 55544
rect 4724 55504 4733 55544
rect 4675 55503 4733 55504
rect 5923 55544 5981 55545
rect 5923 55504 5932 55544
rect 5972 55504 5981 55544
rect 5923 55503 5981 55504
rect 6499 55544 6557 55545
rect 6499 55504 6508 55544
rect 6548 55504 6557 55544
rect 6499 55503 6557 55504
rect 7747 55544 7805 55545
rect 7747 55504 7756 55544
rect 7796 55504 7805 55544
rect 7747 55503 7805 55504
rect 8235 55544 8277 55553
rect 8235 55504 8236 55544
rect 8276 55504 8277 55544
rect 8235 55495 8277 55504
rect 8331 55544 8373 55553
rect 8331 55504 8332 55544
rect 8372 55504 8373 55544
rect 8331 55495 8373 55504
rect 8715 55544 8757 55553
rect 8715 55504 8716 55544
rect 8756 55504 8757 55544
rect 8715 55495 8757 55504
rect 9283 55544 9341 55545
rect 9283 55504 9292 55544
rect 9332 55504 9341 55544
rect 9819 55513 9820 55553
rect 9860 55513 9861 55553
rect 9819 55504 9861 55513
rect 11499 55544 11541 55553
rect 11499 55504 11500 55544
rect 11540 55504 11541 55544
rect 9283 55503 9341 55504
rect 11499 55495 11541 55504
rect 11595 55544 11637 55553
rect 11595 55504 11596 55544
rect 11636 55504 11637 55544
rect 11595 55495 11637 55504
rect 11979 55544 12021 55553
rect 11979 55504 11980 55544
rect 12020 55504 12021 55544
rect 11979 55495 12021 55504
rect 12075 55544 12117 55553
rect 12075 55504 12076 55544
rect 12116 55504 12117 55544
rect 12075 55495 12117 55504
rect 12547 55544 12605 55545
rect 12547 55504 12556 55544
rect 12596 55504 12605 55544
rect 13083 55513 13084 55553
rect 13124 55513 13125 55553
rect 13083 55504 13125 55513
rect 15811 55544 15869 55545
rect 15811 55504 15820 55544
rect 15860 55504 15869 55544
rect 12547 55503 12605 55504
rect 15811 55503 15869 55504
rect 17059 55544 17117 55545
rect 17059 55504 17068 55544
rect 17108 55504 17117 55544
rect 17059 55503 17117 55504
rect 17443 55544 17501 55545
rect 17443 55504 17452 55544
rect 17492 55504 17501 55544
rect 17443 55503 17501 55504
rect 18691 55544 18749 55545
rect 18691 55504 18700 55544
rect 18740 55504 18749 55544
rect 18691 55503 18749 55504
rect 7947 55460 7989 55469
rect 7947 55420 7948 55460
rect 7988 55420 7989 55460
rect 7947 55411 7989 55420
rect 13227 55460 13269 55469
rect 13227 55420 13228 55460
rect 13268 55420 13269 55460
rect 13227 55411 13269 55420
rect 17259 55460 17301 55469
rect 17259 55420 17260 55460
rect 17300 55420 17301 55460
rect 17259 55411 17301 55420
rect 2667 55376 2709 55385
rect 2667 55336 2668 55376
rect 2708 55336 2709 55376
rect 2667 55327 2709 55336
rect 2859 55376 2901 55385
rect 2859 55336 2860 55376
rect 2900 55336 2901 55376
rect 2859 55327 2901 55336
rect 6123 55376 6165 55385
rect 6123 55336 6124 55376
rect 6164 55336 6165 55376
rect 6123 55327 6165 55336
rect 9963 55376 10005 55385
rect 9963 55336 9964 55376
rect 10004 55336 10005 55376
rect 9963 55327 10005 55336
rect 13419 55376 13461 55385
rect 13419 55336 13420 55376
rect 13460 55336 13461 55376
rect 13419 55327 13461 55336
rect 18891 55376 18933 55385
rect 18891 55336 18892 55376
rect 18932 55336 18933 55376
rect 18891 55327 18933 55336
rect 19563 55376 19605 55385
rect 19563 55336 19564 55376
rect 19604 55336 19605 55376
rect 19563 55327 19605 55336
rect 19947 55376 19989 55385
rect 19947 55336 19948 55376
rect 19988 55336 19989 55376
rect 19947 55327 19989 55336
rect 1152 55208 20452 55232
rect 1152 55168 4928 55208
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 5296 55168 20048 55208
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20416 55168 20452 55208
rect 1152 55144 20452 55168
rect 11499 55040 11541 55049
rect 11499 55000 11500 55040
rect 11540 55000 11541 55040
rect 11499 54991 11541 55000
rect 13227 55040 13269 55049
rect 13227 55000 13228 55040
rect 13268 55000 13269 55040
rect 13227 54991 13269 55000
rect 13419 55040 13461 55049
rect 13419 55000 13420 55040
rect 13460 55000 13461 55040
rect 13419 54991 13461 55000
rect 2475 54956 2517 54965
rect 2475 54916 2476 54956
rect 2516 54916 2517 54956
rect 2475 54907 2517 54916
rect 7755 54956 7797 54965
rect 7755 54916 7756 54956
rect 7796 54916 7797 54956
rect 7755 54907 7797 54916
rect 16107 54956 16149 54965
rect 16107 54916 16108 54956
rect 16148 54916 16149 54956
rect 16107 54907 16149 54916
rect 19563 54956 19605 54965
rect 19563 54916 19564 54956
rect 19604 54916 19605 54956
rect 19563 54907 19605 54916
rect 3139 54872 3197 54873
rect 2667 54858 2709 54867
rect 2667 54818 2668 54858
rect 2708 54818 2709 54858
rect 3139 54832 3148 54872
rect 3188 54832 3197 54872
rect 3139 54831 3197 54832
rect 3627 54872 3669 54881
rect 3627 54832 3628 54872
rect 3668 54832 3669 54872
rect 3627 54823 3669 54832
rect 4107 54872 4149 54881
rect 4107 54832 4108 54872
rect 4148 54832 4149 54872
rect 4107 54823 4149 54832
rect 4203 54872 4245 54881
rect 4203 54832 4204 54872
rect 4244 54832 4245 54872
rect 4203 54823 4245 54832
rect 6027 54872 6069 54881
rect 6027 54832 6028 54872
rect 6068 54832 6069 54872
rect 6027 54823 6069 54832
rect 6123 54872 6165 54881
rect 6123 54832 6124 54872
rect 6164 54832 6165 54872
rect 6123 54823 6165 54832
rect 6603 54872 6645 54881
rect 6603 54832 6604 54872
rect 6644 54832 6645 54872
rect 6603 54823 6645 54832
rect 7075 54872 7133 54873
rect 7075 54832 7084 54872
rect 7124 54832 7133 54872
rect 7075 54831 7133 54832
rect 7563 54867 7605 54876
rect 7563 54827 7564 54867
rect 7604 54827 7605 54867
rect 8419 54872 8477 54873
rect 8419 54832 8428 54872
rect 8468 54832 8477 54872
rect 8419 54831 8477 54832
rect 9667 54872 9725 54873
rect 9667 54832 9676 54872
rect 9716 54832 9725 54872
rect 9667 54831 9725 54832
rect 10051 54872 10109 54873
rect 10051 54832 10060 54872
rect 10100 54832 10109 54872
rect 10051 54831 10109 54832
rect 11299 54872 11357 54873
rect 11299 54832 11308 54872
rect 11348 54832 11357 54872
rect 11299 54831 11357 54832
rect 11779 54872 11837 54873
rect 11779 54832 11788 54872
rect 11828 54832 11837 54872
rect 11779 54831 11837 54832
rect 13027 54872 13085 54873
rect 13027 54832 13036 54872
rect 13076 54832 13085 54872
rect 13027 54831 13085 54832
rect 14379 54872 14421 54881
rect 14379 54832 14380 54872
rect 14420 54832 14421 54872
rect 7563 54818 7605 54827
rect 14379 54823 14421 54832
rect 14475 54872 14517 54881
rect 14475 54832 14476 54872
rect 14516 54832 14517 54872
rect 14475 54823 14517 54832
rect 14955 54872 14997 54881
rect 14955 54832 14956 54872
rect 14996 54832 14997 54872
rect 14955 54823 14997 54832
rect 15427 54872 15485 54873
rect 15427 54832 15436 54872
rect 15476 54832 15485 54872
rect 16387 54872 16445 54873
rect 15427 54831 15485 54832
rect 15915 54858 15957 54867
rect 15915 54818 15916 54858
rect 15956 54818 15957 54858
rect 16387 54832 16396 54872
rect 16436 54832 16445 54872
rect 16387 54831 16445 54832
rect 16683 54872 16725 54881
rect 16683 54832 16684 54872
rect 16724 54832 16725 54872
rect 16683 54823 16725 54832
rect 16779 54872 16821 54881
rect 16779 54832 16780 54872
rect 16820 54832 16821 54872
rect 16779 54823 16821 54832
rect 17835 54872 17877 54881
rect 17835 54832 17836 54872
rect 17876 54832 17877 54872
rect 17835 54823 17877 54832
rect 17931 54872 17973 54881
rect 17931 54832 17932 54872
rect 17972 54832 17973 54872
rect 17931 54823 17973 54832
rect 18411 54872 18453 54881
rect 18411 54832 18412 54872
rect 18452 54832 18453 54872
rect 18411 54823 18453 54832
rect 18883 54872 18941 54873
rect 18883 54832 18892 54872
rect 18932 54832 18941 54872
rect 18883 54831 18941 54832
rect 19371 54867 19413 54876
rect 19371 54827 19372 54867
rect 19412 54827 19413 54867
rect 19371 54818 19413 54827
rect 2667 54809 2709 54818
rect 15915 54809 15957 54818
rect 1699 54788 1757 54789
rect 1699 54748 1708 54788
rect 1748 54748 1757 54788
rect 1699 54747 1757 54748
rect 2083 54788 2141 54789
rect 2083 54748 2092 54788
rect 2132 54748 2141 54788
rect 2083 54747 2141 54748
rect 3723 54788 3765 54797
rect 3723 54748 3724 54788
rect 3764 54748 3765 54788
rect 3723 54739 3765 54748
rect 6507 54788 6549 54797
rect 6507 54748 6508 54788
rect 6548 54748 6549 54788
rect 6507 54739 6549 54748
rect 13603 54788 13661 54789
rect 13603 54748 13612 54788
rect 13652 54748 13661 54788
rect 13603 54747 13661 54748
rect 14859 54788 14901 54797
rect 14859 54748 14860 54788
rect 14900 54748 14901 54788
rect 14859 54739 14901 54748
rect 18315 54788 18357 54797
rect 18315 54748 18316 54788
rect 18356 54748 18357 54788
rect 18315 54739 18357 54748
rect 19747 54788 19805 54789
rect 19747 54748 19756 54788
rect 19796 54748 19805 54788
rect 19747 54747 19805 54748
rect 17059 54704 17117 54705
rect 17059 54664 17068 54704
rect 17108 54664 17117 54704
rect 17059 54663 17117 54664
rect 1515 54620 1557 54629
rect 1515 54580 1516 54620
rect 1556 54580 1557 54620
rect 1515 54571 1557 54580
rect 1899 54620 1941 54629
rect 1899 54580 1900 54620
rect 1940 54580 1941 54620
rect 1899 54571 1941 54580
rect 9867 54620 9909 54629
rect 9867 54580 9868 54620
rect 9908 54580 9909 54620
rect 9867 54571 9909 54580
rect 19947 54620 19989 54629
rect 19947 54580 19948 54620
rect 19988 54580 19989 54620
rect 19947 54571 19989 54580
rect 1152 54452 20352 54476
rect 1152 54412 3688 54452
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 4056 54412 18808 54452
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 19176 54412 20352 54452
rect 1152 54388 20352 54412
rect 14667 54284 14709 54293
rect 14667 54244 14668 54284
rect 14708 54244 14709 54284
rect 14667 54235 14709 54244
rect 16299 54284 16341 54293
rect 16299 54244 16300 54284
rect 16340 54244 16341 54284
rect 16299 54235 16341 54244
rect 4011 54200 4053 54209
rect 4011 54160 4012 54200
rect 4052 54160 4053 54200
rect 4011 54151 4053 54160
rect 17835 54200 17877 54209
rect 17835 54160 17836 54200
rect 17876 54160 17877 54200
rect 17835 54151 17877 54160
rect 1699 54116 1757 54117
rect 1699 54076 1708 54116
rect 1748 54076 1757 54116
rect 1699 54075 1757 54076
rect 2083 54116 2141 54117
rect 2083 54076 2092 54116
rect 2132 54076 2141 54116
rect 11395 54116 11453 54117
rect 2083 54075 2141 54076
rect 9627 54074 9669 54083
rect 11395 54076 11404 54116
rect 11444 54076 11453 54116
rect 11395 54075 11453 54076
rect 17635 54116 17693 54117
rect 17635 54076 17644 54116
rect 17684 54076 17693 54116
rect 17635 54075 17693 54076
rect 19651 54116 19709 54117
rect 19651 54076 19660 54116
rect 19700 54076 19709 54116
rect 19651 54075 19709 54076
rect 20035 54116 20093 54117
rect 20035 54076 20044 54116
rect 20084 54076 20093 54116
rect 20035 54075 20093 54076
rect 2563 54032 2621 54033
rect 2563 53992 2572 54032
rect 2612 53992 2621 54032
rect 2563 53991 2621 53992
rect 3811 54032 3869 54033
rect 3811 53992 3820 54032
rect 3860 53992 3869 54032
rect 3811 53991 3869 53992
rect 4387 54032 4445 54033
rect 4387 53992 4396 54032
rect 4436 53992 4445 54032
rect 4387 53991 4445 53992
rect 5635 54032 5693 54033
rect 5635 53992 5644 54032
rect 5684 53992 5693 54032
rect 5635 53991 5693 53992
rect 6307 54032 6365 54033
rect 6307 53992 6316 54032
rect 6356 53992 6365 54032
rect 6307 53991 6365 53992
rect 7555 54032 7613 54033
rect 7555 53992 7564 54032
rect 7604 53992 7613 54032
rect 7555 53991 7613 53992
rect 8043 54032 8085 54041
rect 8043 53992 8044 54032
rect 8084 53992 8085 54032
rect 8043 53983 8085 53992
rect 8139 54032 8181 54041
rect 8139 53992 8140 54032
rect 8180 53992 8181 54032
rect 8139 53983 8181 53992
rect 8523 54032 8565 54041
rect 8523 53992 8524 54032
rect 8564 53992 8565 54032
rect 8523 53983 8565 53992
rect 8619 54032 8661 54041
rect 9627 54034 9628 54074
rect 9668 54034 9669 54074
rect 8619 53992 8620 54032
rect 8660 53992 8661 54032
rect 8619 53983 8661 53992
rect 9091 54032 9149 54033
rect 9091 53992 9100 54032
rect 9140 53992 9149 54032
rect 9627 54025 9669 54034
rect 11587 54032 11645 54033
rect 9091 53991 9149 53992
rect 11587 53992 11596 54032
rect 11636 53992 11645 54032
rect 11587 53991 11645 53992
rect 12835 54032 12893 54033
rect 12835 53992 12844 54032
rect 12884 53992 12893 54032
rect 12835 53991 12893 53992
rect 13219 54032 13277 54033
rect 13219 53992 13228 54032
rect 13268 53992 13277 54032
rect 13219 53991 13277 53992
rect 14467 54032 14525 54033
rect 14467 53992 14476 54032
rect 14516 53992 14525 54032
rect 14467 53991 14525 53992
rect 14851 54032 14909 54033
rect 14851 53992 14860 54032
rect 14900 53992 14909 54032
rect 14851 53991 14909 53992
rect 16099 54032 16157 54033
rect 16099 53992 16108 54032
rect 16148 53992 16157 54032
rect 16099 53991 16157 53992
rect 18019 54032 18077 54033
rect 18019 53992 18028 54032
rect 18068 53992 18077 54032
rect 18019 53991 18077 53992
rect 19267 54032 19325 54033
rect 19267 53992 19276 54032
rect 19316 53992 19325 54032
rect 19267 53991 19325 53992
rect 9771 53948 9813 53957
rect 9771 53908 9772 53948
rect 9812 53908 9813 53948
rect 9771 53899 9813 53908
rect 1515 53864 1557 53873
rect 1515 53824 1516 53864
rect 1556 53824 1557 53864
rect 1515 53815 1557 53824
rect 1899 53864 1941 53873
rect 1899 53824 1900 53864
rect 1940 53824 1941 53864
rect 1899 53815 1941 53824
rect 5835 53864 5877 53873
rect 5835 53824 5836 53864
rect 5876 53824 5877 53864
rect 5835 53815 5877 53824
rect 7755 53864 7797 53873
rect 7755 53824 7756 53864
rect 7796 53824 7797 53864
rect 7755 53815 7797 53824
rect 11211 53864 11253 53873
rect 11211 53824 11212 53864
rect 11252 53824 11253 53864
rect 11211 53815 11253 53824
rect 13035 53864 13077 53873
rect 13035 53824 13036 53864
rect 13076 53824 13077 53864
rect 13035 53815 13077 53824
rect 19467 53864 19509 53873
rect 19467 53824 19468 53864
rect 19508 53824 19509 53864
rect 19467 53815 19509 53824
rect 19851 53864 19893 53873
rect 19851 53824 19852 53864
rect 19892 53824 19893 53864
rect 19851 53815 19893 53824
rect 20235 53864 20277 53873
rect 20235 53824 20236 53864
rect 20276 53824 20277 53864
rect 20235 53815 20277 53824
rect 1152 53696 20452 53720
rect 1152 53656 4928 53696
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 5296 53656 20048 53696
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20416 53656 20452 53696
rect 1152 53632 20452 53656
rect 5739 53528 5781 53537
rect 5739 53488 5740 53528
rect 5780 53488 5781 53528
rect 5739 53479 5781 53488
rect 13323 53528 13365 53537
rect 13323 53488 13324 53528
rect 13364 53488 13365 53528
rect 13323 53479 13365 53488
rect 3531 53444 3573 53453
rect 3531 53404 3532 53444
rect 3572 53404 3573 53444
rect 3531 53395 3573 53404
rect 11307 53444 11349 53453
rect 11307 53404 11308 53444
rect 11348 53404 11349 53444
rect 11307 53395 11349 53404
rect 15435 53444 15477 53453
rect 15435 53404 15436 53444
rect 15476 53404 15477 53444
rect 15435 53395 15477 53404
rect 2083 53360 2141 53361
rect 2083 53320 2092 53360
rect 2132 53320 2141 53360
rect 2083 53319 2141 53320
rect 3331 53360 3389 53361
rect 3331 53320 3340 53360
rect 3380 53320 3389 53360
rect 3331 53319 3389 53320
rect 4011 53360 4053 53369
rect 4011 53320 4012 53360
rect 4052 53320 4053 53360
rect 4011 53311 4053 53320
rect 4107 53360 4149 53369
rect 4107 53320 4108 53360
rect 4148 53320 4149 53360
rect 4107 53311 4149 53320
rect 5059 53360 5117 53361
rect 5059 53320 5068 53360
rect 5108 53320 5117 53360
rect 8227 53360 8285 53361
rect 5059 53319 5117 53320
rect 5595 53350 5637 53359
rect 5595 53310 5596 53350
rect 5636 53310 5637 53350
rect 8227 53320 8236 53360
rect 8276 53320 8285 53360
rect 8227 53319 8285 53320
rect 9475 53360 9533 53361
rect 9475 53320 9484 53360
rect 9524 53320 9533 53360
rect 9475 53319 9533 53320
rect 9859 53360 9917 53361
rect 9859 53320 9868 53360
rect 9908 53320 9917 53360
rect 9859 53319 9917 53320
rect 11107 53360 11165 53361
rect 11107 53320 11116 53360
rect 11156 53320 11165 53360
rect 11107 53319 11165 53320
rect 11595 53360 11637 53369
rect 11595 53320 11596 53360
rect 11636 53320 11637 53360
rect 11595 53311 11637 53320
rect 11691 53360 11733 53369
rect 11691 53320 11692 53360
rect 11732 53320 11733 53360
rect 11691 53311 11733 53320
rect 12075 53360 12117 53369
rect 12075 53320 12076 53360
rect 12116 53320 12117 53360
rect 12075 53311 12117 53320
rect 12643 53360 12701 53361
rect 12643 53320 12652 53360
rect 12692 53320 12701 53360
rect 12643 53319 12701 53320
rect 13131 53355 13173 53364
rect 13131 53315 13132 53355
rect 13172 53315 13173 53355
rect 5595 53301 5637 53310
rect 13131 53306 13173 53315
rect 13707 53360 13749 53369
rect 13707 53320 13708 53360
rect 13748 53320 13749 53360
rect 13707 53311 13749 53320
rect 13803 53360 13845 53369
rect 13803 53320 13804 53360
rect 13844 53320 13845 53360
rect 13803 53311 13845 53320
rect 14187 53360 14229 53369
rect 14187 53320 14188 53360
rect 14228 53320 14229 53360
rect 14187 53311 14229 53320
rect 14755 53360 14813 53361
rect 14755 53320 14764 53360
rect 14804 53320 14813 53360
rect 15619 53360 15677 53361
rect 14755 53319 14813 53320
rect 15243 53346 15285 53355
rect 15243 53306 15244 53346
rect 15284 53306 15285 53346
rect 15619 53320 15628 53360
rect 15668 53320 15677 53360
rect 15619 53319 15677 53320
rect 15907 53360 15965 53361
rect 15907 53320 15916 53360
rect 15956 53320 15965 53360
rect 15907 53319 15965 53320
rect 17155 53360 17213 53361
rect 17155 53320 17164 53360
rect 17204 53320 17213 53360
rect 17155 53319 17213 53320
rect 18307 53360 18365 53361
rect 18307 53320 18316 53360
rect 18356 53320 18365 53360
rect 18307 53319 18365 53320
rect 19555 53360 19613 53361
rect 19555 53320 19564 53360
rect 19604 53320 19613 53360
rect 19555 53319 19613 53320
rect 15243 53297 15285 53306
rect 1507 53276 1565 53277
rect 1507 53236 1516 53276
rect 1556 53236 1565 53276
rect 1507 53235 1565 53236
rect 1891 53276 1949 53277
rect 1891 53236 1900 53276
rect 1940 53236 1949 53276
rect 1891 53235 1949 53236
rect 4491 53276 4533 53285
rect 4491 53236 4492 53276
rect 4532 53236 4533 53276
rect 4491 53227 4533 53236
rect 4587 53276 4629 53285
rect 4587 53236 4588 53276
rect 4628 53236 4629 53276
rect 4587 53227 4629 53236
rect 12171 53276 12213 53285
rect 12171 53236 12172 53276
rect 12212 53236 12213 53276
rect 12171 53227 12213 53236
rect 14283 53276 14325 53285
rect 14283 53236 14284 53276
rect 14324 53236 14325 53276
rect 14283 53227 14325 53236
rect 19939 53276 19997 53277
rect 19939 53236 19948 53276
rect 19988 53236 19997 53276
rect 19939 53235 19997 53236
rect 1323 53108 1365 53117
rect 1323 53068 1324 53108
rect 1364 53068 1365 53108
rect 1323 53059 1365 53068
rect 1707 53108 1749 53117
rect 1707 53068 1708 53108
rect 1748 53068 1749 53108
rect 1707 53059 1749 53068
rect 9675 53108 9717 53117
rect 9675 53068 9676 53108
rect 9716 53068 9717 53108
rect 9675 53059 9717 53068
rect 15723 53108 15765 53117
rect 15723 53068 15724 53108
rect 15764 53068 15765 53108
rect 15723 53059 15765 53068
rect 17355 53108 17397 53117
rect 17355 53068 17356 53108
rect 17396 53068 17397 53108
rect 17355 53059 17397 53068
rect 19755 53108 19797 53117
rect 19755 53068 19756 53108
rect 19796 53068 19797 53108
rect 19755 53059 19797 53068
rect 20139 53108 20181 53117
rect 20139 53068 20140 53108
rect 20180 53068 20181 53108
rect 20139 53059 20181 53068
rect 1152 52940 20352 52964
rect 1152 52900 3688 52940
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 4056 52900 18808 52940
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 19176 52900 20352 52940
rect 1152 52876 20352 52900
rect 14379 52688 14421 52697
rect 14379 52648 14380 52688
rect 14420 52648 14421 52688
rect 14379 52639 14421 52648
rect 15523 52688 15581 52689
rect 15523 52648 15532 52688
rect 15572 52648 15581 52688
rect 15523 52647 15581 52648
rect 17931 52604 17973 52613
rect 17931 52564 17932 52604
rect 17972 52564 17973 52604
rect 17931 52555 17973 52564
rect 18027 52604 18069 52613
rect 18027 52564 18028 52604
rect 18068 52564 18069 52604
rect 18027 52555 18069 52564
rect 19363 52604 19421 52605
rect 19363 52564 19372 52604
rect 19412 52564 19421 52604
rect 19363 52563 19421 52564
rect 19747 52604 19805 52605
rect 19747 52564 19756 52604
rect 19796 52564 19805 52604
rect 19747 52563 19805 52564
rect 9867 52534 9909 52543
rect 1507 52520 1565 52521
rect 1507 52480 1516 52520
rect 1556 52480 1565 52520
rect 1507 52479 1565 52480
rect 2755 52520 2813 52521
rect 2755 52480 2764 52520
rect 2804 52480 2813 52520
rect 2755 52479 2813 52480
rect 3243 52520 3285 52529
rect 3243 52480 3244 52520
rect 3284 52480 3285 52520
rect 3243 52471 3285 52480
rect 3339 52520 3381 52529
rect 3339 52480 3340 52520
rect 3380 52480 3381 52520
rect 3339 52471 3381 52480
rect 3723 52520 3765 52529
rect 3723 52480 3724 52520
rect 3764 52480 3765 52520
rect 3723 52471 3765 52480
rect 3819 52520 3861 52529
rect 4779 52525 4821 52534
rect 3819 52480 3820 52520
rect 3860 52480 3861 52520
rect 3819 52471 3861 52480
rect 4291 52520 4349 52521
rect 4291 52480 4300 52520
rect 4340 52480 4349 52520
rect 4291 52479 4349 52480
rect 4779 52485 4780 52525
rect 4820 52485 4821 52525
rect 4779 52476 4821 52485
rect 6595 52520 6653 52521
rect 6595 52480 6604 52520
rect 6644 52480 6653 52520
rect 6595 52479 6653 52480
rect 7843 52520 7901 52521
rect 7843 52480 7852 52520
rect 7892 52480 7901 52520
rect 7843 52479 7901 52480
rect 8331 52520 8373 52529
rect 8331 52480 8332 52520
rect 8372 52480 8373 52520
rect 8331 52471 8373 52480
rect 8427 52520 8469 52529
rect 8427 52480 8428 52520
rect 8468 52480 8469 52520
rect 8427 52471 8469 52480
rect 8811 52520 8853 52529
rect 8811 52480 8812 52520
rect 8852 52480 8853 52520
rect 8811 52471 8853 52480
rect 8907 52520 8949 52529
rect 8907 52480 8908 52520
rect 8948 52480 8949 52520
rect 8907 52471 8949 52480
rect 9379 52520 9437 52521
rect 9379 52480 9388 52520
rect 9428 52480 9437 52520
rect 9867 52494 9868 52534
rect 9908 52494 9909 52534
rect 18987 52534 19029 52543
rect 9867 52485 9909 52494
rect 12931 52520 12989 52521
rect 9379 52479 9437 52480
rect 12931 52480 12940 52520
rect 12980 52480 12989 52520
rect 12931 52479 12989 52480
rect 14179 52520 14237 52521
rect 14179 52480 14188 52520
rect 14228 52480 14237 52520
rect 14179 52479 14237 52480
rect 14851 52520 14909 52521
rect 14851 52480 14860 52520
rect 14900 52480 14909 52520
rect 14851 52479 14909 52480
rect 15147 52520 15189 52529
rect 15147 52480 15148 52520
rect 15188 52480 15189 52520
rect 15147 52471 15189 52480
rect 15243 52520 15285 52529
rect 15243 52480 15244 52520
rect 15284 52480 15285 52520
rect 15243 52471 15285 52480
rect 15715 52520 15773 52521
rect 15715 52480 15724 52520
rect 15764 52480 15773 52520
rect 15715 52479 15773 52480
rect 16963 52520 17021 52521
rect 16963 52480 16972 52520
rect 17012 52480 17021 52520
rect 16963 52479 17021 52480
rect 17451 52520 17493 52529
rect 17451 52480 17452 52520
rect 17492 52480 17493 52520
rect 17451 52471 17493 52480
rect 17547 52520 17589 52529
rect 17547 52480 17548 52520
rect 17588 52480 17589 52520
rect 17547 52471 17589 52480
rect 18499 52520 18557 52521
rect 18499 52480 18508 52520
rect 18548 52480 18557 52520
rect 18987 52494 18988 52534
rect 19028 52494 19029 52534
rect 18987 52485 19029 52494
rect 18499 52479 18557 52480
rect 2955 52436 2997 52445
rect 2955 52396 2956 52436
rect 2996 52396 2997 52436
rect 2955 52387 2997 52396
rect 4971 52436 5013 52445
rect 4971 52396 4972 52436
rect 5012 52396 5013 52436
rect 4971 52387 5013 52396
rect 8043 52436 8085 52445
rect 8043 52396 8044 52436
rect 8084 52396 8085 52436
rect 8043 52387 8085 52396
rect 10059 52436 10101 52445
rect 10059 52396 10060 52436
rect 10100 52396 10101 52436
rect 10059 52387 10101 52396
rect 17163 52436 17205 52445
rect 17163 52396 17164 52436
rect 17204 52396 17205 52436
rect 17163 52387 17205 52396
rect 19179 52352 19221 52361
rect 19179 52312 19180 52352
rect 19220 52312 19221 52352
rect 19179 52303 19221 52312
rect 19563 52352 19605 52361
rect 19563 52312 19564 52352
rect 19604 52312 19605 52352
rect 19563 52303 19605 52312
rect 19947 52352 19989 52361
rect 19947 52312 19948 52352
rect 19988 52312 19989 52352
rect 19947 52303 19989 52312
rect 1152 52184 20452 52208
rect 1152 52144 4928 52184
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 5296 52144 20048 52184
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20416 52144 20452 52184
rect 1152 52120 20452 52144
rect 4587 52016 4629 52025
rect 4587 51976 4588 52016
rect 4628 51976 4629 52016
rect 4587 51967 4629 51976
rect 6219 52016 6261 52025
rect 6219 51976 6220 52016
rect 6260 51976 6261 52016
rect 6219 51967 6261 51976
rect 13707 52016 13749 52025
rect 13707 51976 13708 52016
rect 13748 51976 13749 52016
rect 13707 51967 13749 51976
rect 8235 51932 8277 51941
rect 8235 51892 8236 51932
rect 8276 51892 8277 51932
rect 8235 51883 8277 51892
rect 11691 51932 11733 51941
rect 11691 51892 11692 51932
rect 11732 51892 11733 51932
rect 11691 51883 11733 51892
rect 16011 51932 16053 51941
rect 16011 51892 16012 51932
rect 16052 51892 16053 51932
rect 16011 51883 16053 51892
rect 19083 51932 19125 51941
rect 19083 51892 19084 51932
rect 19124 51892 19125 51932
rect 19083 51883 19125 51892
rect 16580 51859 16638 51860
rect 1507 51848 1565 51849
rect 1507 51808 1516 51848
rect 1556 51808 1565 51848
rect 1507 51807 1565 51808
rect 2755 51848 2813 51849
rect 2755 51808 2764 51848
rect 2804 51808 2813 51848
rect 2755 51807 2813 51808
rect 3139 51848 3197 51849
rect 3139 51808 3148 51848
rect 3188 51808 3197 51848
rect 3139 51807 3197 51808
rect 4387 51848 4445 51849
rect 4387 51808 4396 51848
rect 4436 51808 4445 51848
rect 4387 51807 4445 51808
rect 4771 51848 4829 51849
rect 4771 51808 4780 51848
rect 4820 51808 4829 51848
rect 4771 51807 4829 51808
rect 6019 51848 6077 51849
rect 6019 51808 6028 51848
rect 6068 51808 6077 51848
rect 6019 51807 6077 51808
rect 6507 51848 6549 51857
rect 6507 51808 6508 51848
rect 6548 51808 6549 51848
rect 6507 51799 6549 51808
rect 6603 51848 6645 51857
rect 6603 51808 6604 51848
rect 6644 51808 6645 51848
rect 6603 51799 6645 51808
rect 6987 51848 7029 51857
rect 6987 51808 6988 51848
rect 7028 51808 7029 51848
rect 6987 51799 7029 51808
rect 7083 51848 7125 51857
rect 7083 51808 7084 51848
rect 7124 51808 7125 51848
rect 7083 51799 7125 51808
rect 7555 51848 7613 51849
rect 7555 51808 7564 51848
rect 7604 51808 7613 51848
rect 9291 51848 9333 51857
rect 7555 51807 7613 51808
rect 8043 51834 8085 51843
rect 8043 51794 8044 51834
rect 8084 51794 8085 51834
rect 9291 51808 9292 51848
rect 9332 51808 9333 51848
rect 9291 51799 9333 51808
rect 9579 51848 9621 51857
rect 9579 51808 9580 51848
rect 9620 51808 9621 51848
rect 9579 51799 9621 51808
rect 9963 51848 10005 51857
rect 9963 51808 9964 51848
rect 10004 51808 10005 51848
rect 9963 51799 10005 51808
rect 10059 51848 10101 51857
rect 10059 51808 10060 51848
rect 10100 51808 10101 51848
rect 10059 51799 10101 51808
rect 10539 51848 10581 51857
rect 10539 51808 10540 51848
rect 10580 51808 10581 51848
rect 10539 51799 10581 51808
rect 11011 51848 11069 51849
rect 11011 51808 11020 51848
rect 11060 51808 11069 51848
rect 12259 51848 12317 51849
rect 11011 51807 11069 51808
rect 11499 51834 11541 51843
rect 8043 51785 8085 51794
rect 11499 51794 11500 51834
rect 11540 51794 11541 51834
rect 12259 51808 12268 51848
rect 12308 51808 12317 51848
rect 12259 51807 12317 51808
rect 13507 51848 13565 51849
rect 13507 51808 13516 51848
rect 13556 51808 13565 51848
rect 13507 51807 13565 51808
rect 14091 51848 14133 51857
rect 14091 51808 14092 51848
rect 14132 51808 14133 51848
rect 14091 51799 14133 51808
rect 14379 51848 14421 51857
rect 14379 51808 14380 51848
rect 14420 51808 14421 51848
rect 14379 51799 14421 51808
rect 14563 51848 14621 51849
rect 14563 51808 14572 51848
rect 14612 51808 14621 51848
rect 14563 51807 14621 51808
rect 15811 51848 15869 51849
rect 15811 51808 15820 51848
rect 15860 51808 15869 51848
rect 15811 51807 15869 51808
rect 16203 51848 16245 51857
rect 16203 51808 16204 51848
rect 16244 51808 16245 51848
rect 16203 51799 16245 51808
rect 16395 51848 16437 51857
rect 16395 51808 16396 51848
rect 16436 51808 16437 51848
rect 16580 51819 16589 51859
rect 16629 51819 16638 51859
rect 16580 51818 16638 51819
rect 16779 51848 16821 51857
rect 16395 51799 16437 51808
rect 16779 51808 16780 51848
rect 16820 51808 16821 51848
rect 16779 51799 16821 51808
rect 17355 51848 17397 51857
rect 17355 51808 17356 51848
rect 17396 51808 17397 51848
rect 17355 51799 17397 51808
rect 17451 51848 17493 51857
rect 17451 51808 17452 51848
rect 17492 51808 17493 51848
rect 17451 51799 17493 51808
rect 17835 51848 17877 51857
rect 17835 51808 17836 51848
rect 17876 51808 17877 51848
rect 17835 51799 17877 51808
rect 17931 51848 17973 51857
rect 17931 51808 17932 51848
rect 17972 51808 17973 51848
rect 17931 51799 17973 51808
rect 18403 51848 18461 51849
rect 18403 51808 18412 51848
rect 18452 51808 18461 51848
rect 18403 51807 18461 51808
rect 18891 51843 18933 51852
rect 18891 51803 18892 51843
rect 18932 51803 18933 51843
rect 18891 51794 18933 51803
rect 11499 51785 11541 51794
rect 8611 51764 8669 51765
rect 8611 51724 8620 51764
rect 8660 51724 8669 51764
rect 8611 51723 8669 51724
rect 10443 51764 10485 51773
rect 10443 51724 10444 51764
rect 10484 51724 10485 51764
rect 10443 51715 10485 51724
rect 14187 51764 14229 51773
rect 14187 51724 14188 51764
rect 14228 51724 14229 51764
rect 14187 51715 14229 51724
rect 16299 51764 16341 51773
rect 16299 51724 16300 51764
rect 16340 51724 16341 51764
rect 16299 51715 16341 51724
rect 19363 51764 19421 51765
rect 19363 51724 19372 51764
rect 19412 51724 19421 51764
rect 19363 51723 19421 51724
rect 19747 51764 19805 51765
rect 19747 51724 19756 51764
rect 19796 51724 19805 51764
rect 19747 51723 19805 51724
rect 2955 51680 2997 51689
rect 2955 51640 2956 51680
rect 2996 51640 2997 51680
rect 2955 51631 2997 51640
rect 19563 51680 19605 51689
rect 19563 51640 19564 51680
rect 19604 51640 19605 51680
rect 19563 51631 19605 51640
rect 19947 51680 19989 51689
rect 19947 51640 19948 51680
rect 19988 51640 19989 51680
rect 19947 51631 19989 51640
rect 8427 51596 8469 51605
rect 8427 51556 8428 51596
rect 8468 51556 8469 51596
rect 8427 51547 8469 51556
rect 9291 51596 9333 51605
rect 9291 51556 9292 51596
rect 9332 51556 9333 51596
rect 9291 51547 9333 51556
rect 16587 51596 16629 51605
rect 16587 51556 16588 51596
rect 16628 51556 16629 51596
rect 16587 51547 16629 51556
rect 1152 51428 20352 51452
rect 1152 51388 3688 51428
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 4056 51388 18808 51428
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 19176 51388 20352 51428
rect 1152 51364 20352 51388
rect 7947 51260 7989 51269
rect 7947 51220 7948 51260
rect 7988 51220 7989 51260
rect 7947 51211 7989 51220
rect 9963 51260 10005 51269
rect 9963 51220 9964 51260
rect 10004 51220 10005 51260
rect 9963 51211 10005 51220
rect 11787 51260 11829 51269
rect 11787 51220 11788 51260
rect 11828 51220 11829 51260
rect 11787 51211 11829 51220
rect 15435 51260 15477 51269
rect 15435 51220 15436 51260
rect 15476 51220 15477 51260
rect 15435 51211 15477 51220
rect 3043 51092 3101 51093
rect 3043 51052 3052 51092
rect 3092 51052 3101 51092
rect 3043 51051 3101 51052
rect 4587 51092 4629 51101
rect 4587 51052 4588 51092
rect 4628 51052 4629 51092
rect 4587 51043 4629 51052
rect 1219 51008 1277 51009
rect 1219 50968 1228 51008
rect 1268 50968 1277 51008
rect 1219 50967 1277 50968
rect 2467 51008 2525 51009
rect 2467 50968 2476 51008
rect 2516 50968 2525 51008
rect 2467 50967 2525 50968
rect 4011 51008 4053 51017
rect 4011 50968 4012 51008
rect 4052 50968 4053 51008
rect 4011 50959 4053 50968
rect 4107 51008 4149 51017
rect 4107 50968 4108 51008
rect 4148 50968 4149 51008
rect 4107 50959 4149 50968
rect 4491 51008 4533 51017
rect 5547 51013 5589 51022
rect 4491 50968 4492 51008
rect 4532 50968 4533 51008
rect 4491 50959 4533 50968
rect 5059 51008 5117 51009
rect 5059 50968 5068 51008
rect 5108 50968 5117 51008
rect 5059 50967 5117 50968
rect 5547 50973 5548 51013
rect 5588 50973 5589 51013
rect 5547 50964 5589 50973
rect 6499 51008 6557 51009
rect 6499 50968 6508 51008
rect 6548 50968 6557 51008
rect 6499 50967 6557 50968
rect 7747 51008 7805 51009
rect 7747 50968 7756 51008
rect 7796 50968 7805 51008
rect 7747 50967 7805 50968
rect 8515 51008 8573 51009
rect 8515 50968 8524 51008
rect 8564 50968 8573 51008
rect 8515 50967 8573 50968
rect 9763 51008 9821 51009
rect 9763 50968 9772 51008
rect 9812 50968 9821 51008
rect 9763 50967 9821 50968
rect 10339 51008 10397 51009
rect 10339 50968 10348 51008
rect 10388 50968 10397 51008
rect 10339 50967 10397 50968
rect 11587 51008 11645 51009
rect 11587 50968 11596 51008
rect 11636 50968 11645 51008
rect 11587 50967 11645 50968
rect 12739 51008 12797 51009
rect 12739 50968 12748 51008
rect 12788 50968 12797 51008
rect 12739 50967 12797 50968
rect 13987 51008 14045 51009
rect 13987 50968 13996 51008
rect 14036 50968 14045 51008
rect 13987 50967 14045 50968
rect 14475 51008 14517 51017
rect 14475 50968 14476 51008
rect 14516 50968 14517 51008
rect 14475 50959 14517 50968
rect 14571 51008 14613 51017
rect 14571 50968 14572 51008
rect 14612 50968 14613 51008
rect 14571 50959 14613 50968
rect 14667 51008 14709 51017
rect 14667 50968 14668 51008
rect 14708 50968 14709 51008
rect 14667 50959 14709 50968
rect 14763 51008 14805 51017
rect 14763 50968 14764 51008
rect 14804 50968 14805 51008
rect 14763 50959 14805 50968
rect 14955 51008 14997 51017
rect 14955 50968 14956 51008
rect 14996 50968 14997 51008
rect 14955 50959 14997 50968
rect 15051 51008 15093 51017
rect 15051 50968 15052 51008
rect 15092 50968 15093 51008
rect 15051 50959 15093 50968
rect 15147 51008 15189 51017
rect 15147 50968 15148 51008
rect 15188 50968 15189 51008
rect 15147 50959 15189 50968
rect 15243 51008 15285 51017
rect 15243 50968 15244 51008
rect 15284 50968 15285 51008
rect 15243 50959 15285 50968
rect 15435 51008 15477 51017
rect 15435 50968 15436 51008
rect 15476 50968 15477 51008
rect 15435 50959 15477 50968
rect 15627 51008 15669 51017
rect 15627 50968 15628 51008
rect 15668 50968 15669 51008
rect 15627 50959 15669 50968
rect 15715 51008 15773 51009
rect 15715 50968 15724 51008
rect 15764 50968 15773 51008
rect 15715 50967 15773 50968
rect 16291 51008 16349 51009
rect 16291 50968 16300 51008
rect 16340 50968 16349 51008
rect 16291 50967 16349 50968
rect 17539 51008 17597 51009
rect 17539 50968 17548 51008
rect 17588 50968 17597 51008
rect 17539 50967 17597 50968
rect 18307 51008 18365 51009
rect 18307 50968 18316 51008
rect 18356 50968 18365 51008
rect 18307 50967 18365 50968
rect 19555 51008 19613 51009
rect 19555 50968 19564 51008
rect 19604 50968 19613 51008
rect 19555 50967 19613 50968
rect 5739 50924 5781 50933
rect 5739 50884 5740 50924
rect 5780 50884 5781 50924
rect 5739 50875 5781 50884
rect 20131 50882 20189 50883
rect 2667 50840 2709 50849
rect 2667 50800 2668 50840
rect 2708 50800 2709 50840
rect 2667 50791 2709 50800
rect 2859 50840 2901 50849
rect 2859 50800 2860 50840
rect 2900 50800 2901 50840
rect 2859 50791 2901 50800
rect 14187 50840 14229 50849
rect 14187 50800 14188 50840
rect 14228 50800 14229 50840
rect 14187 50791 14229 50800
rect 17739 50840 17781 50849
rect 17739 50800 17740 50840
rect 17780 50800 17781 50840
rect 17739 50791 17781 50800
rect 19755 50840 19797 50849
rect 20131 50842 20140 50882
rect 20180 50842 20189 50882
rect 20131 50841 20189 50842
rect 19755 50800 19756 50840
rect 19796 50800 19797 50840
rect 19755 50791 19797 50800
rect 1152 50672 20452 50696
rect 1152 50632 4928 50672
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 5296 50632 20048 50672
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20416 50632 20452 50672
rect 1152 50608 20452 50632
rect 5739 50504 5781 50513
rect 5739 50464 5740 50504
rect 5780 50464 5781 50504
rect 5739 50455 5781 50464
rect 9195 50420 9237 50429
rect 9195 50380 9196 50420
rect 9236 50380 9237 50420
rect 9195 50371 9237 50380
rect 14283 50420 14325 50429
rect 14283 50380 14284 50420
rect 14324 50380 14325 50420
rect 14283 50371 14325 50380
rect 2659 50336 2717 50337
rect 2659 50296 2668 50336
rect 2708 50296 2717 50336
rect 2659 50295 2717 50296
rect 3907 50336 3965 50337
rect 3907 50296 3916 50336
rect 3956 50296 3965 50336
rect 3907 50295 3965 50296
rect 4291 50336 4349 50337
rect 4291 50296 4300 50336
rect 4340 50296 4349 50336
rect 4291 50295 4349 50296
rect 5539 50336 5597 50337
rect 5539 50296 5548 50336
rect 5588 50296 5597 50336
rect 5539 50295 5597 50296
rect 5923 50336 5981 50337
rect 5923 50296 5932 50336
rect 5972 50296 5981 50336
rect 5923 50295 5981 50296
rect 7171 50336 7229 50337
rect 7171 50296 7180 50336
rect 7220 50296 7229 50336
rect 7171 50295 7229 50296
rect 7747 50336 7805 50337
rect 7747 50296 7756 50336
rect 7796 50296 7805 50336
rect 7747 50295 7805 50296
rect 8995 50336 9053 50337
rect 8995 50296 9004 50336
rect 9044 50296 9053 50336
rect 8995 50295 9053 50296
rect 9475 50336 9533 50337
rect 9475 50296 9484 50336
rect 9524 50296 9533 50336
rect 9475 50295 9533 50296
rect 9963 50336 10005 50345
rect 9963 50296 9964 50336
rect 10004 50296 10005 50336
rect 9963 50287 10005 50296
rect 10059 50336 10101 50345
rect 10059 50296 10060 50336
rect 10100 50296 10101 50336
rect 10059 50287 10101 50296
rect 10339 50336 10397 50337
rect 10339 50296 10348 50336
rect 10388 50296 10397 50336
rect 10339 50295 10397 50296
rect 10819 50336 10877 50337
rect 10819 50296 10828 50336
rect 10868 50296 10877 50336
rect 10819 50295 10877 50296
rect 12067 50336 12125 50337
rect 12067 50296 12076 50336
rect 12116 50296 12125 50336
rect 12067 50295 12125 50296
rect 12555 50336 12597 50345
rect 12555 50296 12556 50336
rect 12596 50296 12597 50336
rect 12555 50287 12597 50296
rect 12651 50336 12693 50345
rect 12651 50296 12652 50336
rect 12692 50296 12693 50336
rect 13603 50336 13661 50337
rect 12651 50287 12693 50296
rect 13131 50294 13173 50303
rect 13603 50296 13612 50336
rect 13652 50296 13661 50336
rect 14467 50336 14525 50337
rect 13603 50295 13661 50296
rect 14139 50326 14181 50335
rect 1699 50252 1757 50253
rect 1699 50212 1708 50252
rect 1748 50212 1757 50252
rect 1699 50211 1757 50212
rect 2083 50252 2141 50253
rect 2083 50212 2092 50252
rect 2132 50212 2141 50252
rect 2083 50211 2141 50212
rect 2467 50252 2525 50253
rect 2467 50212 2476 50252
rect 2516 50212 2525 50252
rect 2467 50211 2525 50212
rect 13035 50252 13077 50261
rect 13035 50212 13036 50252
rect 13076 50212 13077 50252
rect 13131 50254 13132 50294
rect 13172 50254 13173 50294
rect 14139 50286 14140 50326
rect 14180 50286 14181 50326
rect 14467 50296 14476 50336
rect 14516 50296 14525 50336
rect 14467 50295 14525 50296
rect 15715 50336 15773 50337
rect 15715 50296 15724 50336
rect 15764 50296 15773 50336
rect 15715 50295 15773 50296
rect 16099 50336 16157 50337
rect 16099 50296 16108 50336
rect 16148 50296 16157 50336
rect 17923 50336 17981 50337
rect 16099 50295 16157 50296
rect 17347 50315 17405 50316
rect 14139 50277 14181 50286
rect 17347 50275 17356 50315
rect 17396 50275 17405 50315
rect 17923 50296 17932 50336
rect 17972 50296 17981 50336
rect 17923 50295 17981 50296
rect 19171 50336 19229 50337
rect 19171 50296 19180 50336
rect 19220 50296 19229 50336
rect 19171 50295 19229 50296
rect 17347 50274 17405 50275
rect 13131 50245 13173 50254
rect 19363 50252 19421 50253
rect 13035 50203 13077 50212
rect 19363 50212 19372 50252
rect 19412 50212 19421 50252
rect 19363 50211 19421 50212
rect 12267 50168 12309 50177
rect 12267 50128 12268 50168
rect 12308 50128 12309 50168
rect 12267 50119 12309 50128
rect 19563 50168 19605 50177
rect 19563 50128 19564 50168
rect 19604 50128 19605 50168
rect 19563 50119 19605 50128
rect 19947 50168 19989 50177
rect 19947 50128 19948 50168
rect 19988 50128 19989 50168
rect 19947 50119 19989 50128
rect 1515 50084 1557 50093
rect 1515 50044 1516 50084
rect 1556 50044 1557 50084
rect 1515 50035 1557 50044
rect 1899 50084 1941 50093
rect 1899 50044 1900 50084
rect 1940 50044 1941 50084
rect 1899 50035 1941 50044
rect 2283 50084 2325 50093
rect 2283 50044 2284 50084
rect 2324 50044 2325 50084
rect 2283 50035 2325 50044
rect 4107 50084 4149 50093
rect 4107 50044 4108 50084
rect 4148 50044 4149 50084
rect 4107 50035 4149 50044
rect 7371 50084 7413 50093
rect 7371 50044 7372 50084
rect 7412 50044 7413 50084
rect 7371 50035 7413 50044
rect 9387 50084 9429 50093
rect 9387 50044 9388 50084
rect 9428 50044 9429 50084
rect 9387 50035 9429 50044
rect 9667 50084 9725 50085
rect 9667 50044 9676 50084
rect 9716 50044 9725 50084
rect 9667 50043 9725 50044
rect 15915 50084 15957 50093
rect 15915 50044 15916 50084
rect 15956 50044 15957 50084
rect 15915 50035 15957 50044
rect 17547 50084 17589 50093
rect 17547 50044 17548 50084
rect 17588 50044 17589 50084
rect 17547 50035 17589 50044
rect 17739 50084 17781 50093
rect 17739 50044 17740 50084
rect 17780 50044 17781 50084
rect 17739 50035 17781 50044
rect 1152 49916 20352 49940
rect 1152 49876 3688 49916
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 4056 49876 18808 49916
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 19176 49876 20352 49916
rect 1152 49852 20352 49876
rect 8139 49748 8181 49757
rect 8139 49708 8140 49748
rect 8180 49708 8181 49748
rect 8139 49699 8181 49708
rect 8907 49580 8949 49589
rect 8907 49540 8908 49580
rect 8948 49540 8949 49580
rect 8907 49531 8949 49540
rect 9003 49580 9045 49589
rect 9003 49540 9004 49580
rect 9044 49540 9045 49580
rect 9003 49531 9045 49540
rect 18603 49580 18645 49589
rect 18603 49540 18604 49580
rect 18644 49540 18645 49580
rect 18603 49531 18645 49540
rect 19611 49538 19653 49547
rect 4299 49510 4341 49519
rect 2763 49496 2805 49505
rect 2763 49456 2764 49496
rect 2804 49456 2805 49496
rect 2763 49447 2805 49456
rect 2859 49496 2901 49505
rect 2859 49456 2860 49496
rect 2900 49456 2901 49496
rect 2859 49447 2901 49456
rect 3243 49496 3285 49505
rect 3243 49456 3244 49496
rect 3284 49456 3285 49496
rect 3243 49447 3285 49456
rect 3339 49496 3381 49505
rect 3339 49456 3340 49496
rect 3380 49456 3381 49496
rect 3339 49447 3381 49456
rect 3811 49496 3869 49497
rect 3811 49456 3820 49496
rect 3860 49456 3869 49496
rect 4299 49470 4300 49510
rect 4340 49470 4341 49510
rect 9963 49510 10005 49519
rect 4299 49461 4341 49470
rect 4675 49496 4733 49497
rect 3811 49455 3869 49456
rect 4675 49456 4684 49496
rect 4724 49456 4733 49496
rect 4675 49455 4733 49456
rect 5923 49496 5981 49497
rect 5923 49456 5932 49496
rect 5972 49456 5981 49496
rect 5923 49455 5981 49456
rect 6691 49496 6749 49497
rect 6691 49456 6700 49496
rect 6740 49456 6749 49496
rect 6691 49455 6749 49456
rect 7939 49496 7997 49497
rect 7939 49456 7948 49496
rect 7988 49456 7997 49496
rect 7939 49455 7997 49456
rect 8427 49496 8469 49505
rect 8427 49456 8428 49496
rect 8468 49456 8469 49496
rect 8427 49447 8469 49456
rect 8523 49496 8565 49505
rect 8523 49456 8524 49496
rect 8564 49456 8565 49496
rect 8523 49447 8565 49456
rect 9475 49496 9533 49497
rect 9475 49456 9484 49496
rect 9524 49456 9533 49496
rect 9963 49470 9964 49510
rect 10004 49470 10005 49510
rect 9963 49461 10005 49470
rect 10347 49496 10389 49505
rect 9475 49455 9533 49456
rect 10347 49456 10348 49496
rect 10388 49456 10389 49496
rect 10347 49447 10389 49456
rect 10443 49496 10485 49505
rect 10443 49456 10444 49496
rect 10484 49456 10485 49496
rect 10443 49447 10485 49456
rect 10539 49504 10581 49513
rect 14523 49505 14565 49514
rect 10539 49464 10540 49504
rect 10580 49464 10581 49504
rect 10539 49455 10581 49464
rect 10827 49496 10869 49505
rect 10827 49456 10828 49496
rect 10868 49456 10869 49496
rect 10827 49447 10869 49456
rect 11019 49496 11061 49505
rect 11019 49456 11020 49496
rect 11060 49456 11061 49496
rect 11019 49447 11061 49456
rect 11203 49496 11261 49497
rect 11203 49456 11212 49496
rect 11252 49456 11261 49496
rect 11203 49455 11261 49456
rect 12451 49496 12509 49497
rect 12451 49456 12460 49496
rect 12500 49456 12509 49496
rect 12451 49455 12509 49456
rect 12939 49496 12981 49505
rect 12939 49456 12940 49496
rect 12980 49456 12981 49496
rect 12939 49447 12981 49456
rect 13035 49496 13077 49505
rect 13035 49456 13036 49496
rect 13076 49456 13077 49496
rect 13035 49447 13077 49456
rect 13419 49496 13461 49505
rect 13419 49456 13420 49496
rect 13460 49456 13461 49496
rect 13419 49447 13461 49456
rect 13515 49496 13557 49505
rect 13515 49456 13516 49496
rect 13556 49456 13557 49496
rect 13515 49447 13557 49456
rect 13987 49496 14045 49497
rect 13987 49456 13996 49496
rect 14036 49456 14045 49496
rect 14523 49465 14524 49505
rect 14564 49465 14565 49505
rect 14523 49456 14565 49465
rect 15043 49496 15101 49497
rect 15043 49456 15052 49496
rect 15092 49456 15101 49496
rect 13987 49455 14045 49456
rect 15043 49455 15101 49456
rect 16291 49496 16349 49497
rect 16291 49456 16300 49496
rect 16340 49456 16349 49496
rect 16291 49455 16349 49456
rect 18027 49496 18069 49505
rect 18027 49456 18028 49496
rect 18068 49456 18069 49496
rect 18027 49447 18069 49456
rect 18123 49496 18165 49505
rect 18123 49456 18124 49496
rect 18164 49456 18165 49496
rect 18123 49447 18165 49456
rect 18507 49496 18549 49505
rect 19611 49498 19612 49538
rect 19652 49498 19653 49538
rect 18507 49456 18508 49496
rect 18548 49456 18549 49496
rect 18507 49447 18549 49456
rect 19075 49496 19133 49497
rect 19075 49456 19084 49496
rect 19124 49456 19133 49496
rect 19611 49489 19653 49498
rect 19075 49455 19133 49456
rect 10155 49412 10197 49421
rect 10155 49372 10156 49412
rect 10196 49372 10197 49412
rect 10155 49363 10197 49372
rect 12651 49412 12693 49421
rect 12651 49372 12652 49412
rect 12692 49372 12693 49412
rect 12651 49363 12693 49372
rect 14859 49412 14901 49421
rect 14859 49372 14860 49412
rect 14900 49372 14901 49412
rect 14859 49363 14901 49372
rect 4491 49328 4533 49337
rect 4491 49288 4492 49328
rect 4532 49288 4533 49328
rect 4491 49279 4533 49288
rect 6123 49328 6165 49337
rect 6123 49288 6124 49328
rect 6164 49288 6165 49328
rect 6123 49279 6165 49288
rect 10627 49328 10685 49329
rect 10627 49288 10636 49328
rect 10676 49288 10685 49328
rect 10627 49287 10685 49288
rect 10923 49328 10965 49337
rect 10923 49288 10924 49328
rect 10964 49288 10965 49328
rect 10923 49279 10965 49288
rect 14667 49328 14709 49337
rect 14667 49288 14668 49328
rect 14708 49288 14709 49328
rect 14667 49279 14709 49288
rect 19755 49286 19797 49295
rect 19755 49246 19756 49286
rect 19796 49246 19797 49286
rect 19755 49237 19797 49246
rect 1152 49160 20452 49184
rect 1152 49120 4928 49160
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 5296 49120 20048 49160
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20416 49120 20452 49160
rect 1152 49096 20452 49120
rect 1899 48992 1941 49001
rect 1899 48952 1900 48992
rect 1940 48952 1941 48992
rect 1899 48943 1941 48952
rect 9867 48992 9909 49001
rect 9867 48952 9868 48992
rect 9908 48952 9909 48992
rect 9867 48943 9909 48952
rect 10339 48992 10397 48993
rect 10339 48952 10348 48992
rect 10388 48952 10397 48992
rect 10339 48951 10397 48952
rect 7659 48908 7701 48917
rect 7659 48868 7660 48908
rect 7700 48868 7701 48908
rect 7659 48859 7701 48868
rect 17259 48908 17301 48917
rect 17259 48868 17260 48908
rect 17300 48868 17301 48908
rect 17259 48859 17301 48868
rect 19755 48908 19797 48917
rect 19755 48868 19756 48908
rect 19796 48868 19797 48908
rect 19755 48859 19797 48868
rect 2563 48824 2621 48825
rect 2563 48784 2572 48824
rect 2612 48784 2621 48824
rect 2563 48783 2621 48784
rect 3811 48824 3869 48825
rect 3811 48784 3820 48824
rect 3860 48784 3869 48824
rect 3811 48783 3869 48784
rect 4195 48824 4253 48825
rect 4195 48784 4204 48824
rect 4244 48784 4253 48824
rect 4195 48783 4253 48784
rect 5443 48824 5501 48825
rect 5443 48784 5452 48824
rect 5492 48784 5501 48824
rect 5443 48783 5501 48784
rect 5931 48824 5973 48833
rect 5931 48784 5932 48824
rect 5972 48784 5973 48824
rect 5931 48775 5973 48784
rect 6027 48824 6069 48833
rect 6027 48784 6028 48824
rect 6068 48784 6069 48824
rect 6027 48775 6069 48784
rect 6507 48824 6549 48833
rect 6507 48784 6508 48824
rect 6548 48784 6549 48824
rect 6507 48775 6549 48784
rect 6979 48824 7037 48825
rect 6979 48784 6988 48824
rect 7028 48784 7037 48824
rect 6979 48783 7037 48784
rect 7467 48819 7509 48828
rect 7467 48779 7468 48819
rect 7508 48779 7509 48819
rect 7939 48824 7997 48825
rect 7939 48784 7948 48824
rect 7988 48784 7997 48824
rect 7939 48783 7997 48784
rect 8043 48824 8085 48833
rect 8043 48784 8044 48824
rect 8084 48784 8085 48824
rect 7467 48770 7509 48779
rect 8043 48775 8085 48784
rect 8235 48824 8277 48833
rect 8235 48784 8236 48824
rect 8276 48784 8277 48824
rect 8235 48775 8277 48784
rect 8419 48824 8477 48825
rect 8419 48784 8428 48824
rect 8468 48784 8477 48824
rect 8419 48783 8477 48784
rect 9667 48824 9725 48825
rect 9667 48784 9676 48824
rect 9716 48784 9725 48824
rect 9667 48783 9725 48784
rect 10059 48824 10101 48833
rect 10059 48784 10060 48824
rect 10100 48784 10101 48824
rect 10059 48775 10101 48784
rect 10155 48824 10197 48833
rect 10155 48784 10156 48824
rect 10196 48784 10197 48824
rect 10155 48775 10197 48784
rect 10251 48824 10293 48833
rect 10251 48784 10252 48824
rect 10292 48784 10293 48824
rect 10251 48775 10293 48784
rect 10627 48824 10685 48825
rect 10627 48784 10636 48824
rect 10676 48784 10685 48824
rect 10627 48783 10685 48784
rect 11875 48824 11933 48825
rect 11875 48784 11884 48824
rect 11924 48784 11933 48824
rect 11875 48783 11933 48784
rect 13123 48824 13181 48825
rect 13123 48784 13132 48824
rect 13172 48784 13181 48824
rect 13123 48783 13181 48784
rect 14371 48824 14429 48825
rect 14371 48784 14380 48824
rect 14420 48784 14429 48824
rect 14371 48783 14429 48784
rect 15531 48824 15573 48833
rect 15531 48784 15532 48824
rect 15572 48784 15573 48824
rect 15531 48775 15573 48784
rect 15627 48824 15669 48833
rect 15627 48784 15628 48824
rect 15668 48784 15669 48824
rect 15627 48775 15669 48784
rect 16107 48824 16149 48833
rect 16107 48784 16108 48824
rect 16148 48784 16149 48824
rect 16107 48775 16149 48784
rect 16579 48824 16637 48825
rect 16579 48784 16588 48824
rect 16628 48784 16637 48824
rect 18027 48824 18069 48833
rect 16579 48783 16637 48784
rect 17115 48814 17157 48823
rect 17115 48774 17116 48814
rect 17156 48774 17157 48814
rect 18027 48784 18028 48824
rect 18068 48784 18069 48824
rect 18027 48775 18069 48784
rect 18123 48824 18165 48833
rect 18123 48784 18124 48824
rect 18164 48784 18165 48824
rect 18123 48775 18165 48784
rect 18507 48824 18549 48833
rect 18507 48784 18508 48824
rect 18548 48784 18549 48824
rect 18507 48775 18549 48784
rect 18603 48824 18645 48833
rect 18603 48784 18604 48824
rect 18644 48784 18645 48824
rect 18603 48775 18645 48784
rect 19075 48824 19133 48825
rect 19075 48784 19084 48824
rect 19124 48784 19133 48824
rect 19075 48783 19133 48784
rect 19611 48814 19653 48823
rect 17115 48765 17157 48774
rect 19611 48774 19612 48814
rect 19652 48774 19653 48814
rect 19611 48765 19653 48774
rect 1699 48740 1757 48741
rect 1699 48700 1708 48740
rect 1748 48700 1757 48740
rect 1699 48699 1757 48700
rect 2083 48740 2141 48741
rect 2083 48700 2092 48740
rect 2132 48700 2141 48740
rect 2083 48699 2141 48700
rect 6411 48740 6453 48749
rect 6411 48700 6412 48740
rect 6452 48700 6453 48740
rect 6411 48691 6453 48700
rect 16011 48740 16053 48749
rect 16011 48700 16012 48740
rect 16052 48700 16053 48740
rect 16011 48691 16053 48700
rect 1515 48572 1557 48581
rect 1515 48532 1516 48572
rect 1556 48532 1557 48572
rect 1515 48523 1557 48532
rect 4011 48572 4053 48581
rect 4011 48532 4012 48572
rect 4052 48532 4053 48572
rect 4011 48523 4053 48532
rect 5643 48572 5685 48581
rect 5643 48532 5644 48572
rect 5684 48532 5685 48572
rect 5643 48523 5685 48532
rect 8235 48572 8277 48581
rect 8235 48532 8236 48572
rect 8276 48532 8277 48572
rect 8235 48523 8277 48532
rect 12075 48572 12117 48581
rect 12075 48532 12076 48572
rect 12116 48532 12117 48572
rect 12075 48523 12117 48532
rect 14571 48572 14613 48581
rect 14571 48532 14572 48572
rect 14612 48532 14613 48572
rect 14571 48523 14613 48532
rect 1152 48404 20352 48428
rect 1152 48364 3688 48404
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 4056 48364 18808 48404
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 19176 48364 20352 48404
rect 1152 48340 20352 48364
rect 1515 48236 1557 48245
rect 1515 48196 1516 48236
rect 1556 48196 1557 48236
rect 1515 48187 1557 48196
rect 1699 48068 1757 48069
rect 1699 48028 1708 48068
rect 1748 48028 1757 48068
rect 1699 48027 1757 48028
rect 2083 48068 2141 48069
rect 2083 48028 2092 48068
rect 2132 48028 2141 48068
rect 2083 48027 2141 48028
rect 2467 48068 2525 48069
rect 2467 48028 2476 48068
rect 2516 48028 2525 48068
rect 2467 48027 2525 48028
rect 3339 48068 3381 48077
rect 3339 48028 3340 48068
rect 3380 48028 3381 48068
rect 3339 48019 3381 48028
rect 8715 48068 8757 48077
rect 8715 48028 8716 48068
rect 8756 48028 8757 48068
rect 8715 48019 8757 48028
rect 10243 48026 10301 48027
rect 4299 47998 4341 48007
rect 2763 47984 2805 47993
rect 2763 47944 2764 47984
rect 2804 47944 2805 47984
rect 2763 47935 2805 47944
rect 2859 47984 2901 47993
rect 2859 47944 2860 47984
rect 2900 47944 2901 47984
rect 2859 47935 2901 47944
rect 3243 47984 3285 47993
rect 3243 47944 3244 47984
rect 3284 47944 3285 47984
rect 3243 47935 3285 47944
rect 3811 47984 3869 47985
rect 3811 47944 3820 47984
rect 3860 47944 3869 47984
rect 4299 47958 4300 47998
rect 4340 47958 4341 47998
rect 4299 47949 4341 47958
rect 4771 47984 4829 47985
rect 3811 47943 3869 47944
rect 4771 47944 4780 47984
rect 4820 47944 4829 47984
rect 4771 47943 4829 47944
rect 6019 47984 6077 47985
rect 6019 47944 6028 47984
rect 6068 47944 6077 47984
rect 6019 47943 6077 47944
rect 6403 47984 6461 47985
rect 6403 47944 6412 47984
rect 6452 47944 6461 47984
rect 6403 47943 6461 47944
rect 7651 47984 7709 47985
rect 7651 47944 7660 47984
rect 7700 47944 7709 47984
rect 7651 47943 7709 47944
rect 8619 47984 8661 47993
rect 8619 47944 8620 47984
rect 8660 47944 8661 47984
rect 8619 47935 8661 47944
rect 8811 47984 8853 47993
rect 10243 47986 10252 48026
rect 10292 47986 10301 48026
rect 14283 47998 14325 48007
rect 10243 47985 10301 47986
rect 8811 47944 8812 47984
rect 8852 47944 8853 47984
rect 8811 47935 8853 47944
rect 8995 47984 9053 47985
rect 8995 47944 9004 47984
rect 9044 47944 9053 47984
rect 8995 47943 9053 47944
rect 11011 47984 11069 47985
rect 11011 47944 11020 47984
rect 11060 47944 11069 47984
rect 11011 47943 11069 47944
rect 12259 47984 12317 47985
rect 12259 47944 12268 47984
rect 12308 47944 12317 47984
rect 12259 47943 12317 47944
rect 12747 47984 12789 47993
rect 12747 47944 12748 47984
rect 12788 47944 12789 47984
rect 12747 47935 12789 47944
rect 12843 47984 12885 47993
rect 12843 47944 12844 47984
rect 12884 47944 12885 47984
rect 12843 47935 12885 47944
rect 13227 47984 13269 47993
rect 13227 47944 13228 47984
rect 13268 47944 13269 47984
rect 13227 47935 13269 47944
rect 13323 47984 13365 47993
rect 13323 47944 13324 47984
rect 13364 47944 13365 47984
rect 13323 47935 13365 47944
rect 13795 47984 13853 47985
rect 13795 47944 13804 47984
rect 13844 47944 13853 47984
rect 14283 47958 14284 47998
rect 14324 47958 14325 47998
rect 14283 47949 14325 47958
rect 14659 47984 14717 47985
rect 13795 47943 13853 47944
rect 14659 47944 14668 47984
rect 14708 47944 14717 47984
rect 14659 47943 14717 47944
rect 15907 47984 15965 47985
rect 15907 47944 15916 47984
rect 15956 47944 15965 47984
rect 15907 47943 15965 47944
rect 16483 47984 16541 47985
rect 16483 47944 16492 47984
rect 16532 47944 16541 47984
rect 16483 47943 16541 47944
rect 17731 47984 17789 47985
rect 17731 47944 17740 47984
rect 17780 47944 17789 47984
rect 17731 47943 17789 47944
rect 18115 47984 18173 47985
rect 18115 47944 18124 47984
rect 18164 47944 18173 47984
rect 18115 47943 18173 47944
rect 19363 47984 19421 47985
rect 19363 47944 19372 47984
rect 19412 47944 19421 47984
rect 19363 47943 19421 47944
rect 4491 47900 4533 47909
rect 4491 47860 4492 47900
rect 4532 47860 4533 47900
rect 4491 47851 4533 47860
rect 12459 47900 12501 47909
rect 12459 47860 12460 47900
rect 12500 47860 12501 47900
rect 12459 47851 12501 47860
rect 1899 47816 1941 47825
rect 1899 47776 1900 47816
rect 1940 47776 1941 47816
rect 1899 47767 1941 47776
rect 2283 47816 2325 47825
rect 2283 47776 2284 47816
rect 2324 47776 2325 47816
rect 2283 47767 2325 47776
rect 6219 47816 6261 47825
rect 6219 47776 6220 47816
rect 6260 47776 6261 47816
rect 6219 47767 6261 47776
rect 7851 47816 7893 47825
rect 7851 47776 7852 47816
rect 7892 47776 7893 47816
rect 7851 47767 7893 47776
rect 10443 47816 10485 47825
rect 10443 47776 10444 47816
rect 10484 47776 10485 47816
rect 10443 47767 10485 47776
rect 14475 47816 14517 47825
rect 14475 47776 14476 47816
rect 14516 47776 14517 47816
rect 14475 47767 14517 47776
rect 16107 47816 16149 47825
rect 16107 47776 16108 47816
rect 16148 47776 16149 47816
rect 16107 47767 16149 47776
rect 16299 47816 16341 47825
rect 16299 47776 16300 47816
rect 16340 47776 16341 47816
rect 16299 47767 16341 47776
rect 17931 47816 17973 47825
rect 17931 47776 17932 47816
rect 17972 47776 17973 47816
rect 17931 47767 17973 47776
rect 1152 47648 20452 47672
rect 1152 47608 4928 47648
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 5296 47608 20048 47648
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20416 47608 20452 47648
rect 1152 47584 20452 47608
rect 7947 47480 7989 47489
rect 7947 47440 7948 47480
rect 7988 47440 7989 47480
rect 7947 47431 7989 47440
rect 12075 47480 12117 47489
rect 12075 47440 12076 47480
rect 12116 47440 12117 47480
rect 12075 47431 12117 47440
rect 3339 47396 3381 47405
rect 3339 47356 3340 47396
rect 3380 47356 3381 47396
rect 3339 47347 3381 47356
rect 5547 47396 5589 47405
rect 5547 47356 5548 47396
rect 5588 47356 5589 47396
rect 5547 47347 5589 47356
rect 17163 47396 17205 47405
rect 17163 47356 17164 47396
rect 17204 47356 17205 47396
rect 17163 47347 17205 47356
rect 20043 47396 20085 47405
rect 20043 47356 20044 47396
rect 20084 47356 20085 47396
rect 20043 47347 20085 47356
rect 1891 47312 1949 47313
rect 1891 47272 1900 47312
rect 1940 47272 1949 47312
rect 1891 47271 1949 47272
rect 3139 47312 3197 47313
rect 3139 47272 3148 47312
rect 3188 47272 3197 47312
rect 3139 47271 3197 47272
rect 3819 47312 3861 47321
rect 3819 47272 3820 47312
rect 3860 47272 3861 47312
rect 3819 47263 3861 47272
rect 3915 47312 3957 47321
rect 3915 47272 3916 47312
rect 3956 47272 3957 47312
rect 3915 47263 3957 47272
rect 4299 47312 4341 47321
rect 4299 47272 4300 47312
rect 4340 47272 4341 47312
rect 4299 47263 4341 47272
rect 4395 47312 4437 47321
rect 4395 47272 4396 47312
rect 4436 47272 4437 47312
rect 4395 47263 4437 47272
rect 4867 47312 4925 47313
rect 4867 47272 4876 47312
rect 4916 47272 4925 47312
rect 6219 47312 6261 47321
rect 4867 47271 4925 47272
rect 5403 47302 5445 47311
rect 5403 47262 5404 47302
rect 5444 47262 5445 47302
rect 6219 47272 6220 47312
rect 6260 47272 6261 47312
rect 6219 47263 6261 47272
rect 6315 47312 6357 47321
rect 6315 47272 6316 47312
rect 6356 47272 6357 47312
rect 6315 47263 6357 47272
rect 6699 47312 6741 47321
rect 6699 47272 6700 47312
rect 6740 47272 6741 47312
rect 6699 47263 6741 47272
rect 6795 47312 6837 47321
rect 6795 47272 6796 47312
rect 6836 47272 6837 47312
rect 6795 47263 6837 47272
rect 7267 47312 7325 47313
rect 7267 47272 7276 47312
rect 7316 47272 7325 47312
rect 8515 47312 8573 47313
rect 7267 47271 7325 47272
rect 7803 47302 7845 47311
rect 5403 47253 5445 47262
rect 7803 47262 7804 47302
rect 7844 47262 7845 47302
rect 8515 47272 8524 47312
rect 8564 47272 8573 47312
rect 8515 47271 8573 47272
rect 9763 47312 9821 47313
rect 9763 47272 9772 47312
rect 9812 47272 9821 47312
rect 9763 47271 9821 47272
rect 10347 47312 10389 47321
rect 10347 47272 10348 47312
rect 10388 47272 10389 47312
rect 10347 47263 10389 47272
rect 10443 47312 10485 47321
rect 10443 47272 10444 47312
rect 10484 47272 10485 47312
rect 10443 47263 10485 47272
rect 10923 47312 10965 47321
rect 10923 47272 10924 47312
rect 10964 47272 10965 47312
rect 10923 47263 10965 47272
rect 11395 47312 11453 47313
rect 11395 47272 11404 47312
rect 11444 47272 11453 47312
rect 12931 47312 12989 47313
rect 11395 47271 11453 47272
rect 11931 47302 11973 47311
rect 7803 47253 7845 47262
rect 11931 47262 11932 47302
rect 11972 47262 11973 47302
rect 12931 47272 12940 47312
rect 12980 47272 12989 47312
rect 12931 47271 12989 47272
rect 14179 47312 14237 47313
rect 14179 47272 14188 47312
rect 14228 47272 14237 47312
rect 14179 47271 14237 47272
rect 15435 47312 15477 47321
rect 15435 47272 15436 47312
rect 15476 47272 15477 47312
rect 15435 47263 15477 47272
rect 15531 47312 15573 47321
rect 15531 47272 15532 47312
rect 15572 47272 15573 47312
rect 15531 47263 15573 47272
rect 15915 47312 15957 47321
rect 15915 47272 15916 47312
rect 15956 47272 15957 47312
rect 15915 47263 15957 47272
rect 16011 47312 16053 47321
rect 16011 47272 16012 47312
rect 16052 47272 16053 47312
rect 16011 47263 16053 47272
rect 16483 47312 16541 47313
rect 16483 47272 16492 47312
rect 16532 47272 16541 47312
rect 16483 47271 16541 47272
rect 16971 47307 17013 47316
rect 16971 47267 16972 47307
rect 17012 47267 17013 47307
rect 11931 47253 11973 47262
rect 16971 47258 17013 47267
rect 18315 47312 18357 47321
rect 18315 47272 18316 47312
rect 18356 47272 18357 47312
rect 18315 47263 18357 47272
rect 18411 47312 18453 47321
rect 18411 47272 18412 47312
rect 18452 47272 18453 47312
rect 18411 47263 18453 47272
rect 18795 47312 18837 47321
rect 18795 47272 18796 47312
rect 18836 47272 18837 47312
rect 18795 47263 18837 47272
rect 18891 47312 18933 47321
rect 18891 47272 18892 47312
rect 18932 47272 18933 47312
rect 18891 47263 18933 47272
rect 19363 47312 19421 47313
rect 19363 47272 19372 47312
rect 19412 47272 19421 47312
rect 19363 47271 19421 47272
rect 19851 47298 19893 47307
rect 19851 47258 19852 47298
rect 19892 47258 19893 47298
rect 19851 47249 19893 47258
rect 1699 47228 1757 47229
rect 1699 47188 1708 47228
rect 1748 47188 1757 47228
rect 1699 47187 1757 47188
rect 10827 47228 10869 47237
rect 10827 47188 10828 47228
rect 10868 47188 10869 47228
rect 10827 47179 10869 47188
rect 1515 47060 1557 47069
rect 1515 47020 1516 47060
rect 1556 47020 1557 47060
rect 1515 47011 1557 47020
rect 9963 47060 10005 47069
rect 9963 47020 9964 47060
rect 10004 47020 10005 47060
rect 9963 47011 10005 47020
rect 14379 47060 14421 47069
rect 14379 47020 14380 47060
rect 14420 47020 14421 47060
rect 14379 47011 14421 47020
rect 1152 46892 20352 46916
rect 1152 46852 3688 46892
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 4056 46852 18808 46892
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 19176 46852 20352 46892
rect 1152 46828 20352 46852
rect 2667 46640 2709 46649
rect 2667 46600 2668 46640
rect 2708 46600 2709 46640
rect 2667 46591 2709 46600
rect 3043 46556 3101 46557
rect 3043 46516 3052 46556
rect 3092 46516 3101 46556
rect 3043 46515 3101 46516
rect 3427 46556 3485 46557
rect 3427 46516 3436 46556
rect 3476 46516 3485 46556
rect 3427 46515 3485 46516
rect 8715 46556 8757 46565
rect 8715 46516 8716 46556
rect 8756 46516 8757 46556
rect 18891 46556 18933 46565
rect 8715 46507 8757 46516
rect 9723 46514 9765 46523
rect 1219 46472 1277 46473
rect 1219 46432 1228 46472
rect 1268 46432 1277 46472
rect 1219 46431 1277 46432
rect 2467 46472 2525 46473
rect 2467 46432 2476 46472
rect 2516 46432 2525 46472
rect 2467 46431 2525 46432
rect 4099 46472 4157 46473
rect 4099 46432 4108 46472
rect 4148 46432 4157 46472
rect 4099 46431 4157 46432
rect 5347 46472 5405 46473
rect 5347 46432 5356 46472
rect 5396 46432 5405 46472
rect 5347 46431 5405 46432
rect 6403 46472 6461 46473
rect 6403 46432 6412 46472
rect 6452 46432 6461 46472
rect 6403 46431 6461 46432
rect 7651 46472 7709 46473
rect 7651 46432 7660 46472
rect 7700 46432 7709 46472
rect 7651 46431 7709 46432
rect 8139 46472 8181 46481
rect 8139 46432 8140 46472
rect 8180 46432 8181 46472
rect 8139 46423 8181 46432
rect 8235 46472 8277 46481
rect 8235 46432 8236 46472
rect 8276 46432 8277 46472
rect 8235 46423 8277 46432
rect 8619 46472 8661 46481
rect 9723 46474 9724 46514
rect 9764 46474 9765 46514
rect 18891 46516 18892 46556
rect 18932 46516 18933 46556
rect 18891 46507 18933 46516
rect 18987 46556 19029 46565
rect 18987 46516 18988 46556
rect 19028 46516 19029 46556
rect 18987 46507 19029 46516
rect 14187 46486 14229 46495
rect 8619 46432 8620 46472
rect 8660 46432 8661 46472
rect 8619 46423 8661 46432
rect 9187 46472 9245 46473
rect 9187 46432 9196 46472
rect 9236 46432 9245 46472
rect 9723 46465 9765 46474
rect 10915 46472 10973 46473
rect 9187 46431 9245 46432
rect 10915 46432 10924 46472
rect 10964 46432 10973 46472
rect 10915 46431 10973 46432
rect 12163 46472 12221 46473
rect 12163 46432 12172 46472
rect 12212 46432 12221 46472
rect 12163 46431 12221 46432
rect 12651 46472 12693 46481
rect 12651 46432 12652 46472
rect 12692 46432 12693 46472
rect 12651 46423 12693 46432
rect 12747 46472 12789 46481
rect 12747 46432 12748 46472
rect 12788 46432 12789 46472
rect 12747 46423 12789 46432
rect 13131 46472 13173 46481
rect 13131 46432 13132 46472
rect 13172 46432 13173 46472
rect 13131 46423 13173 46432
rect 13227 46472 13269 46481
rect 13227 46432 13228 46472
rect 13268 46432 13269 46472
rect 13227 46423 13269 46432
rect 13699 46472 13757 46473
rect 13699 46432 13708 46472
rect 13748 46432 13757 46472
rect 14187 46446 14188 46486
rect 14228 46446 14229 46486
rect 14187 46437 14229 46446
rect 15715 46472 15773 46473
rect 13699 46431 13757 46432
rect 15715 46432 15724 46472
rect 15764 46432 15773 46472
rect 15715 46431 15773 46432
rect 16963 46472 17021 46473
rect 16963 46432 16972 46472
rect 17012 46432 17021 46472
rect 16963 46431 17021 46432
rect 18411 46472 18453 46481
rect 18411 46432 18412 46472
rect 18452 46432 18453 46472
rect 18411 46423 18453 46432
rect 18507 46472 18549 46481
rect 19947 46477 19989 46486
rect 18507 46432 18508 46472
rect 18548 46432 18549 46472
rect 18507 46423 18549 46432
rect 19459 46472 19517 46473
rect 19459 46432 19468 46472
rect 19508 46432 19517 46472
rect 19459 46431 19517 46432
rect 19947 46437 19948 46477
rect 19988 46437 19989 46477
rect 19947 46428 19989 46437
rect 7851 46388 7893 46397
rect 7851 46348 7852 46388
rect 7892 46348 7893 46388
rect 7851 46339 7893 46348
rect 9867 46388 9909 46397
rect 9867 46348 9868 46388
rect 9908 46348 9909 46388
rect 9867 46339 9909 46348
rect 12363 46388 12405 46397
rect 12363 46348 12364 46388
rect 12404 46348 12405 46388
rect 12363 46339 12405 46348
rect 14379 46388 14421 46397
rect 14379 46348 14380 46388
rect 14420 46348 14421 46388
rect 14379 46339 14421 46348
rect 2859 46304 2901 46313
rect 2859 46264 2860 46304
rect 2900 46264 2901 46304
rect 2859 46255 2901 46264
rect 3243 46304 3285 46313
rect 3243 46264 3244 46304
rect 3284 46264 3285 46304
rect 3243 46255 3285 46264
rect 5547 46304 5589 46313
rect 5547 46264 5548 46304
rect 5588 46264 5589 46304
rect 5547 46255 5589 46264
rect 17163 46304 17205 46313
rect 17163 46264 17164 46304
rect 17204 46264 17205 46304
rect 17163 46255 17205 46264
rect 20139 46304 20181 46313
rect 20139 46264 20140 46304
rect 20180 46264 20181 46304
rect 20139 46255 20181 46264
rect 1152 46136 20452 46160
rect 1152 46096 4928 46136
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 5296 46096 20048 46136
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20416 46096 20452 46136
rect 1152 46072 20452 46096
rect 2283 45968 2325 45977
rect 2283 45928 2284 45968
rect 2324 45928 2325 45968
rect 2283 45919 2325 45928
rect 18891 45968 18933 45977
rect 18891 45928 18892 45968
rect 18932 45928 18933 45968
rect 18891 45919 18933 45928
rect 4387 45800 4445 45801
rect 4387 45760 4396 45800
rect 4436 45760 4445 45800
rect 4387 45759 4445 45760
rect 5635 45800 5693 45801
rect 5635 45760 5644 45800
rect 5684 45760 5693 45800
rect 5635 45759 5693 45760
rect 8707 45800 8765 45801
rect 8707 45760 8716 45800
rect 8756 45760 8765 45800
rect 8707 45759 8765 45760
rect 9955 45800 10013 45801
rect 9955 45760 9964 45800
rect 10004 45760 10013 45800
rect 9955 45759 10013 45760
rect 10339 45800 10397 45801
rect 10339 45760 10348 45800
rect 10388 45760 10397 45800
rect 10339 45759 10397 45760
rect 11587 45800 11645 45801
rect 11587 45760 11596 45800
rect 11636 45760 11645 45800
rect 11587 45759 11645 45760
rect 14947 45800 15005 45801
rect 14947 45760 14956 45800
rect 14996 45760 15005 45800
rect 14947 45759 15005 45760
rect 15811 45800 15869 45801
rect 15811 45760 15820 45800
rect 15860 45760 15869 45800
rect 15811 45759 15869 45760
rect 17059 45800 17117 45801
rect 17059 45760 17068 45800
rect 17108 45760 17117 45800
rect 17059 45759 17117 45760
rect 17443 45800 17501 45801
rect 17443 45760 17452 45800
rect 17492 45760 17501 45800
rect 17443 45759 17501 45760
rect 18691 45800 18749 45801
rect 18691 45760 18700 45800
rect 18740 45760 18749 45800
rect 18691 45759 18749 45760
rect 13699 45758 13757 45759
rect 13699 45718 13708 45758
rect 13748 45718 13757 45758
rect 13699 45717 13757 45718
rect 1699 45716 1757 45717
rect 1699 45676 1708 45716
rect 1748 45676 1757 45716
rect 1699 45675 1757 45676
rect 2083 45716 2141 45717
rect 2083 45676 2092 45716
rect 2132 45676 2141 45716
rect 2083 45675 2141 45676
rect 2467 45716 2525 45717
rect 2467 45676 2476 45716
rect 2516 45676 2525 45716
rect 2467 45675 2525 45676
rect 2851 45716 2909 45717
rect 2851 45676 2860 45716
rect 2900 45676 2909 45716
rect 2851 45675 2909 45676
rect 19363 45716 19421 45717
rect 19363 45676 19372 45716
rect 19412 45676 19421 45716
rect 19363 45675 19421 45676
rect 19747 45716 19805 45717
rect 19747 45676 19756 45716
rect 19796 45676 19805 45716
rect 19747 45675 19805 45676
rect 1515 45548 1557 45557
rect 1515 45508 1516 45548
rect 1556 45508 1557 45548
rect 1515 45499 1557 45508
rect 1899 45548 1941 45557
rect 1899 45508 1900 45548
rect 1940 45508 1941 45548
rect 1899 45499 1941 45508
rect 2667 45548 2709 45557
rect 2667 45508 2668 45548
rect 2708 45508 2709 45548
rect 2667 45499 2709 45508
rect 5835 45548 5877 45557
rect 5835 45508 5836 45548
rect 5876 45508 5877 45548
rect 5835 45499 5877 45508
rect 10155 45548 10197 45557
rect 10155 45508 10156 45548
rect 10196 45508 10197 45548
rect 10155 45499 10197 45508
rect 11787 45548 11829 45557
rect 11787 45508 11788 45548
rect 11828 45508 11829 45548
rect 11787 45499 11829 45508
rect 15147 45548 15189 45557
rect 15147 45508 15148 45548
rect 15188 45508 15189 45548
rect 15147 45499 15189 45508
rect 17259 45548 17301 45557
rect 17259 45508 17260 45548
rect 17300 45508 17301 45548
rect 17259 45499 17301 45508
rect 19563 45548 19605 45557
rect 19563 45508 19564 45548
rect 19604 45508 19605 45548
rect 19563 45499 19605 45508
rect 19947 45548 19989 45557
rect 19947 45508 19948 45548
rect 19988 45508 19989 45548
rect 19947 45499 19989 45508
rect 1152 45380 20352 45404
rect 1152 45340 3688 45380
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 4056 45340 18808 45380
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 19176 45340 20352 45380
rect 1152 45316 20352 45340
rect 18315 45212 18357 45221
rect 18315 45172 18316 45212
rect 18356 45172 18357 45212
rect 18315 45163 18357 45172
rect 19947 45212 19989 45221
rect 19947 45172 19948 45212
rect 19988 45172 19989 45212
rect 19947 45163 19989 45172
rect 1411 45044 1469 45045
rect 1411 45004 1420 45044
rect 1460 45004 1469 45044
rect 1411 45003 1469 45004
rect 1795 45044 1853 45045
rect 1795 45004 1804 45044
rect 1844 45004 1853 45044
rect 1795 45003 1853 45004
rect 4203 45044 4245 45053
rect 4203 45004 4204 45044
rect 4244 45004 4245 45044
rect 4203 44995 4245 45004
rect 4299 45044 4341 45053
rect 4299 45004 4300 45044
rect 4340 45004 4341 45044
rect 8427 45044 8469 45053
rect 4299 44995 4341 45004
rect 5307 45002 5349 45011
rect 1987 44960 2045 44961
rect 1987 44920 1996 44960
rect 2036 44920 2045 44960
rect 1987 44919 2045 44920
rect 3235 44960 3293 44961
rect 3235 44920 3244 44960
rect 3284 44920 3293 44960
rect 3235 44919 3293 44920
rect 3723 44960 3765 44969
rect 3723 44920 3724 44960
rect 3764 44920 3765 44960
rect 3723 44911 3765 44920
rect 3819 44960 3861 44969
rect 5307 44962 5308 45002
rect 5348 44962 5349 45002
rect 8427 45004 8428 45044
rect 8468 45004 8469 45044
rect 8427 44995 8469 45004
rect 10731 45044 10773 45053
rect 10731 45004 10732 45044
rect 10772 45004 10773 45044
rect 15915 45044 15957 45053
rect 10731 44995 10773 45004
rect 11739 45002 11781 45011
rect 9435 44969 9477 44978
rect 3819 44920 3820 44960
rect 3860 44920 3861 44960
rect 3819 44911 3861 44920
rect 4771 44960 4829 44961
rect 4771 44920 4780 44960
rect 4820 44920 4829 44960
rect 5307 44953 5349 44962
rect 6115 44960 6173 44961
rect 4771 44919 4829 44920
rect 6115 44920 6124 44960
rect 6164 44920 6173 44960
rect 6115 44919 6173 44920
rect 7363 44960 7421 44961
rect 7363 44920 7372 44960
rect 7412 44920 7421 44960
rect 7363 44919 7421 44920
rect 7851 44960 7893 44969
rect 7851 44920 7852 44960
rect 7892 44920 7893 44960
rect 7851 44911 7893 44920
rect 7947 44960 7989 44969
rect 7947 44920 7948 44960
rect 7988 44920 7989 44960
rect 7947 44911 7989 44920
rect 8331 44960 8373 44969
rect 8331 44920 8332 44960
rect 8372 44920 8373 44960
rect 8331 44911 8373 44920
rect 8899 44960 8957 44961
rect 8899 44920 8908 44960
rect 8948 44920 8957 44960
rect 9435 44929 9436 44969
rect 9476 44929 9477 44969
rect 9435 44920 9477 44929
rect 10155 44960 10197 44969
rect 10155 44920 10156 44960
rect 10196 44920 10197 44960
rect 8899 44919 8957 44920
rect 10155 44911 10197 44920
rect 10251 44960 10293 44969
rect 10251 44920 10252 44960
rect 10292 44920 10293 44960
rect 10251 44911 10293 44920
rect 10635 44960 10677 44969
rect 11739 44962 11740 45002
rect 11780 44962 11781 45002
rect 15915 45004 15916 45044
rect 15956 45004 15957 45044
rect 15915 44995 15957 45004
rect 16011 45044 16053 45053
rect 16011 45004 16012 45044
rect 16052 45004 16053 45044
rect 18115 45044 18173 45045
rect 16011 44995 16053 45004
rect 17019 45002 17061 45011
rect 18115 45004 18124 45044
rect 18164 45004 18173 45044
rect 18115 45003 18173 45004
rect 10635 44920 10636 44960
rect 10676 44920 10677 44960
rect 10635 44911 10677 44920
rect 11203 44960 11261 44961
rect 11203 44920 11212 44960
rect 11252 44920 11261 44960
rect 11739 44953 11781 44962
rect 12163 44960 12221 44961
rect 11203 44919 11261 44920
rect 12163 44920 12172 44960
rect 12212 44920 12221 44960
rect 12163 44919 12221 44920
rect 13411 44960 13469 44961
rect 13411 44920 13420 44960
rect 13460 44920 13469 44960
rect 13411 44919 13469 44920
rect 15435 44960 15477 44969
rect 15435 44920 15436 44960
rect 15476 44920 15477 44960
rect 15435 44911 15477 44920
rect 15531 44960 15573 44969
rect 17019 44962 17020 45002
rect 17060 44962 17061 45002
rect 15531 44920 15532 44960
rect 15572 44920 15573 44960
rect 15531 44911 15573 44920
rect 16483 44960 16541 44961
rect 16483 44920 16492 44960
rect 16532 44920 16541 44960
rect 17019 44953 17061 44962
rect 18499 44960 18557 44961
rect 16483 44919 16541 44920
rect 18499 44920 18508 44960
rect 18548 44920 18557 44960
rect 18499 44919 18557 44920
rect 19747 44960 19805 44961
rect 19747 44920 19756 44960
rect 19796 44920 19805 44960
rect 19747 44919 19805 44920
rect 5451 44876 5493 44885
rect 5451 44836 5452 44876
rect 5492 44836 5493 44876
rect 5451 44827 5493 44836
rect 7563 44876 7605 44885
rect 7563 44836 7564 44876
rect 7604 44836 7605 44876
rect 7563 44827 7605 44836
rect 9579 44876 9621 44885
rect 9579 44836 9580 44876
rect 9620 44836 9621 44876
rect 9579 44827 9621 44836
rect 1227 44792 1269 44801
rect 1227 44752 1228 44792
rect 1268 44752 1269 44792
rect 1227 44743 1269 44752
rect 1611 44792 1653 44801
rect 1611 44752 1612 44792
rect 1652 44752 1653 44792
rect 1611 44743 1653 44752
rect 3435 44792 3477 44801
rect 3435 44752 3436 44792
rect 3476 44752 3477 44792
rect 3435 44743 3477 44752
rect 11883 44792 11925 44801
rect 11883 44752 11884 44792
rect 11924 44752 11925 44792
rect 11883 44743 11925 44752
rect 13611 44792 13653 44801
rect 13611 44752 13612 44792
rect 13652 44752 13653 44792
rect 13611 44743 13653 44752
rect 17163 44792 17205 44801
rect 17163 44752 17164 44792
rect 17204 44752 17205 44792
rect 17163 44743 17205 44752
rect 1152 44624 20452 44648
rect 1152 44584 4928 44624
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 5296 44584 20048 44624
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20416 44584 20452 44624
rect 1152 44560 20452 44584
rect 9579 44456 9621 44465
rect 9579 44416 9580 44456
rect 9620 44416 9621 44456
rect 9579 44407 9621 44416
rect 17163 44456 17205 44465
rect 17163 44416 17164 44456
rect 17204 44416 17205 44456
rect 17163 44407 17205 44416
rect 17931 44456 17973 44465
rect 17931 44416 17932 44456
rect 17972 44416 17973 44456
rect 17931 44407 17973 44416
rect 18315 44456 18357 44465
rect 18315 44416 18316 44456
rect 18356 44416 18357 44456
rect 18315 44407 18357 44416
rect 20043 44456 20085 44465
rect 20043 44416 20044 44456
rect 20084 44416 20085 44456
rect 20043 44407 20085 44416
rect 5547 44372 5589 44381
rect 5547 44332 5548 44372
rect 5588 44332 5589 44372
rect 5547 44323 5589 44332
rect 11691 44372 11733 44381
rect 11691 44332 11692 44372
rect 11732 44332 11733 44372
rect 11691 44323 11733 44332
rect 13707 44372 13749 44381
rect 13707 44332 13708 44372
rect 13748 44332 13749 44372
rect 13707 44323 13749 44332
rect 1987 44288 2045 44289
rect 1987 44248 1996 44288
rect 2036 44248 2045 44288
rect 1987 44247 2045 44248
rect 3235 44288 3293 44289
rect 3235 44248 3244 44288
rect 3284 44248 3293 44288
rect 3235 44247 3293 44248
rect 3819 44288 3861 44297
rect 3819 44248 3820 44288
rect 3860 44248 3861 44288
rect 3819 44239 3861 44248
rect 3915 44288 3957 44297
rect 3915 44248 3916 44288
rect 3956 44248 3957 44288
rect 3915 44239 3957 44248
rect 4299 44288 4341 44297
rect 4299 44248 4300 44288
rect 4340 44248 4341 44288
rect 4299 44239 4341 44248
rect 4395 44288 4437 44297
rect 4395 44248 4396 44288
rect 4436 44248 4437 44288
rect 4395 44239 4437 44248
rect 4867 44288 4925 44289
rect 4867 44248 4876 44288
rect 4916 44248 4925 44288
rect 6403 44288 6461 44289
rect 4867 44247 4925 44248
rect 5403 44278 5445 44287
rect 5403 44238 5404 44278
rect 5444 44238 5445 44278
rect 6403 44248 6412 44288
rect 6452 44248 6461 44288
rect 6403 44247 6461 44248
rect 7651 44288 7709 44289
rect 7651 44248 7660 44288
rect 7700 44248 7709 44288
rect 7651 44247 7709 44248
rect 8131 44288 8189 44289
rect 8131 44248 8140 44288
rect 8180 44248 8189 44288
rect 8131 44247 8189 44248
rect 9379 44288 9437 44289
rect 9379 44248 9388 44288
rect 9428 44248 9437 44288
rect 9379 44247 9437 44248
rect 10243 44288 10301 44289
rect 10243 44248 10252 44288
rect 10292 44248 10301 44288
rect 10243 44247 10301 44248
rect 11491 44288 11549 44289
rect 11491 44248 11500 44288
rect 11540 44248 11549 44288
rect 11491 44247 11549 44248
rect 11979 44288 12021 44297
rect 11979 44248 11980 44288
rect 12020 44248 12021 44288
rect 11979 44239 12021 44248
rect 12075 44288 12117 44297
rect 12075 44248 12076 44288
rect 12116 44248 12117 44288
rect 12075 44239 12117 44248
rect 12555 44288 12597 44297
rect 12555 44248 12556 44288
rect 12596 44248 12597 44288
rect 12555 44239 12597 44248
rect 13027 44288 13085 44289
rect 13027 44248 13036 44288
rect 13076 44248 13085 44288
rect 15531 44288 15573 44297
rect 13027 44247 13085 44248
rect 13563 44278 13605 44287
rect 5403 44229 5445 44238
rect 13563 44238 13564 44278
rect 13604 44238 13605 44278
rect 13563 44229 13605 44238
rect 15435 44269 15477 44278
rect 15435 44229 15436 44269
rect 15476 44229 15477 44269
rect 15531 44248 15532 44288
rect 15572 44248 15573 44288
rect 15531 44239 15573 44248
rect 15915 44288 15957 44297
rect 15915 44248 15916 44288
rect 15956 44248 15957 44288
rect 15915 44239 15957 44248
rect 16011 44288 16053 44297
rect 16011 44248 16012 44288
rect 16052 44248 16053 44288
rect 16011 44239 16053 44248
rect 16483 44288 16541 44289
rect 16483 44248 16492 44288
rect 16532 44248 16541 44288
rect 16483 44247 16541 44248
rect 16971 44283 17013 44292
rect 16971 44243 16972 44283
rect 17012 44243 17013 44283
rect 18595 44288 18653 44289
rect 18595 44248 18604 44288
rect 18644 44248 18653 44288
rect 18595 44247 18653 44248
rect 19843 44288 19901 44289
rect 19843 44248 19852 44288
rect 19892 44248 19901 44288
rect 19843 44247 19901 44248
rect 16971 44234 17013 44243
rect 15435 44220 15477 44229
rect 1795 44204 1853 44205
rect 1795 44164 1804 44204
rect 1844 44164 1853 44204
rect 1795 44163 1853 44164
rect 12459 44204 12501 44213
rect 12459 44164 12460 44204
rect 12500 44164 12501 44204
rect 12459 44155 12501 44164
rect 15139 44204 15197 44205
rect 15139 44164 15148 44204
rect 15188 44164 15197 44204
rect 15139 44163 15197 44164
rect 17731 44204 17789 44205
rect 17731 44164 17740 44204
rect 17780 44164 17789 44204
rect 17731 44163 17789 44164
rect 18115 44204 18173 44205
rect 18115 44164 18124 44204
rect 18164 44164 18173 44204
rect 18115 44163 18173 44164
rect 3435 44120 3477 44129
rect 3435 44080 3436 44120
rect 3476 44080 3477 44120
rect 3435 44071 3477 44080
rect 14955 44120 14997 44129
rect 14955 44080 14956 44120
rect 14996 44080 14997 44120
rect 14955 44071 14997 44080
rect 1611 44036 1653 44045
rect 1611 43996 1612 44036
rect 1652 43996 1653 44036
rect 1611 43987 1653 43996
rect 7851 44036 7893 44045
rect 7851 43996 7852 44036
rect 7892 43996 7893 44036
rect 7851 43987 7893 43996
rect 1152 43868 20352 43892
rect 1152 43828 3688 43868
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 4056 43828 18808 43868
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 19176 43828 20352 43868
rect 1152 43804 20352 43828
rect 15243 43700 15285 43709
rect 15243 43660 15244 43700
rect 15284 43660 15285 43700
rect 15243 43651 15285 43660
rect 17739 43700 17781 43709
rect 17739 43660 17740 43700
rect 17780 43660 17781 43700
rect 17739 43651 17781 43660
rect 18795 43700 18837 43709
rect 18795 43660 18796 43700
rect 18836 43660 18837 43700
rect 18795 43651 18837 43660
rect 19563 43700 19605 43709
rect 19563 43660 19564 43700
rect 19604 43660 19605 43700
rect 19563 43651 19605 43660
rect 19947 43700 19989 43709
rect 19947 43660 19948 43700
rect 19988 43660 19989 43700
rect 19947 43651 19989 43660
rect 13131 43616 13173 43625
rect 13131 43576 13132 43616
rect 13172 43576 13173 43616
rect 13131 43567 13173 43576
rect 11875 43532 11933 43533
rect 11875 43492 11884 43532
rect 11924 43492 11933 43532
rect 11875 43491 11933 43492
rect 13315 43532 13373 43533
rect 13315 43492 13324 43532
rect 13364 43492 13373 43532
rect 13315 43491 13373 43492
rect 17539 43532 17597 43533
rect 17539 43492 17548 43532
rect 17588 43492 17597 43532
rect 17539 43491 17597 43492
rect 17923 43532 17981 43533
rect 17923 43492 17932 43532
rect 17972 43492 17981 43532
rect 17923 43491 17981 43492
rect 18595 43532 18653 43533
rect 18595 43492 18604 43532
rect 18644 43492 18653 43532
rect 18595 43491 18653 43492
rect 18979 43532 19037 43533
rect 18979 43492 18988 43532
rect 19028 43492 19037 43532
rect 18979 43491 19037 43492
rect 19363 43532 19421 43533
rect 19363 43492 19372 43532
rect 19412 43492 19421 43532
rect 19363 43491 19421 43492
rect 19747 43532 19805 43533
rect 19747 43492 19756 43532
rect 19796 43492 19805 43532
rect 19747 43491 19805 43492
rect 2179 43448 2237 43449
rect 2179 43408 2188 43448
rect 2228 43408 2237 43448
rect 2179 43407 2237 43408
rect 3427 43448 3485 43449
rect 3427 43408 3436 43448
rect 3476 43408 3485 43448
rect 3427 43407 3485 43408
rect 3811 43448 3869 43449
rect 3811 43408 3820 43448
rect 3860 43408 3869 43448
rect 3811 43407 3869 43408
rect 3915 43448 3957 43457
rect 3915 43408 3916 43448
rect 3956 43408 3957 43448
rect 3915 43399 3957 43408
rect 4107 43448 4149 43457
rect 4107 43408 4108 43448
rect 4148 43408 4149 43448
rect 4107 43399 4149 43408
rect 6411 43448 6453 43457
rect 6411 43408 6412 43448
rect 6452 43408 6453 43448
rect 6411 43399 6453 43408
rect 6595 43448 6653 43449
rect 6595 43408 6604 43448
rect 6644 43408 6653 43448
rect 6595 43407 6653 43408
rect 6787 43448 6845 43449
rect 6787 43408 6796 43448
rect 6836 43408 6845 43448
rect 6787 43407 6845 43408
rect 6891 43448 6933 43457
rect 6891 43408 6892 43448
rect 6932 43408 6933 43448
rect 6891 43399 6933 43408
rect 7083 43448 7125 43457
rect 7083 43408 7084 43448
rect 7124 43408 7125 43448
rect 7083 43399 7125 43408
rect 7275 43448 7317 43457
rect 7275 43408 7276 43448
rect 7316 43408 7317 43448
rect 7275 43399 7317 43408
rect 7371 43448 7413 43457
rect 7371 43408 7372 43448
rect 7412 43408 7413 43448
rect 7371 43399 7413 43408
rect 7747 43448 7805 43449
rect 7747 43408 7756 43448
rect 7796 43408 7805 43448
rect 7747 43407 7805 43408
rect 7851 43448 7893 43457
rect 7851 43408 7852 43448
rect 7892 43408 7893 43448
rect 7851 43399 7893 43408
rect 8043 43448 8085 43457
rect 8043 43408 8044 43448
rect 8084 43408 8085 43448
rect 8043 43399 8085 43408
rect 8235 43448 8277 43457
rect 8235 43408 8236 43448
rect 8276 43408 8277 43448
rect 8235 43399 8277 43408
rect 8323 43448 8381 43449
rect 8323 43408 8332 43448
rect 8372 43408 8381 43448
rect 8323 43407 8381 43408
rect 9379 43448 9437 43449
rect 9379 43408 9388 43448
rect 9428 43408 9437 43448
rect 9379 43407 9437 43408
rect 13795 43448 13853 43449
rect 13795 43408 13804 43448
rect 13844 43408 13853 43448
rect 13795 43407 13853 43408
rect 15043 43448 15101 43449
rect 15043 43408 15052 43448
rect 15092 43408 15101 43448
rect 15043 43407 15101 43408
rect 6507 43364 6549 43373
rect 6507 43324 6508 43364
rect 6548 43324 6549 43364
rect 6507 43315 6549 43324
rect 3627 43280 3669 43289
rect 3627 43240 3628 43280
rect 3668 43240 3669 43280
rect 3627 43231 3669 43240
rect 4003 43280 4061 43281
rect 4003 43240 4012 43280
rect 4052 43240 4061 43280
rect 4003 43239 4061 43240
rect 6979 43280 7037 43281
rect 6979 43240 6988 43280
rect 7028 43240 7037 43280
rect 6979 43239 7037 43240
rect 7555 43280 7613 43281
rect 7555 43240 7564 43280
rect 7604 43240 7613 43280
rect 7555 43239 7613 43240
rect 8131 43280 8189 43281
rect 8131 43240 8140 43280
rect 8180 43240 8189 43280
rect 8131 43239 8189 43240
rect 9291 43280 9333 43289
rect 9291 43240 9292 43280
rect 9332 43240 9333 43280
rect 9291 43231 9333 43240
rect 11691 43280 11733 43289
rect 11691 43240 11692 43280
rect 11732 43240 11733 43280
rect 11691 43231 11733 43240
rect 18123 43280 18165 43289
rect 18123 43240 18124 43280
rect 18164 43240 18165 43280
rect 18123 43231 18165 43240
rect 19179 43280 19221 43289
rect 19179 43240 19180 43280
rect 19220 43240 19221 43280
rect 19179 43231 19221 43240
rect 1152 43112 20452 43136
rect 1152 43072 4928 43112
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 5296 43072 20048 43112
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20416 43072 20452 43112
rect 1152 43048 20452 43072
rect 8515 42944 8573 42945
rect 8515 42904 8524 42944
rect 8564 42904 8573 42944
rect 8515 42903 8573 42904
rect 17355 42944 17397 42953
rect 17355 42904 17356 42944
rect 17396 42904 17397 42944
rect 17355 42895 17397 42904
rect 4779 42860 4821 42869
rect 4779 42820 4780 42860
rect 4820 42820 4821 42860
rect 4779 42811 4821 42820
rect 9483 42860 9525 42869
rect 9483 42820 9484 42860
rect 9524 42820 9525 42860
rect 9483 42811 9525 42820
rect 4203 42797 4245 42806
rect 2763 42776 2805 42785
rect 2763 42736 2764 42776
rect 2804 42736 2805 42776
rect 2763 42727 2805 42736
rect 2955 42776 2997 42785
rect 2955 42736 2956 42776
rect 2996 42736 2997 42776
rect 2955 42727 2997 42736
rect 3043 42776 3101 42777
rect 3043 42736 3052 42776
rect 3092 42736 3101 42776
rect 3043 42735 3101 42736
rect 3243 42776 3285 42785
rect 3243 42736 3244 42776
rect 3284 42736 3285 42776
rect 3243 42727 3285 42736
rect 3435 42776 3477 42785
rect 3435 42736 3436 42776
rect 3476 42736 3477 42776
rect 3435 42727 3477 42736
rect 3531 42776 3573 42785
rect 3531 42736 3532 42776
rect 3572 42736 3573 42776
rect 3531 42727 3573 42736
rect 3723 42776 3765 42785
rect 3723 42736 3724 42776
rect 3764 42736 3765 42776
rect 3723 42727 3765 42736
rect 3819 42776 3861 42785
rect 3819 42736 3820 42776
rect 3860 42736 3861 42776
rect 3819 42727 3861 42736
rect 3915 42776 3957 42785
rect 3915 42736 3916 42776
rect 3956 42736 3957 42776
rect 3915 42727 3957 42736
rect 4011 42776 4053 42785
rect 4011 42736 4012 42776
rect 4052 42736 4053 42776
rect 4203 42757 4204 42797
rect 4244 42757 4245 42797
rect 4203 42748 4245 42757
rect 4299 42797 4341 42806
rect 4299 42757 4300 42797
rect 4340 42757 4341 42797
rect 4299 42748 4341 42757
rect 4395 42776 4437 42785
rect 4011 42727 4053 42736
rect 4395 42736 4396 42776
rect 4436 42736 4437 42776
rect 4395 42727 4437 42736
rect 4491 42776 4533 42785
rect 4491 42736 4492 42776
rect 4532 42736 4533 42776
rect 4491 42727 4533 42736
rect 4675 42776 4733 42777
rect 4675 42736 4684 42776
rect 4724 42736 4733 42776
rect 4675 42735 4733 42736
rect 4875 42776 4917 42785
rect 4875 42736 4876 42776
rect 4916 42736 4917 42776
rect 4875 42727 4917 42736
rect 5251 42776 5309 42777
rect 5251 42736 5260 42776
rect 5300 42736 5309 42776
rect 5251 42735 5309 42736
rect 6499 42776 6557 42777
rect 6499 42736 6508 42776
rect 6548 42736 6557 42776
rect 6499 42735 6557 42736
rect 7371 42776 7413 42785
rect 7371 42736 7372 42776
rect 7412 42736 7413 42776
rect 7371 42727 7413 42736
rect 7747 42776 7805 42777
rect 7747 42736 7756 42776
rect 7796 42736 7805 42776
rect 7747 42735 7805 42736
rect 8139 42776 8181 42785
rect 8139 42736 8140 42776
rect 8180 42736 8181 42776
rect 8139 42727 8181 42736
rect 8323 42776 8381 42777
rect 8323 42736 8332 42776
rect 8372 42736 8381 42776
rect 8323 42735 8381 42736
rect 8419 42776 8477 42777
rect 8419 42736 8428 42776
rect 8468 42736 8477 42776
rect 8419 42735 8477 42736
rect 8619 42776 8661 42785
rect 8619 42736 8620 42776
rect 8660 42736 8661 42776
rect 8619 42727 8661 42736
rect 8715 42776 8757 42785
rect 8715 42736 8716 42776
rect 8756 42736 8757 42776
rect 9099 42776 9141 42785
rect 8715 42727 8757 42736
rect 8872 42761 8914 42770
rect 8872 42721 8873 42761
rect 8913 42721 8914 42761
rect 9099 42736 9100 42776
rect 9140 42736 9141 42776
rect 9099 42727 9141 42736
rect 9283 42776 9341 42777
rect 9283 42736 9292 42776
rect 9332 42736 9341 42776
rect 9283 42735 9341 42736
rect 9667 42776 9725 42777
rect 9667 42736 9676 42776
rect 9716 42736 9725 42776
rect 9667 42735 9725 42736
rect 10915 42776 10973 42777
rect 10915 42736 10924 42776
rect 10964 42736 10973 42776
rect 10915 42735 10973 42736
rect 11491 42776 11549 42777
rect 11491 42736 11500 42776
rect 11540 42736 11549 42776
rect 11491 42735 11549 42736
rect 12739 42776 12797 42777
rect 12739 42736 12748 42776
rect 12788 42736 12797 42776
rect 12739 42735 12797 42736
rect 13123 42776 13181 42777
rect 13123 42736 13132 42776
rect 13172 42736 13181 42776
rect 13123 42735 13181 42736
rect 14371 42776 14429 42777
rect 14371 42736 14380 42776
rect 14420 42736 14429 42776
rect 14371 42735 14429 42736
rect 8872 42712 8914 42721
rect 7851 42692 7893 42701
rect 7851 42652 7852 42692
rect 7892 42652 7893 42692
rect 7851 42643 7893 42652
rect 8043 42692 8085 42701
rect 8043 42652 8044 42692
rect 8084 42652 8085 42692
rect 8043 42643 8085 42652
rect 14947 42692 15005 42693
rect 14947 42652 14956 42692
rect 14996 42652 15005 42692
rect 14947 42651 15005 42652
rect 16099 42692 16157 42693
rect 16099 42652 16108 42692
rect 16148 42652 16157 42692
rect 16099 42651 16157 42652
rect 16579 42692 16637 42693
rect 16579 42652 16588 42692
rect 16628 42652 16637 42692
rect 16579 42651 16637 42652
rect 17155 42692 17213 42693
rect 17155 42652 17164 42692
rect 17204 42652 17213 42692
rect 17155 42651 17213 42652
rect 17731 42692 17789 42693
rect 17731 42652 17740 42692
rect 17780 42652 17789 42692
rect 17731 42651 17789 42652
rect 18115 42692 18173 42693
rect 18115 42652 18124 42692
rect 18164 42652 18173 42692
rect 18115 42651 18173 42652
rect 18787 42692 18845 42693
rect 18787 42652 18796 42692
rect 18836 42652 18845 42692
rect 18787 42651 18845 42652
rect 19363 42692 19421 42693
rect 19363 42652 19372 42692
rect 19412 42652 19421 42692
rect 19363 42651 19421 42652
rect 19747 42692 19805 42693
rect 19747 42652 19756 42692
rect 19796 42652 19805 42692
rect 19747 42651 19805 42652
rect 3339 42608 3381 42617
rect 3339 42568 3340 42608
rect 3380 42568 3381 42608
rect 3339 42559 3381 42568
rect 6987 42608 7029 42617
rect 6987 42568 6988 42608
rect 7028 42568 7029 42608
rect 6987 42559 7029 42568
rect 7371 42608 7413 42617
rect 7371 42568 7372 42608
rect 7412 42568 7413 42608
rect 7371 42559 7413 42568
rect 7947 42608 7989 42617
rect 7947 42568 7948 42608
rect 7988 42568 7989 42608
rect 7947 42559 7989 42568
rect 9195 42608 9237 42617
rect 9195 42568 9196 42608
rect 9236 42568 9237 42608
rect 9195 42559 9237 42568
rect 15147 42608 15189 42617
rect 15147 42568 15148 42608
rect 15188 42568 15189 42608
rect 15147 42559 15189 42568
rect 16299 42608 16341 42617
rect 16299 42568 16300 42608
rect 16340 42568 16341 42608
rect 16299 42559 16341 42568
rect 16779 42608 16821 42617
rect 16779 42568 16780 42608
rect 16820 42568 16821 42608
rect 16779 42559 16821 42568
rect 17931 42608 17973 42617
rect 17931 42568 17932 42608
rect 17972 42568 17973 42608
rect 17931 42559 17973 42568
rect 18315 42608 18357 42617
rect 18315 42568 18316 42608
rect 18356 42568 18357 42608
rect 18315 42559 18357 42568
rect 18987 42608 19029 42617
rect 18987 42568 18988 42608
rect 19028 42568 19029 42608
rect 18987 42559 19029 42568
rect 19563 42608 19605 42617
rect 19563 42568 19564 42608
rect 19604 42568 19605 42608
rect 19563 42559 19605 42568
rect 2763 42524 2805 42533
rect 2763 42484 2764 42524
rect 2804 42484 2805 42524
rect 2763 42475 2805 42484
rect 6699 42524 6741 42533
rect 6699 42484 6700 42524
rect 6740 42484 6741 42524
rect 6699 42475 6741 42484
rect 7563 42524 7605 42533
rect 7563 42484 7564 42524
rect 7604 42484 7605 42524
rect 7563 42475 7605 42484
rect 12939 42524 12981 42533
rect 12939 42484 12940 42524
rect 12980 42484 12981 42524
rect 12939 42475 12981 42484
rect 14571 42524 14613 42533
rect 14571 42484 14572 42524
rect 14612 42484 14613 42524
rect 14571 42475 14613 42484
rect 19947 42524 19989 42533
rect 19947 42484 19948 42524
rect 19988 42484 19989 42524
rect 19947 42475 19989 42484
rect 1152 42356 20352 42380
rect 1152 42316 3688 42356
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 4056 42316 18808 42356
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 19176 42316 20352 42356
rect 1152 42292 20352 42316
rect 15147 42188 15189 42197
rect 15147 42148 15148 42188
rect 15188 42148 15189 42188
rect 15147 42139 15189 42148
rect 17835 42188 17877 42197
rect 17835 42148 17836 42188
rect 17876 42148 17877 42188
rect 17835 42139 17877 42148
rect 18219 42188 18261 42197
rect 18219 42148 18220 42188
rect 18260 42148 18261 42188
rect 18219 42139 18261 42148
rect 18603 42188 18645 42197
rect 18603 42148 18604 42188
rect 18644 42148 18645 42188
rect 18603 42139 18645 42148
rect 18987 42188 19029 42197
rect 18987 42148 18988 42188
rect 19028 42148 19029 42188
rect 18987 42139 19029 42148
rect 19371 42188 19413 42197
rect 19371 42148 19372 42188
rect 19412 42148 19413 42188
rect 19371 42139 19413 42148
rect 20139 42188 20181 42197
rect 20139 42148 20140 42188
rect 20180 42148 20181 42188
rect 20139 42139 20181 42148
rect 3523 42104 3581 42105
rect 3523 42064 3532 42104
rect 3572 42064 3581 42104
rect 3523 42063 3581 42064
rect 4099 42104 4157 42105
rect 4099 42064 4108 42104
rect 4148 42064 4157 42104
rect 4099 42063 4157 42064
rect 4395 42104 4437 42113
rect 4395 42064 4396 42104
rect 4436 42064 4437 42104
rect 4395 42055 4437 42064
rect 14947 42020 15005 42021
rect 14947 41980 14956 42020
rect 14996 41980 15005 42020
rect 14947 41979 15005 41980
rect 17635 42020 17693 42021
rect 17635 41980 17644 42020
rect 17684 41980 17693 42020
rect 17635 41979 17693 41980
rect 18019 42020 18077 42021
rect 18019 41980 18028 42020
rect 18068 41980 18077 42020
rect 18019 41979 18077 41980
rect 18403 42020 18461 42021
rect 18403 41980 18412 42020
rect 18452 41980 18461 42020
rect 18403 41979 18461 41980
rect 18787 42020 18845 42021
rect 18787 41980 18796 42020
rect 18836 41980 18845 42020
rect 18787 41979 18845 41980
rect 19171 42020 19229 42021
rect 19171 41980 19180 42020
rect 19220 41980 19229 42020
rect 19171 41979 19229 41980
rect 19555 42020 19613 42021
rect 19555 41980 19564 42020
rect 19604 41980 19613 42020
rect 19555 41979 19613 41980
rect 19939 42020 19997 42021
rect 19939 41980 19948 42020
rect 19988 41980 19997 42020
rect 19939 41979 19997 41980
rect 6891 41946 6933 41955
rect 1219 41936 1277 41937
rect 1219 41896 1228 41936
rect 1268 41896 1277 41936
rect 1219 41895 1277 41896
rect 2467 41936 2525 41937
rect 2467 41896 2476 41936
rect 2516 41896 2525 41936
rect 2467 41895 2525 41896
rect 2859 41936 2901 41945
rect 2859 41896 2860 41936
rect 2900 41896 2901 41936
rect 2859 41887 2901 41896
rect 3051 41936 3093 41945
rect 3051 41896 3052 41936
rect 3092 41896 3093 41936
rect 3051 41887 3093 41896
rect 3139 41936 3197 41937
rect 3139 41896 3148 41936
rect 3188 41896 3197 41936
rect 3139 41895 3197 41896
rect 3339 41936 3381 41945
rect 3339 41896 3340 41936
rect 3380 41896 3381 41936
rect 3339 41887 3381 41896
rect 3531 41936 3573 41945
rect 3531 41896 3532 41936
rect 3572 41896 3573 41936
rect 3531 41887 3573 41896
rect 3627 41936 3669 41945
rect 3627 41896 3628 41936
rect 3668 41896 3669 41936
rect 3627 41887 3669 41896
rect 3819 41936 3861 41945
rect 3819 41896 3820 41936
rect 3860 41896 3861 41936
rect 3819 41887 3861 41896
rect 4011 41936 4053 41945
rect 4011 41896 4012 41936
rect 4052 41896 4053 41936
rect 4011 41887 4053 41896
rect 4107 41936 4149 41945
rect 4107 41896 4108 41936
rect 4148 41896 4149 41936
rect 4107 41887 4149 41896
rect 4587 41936 4629 41945
rect 4587 41896 4588 41936
rect 4628 41896 4629 41936
rect 4587 41887 4629 41896
rect 4683 41936 4725 41945
rect 4683 41896 4684 41936
rect 4724 41896 4725 41936
rect 4683 41887 4725 41896
rect 4779 41936 4821 41945
rect 4779 41896 4780 41936
rect 4820 41896 4821 41936
rect 4779 41887 4821 41896
rect 4875 41936 4917 41945
rect 4875 41896 4876 41936
rect 4916 41896 4917 41936
rect 4875 41887 4917 41896
rect 5251 41936 5309 41937
rect 5251 41896 5260 41936
rect 5300 41896 5309 41936
rect 5251 41895 5309 41896
rect 6499 41936 6557 41937
rect 6499 41896 6508 41936
rect 6548 41896 6557 41936
rect 6891 41906 6892 41946
rect 6932 41906 6933 41946
rect 14571 41950 14613 41959
rect 6891 41897 6933 41906
rect 6987 41936 7029 41945
rect 6499 41895 6557 41896
rect 6987 41896 6988 41936
rect 7028 41896 7029 41936
rect 6987 41887 7029 41896
rect 7363 41936 7421 41937
rect 7363 41896 7372 41936
rect 7412 41896 7421 41936
rect 7363 41895 7421 41896
rect 7563 41936 7605 41945
rect 7563 41896 7564 41936
rect 7604 41896 7605 41936
rect 7563 41887 7605 41896
rect 7651 41936 7709 41937
rect 7651 41896 7660 41936
rect 7700 41896 7709 41936
rect 7651 41895 7709 41896
rect 8043 41936 8085 41945
rect 8043 41896 8044 41936
rect 8084 41896 8085 41936
rect 8043 41887 8085 41896
rect 8139 41936 8181 41945
rect 8139 41896 8140 41936
rect 8180 41896 8181 41936
rect 8139 41887 8181 41896
rect 8811 41936 8853 41945
rect 8811 41896 8812 41936
rect 8852 41896 8853 41936
rect 8811 41887 8853 41896
rect 8907 41936 8949 41945
rect 8907 41896 8908 41936
rect 8948 41896 8949 41936
rect 8907 41887 8949 41896
rect 9195 41936 9237 41945
rect 9195 41896 9196 41936
rect 9236 41896 9237 41936
rect 9195 41887 9237 41896
rect 9291 41936 9333 41945
rect 9291 41896 9292 41936
rect 9332 41896 9333 41936
rect 9291 41887 9333 41896
rect 9387 41936 9429 41945
rect 9387 41896 9388 41936
rect 9428 41896 9429 41936
rect 9387 41887 9429 41896
rect 9859 41936 9917 41937
rect 9859 41896 9868 41936
rect 9908 41896 9917 41936
rect 9859 41895 9917 41896
rect 11107 41936 11165 41937
rect 11107 41896 11116 41936
rect 11156 41896 11165 41936
rect 11107 41895 11165 41896
rect 11299 41936 11357 41937
rect 11299 41896 11308 41936
rect 11348 41896 11357 41936
rect 11299 41895 11357 41896
rect 12547 41936 12605 41937
rect 12547 41896 12556 41936
rect 12596 41896 12605 41936
rect 12547 41895 12605 41896
rect 13035 41936 13077 41945
rect 13035 41896 13036 41936
rect 13076 41896 13077 41936
rect 13035 41887 13077 41896
rect 13131 41936 13173 41945
rect 13131 41896 13132 41936
rect 13172 41896 13173 41936
rect 13131 41887 13173 41896
rect 13515 41936 13557 41945
rect 13515 41896 13516 41936
rect 13556 41896 13557 41936
rect 13515 41887 13557 41896
rect 13611 41936 13653 41945
rect 13611 41896 13612 41936
rect 13652 41896 13653 41936
rect 13611 41887 13653 41896
rect 14083 41936 14141 41937
rect 14083 41896 14092 41936
rect 14132 41896 14141 41936
rect 14571 41910 14572 41950
rect 14612 41910 14613 41950
rect 17307 41945 17349 41954
rect 14571 41901 14613 41910
rect 15723 41936 15765 41945
rect 14083 41895 14141 41896
rect 15723 41896 15724 41936
rect 15764 41896 15765 41936
rect 15723 41887 15765 41896
rect 15819 41936 15861 41945
rect 15819 41896 15820 41936
rect 15860 41896 15861 41936
rect 15819 41887 15861 41896
rect 16203 41936 16245 41945
rect 16203 41896 16204 41936
rect 16244 41896 16245 41936
rect 16203 41887 16245 41896
rect 16299 41936 16341 41945
rect 16299 41896 16300 41936
rect 16340 41896 16341 41936
rect 16299 41887 16341 41896
rect 16771 41936 16829 41937
rect 16771 41896 16780 41936
rect 16820 41896 16829 41936
rect 17307 41905 17308 41945
rect 17348 41905 17349 41945
rect 17307 41896 17349 41905
rect 16771 41895 16829 41896
rect 2955 41852 2997 41861
rect 2955 41812 2956 41852
rect 2996 41812 2997 41852
rect 2955 41803 2997 41812
rect 6699 41852 6741 41861
rect 6699 41812 6700 41852
rect 6740 41812 6741 41852
rect 6699 41803 6741 41812
rect 8227 41852 8285 41853
rect 8227 41812 8236 41852
rect 8276 41812 8285 41852
rect 8227 41811 8285 41812
rect 14763 41852 14805 41861
rect 14763 41812 14764 41852
rect 14804 41812 14805 41852
rect 14763 41803 14805 41812
rect 17451 41852 17493 41861
rect 17451 41812 17452 41852
rect 17492 41812 17493 41852
rect 17451 41803 17493 41812
rect 2667 41768 2709 41777
rect 2667 41728 2668 41768
rect 2708 41728 2709 41768
rect 2667 41719 2709 41728
rect 7171 41768 7229 41769
rect 7171 41728 7180 41768
rect 7220 41728 7229 41768
rect 7171 41727 7229 41728
rect 7851 41768 7893 41777
rect 7851 41728 7852 41768
rect 7892 41728 7893 41768
rect 7851 41719 7893 41728
rect 8323 41768 8381 41769
rect 8323 41728 8332 41768
rect 8372 41728 8381 41768
rect 8323 41727 8381 41728
rect 8427 41768 8469 41777
rect 8427 41728 8428 41768
rect 8468 41728 8469 41768
rect 8427 41719 8469 41728
rect 8611 41768 8669 41769
rect 8611 41728 8620 41768
rect 8660 41728 8669 41768
rect 8611 41727 8669 41728
rect 9475 41768 9533 41769
rect 9475 41728 9484 41768
rect 9524 41728 9533 41768
rect 9475 41727 9533 41728
rect 9675 41768 9717 41777
rect 9675 41728 9676 41768
rect 9716 41728 9717 41768
rect 9675 41719 9717 41728
rect 12747 41768 12789 41777
rect 12747 41728 12748 41768
rect 12788 41728 12789 41768
rect 12747 41719 12789 41728
rect 19755 41768 19797 41777
rect 19755 41728 19756 41768
rect 19796 41728 19797 41768
rect 19755 41719 19797 41728
rect 1152 41600 20452 41624
rect 1152 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20452 41600
rect 1152 41536 20452 41560
rect 2955 41432 2997 41441
rect 2955 41392 2956 41432
rect 2996 41392 2997 41432
rect 2955 41383 2997 41392
rect 4395 41432 4437 41441
rect 4395 41392 4396 41432
rect 4436 41392 4437 41432
rect 4395 41383 4437 41392
rect 6507 41432 6549 41441
rect 6507 41392 6508 41432
rect 6548 41392 6549 41432
rect 6507 41383 6549 41392
rect 8035 41432 8093 41433
rect 8035 41392 8044 41432
rect 8084 41392 8093 41432
rect 8035 41391 8093 41392
rect 8523 41432 8565 41441
rect 8523 41392 8524 41432
rect 8564 41392 8565 41432
rect 8523 41383 8565 41392
rect 9291 41432 9333 41441
rect 9291 41392 9292 41432
rect 9332 41392 9333 41432
rect 9291 41383 9333 41392
rect 10251 41432 10293 41441
rect 10251 41392 10252 41432
rect 10292 41392 10293 41432
rect 10251 41383 10293 41392
rect 15627 41432 15669 41441
rect 15627 41392 15628 41432
rect 15668 41392 15669 41432
rect 15627 41383 15669 41392
rect 17355 41432 17397 41441
rect 17355 41392 17356 41432
rect 17396 41392 17397 41432
rect 17355 41383 17397 41392
rect 19747 41432 19805 41433
rect 19747 41392 19756 41432
rect 19796 41392 19805 41432
rect 19747 41391 19805 41392
rect 20235 41432 20277 41441
rect 20235 41392 20236 41432
rect 20276 41392 20277 41432
rect 20235 41383 20277 41392
rect 7939 41348 7997 41349
rect 7939 41308 7948 41348
rect 7988 41308 7997 41348
rect 7939 41307 7997 41308
rect 10731 41348 10773 41357
rect 10731 41308 10732 41348
rect 10772 41308 10773 41348
rect 10731 41299 10773 41308
rect 11115 41285 11157 41294
rect 1219 41264 1277 41265
rect 1219 41224 1228 41264
rect 1268 41224 1277 41264
rect 1219 41223 1277 41224
rect 2467 41264 2525 41265
rect 2467 41224 2476 41264
rect 2516 41224 2525 41264
rect 2467 41223 2525 41224
rect 2851 41264 2909 41265
rect 2851 41224 2860 41264
rect 2900 41224 2909 41264
rect 2851 41223 2909 41224
rect 3147 41264 3189 41273
rect 3147 41224 3148 41264
rect 3188 41224 3189 41264
rect 3147 41215 3189 41224
rect 3339 41264 3381 41273
rect 3339 41224 3340 41264
rect 3380 41224 3381 41264
rect 3339 41215 3381 41224
rect 3435 41264 3477 41273
rect 3435 41224 3436 41264
rect 3476 41224 3477 41264
rect 3435 41215 3477 41224
rect 3619 41264 3677 41265
rect 3619 41224 3628 41264
rect 3668 41224 3677 41264
rect 3619 41223 3677 41224
rect 4011 41264 4053 41273
rect 4011 41224 4012 41264
rect 4052 41224 4053 41264
rect 4011 41215 4053 41224
rect 4203 41264 4245 41273
rect 4203 41224 4204 41264
rect 4244 41224 4245 41264
rect 4203 41215 4245 41224
rect 4306 41263 4348 41272
rect 4306 41223 4307 41263
rect 4347 41223 4348 41263
rect 4306 41214 4348 41223
rect 4491 41264 4533 41273
rect 4491 41224 4492 41264
rect 4532 41224 4533 41264
rect 4491 41215 4533 41224
rect 4675 41264 4733 41265
rect 4675 41224 4684 41264
rect 4724 41224 4733 41264
rect 4675 41223 4733 41224
rect 4779 41264 4821 41273
rect 4779 41224 4780 41264
rect 4820 41224 4821 41264
rect 4779 41215 4821 41224
rect 4875 41264 4917 41273
rect 4875 41224 4876 41264
rect 4916 41224 4917 41264
rect 4875 41215 4917 41224
rect 5059 41264 5117 41265
rect 5059 41224 5068 41264
rect 5108 41224 5117 41264
rect 5059 41223 5117 41224
rect 6307 41264 6365 41265
rect 6307 41224 6316 41264
rect 6356 41224 6365 41264
rect 6307 41223 6365 41224
rect 6691 41264 6749 41265
rect 6691 41224 6700 41264
rect 6740 41224 6749 41264
rect 6691 41223 6749 41224
rect 6987 41264 7029 41273
rect 6987 41224 6988 41264
rect 7028 41224 7029 41264
rect 6987 41215 7029 41224
rect 7363 41264 7421 41265
rect 7363 41224 7372 41264
rect 7412 41224 7421 41264
rect 7363 41223 7421 41224
rect 7755 41264 7797 41273
rect 7755 41224 7756 41264
rect 7796 41224 7797 41264
rect 7265 41222 7323 41223
rect 3723 41180 3765 41189
rect 3723 41140 3724 41180
rect 3764 41140 3765 41180
rect 3723 41131 3765 41140
rect 3915 41180 3957 41189
rect 3915 41140 3916 41180
rect 3956 41140 3957 41180
rect 3915 41131 3957 41140
rect 6795 41180 6837 41189
rect 6795 41140 6796 41180
rect 6836 41140 6837 41180
rect 6795 41131 6837 41140
rect 7083 41180 7125 41189
rect 7265 41182 7274 41222
rect 7314 41182 7323 41222
rect 7755 41215 7797 41224
rect 7851 41264 7893 41273
rect 7851 41224 7852 41264
rect 7892 41224 7893 41264
rect 7851 41215 7893 41224
rect 8331 41264 8373 41273
rect 8331 41224 8332 41264
rect 8372 41224 8373 41264
rect 8331 41215 8373 41224
rect 8427 41264 8469 41273
rect 8427 41224 8428 41264
rect 8468 41224 8469 41264
rect 8427 41215 8469 41224
rect 8619 41264 8661 41273
rect 8619 41224 8620 41264
rect 8660 41224 8661 41264
rect 8619 41215 8661 41224
rect 8811 41264 8853 41273
rect 8811 41224 8812 41264
rect 8852 41224 8853 41264
rect 8811 41215 8853 41224
rect 8907 41264 8949 41273
rect 8907 41224 8908 41264
rect 8948 41224 8949 41264
rect 8907 41215 8949 41224
rect 9003 41264 9045 41273
rect 9003 41224 9004 41264
rect 9044 41224 9045 41264
rect 9003 41215 9045 41224
rect 9099 41264 9141 41273
rect 9099 41224 9100 41264
rect 9140 41224 9141 41264
rect 9099 41215 9141 41224
rect 9283 41264 9341 41265
rect 9283 41224 9292 41264
rect 9332 41224 9341 41264
rect 9283 41223 9341 41224
rect 9483 41264 9525 41273
rect 9483 41224 9484 41264
rect 9524 41224 9525 41264
rect 9483 41215 9525 41224
rect 9571 41264 9629 41265
rect 9571 41224 9580 41264
rect 9620 41224 9629 41264
rect 9571 41223 9629 41224
rect 9867 41264 9909 41273
rect 9867 41224 9868 41264
rect 9908 41224 9909 41264
rect 9867 41215 9909 41224
rect 9963 41264 10005 41273
rect 9963 41224 9964 41264
rect 10004 41224 10005 41264
rect 9963 41215 10005 41224
rect 10059 41264 10101 41273
rect 10059 41224 10060 41264
rect 10100 41224 10101 41264
rect 10059 41215 10101 41224
rect 10443 41264 10485 41273
rect 10443 41224 10444 41264
rect 10484 41224 10485 41264
rect 10443 41215 10485 41224
rect 10539 41264 10581 41273
rect 10539 41224 10540 41264
rect 10580 41224 10581 41264
rect 10539 41215 10581 41224
rect 10635 41264 10677 41273
rect 10635 41224 10636 41264
rect 10676 41224 10677 41264
rect 10635 41215 10677 41224
rect 10923 41264 10965 41273
rect 10923 41224 10924 41264
rect 10964 41224 10965 41264
rect 10923 41215 10965 41224
rect 11019 41264 11061 41273
rect 11019 41224 11020 41264
rect 11060 41224 11061 41264
rect 11115 41245 11116 41285
rect 11156 41245 11157 41285
rect 11115 41236 11157 41245
rect 11211 41264 11253 41273
rect 11019 41215 11061 41224
rect 11211 41224 11212 41264
rect 11252 41224 11253 41264
rect 11211 41215 11253 41224
rect 13227 41264 13269 41273
rect 13227 41224 13228 41264
rect 13268 41224 13269 41264
rect 13227 41215 13269 41224
rect 13419 41264 13461 41273
rect 13419 41224 13420 41264
rect 13460 41224 13461 41264
rect 13419 41215 13461 41224
rect 13611 41264 13653 41273
rect 13611 41224 13612 41264
rect 13652 41224 13653 41264
rect 13611 41215 13653 41224
rect 13803 41264 13845 41273
rect 13803 41224 13804 41264
rect 13844 41224 13845 41264
rect 13803 41215 13845 41224
rect 13891 41264 13949 41265
rect 13891 41224 13900 41264
rect 13940 41224 13949 41264
rect 13891 41223 13949 41224
rect 14179 41264 14237 41265
rect 14179 41224 14188 41264
rect 14228 41224 14237 41264
rect 14179 41223 14237 41224
rect 15427 41264 15485 41265
rect 15427 41224 15436 41264
rect 15476 41224 15485 41264
rect 15427 41223 15485 41224
rect 15907 41264 15965 41265
rect 15907 41224 15916 41264
rect 15956 41224 15965 41264
rect 15907 41223 15965 41224
rect 17155 41264 17213 41265
rect 17155 41224 17164 41264
rect 17204 41224 17213 41264
rect 17155 41223 17213 41224
rect 17923 41264 17981 41265
rect 17923 41224 17932 41264
rect 17972 41224 17981 41264
rect 17923 41223 17981 41224
rect 19171 41264 19229 41265
rect 19171 41224 19180 41264
rect 19220 41224 19229 41264
rect 19171 41223 19229 41224
rect 19555 41264 19613 41265
rect 19555 41224 19564 41264
rect 19604 41224 19613 41264
rect 19851 41264 19893 41273
rect 19555 41223 19613 41224
rect 19651 41250 19709 41251
rect 19651 41210 19660 41250
rect 19700 41210 19709 41250
rect 19851 41224 19852 41264
rect 19892 41224 19893 41264
rect 19851 41215 19893 41224
rect 19651 41209 19709 41210
rect 7265 41181 7323 41182
rect 7083 41140 7084 41180
rect 7124 41140 7125 41180
rect 7083 41131 7125 41140
rect 17539 41180 17597 41181
rect 17539 41140 17548 41180
rect 17588 41140 17597 41180
rect 17539 41139 17597 41140
rect 20035 41180 20093 41181
rect 20035 41140 20044 41180
rect 20084 41140 20093 41180
rect 20035 41139 20093 41140
rect 2667 41096 2709 41105
rect 2667 41056 2668 41096
rect 2708 41056 2709 41096
rect 2667 41047 2709 41056
rect 3427 41096 3485 41097
rect 3427 41056 3436 41096
rect 3476 41056 3485 41096
rect 3427 41055 3485 41056
rect 3819 41096 3861 41105
rect 3819 41056 3820 41096
rect 3860 41056 3861 41096
rect 3819 41047 3861 41056
rect 7179 41054 7221 41063
rect 2955 41012 2997 41021
rect 2955 40972 2956 41012
rect 2996 40972 2997 41012
rect 7179 41014 7180 41054
rect 7220 41014 7221 41054
rect 7179 41005 7221 41014
rect 8043 41012 8085 41021
rect 2955 40963 2997 40972
rect 8043 40972 8044 41012
rect 8084 40972 8085 41012
rect 8043 40963 8085 40972
rect 13419 41012 13461 41021
rect 13419 40972 13420 41012
rect 13460 40972 13461 41012
rect 13419 40963 13461 40972
rect 13611 41012 13653 41021
rect 13611 40972 13612 41012
rect 13652 40972 13653 41012
rect 13611 40963 13653 40972
rect 17739 41012 17781 41021
rect 17739 40972 17740 41012
rect 17780 40972 17781 41012
rect 17739 40963 17781 40972
rect 19371 41012 19413 41021
rect 19371 40972 19372 41012
rect 19412 40972 19413 41012
rect 19371 40963 19413 40972
rect 1152 40844 20352 40868
rect 1152 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 20352 40844
rect 1152 40780 20352 40804
rect 6219 40676 6261 40685
rect 6219 40636 6220 40676
rect 6260 40636 6261 40676
rect 6219 40627 6261 40636
rect 6987 40676 7029 40685
rect 6987 40636 6988 40676
rect 7028 40636 7029 40676
rect 6987 40627 7029 40636
rect 7179 40676 7221 40685
rect 7179 40636 7180 40676
rect 7220 40636 7221 40676
rect 7179 40627 7221 40636
rect 8139 40676 8181 40685
rect 8139 40636 8140 40676
rect 8180 40636 8181 40676
rect 8139 40627 8181 40636
rect 8331 40676 8373 40685
rect 8331 40636 8332 40676
rect 8372 40636 8373 40676
rect 8331 40627 8373 40636
rect 13323 40676 13365 40685
rect 13323 40636 13324 40676
rect 13364 40636 13365 40676
rect 13323 40627 13365 40636
rect 15435 40676 15477 40685
rect 15435 40636 15436 40676
rect 15476 40636 15477 40676
rect 15435 40627 15477 40636
rect 4971 40592 5013 40601
rect 4971 40552 4972 40592
rect 5012 40552 5013 40592
rect 4971 40543 5013 40552
rect 6019 40592 6077 40593
rect 6019 40552 6028 40592
rect 6068 40552 6077 40592
rect 6019 40551 6077 40552
rect 6795 40592 6837 40601
rect 6795 40552 6796 40592
rect 6836 40552 6837 40592
rect 6795 40543 6837 40552
rect 9099 40592 9141 40601
rect 9099 40552 9100 40592
rect 9140 40552 9141 40592
rect 9099 40543 9141 40552
rect 9771 40592 9813 40601
rect 9771 40552 9772 40592
rect 9812 40552 9813 40592
rect 9771 40543 9813 40552
rect 3051 40508 3093 40517
rect 3051 40468 3052 40508
rect 3092 40468 3093 40508
rect 3051 40459 3093 40468
rect 7275 40508 7317 40517
rect 7275 40468 7276 40508
rect 7316 40468 7317 40508
rect 7275 40459 7317 40468
rect 9675 40508 9717 40517
rect 9675 40468 9676 40508
rect 9716 40468 9717 40508
rect 9675 40459 9717 40468
rect 9867 40508 9909 40517
rect 9867 40468 9868 40508
rect 9908 40468 9909 40508
rect 9867 40459 9909 40468
rect 16203 40508 16245 40517
rect 16203 40468 16204 40508
rect 16244 40468 16245 40508
rect 11491 40466 11549 40467
rect 4107 40438 4149 40447
rect 2187 40424 2229 40433
rect 2187 40384 2188 40424
rect 2228 40384 2229 40424
rect 2187 40375 2229 40384
rect 2283 40424 2325 40433
rect 2283 40384 2284 40424
rect 2324 40384 2325 40424
rect 2283 40375 2325 40384
rect 2571 40424 2613 40433
rect 2571 40384 2572 40424
rect 2612 40384 2613 40424
rect 2571 40375 2613 40384
rect 2667 40424 2709 40433
rect 2667 40384 2668 40424
rect 2708 40384 2709 40424
rect 2667 40375 2709 40384
rect 3147 40424 3189 40433
rect 3147 40384 3148 40424
rect 3188 40384 3189 40424
rect 3147 40375 3189 40384
rect 3619 40424 3677 40425
rect 3619 40384 3628 40424
rect 3668 40384 3677 40424
rect 4107 40398 4108 40438
rect 4148 40398 4149 40438
rect 7172 40441 7214 40450
rect 4107 40389 4149 40398
rect 4491 40424 4533 40433
rect 3619 40383 3677 40384
rect 4491 40384 4492 40424
rect 4532 40384 4533 40424
rect 4491 40375 4533 40384
rect 4587 40424 4629 40433
rect 4587 40384 4588 40424
rect 4628 40384 4629 40424
rect 4587 40375 4629 40384
rect 4683 40424 4725 40433
rect 4683 40384 4684 40424
rect 4724 40384 4725 40424
rect 4683 40375 4725 40384
rect 4779 40424 4821 40433
rect 4779 40384 4780 40424
rect 4820 40384 4821 40424
rect 4779 40375 4821 40384
rect 4971 40424 5013 40433
rect 4971 40384 4972 40424
rect 5012 40384 5013 40424
rect 4971 40375 5013 40384
rect 5259 40424 5301 40433
rect 5259 40384 5260 40424
rect 5300 40384 5301 40424
rect 5259 40375 5301 40384
rect 5827 40424 5885 40425
rect 5827 40384 5836 40424
rect 5876 40384 5885 40424
rect 5827 40383 5885 40384
rect 6219 40424 6261 40433
rect 6219 40384 6220 40424
rect 6260 40384 6261 40424
rect 6219 40375 6261 40384
rect 6411 40424 6453 40433
rect 6411 40384 6412 40424
rect 6452 40384 6453 40424
rect 6411 40375 6453 40384
rect 6499 40424 6557 40425
rect 6499 40384 6508 40424
rect 6548 40384 6557 40424
rect 6499 40383 6557 40384
rect 6795 40424 6837 40433
rect 6795 40384 6796 40424
rect 6836 40384 6837 40424
rect 7172 40401 7173 40441
rect 7213 40401 7214 40441
rect 7172 40392 7214 40401
rect 7467 40424 7509 40433
rect 6795 40375 6837 40384
rect 7467 40384 7468 40424
rect 7508 40384 7509 40424
rect 7467 40375 7509 40384
rect 7843 40424 7901 40425
rect 7843 40384 7852 40424
rect 7892 40384 7901 40424
rect 7843 40383 7901 40384
rect 7947 40424 7989 40433
rect 7947 40384 7948 40424
rect 7988 40384 7989 40424
rect 7947 40375 7989 40384
rect 8131 40424 8189 40425
rect 8131 40384 8140 40424
rect 8180 40384 8189 40424
rect 8131 40383 8189 40384
rect 8331 40424 8373 40433
rect 8331 40384 8332 40424
rect 8372 40384 8373 40424
rect 8331 40375 8373 40384
rect 8523 40424 8565 40433
rect 8523 40384 8524 40424
rect 8564 40384 8565 40424
rect 8523 40375 8565 40384
rect 8611 40424 8669 40425
rect 8611 40384 8620 40424
rect 8660 40384 8669 40424
rect 8611 40383 8669 40384
rect 8907 40424 8949 40433
rect 8907 40384 8908 40424
rect 8948 40384 8949 40424
rect 8907 40375 8949 40384
rect 9099 40424 9141 40433
rect 9099 40384 9100 40424
rect 9140 40384 9141 40424
rect 9099 40375 9141 40384
rect 9579 40424 9621 40433
rect 9579 40384 9580 40424
rect 9620 40384 9621 40424
rect 9579 40375 9621 40384
rect 9955 40424 10013 40425
rect 9955 40384 9964 40424
rect 10004 40384 10013 40424
rect 9955 40383 10013 40384
rect 10155 40424 10197 40433
rect 10155 40384 10156 40424
rect 10196 40384 10197 40424
rect 10155 40375 10197 40384
rect 10251 40424 10293 40433
rect 10251 40384 10252 40424
rect 10292 40384 10293 40424
rect 10251 40375 10293 40384
rect 10347 40424 10389 40433
rect 10347 40384 10348 40424
rect 10388 40384 10389 40424
rect 10347 40375 10389 40384
rect 10443 40424 10485 40433
rect 10443 40384 10444 40424
rect 10484 40384 10485 40424
rect 10443 40375 10485 40384
rect 10627 40424 10685 40425
rect 10627 40384 10636 40424
rect 10676 40384 10685 40424
rect 10627 40383 10685 40384
rect 10827 40424 10869 40433
rect 11491 40426 11500 40466
rect 11540 40426 11549 40466
rect 16203 40459 16245 40468
rect 11491 40425 11549 40426
rect 10827 40384 10828 40424
rect 10868 40384 10869 40424
rect 10827 40375 10869 40384
rect 12739 40424 12797 40425
rect 12739 40384 12748 40424
rect 12788 40384 12797 40424
rect 12739 40383 12797 40384
rect 13323 40424 13365 40433
rect 13323 40384 13324 40424
rect 13364 40384 13365 40424
rect 13323 40375 13365 40384
rect 13515 40424 13557 40433
rect 13515 40384 13516 40424
rect 13556 40384 13557 40424
rect 13515 40375 13557 40384
rect 13603 40424 13661 40425
rect 13603 40384 13612 40424
rect 13652 40384 13661 40424
rect 13603 40383 13661 40384
rect 13987 40424 14045 40425
rect 13987 40384 13996 40424
rect 14036 40384 14045 40424
rect 13987 40383 14045 40384
rect 15235 40424 15293 40425
rect 15235 40384 15244 40424
rect 15284 40384 15293 40424
rect 15235 40383 15293 40384
rect 15723 40424 15765 40433
rect 15723 40384 15724 40424
rect 15764 40384 15765 40424
rect 15723 40375 15765 40384
rect 15819 40424 15861 40433
rect 15819 40384 15820 40424
rect 15860 40384 15861 40424
rect 15819 40375 15861 40384
rect 16299 40424 16341 40433
rect 17259 40429 17301 40438
rect 16299 40384 16300 40424
rect 16340 40384 16341 40424
rect 16299 40375 16341 40384
rect 16771 40424 16829 40425
rect 16771 40384 16780 40424
rect 16820 40384 16829 40424
rect 16771 40383 16829 40384
rect 17259 40389 17260 40429
rect 17300 40389 17301 40429
rect 17259 40380 17301 40389
rect 18211 40424 18269 40425
rect 18211 40384 18220 40424
rect 18260 40384 18269 40424
rect 18211 40383 18269 40384
rect 19459 40424 19517 40425
rect 19459 40384 19468 40424
rect 19508 40384 19517 40424
rect 19459 40383 19517 40384
rect 19851 40424 19893 40433
rect 19851 40384 19852 40424
rect 19892 40384 19893 40424
rect 19851 40375 19893 40384
rect 19947 40424 19989 40433
rect 19947 40384 19948 40424
rect 19988 40384 19989 40424
rect 19947 40375 19989 40384
rect 20043 40424 20085 40433
rect 20043 40384 20044 40424
rect 20084 40384 20085 40424
rect 20043 40375 20085 40384
rect 20139 40424 20181 40433
rect 20139 40384 20140 40424
rect 20180 40384 20181 40424
rect 20139 40375 20181 40384
rect 4299 40340 4341 40349
rect 4299 40300 4300 40340
rect 4340 40300 4341 40340
rect 4299 40291 4341 40300
rect 10731 40340 10773 40349
rect 10731 40300 10732 40340
rect 10772 40300 10773 40340
rect 10731 40291 10773 40300
rect 17451 40340 17493 40349
rect 17451 40300 17452 40340
rect 17492 40300 17493 40340
rect 17451 40291 17493 40300
rect 1987 40256 2045 40257
rect 1987 40216 1996 40256
rect 2036 40216 2045 40256
rect 1987 40215 2045 40216
rect 5731 40256 5789 40257
rect 5731 40216 5740 40256
rect 5780 40216 5789 40256
rect 5731 40215 5789 40216
rect 9283 40256 9341 40257
rect 9283 40216 9292 40256
rect 9332 40216 9341 40256
rect 9283 40215 9341 40216
rect 12939 40256 12981 40265
rect 12939 40216 12940 40256
rect 12980 40216 12981 40256
rect 12939 40207 12981 40216
rect 19659 40256 19701 40265
rect 19659 40216 19660 40256
rect 19700 40216 19701 40256
rect 19659 40207 19701 40216
rect 1152 40088 20452 40112
rect 1152 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20452 40088
rect 1152 40024 20452 40048
rect 2571 39920 2613 39929
rect 2571 39880 2572 39920
rect 2612 39880 2613 39920
rect 2571 39871 2613 39880
rect 6699 39920 6741 39929
rect 6699 39880 6700 39920
rect 6740 39880 6741 39920
rect 6699 39871 6741 39880
rect 9003 39920 9045 39929
rect 9003 39880 9004 39920
rect 9044 39880 9045 39920
rect 9003 39871 9045 39880
rect 14467 39920 14525 39921
rect 14467 39880 14476 39920
rect 14516 39880 14525 39920
rect 14467 39879 14525 39880
rect 15427 39920 15485 39921
rect 15427 39880 15436 39920
rect 15476 39880 15485 39920
rect 15427 39879 15485 39880
rect 17163 39920 17205 39929
rect 17163 39880 17164 39920
rect 17204 39880 17205 39920
rect 17163 39871 17205 39880
rect 19851 39920 19893 39929
rect 19851 39880 19852 39920
rect 19892 39880 19893 39920
rect 19851 39871 19893 39880
rect 4971 39836 5013 39845
rect 4971 39796 4972 39836
rect 5012 39796 5013 39836
rect 4971 39787 5013 39796
rect 9771 39836 9813 39845
rect 9771 39796 9772 39836
rect 9812 39796 9813 39836
rect 9771 39787 9813 39796
rect 12747 39836 12789 39845
rect 12747 39796 12748 39836
rect 12788 39796 12789 39836
rect 12747 39787 12789 39796
rect 13707 39836 13749 39845
rect 13707 39796 13708 39836
rect 13748 39796 13749 39836
rect 13611 39779 13653 39788
rect 13707 39787 13749 39796
rect 2467 39752 2525 39753
rect 2467 39712 2476 39752
rect 2516 39712 2525 39752
rect 2467 39711 2525 39712
rect 2755 39752 2813 39753
rect 2755 39712 2764 39752
rect 2804 39712 2813 39752
rect 2755 39711 2813 39712
rect 4003 39752 4061 39753
rect 4003 39712 4012 39752
rect 4052 39712 4061 39752
rect 4003 39711 4061 39712
rect 4395 39752 4437 39761
rect 4395 39712 4396 39752
rect 4436 39712 4437 39752
rect 4395 39703 4437 39712
rect 4491 39752 4533 39761
rect 4491 39712 4492 39752
rect 4532 39712 4533 39752
rect 4491 39703 4533 39712
rect 4587 39752 4629 39761
rect 4587 39712 4588 39752
rect 4628 39712 4629 39752
rect 4587 39703 4629 39712
rect 4683 39752 4725 39761
rect 4683 39712 4684 39752
rect 4724 39712 4725 39752
rect 4683 39703 4725 39712
rect 4867 39752 4925 39753
rect 4867 39712 4876 39752
rect 4916 39712 4925 39752
rect 4867 39711 4925 39712
rect 5067 39752 5109 39761
rect 5067 39712 5068 39752
rect 5108 39712 5109 39752
rect 5067 39703 5109 39712
rect 5251 39752 5309 39753
rect 5251 39712 5260 39752
rect 5300 39712 5309 39752
rect 5251 39711 5309 39712
rect 6499 39752 6557 39753
rect 6499 39712 6508 39752
rect 6548 39712 6557 39752
rect 6499 39711 6557 39712
rect 6883 39752 6941 39753
rect 6883 39712 6892 39752
rect 6932 39712 6941 39752
rect 6883 39711 6941 39712
rect 7275 39752 7317 39761
rect 7275 39712 7276 39752
rect 7316 39712 7317 39752
rect 7275 39703 7317 39712
rect 7371 39752 7413 39761
rect 7371 39712 7372 39752
rect 7412 39712 7413 39752
rect 7371 39703 7413 39712
rect 7755 39752 7797 39761
rect 7755 39712 7756 39752
rect 7796 39712 7797 39752
rect 7755 39703 7797 39712
rect 7851 39752 7893 39761
rect 7851 39712 7852 39752
rect 7892 39712 7893 39752
rect 7851 39703 7893 39712
rect 8323 39752 8381 39753
rect 8323 39712 8332 39752
rect 8372 39712 8381 39752
rect 9379 39752 9437 39753
rect 8323 39711 8381 39712
rect 8811 39738 8853 39747
rect 8811 39698 8812 39738
rect 8852 39698 8853 39738
rect 9379 39712 9388 39752
rect 9428 39712 9437 39752
rect 9379 39711 9437 39712
rect 9675 39752 9717 39761
rect 9675 39712 9676 39752
rect 9716 39712 9717 39752
rect 9675 39703 9717 39712
rect 10347 39752 10389 39761
rect 10347 39712 10348 39752
rect 10388 39712 10389 39752
rect 10347 39703 10389 39712
rect 10539 39752 10581 39761
rect 10539 39712 10540 39752
rect 10580 39712 10581 39752
rect 10539 39703 10581 39712
rect 10627 39752 10685 39753
rect 10627 39712 10636 39752
rect 10676 39712 10685 39752
rect 10627 39711 10685 39712
rect 11299 39752 11357 39753
rect 11299 39712 11308 39752
rect 11348 39712 11357 39752
rect 11299 39711 11357 39712
rect 12547 39752 12605 39753
rect 12547 39712 12556 39752
rect 12596 39712 12605 39752
rect 12547 39711 12605 39712
rect 12931 39752 12989 39753
rect 12931 39712 12940 39752
rect 12980 39712 12989 39752
rect 12931 39711 12989 39712
rect 13315 39752 13373 39753
rect 13315 39712 13324 39752
rect 13364 39712 13373 39752
rect 13611 39739 13612 39779
rect 13652 39739 13653 39779
rect 18123 39772 18165 39781
rect 13611 39730 13653 39739
rect 14187 39752 14229 39761
rect 13315 39711 13373 39712
rect 14187 39712 14188 39752
rect 14228 39712 14229 39752
rect 14187 39703 14229 39712
rect 14283 39752 14325 39761
rect 14283 39712 14284 39752
rect 14324 39712 14325 39752
rect 14283 39703 14325 39712
rect 14379 39752 14421 39761
rect 14379 39712 14380 39752
rect 14420 39712 14421 39752
rect 14379 39703 14421 39712
rect 14667 39752 14709 39761
rect 14667 39712 14668 39752
rect 14708 39712 14709 39752
rect 14667 39703 14709 39712
rect 14763 39752 14805 39761
rect 14763 39712 14764 39752
rect 14804 39712 14805 39752
rect 14763 39703 14805 39712
rect 14859 39752 14901 39761
rect 14859 39712 14860 39752
rect 14900 39712 14901 39752
rect 14859 39703 14901 39712
rect 14955 39752 14997 39761
rect 14955 39712 14956 39752
rect 14996 39712 14997 39752
rect 14955 39703 14997 39712
rect 15147 39752 15189 39761
rect 15147 39712 15148 39752
rect 15188 39712 15189 39752
rect 15147 39703 15189 39712
rect 15243 39752 15285 39761
rect 15243 39712 15244 39752
rect 15284 39712 15285 39752
rect 15243 39703 15285 39712
rect 15339 39752 15381 39761
rect 15339 39712 15340 39752
rect 15380 39712 15381 39752
rect 15339 39703 15381 39712
rect 15715 39752 15773 39753
rect 15715 39712 15724 39752
rect 15764 39712 15773 39752
rect 15715 39711 15773 39712
rect 16963 39752 17021 39753
rect 16963 39712 16972 39752
rect 17012 39712 17021 39752
rect 18123 39732 18124 39772
rect 18164 39732 18165 39772
rect 18123 39723 18165 39732
rect 18219 39752 18261 39761
rect 16963 39711 17021 39712
rect 18219 39712 18220 39752
rect 18260 39712 18261 39752
rect 18219 39703 18261 39712
rect 19171 39752 19229 39753
rect 19171 39712 19180 39752
rect 19220 39712 19229 39752
rect 19171 39711 19229 39712
rect 19659 39747 19701 39756
rect 19659 39707 19660 39747
rect 19700 39707 19701 39747
rect 19659 39698 19701 39707
rect 8811 39689 8853 39698
rect 18603 39668 18645 39677
rect 18603 39628 18604 39668
rect 18644 39628 18645 39668
rect 18603 39619 18645 39628
rect 18699 39668 18741 39677
rect 18699 39628 18700 39668
rect 18740 39628 18741 39668
rect 18699 39619 18741 39628
rect 6987 39584 7029 39593
rect 6987 39544 6988 39584
rect 7028 39544 7029 39584
rect 6987 39535 7029 39544
rect 10051 39584 10109 39585
rect 10051 39544 10060 39584
rect 10100 39544 10109 39584
rect 10051 39543 10109 39544
rect 4203 39500 4245 39509
rect 4203 39460 4204 39500
rect 4244 39460 4245 39500
rect 4203 39451 4245 39460
rect 10347 39500 10389 39509
rect 10347 39460 10348 39500
rect 10388 39460 10389 39500
rect 10347 39451 10389 39460
rect 13035 39500 13077 39509
rect 13035 39460 13036 39500
rect 13076 39460 13077 39500
rect 13035 39451 13077 39460
rect 13987 39500 14045 39501
rect 13987 39460 13996 39500
rect 14036 39460 14045 39500
rect 13987 39459 14045 39460
rect 1152 39332 20352 39356
rect 1152 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 20352 39332
rect 1152 39268 20352 39292
rect 12555 39164 12597 39173
rect 12555 39124 12556 39164
rect 12596 39124 12597 39164
rect 12555 39115 12597 39124
rect 14083 39164 14141 39165
rect 14083 39124 14092 39164
rect 14132 39124 14141 39164
rect 14083 39123 14141 39124
rect 17739 39164 17781 39173
rect 17739 39124 17740 39164
rect 17780 39124 17781 39164
rect 17739 39115 17781 39124
rect 9771 39080 9813 39089
rect 9771 39040 9772 39080
rect 9812 39040 9813 39080
rect 9771 39031 9813 39040
rect 12267 39080 12309 39089
rect 12267 39040 12268 39080
rect 12308 39040 12309 39080
rect 12267 39031 12309 39040
rect 3627 38996 3669 39005
rect 3627 38956 3628 38996
rect 3668 38956 3669 38996
rect 3627 38947 3669 38956
rect 5739 38996 5781 39005
rect 5739 38956 5740 38996
rect 5780 38956 5781 38996
rect 5739 38947 5781 38956
rect 7755 38996 7797 39005
rect 7755 38956 7756 38996
rect 7796 38956 7797 38996
rect 7755 38947 7797 38956
rect 4587 38926 4629 38935
rect 3051 38912 3093 38921
rect 3051 38872 3052 38912
rect 3092 38872 3093 38912
rect 3051 38863 3093 38872
rect 3147 38912 3189 38921
rect 3147 38872 3148 38912
rect 3188 38872 3189 38912
rect 3147 38863 3189 38872
rect 3531 38912 3573 38921
rect 3531 38872 3532 38912
rect 3572 38872 3573 38912
rect 3531 38863 3573 38872
rect 4099 38912 4157 38913
rect 4099 38872 4108 38912
rect 4148 38872 4157 38912
rect 4587 38886 4588 38926
rect 4628 38886 4629 38926
rect 6843 38921 6885 38930
rect 8811 38926 8853 38935
rect 4587 38877 4629 38886
rect 5259 38912 5301 38921
rect 4099 38871 4157 38872
rect 5259 38872 5260 38912
rect 5300 38872 5301 38912
rect 5259 38863 5301 38872
rect 5355 38912 5397 38921
rect 5355 38872 5356 38912
rect 5396 38872 5397 38912
rect 5355 38863 5397 38872
rect 5835 38912 5877 38921
rect 5835 38872 5836 38912
rect 5876 38872 5877 38912
rect 5835 38863 5877 38872
rect 6307 38912 6365 38913
rect 6307 38872 6316 38912
rect 6356 38872 6365 38912
rect 6843 38881 6844 38921
rect 6884 38881 6885 38921
rect 6843 38872 6885 38881
rect 7275 38912 7317 38921
rect 7275 38872 7276 38912
rect 7316 38872 7317 38912
rect 6307 38871 6365 38872
rect 7275 38863 7317 38872
rect 7371 38912 7413 38921
rect 7371 38872 7372 38912
rect 7412 38872 7413 38912
rect 7371 38863 7413 38872
rect 7851 38912 7893 38921
rect 7851 38872 7852 38912
rect 7892 38872 7893 38912
rect 7851 38863 7893 38872
rect 8323 38912 8381 38913
rect 8323 38872 8332 38912
rect 8372 38872 8381 38912
rect 8811 38886 8812 38926
rect 8852 38886 8853 38926
rect 8811 38877 8853 38886
rect 9579 38912 9621 38921
rect 8323 38871 8381 38872
rect 9579 38872 9580 38912
rect 9620 38872 9621 38912
rect 9579 38863 9621 38872
rect 9771 38912 9813 38921
rect 9771 38872 9772 38912
rect 9812 38872 9813 38912
rect 9771 38863 9813 38872
rect 9955 38912 10013 38913
rect 9955 38872 9964 38912
rect 10004 38872 10013 38912
rect 9955 38871 10013 38872
rect 11203 38912 11261 38913
rect 11203 38872 11212 38912
rect 11252 38872 11261 38912
rect 11203 38871 11261 38872
rect 11787 38912 11829 38921
rect 11787 38872 11788 38912
rect 11828 38872 11829 38912
rect 11787 38863 11829 38872
rect 11883 38912 11925 38921
rect 11883 38872 11884 38912
rect 11924 38872 11925 38912
rect 11883 38863 11925 38872
rect 11979 38912 12021 38921
rect 11979 38872 11980 38912
rect 12020 38872 12021 38912
rect 11979 38863 12021 38872
rect 12355 38912 12413 38913
rect 12355 38872 12364 38912
rect 12404 38872 12413 38912
rect 12355 38871 12413 38872
rect 12643 38912 12701 38913
rect 12643 38872 12652 38912
rect 12692 38872 12701 38912
rect 12643 38871 12701 38872
rect 12843 38912 12885 38921
rect 12843 38872 12844 38912
rect 12884 38872 12885 38912
rect 12843 38863 12885 38872
rect 12939 38912 12981 38921
rect 12939 38872 12940 38912
rect 12980 38872 12981 38912
rect 12939 38863 12981 38872
rect 13035 38912 13077 38921
rect 13035 38872 13036 38912
rect 13076 38872 13077 38912
rect 13035 38863 13077 38872
rect 13131 38912 13173 38921
rect 13131 38872 13132 38912
rect 13172 38872 13173 38912
rect 13131 38863 13173 38872
rect 13411 38912 13469 38913
rect 13411 38872 13420 38912
rect 13460 38872 13469 38912
rect 13411 38871 13469 38872
rect 13707 38912 13749 38921
rect 13707 38872 13708 38912
rect 13748 38872 13749 38912
rect 13707 38863 13749 38872
rect 14275 38912 14333 38913
rect 14275 38872 14284 38912
rect 14324 38872 14333 38912
rect 14275 38871 14333 38872
rect 14379 38912 14421 38921
rect 14379 38872 14380 38912
rect 14420 38872 14421 38912
rect 14379 38863 14421 38872
rect 14571 38912 14613 38921
rect 14571 38872 14572 38912
rect 14612 38872 14613 38912
rect 14571 38863 14613 38872
rect 16291 38912 16349 38913
rect 16291 38872 16300 38912
rect 16340 38872 16349 38912
rect 16291 38871 16349 38872
rect 17539 38912 17597 38913
rect 17539 38872 17548 38912
rect 17588 38872 17597 38912
rect 17539 38871 17597 38872
rect 18411 38912 18453 38921
rect 18411 38872 18412 38912
rect 18452 38872 18453 38912
rect 18411 38863 18453 38872
rect 18507 38912 18549 38921
rect 18507 38872 18508 38912
rect 18548 38872 18549 38912
rect 18507 38863 18549 38872
rect 18891 38912 18933 38921
rect 18891 38872 18892 38912
rect 18932 38872 18933 38912
rect 18891 38863 18933 38872
rect 18987 38912 19029 38921
rect 19947 38917 19989 38926
rect 18987 38872 18988 38912
rect 19028 38872 19029 38912
rect 18987 38863 19029 38872
rect 19459 38912 19517 38913
rect 19459 38872 19468 38912
rect 19508 38872 19517 38912
rect 19459 38871 19517 38872
rect 19947 38877 19948 38917
rect 19988 38877 19989 38917
rect 19947 38868 19989 38877
rect 6987 38828 7029 38837
rect 6987 38788 6988 38828
rect 7028 38788 7029 38828
rect 6987 38779 7029 38788
rect 9003 38828 9045 38837
rect 9003 38788 9004 38828
rect 9044 38788 9045 38828
rect 9003 38779 9045 38788
rect 13803 38828 13845 38837
rect 13803 38788 13804 38828
rect 13844 38788 13845 38828
rect 13803 38779 13845 38788
rect 14475 38828 14517 38837
rect 14475 38788 14476 38828
rect 14516 38788 14517 38828
rect 14475 38779 14517 38788
rect 20139 38828 20181 38837
rect 20139 38788 20140 38828
rect 20180 38788 20181 38828
rect 20139 38779 20181 38788
rect 2667 38744 2709 38753
rect 2667 38704 2668 38744
rect 2708 38704 2709 38744
rect 2667 38695 2709 38704
rect 4779 38744 4821 38753
rect 4779 38704 4780 38744
rect 4820 38704 4821 38744
rect 4779 38695 4821 38704
rect 11403 38744 11445 38753
rect 11403 38704 11404 38744
rect 11444 38704 11445 38744
rect 11403 38695 11445 38704
rect 11595 38744 11637 38753
rect 11595 38704 11596 38744
rect 11636 38704 11637 38744
rect 11595 38695 11637 38704
rect 1152 38576 20452 38600
rect 1152 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20452 38576
rect 1152 38512 20452 38536
rect 2667 38408 2709 38417
rect 2667 38368 2668 38408
rect 2708 38368 2709 38408
rect 2667 38359 2709 38368
rect 3043 38408 3101 38409
rect 3043 38368 3052 38408
rect 3092 38368 3101 38408
rect 3043 38367 3101 38368
rect 5355 38408 5397 38417
rect 5355 38368 5356 38408
rect 5396 38368 5397 38408
rect 5355 38359 5397 38368
rect 6987 38408 7029 38417
rect 6987 38368 6988 38408
rect 7028 38368 7029 38408
rect 6987 38359 7029 38368
rect 10731 38408 10773 38417
rect 10731 38368 10732 38408
rect 10772 38368 10773 38408
rect 10731 38359 10773 38368
rect 18891 38408 18933 38417
rect 18891 38368 18892 38408
rect 18932 38368 18933 38408
rect 18891 38359 18933 38368
rect 19563 38408 19605 38417
rect 19563 38368 19564 38408
rect 19604 38368 19605 38408
rect 19563 38359 19605 38368
rect 17259 38324 17301 38333
rect 17259 38284 17260 38324
rect 17300 38284 17301 38324
rect 17259 38275 17301 38284
rect 1219 38240 1277 38241
rect 1219 38200 1228 38240
rect 1268 38200 1277 38240
rect 1219 38199 1277 38200
rect 2467 38240 2525 38241
rect 2467 38200 2476 38240
rect 2516 38200 2525 38240
rect 2467 38199 2525 38200
rect 3907 38240 3965 38241
rect 3907 38200 3916 38240
rect 3956 38200 3965 38240
rect 3907 38199 3965 38200
rect 5155 38240 5213 38241
rect 5155 38200 5164 38240
rect 5204 38200 5213 38240
rect 5155 38199 5213 38200
rect 5539 38240 5597 38241
rect 5539 38200 5548 38240
rect 5588 38200 5597 38240
rect 5539 38199 5597 38200
rect 6787 38240 6845 38241
rect 6787 38200 6796 38240
rect 6836 38200 6845 38240
rect 6787 38199 6845 38200
rect 9283 38240 9341 38241
rect 9283 38200 9292 38240
rect 9332 38200 9341 38240
rect 9283 38199 9341 38200
rect 10531 38240 10589 38241
rect 10531 38200 10540 38240
rect 10580 38200 10589 38240
rect 10531 38199 10589 38200
rect 11115 38240 11157 38249
rect 11115 38200 11116 38240
rect 11156 38200 11157 38240
rect 11115 38191 11157 38200
rect 11211 38240 11253 38249
rect 11211 38200 11212 38240
rect 11252 38200 11253 38240
rect 11211 38191 11253 38200
rect 11307 38240 11349 38249
rect 11307 38200 11308 38240
rect 11348 38200 11349 38240
rect 11307 38191 11349 38200
rect 11403 38240 11445 38249
rect 11403 38200 11404 38240
rect 11444 38200 11445 38240
rect 11403 38191 11445 38200
rect 12643 38240 12701 38241
rect 12643 38200 12652 38240
rect 12692 38200 12701 38240
rect 12643 38199 12701 38200
rect 13891 38240 13949 38241
rect 13891 38200 13900 38240
rect 13940 38200 13949 38240
rect 13891 38199 13949 38200
rect 15531 38240 15573 38249
rect 15531 38200 15532 38240
rect 15572 38200 15573 38240
rect 15531 38191 15573 38200
rect 15627 38240 15669 38249
rect 15627 38200 15628 38240
rect 15668 38200 15669 38240
rect 15627 38191 15669 38200
rect 16107 38240 16149 38249
rect 16107 38200 16108 38240
rect 16148 38200 16149 38240
rect 16107 38191 16149 38200
rect 16579 38240 16637 38241
rect 16579 38200 16588 38240
rect 16628 38200 16637 38240
rect 17443 38240 17501 38241
rect 16579 38199 16637 38200
rect 17115 38198 17157 38207
rect 17443 38200 17452 38240
rect 17492 38200 17501 38240
rect 17443 38199 17501 38200
rect 18691 38240 18749 38241
rect 18691 38200 18700 38240
rect 18740 38200 18749 38240
rect 18691 38199 18749 38200
rect 16011 38156 16053 38165
rect 16011 38116 16012 38156
rect 16052 38116 16053 38156
rect 17115 38158 17116 38198
rect 17156 38158 17157 38198
rect 17115 38149 17157 38158
rect 19363 38156 19421 38157
rect 16011 38107 16053 38116
rect 19363 38116 19372 38156
rect 19412 38116 19421 38156
rect 19363 38115 19421 38116
rect 19747 38156 19805 38157
rect 19747 38116 19756 38156
rect 19796 38116 19805 38156
rect 19747 38115 19805 38116
rect 2955 38072 2997 38081
rect 2955 38032 2956 38072
rect 2996 38032 2997 38072
rect 2955 38023 2997 38032
rect 14091 38072 14133 38081
rect 14091 38032 14092 38072
rect 14132 38032 14133 38072
rect 14091 38023 14133 38032
rect 19947 38072 19989 38081
rect 19947 38032 19948 38072
rect 19988 38032 19989 38072
rect 19947 38023 19989 38032
rect 1152 37820 20352 37844
rect 1152 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 20352 37820
rect 1152 37756 20352 37780
rect 2667 37652 2709 37661
rect 2667 37612 2668 37652
rect 2708 37612 2709 37652
rect 2667 37603 2709 37612
rect 15723 37652 15765 37661
rect 15723 37612 15724 37652
rect 15764 37612 15765 37652
rect 15723 37603 15765 37612
rect 17355 37652 17397 37661
rect 17355 37612 17356 37652
rect 17396 37612 17397 37652
rect 17355 37603 17397 37612
rect 19947 37652 19989 37661
rect 19947 37612 19948 37652
rect 19988 37612 19989 37652
rect 19947 37603 19989 37612
rect 3003 37409 3045 37418
rect 13803 37414 13845 37423
rect 1219 37400 1277 37401
rect 1219 37360 1228 37400
rect 1268 37360 1277 37400
rect 1219 37359 1277 37360
rect 2467 37400 2525 37401
rect 2467 37360 2476 37400
rect 2516 37360 2525 37400
rect 3003 37369 3004 37409
rect 3044 37369 3045 37409
rect 3003 37360 3045 37369
rect 3523 37400 3581 37401
rect 3523 37360 3532 37400
rect 3572 37360 3581 37400
rect 2467 37359 2525 37360
rect 3523 37359 3581 37360
rect 4011 37400 4053 37409
rect 4011 37360 4012 37400
rect 4052 37360 4053 37400
rect 4011 37351 4053 37360
rect 4107 37400 4149 37409
rect 4107 37360 4108 37400
rect 4148 37360 4149 37400
rect 4107 37351 4149 37360
rect 4491 37400 4533 37409
rect 4491 37360 4492 37400
rect 4532 37360 4533 37400
rect 4491 37351 4533 37360
rect 4587 37400 4629 37409
rect 4587 37360 4588 37400
rect 4628 37360 4629 37400
rect 4587 37351 4629 37360
rect 5443 37400 5501 37401
rect 5443 37360 5452 37400
rect 5492 37360 5501 37400
rect 5443 37359 5501 37360
rect 5739 37400 5781 37409
rect 5739 37360 5740 37400
rect 5780 37360 5781 37400
rect 5739 37351 5781 37360
rect 5835 37400 5877 37409
rect 5835 37360 5836 37400
rect 5876 37360 5877 37400
rect 5835 37351 5877 37360
rect 5931 37400 5973 37409
rect 5931 37360 5932 37400
rect 5972 37360 5973 37400
rect 5931 37351 5973 37360
rect 6027 37400 6069 37409
rect 6027 37360 6028 37400
rect 6068 37360 6069 37400
rect 6027 37351 6069 37360
rect 6315 37400 6357 37409
rect 6315 37360 6316 37400
rect 6356 37360 6357 37400
rect 6315 37351 6357 37360
rect 6411 37400 6453 37409
rect 6411 37360 6412 37400
rect 6452 37360 6453 37400
rect 6411 37351 6453 37360
rect 6507 37400 6549 37409
rect 6507 37360 6508 37400
rect 6548 37360 6549 37400
rect 6507 37351 6549 37360
rect 6691 37400 6749 37401
rect 6691 37360 6700 37400
rect 6740 37360 6749 37400
rect 6691 37359 6749 37360
rect 7939 37400 7997 37401
rect 7939 37360 7948 37400
rect 7988 37360 7997 37400
rect 7939 37359 7997 37360
rect 8323 37400 8381 37401
rect 8323 37360 8332 37400
rect 8372 37360 8381 37400
rect 8323 37359 8381 37360
rect 9571 37400 9629 37401
rect 9571 37360 9580 37400
rect 9620 37360 9629 37400
rect 9571 37359 9629 37360
rect 10531 37400 10589 37401
rect 10531 37360 10540 37400
rect 10580 37360 10589 37400
rect 10531 37359 10589 37360
rect 11779 37400 11837 37401
rect 11779 37360 11788 37400
rect 11828 37360 11837 37400
rect 11779 37359 11837 37360
rect 12267 37400 12309 37409
rect 12267 37360 12268 37400
rect 12308 37360 12309 37400
rect 12267 37351 12309 37360
rect 12363 37400 12405 37409
rect 12363 37360 12364 37400
rect 12404 37360 12405 37400
rect 12363 37351 12405 37360
rect 12747 37400 12789 37409
rect 12747 37360 12748 37400
rect 12788 37360 12789 37400
rect 12747 37351 12789 37360
rect 12843 37400 12885 37409
rect 12843 37360 12844 37400
rect 12884 37360 12885 37400
rect 12843 37351 12885 37360
rect 13315 37400 13373 37401
rect 13315 37360 13324 37400
rect 13364 37360 13373 37400
rect 13803 37374 13804 37414
rect 13844 37374 13845 37414
rect 13803 37365 13845 37374
rect 14275 37400 14333 37401
rect 13315 37359 13373 37360
rect 14275 37360 14284 37400
rect 14324 37360 14333 37400
rect 14275 37359 14333 37360
rect 15523 37400 15581 37401
rect 15523 37360 15532 37400
rect 15572 37360 15581 37400
rect 15523 37359 15581 37360
rect 15907 37400 15965 37401
rect 15907 37360 15916 37400
rect 15956 37360 15965 37400
rect 15907 37359 15965 37360
rect 17155 37400 17213 37401
rect 17155 37360 17164 37400
rect 17204 37360 17213 37400
rect 17155 37359 17213 37360
rect 18499 37400 18557 37401
rect 18499 37360 18508 37400
rect 18548 37360 18557 37400
rect 18499 37359 18557 37360
rect 19747 37400 19805 37401
rect 19747 37360 19756 37400
rect 19796 37360 19805 37400
rect 19747 37359 19805 37360
rect 13995 37316 14037 37325
rect 13995 37276 13996 37316
rect 14036 37276 14037 37316
rect 13995 37267 14037 37276
rect 2859 37232 2901 37241
rect 2859 37192 2860 37232
rect 2900 37192 2901 37232
rect 2859 37183 2901 37192
rect 5547 37232 5589 37241
rect 5547 37192 5548 37232
rect 5588 37192 5589 37232
rect 5547 37183 5589 37192
rect 6211 37232 6269 37233
rect 6211 37192 6220 37232
rect 6260 37192 6269 37232
rect 6211 37191 6269 37192
rect 8139 37232 8181 37241
rect 8139 37192 8140 37232
rect 8180 37192 8181 37232
rect 8139 37183 8181 37192
rect 9771 37232 9813 37241
rect 9771 37192 9772 37232
rect 9812 37192 9813 37232
rect 9771 37183 9813 37192
rect 11979 37232 12021 37241
rect 11979 37192 11980 37232
rect 12020 37192 12021 37232
rect 11979 37183 12021 37192
rect 1152 37064 20452 37088
rect 1152 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20452 37064
rect 1152 37000 20452 37024
rect 2667 36896 2709 36905
rect 2667 36856 2668 36896
rect 2708 36856 2709 36896
rect 2667 36847 2709 36856
rect 4299 36896 4341 36905
rect 4299 36856 4300 36896
rect 4340 36856 4341 36896
rect 4299 36847 4341 36856
rect 5931 36896 5973 36905
rect 5931 36856 5932 36896
rect 5972 36856 5973 36896
rect 5931 36847 5973 36856
rect 6787 36896 6845 36897
rect 6787 36856 6796 36896
rect 6836 36856 6845 36896
rect 6787 36855 6845 36856
rect 7659 36896 7701 36905
rect 7659 36856 7660 36896
rect 7700 36856 7701 36896
rect 7659 36847 7701 36856
rect 10059 36896 10101 36905
rect 10059 36856 10060 36896
rect 10100 36856 10101 36896
rect 10059 36847 10101 36856
rect 12267 36896 12309 36905
rect 12267 36856 12268 36896
rect 12308 36856 12309 36896
rect 12267 36847 12309 36856
rect 14475 36896 14517 36905
rect 14475 36856 14476 36896
rect 14516 36856 14517 36896
rect 14475 36847 14517 36856
rect 6219 36812 6261 36821
rect 6219 36772 6220 36812
rect 6260 36772 6261 36812
rect 6219 36763 6261 36772
rect 17355 36812 17397 36821
rect 17355 36772 17356 36812
rect 17396 36772 17397 36812
rect 17355 36763 17397 36772
rect 20043 36812 20085 36821
rect 20043 36772 20044 36812
rect 20084 36772 20085 36812
rect 20043 36763 20085 36772
rect 1219 36728 1277 36729
rect 1219 36688 1228 36728
rect 1268 36688 1277 36728
rect 1219 36687 1277 36688
rect 2467 36728 2525 36729
rect 2467 36688 2476 36728
rect 2516 36688 2525 36728
rect 2467 36687 2525 36688
rect 2851 36728 2909 36729
rect 2851 36688 2860 36728
rect 2900 36688 2909 36728
rect 2851 36687 2909 36688
rect 4099 36728 4157 36729
rect 4099 36688 4108 36728
rect 4148 36688 4157 36728
rect 4099 36687 4157 36688
rect 4483 36728 4541 36729
rect 4483 36688 4492 36728
rect 4532 36688 4541 36728
rect 4483 36687 4541 36688
rect 5731 36728 5789 36729
rect 5731 36688 5740 36728
rect 5780 36688 5789 36728
rect 5731 36687 5789 36688
rect 6123 36728 6165 36737
rect 6123 36688 6124 36728
rect 6164 36688 6165 36728
rect 6123 36679 6165 36688
rect 6315 36728 6357 36737
rect 6315 36688 6316 36728
rect 6356 36688 6357 36728
rect 6595 36728 6653 36729
rect 6315 36679 6357 36688
rect 6403 36709 6461 36710
rect 6403 36669 6412 36709
rect 6452 36669 6461 36709
rect 6595 36688 6604 36728
rect 6644 36688 6653 36728
rect 6595 36687 6653 36688
rect 6699 36728 6741 36737
rect 6699 36688 6700 36728
rect 6740 36688 6741 36728
rect 6699 36679 6741 36688
rect 6891 36728 6933 36737
rect 6891 36688 6892 36728
rect 6932 36688 6933 36728
rect 6891 36679 6933 36688
rect 7083 36728 7125 36737
rect 7083 36688 7084 36728
rect 7124 36688 7125 36728
rect 7083 36679 7125 36688
rect 7275 36728 7317 36737
rect 7275 36688 7276 36728
rect 7316 36688 7317 36728
rect 7275 36679 7317 36688
rect 7363 36728 7421 36729
rect 7363 36688 7372 36728
rect 7412 36688 7421 36728
rect 7363 36687 7421 36688
rect 7563 36728 7605 36737
rect 7563 36688 7564 36728
rect 7604 36688 7605 36728
rect 7563 36679 7605 36688
rect 7755 36728 7797 36737
rect 7755 36688 7756 36728
rect 7796 36688 7797 36728
rect 7755 36679 7797 36688
rect 8331 36728 8373 36737
rect 8331 36688 8332 36728
rect 8372 36688 8373 36728
rect 8331 36679 8373 36688
rect 8427 36728 8469 36737
rect 8427 36688 8428 36728
rect 8468 36688 8469 36728
rect 8427 36679 8469 36688
rect 9379 36728 9437 36729
rect 9379 36688 9388 36728
rect 9428 36688 9437 36728
rect 9379 36687 9437 36688
rect 9867 36723 9909 36732
rect 9867 36683 9868 36723
rect 9908 36683 9909 36723
rect 10819 36728 10877 36729
rect 10819 36688 10828 36728
rect 10868 36688 10877 36728
rect 10819 36687 10877 36688
rect 12067 36728 12125 36729
rect 12067 36688 12076 36728
rect 12116 36688 12125 36728
rect 12067 36687 12125 36688
rect 12747 36728 12789 36737
rect 12747 36688 12748 36728
rect 12788 36688 12789 36728
rect 9867 36674 9909 36683
rect 12747 36679 12789 36688
rect 12843 36728 12885 36737
rect 12843 36688 12844 36728
rect 12884 36688 12885 36728
rect 12843 36679 12885 36688
rect 13795 36728 13853 36729
rect 13795 36688 13804 36728
rect 13844 36688 13853 36728
rect 15627 36728 15669 36737
rect 13795 36687 13853 36688
rect 14331 36686 14373 36695
rect 6403 36668 6461 36669
rect 8811 36644 8853 36653
rect 8811 36604 8812 36644
rect 8852 36604 8853 36644
rect 8811 36595 8853 36604
rect 8907 36644 8949 36653
rect 8907 36604 8908 36644
rect 8948 36604 8949 36644
rect 8907 36595 8949 36604
rect 13227 36644 13269 36653
rect 13227 36604 13228 36644
rect 13268 36604 13269 36644
rect 13227 36595 13269 36604
rect 13323 36644 13365 36653
rect 13323 36604 13324 36644
rect 13364 36604 13365 36644
rect 14331 36646 14332 36686
rect 14372 36646 14373 36686
rect 15627 36688 15628 36728
rect 15668 36688 15669 36728
rect 15627 36679 15669 36688
rect 15723 36728 15765 36737
rect 15723 36688 15724 36728
rect 15764 36688 15765 36728
rect 15723 36679 15765 36688
rect 16675 36728 16733 36729
rect 16675 36688 16684 36728
rect 16724 36688 16733 36728
rect 18315 36728 18357 36737
rect 16675 36687 16733 36688
rect 17163 36714 17205 36723
rect 17163 36674 17164 36714
rect 17204 36674 17205 36714
rect 18315 36688 18316 36728
rect 18356 36688 18357 36728
rect 18315 36679 18357 36688
rect 18411 36728 18453 36737
rect 18411 36688 18412 36728
rect 18452 36688 18453 36728
rect 18411 36679 18453 36688
rect 18891 36728 18933 36737
rect 18891 36688 18892 36728
rect 18932 36688 18933 36728
rect 18891 36679 18933 36688
rect 19363 36728 19421 36729
rect 19363 36688 19372 36728
rect 19412 36688 19421 36728
rect 19363 36687 19421 36688
rect 19851 36714 19893 36723
rect 17163 36665 17205 36674
rect 19851 36674 19852 36714
rect 19892 36674 19893 36714
rect 19851 36665 19893 36674
rect 14331 36637 14373 36646
rect 16107 36644 16149 36653
rect 13323 36595 13365 36604
rect 16107 36604 16108 36644
rect 16148 36604 16149 36644
rect 16107 36595 16149 36604
rect 16203 36644 16245 36653
rect 16203 36604 16204 36644
rect 16244 36604 16245 36644
rect 16203 36595 16245 36604
rect 18795 36644 18837 36653
rect 18795 36604 18796 36644
rect 18836 36604 18837 36644
rect 18795 36595 18837 36604
rect 7083 36560 7125 36569
rect 7083 36520 7084 36560
rect 7124 36520 7125 36560
rect 7083 36511 7125 36520
rect 1152 36308 20352 36332
rect 1152 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 20352 36308
rect 1152 36244 20352 36268
rect 2667 36140 2709 36149
rect 2667 36100 2668 36140
rect 2708 36100 2709 36140
rect 2667 36091 2709 36100
rect 5451 36140 5493 36149
rect 5451 36100 5452 36140
rect 5492 36100 5493 36140
rect 5451 36091 5493 36100
rect 6979 36140 7037 36141
rect 6979 36100 6988 36140
rect 7028 36100 7037 36140
rect 6979 36099 7037 36100
rect 9195 36140 9237 36149
rect 9195 36100 9196 36140
rect 9236 36100 9237 36140
rect 9195 36091 9237 36100
rect 18315 36140 18357 36149
rect 18315 36100 18316 36140
rect 18356 36100 18357 36140
rect 18315 36091 18357 36100
rect 19947 36140 19989 36149
rect 19947 36100 19948 36140
rect 19988 36100 19989 36140
rect 19947 36091 19989 36100
rect 11067 35897 11109 35906
rect 1219 35888 1277 35889
rect 1219 35848 1228 35888
rect 1268 35848 1277 35888
rect 1219 35847 1277 35848
rect 2467 35888 2525 35889
rect 2467 35848 2476 35888
rect 2516 35848 2525 35888
rect 2467 35847 2525 35848
rect 4003 35888 4061 35889
rect 4003 35848 4012 35888
rect 4052 35848 4061 35888
rect 4003 35847 4061 35848
rect 5251 35888 5309 35889
rect 5251 35848 5260 35888
rect 5300 35848 5309 35888
rect 5251 35847 5309 35848
rect 5739 35888 5781 35897
rect 5739 35848 5740 35888
rect 5780 35848 5781 35888
rect 5739 35839 5781 35848
rect 5835 35888 5877 35897
rect 5835 35848 5836 35888
rect 5876 35848 5877 35888
rect 5835 35839 5877 35848
rect 5931 35888 5973 35897
rect 5931 35848 5932 35888
rect 5972 35848 5973 35888
rect 5931 35839 5973 35848
rect 6027 35888 6069 35897
rect 6027 35848 6028 35888
rect 6068 35848 6069 35888
rect 6027 35839 6069 35848
rect 6307 35888 6365 35889
rect 6307 35848 6316 35888
rect 6356 35848 6365 35888
rect 6307 35847 6365 35848
rect 6603 35888 6645 35897
rect 6603 35848 6604 35888
rect 6644 35848 6645 35888
rect 6603 35839 6645 35848
rect 7171 35888 7229 35889
rect 7171 35848 7180 35888
rect 7220 35848 7229 35888
rect 7171 35847 7229 35848
rect 7275 35888 7317 35897
rect 7275 35848 7276 35888
rect 7316 35848 7317 35888
rect 7275 35839 7317 35848
rect 7459 35888 7517 35889
rect 7459 35848 7468 35888
rect 7508 35848 7517 35888
rect 7459 35847 7517 35848
rect 7563 35888 7605 35897
rect 7563 35848 7564 35888
rect 7604 35848 7605 35888
rect 7563 35839 7605 35848
rect 7747 35888 7805 35889
rect 7747 35848 7756 35888
rect 7796 35848 7805 35888
rect 7747 35847 7805 35848
rect 8995 35888 9053 35889
rect 8995 35848 9004 35888
rect 9044 35848 9053 35888
rect 8995 35847 9053 35848
rect 9483 35888 9525 35897
rect 9483 35848 9484 35888
rect 9524 35848 9525 35888
rect 9483 35839 9525 35848
rect 9579 35888 9621 35897
rect 9579 35848 9580 35888
rect 9620 35848 9621 35888
rect 9579 35839 9621 35848
rect 9963 35888 10005 35897
rect 9963 35848 9964 35888
rect 10004 35848 10005 35888
rect 9963 35839 10005 35848
rect 10059 35888 10101 35897
rect 10059 35848 10060 35888
rect 10100 35848 10101 35888
rect 10059 35839 10101 35848
rect 10531 35888 10589 35889
rect 10531 35848 10540 35888
rect 10580 35848 10589 35888
rect 11067 35857 11068 35897
rect 11108 35857 11109 35897
rect 11067 35848 11109 35857
rect 11395 35888 11453 35889
rect 11395 35848 11404 35888
rect 11444 35848 11453 35888
rect 10531 35847 10589 35848
rect 11395 35847 11453 35848
rect 12643 35888 12701 35889
rect 12643 35848 12652 35888
rect 12692 35848 12701 35888
rect 12643 35847 12701 35848
rect 13411 35888 13469 35889
rect 13411 35848 13420 35888
rect 13460 35848 13469 35888
rect 13411 35847 13469 35848
rect 14659 35888 14717 35889
rect 14659 35848 14668 35888
rect 14708 35848 14717 35888
rect 14659 35847 14717 35848
rect 15043 35888 15101 35889
rect 15043 35848 15052 35888
rect 15092 35848 15101 35888
rect 15043 35847 15101 35848
rect 16291 35888 16349 35889
rect 16291 35848 16300 35888
rect 16340 35848 16349 35888
rect 16291 35847 16349 35848
rect 16867 35888 16925 35889
rect 16867 35848 16876 35888
rect 16916 35848 16925 35888
rect 16867 35847 16925 35848
rect 18115 35888 18173 35889
rect 18115 35848 18124 35888
rect 18164 35848 18173 35888
rect 18115 35847 18173 35848
rect 18499 35888 18557 35889
rect 18499 35848 18508 35888
rect 18548 35848 18557 35888
rect 18499 35847 18557 35848
rect 19747 35888 19805 35889
rect 19747 35848 19756 35888
rect 19796 35848 19805 35888
rect 19747 35847 19805 35848
rect 6699 35804 6741 35813
rect 6699 35764 6700 35804
rect 6740 35764 6741 35804
rect 6699 35755 6741 35764
rect 11211 35804 11253 35813
rect 11211 35764 11212 35804
rect 11252 35764 11253 35804
rect 11211 35755 11253 35764
rect 5451 35720 5493 35729
rect 5451 35680 5452 35720
rect 5492 35680 5493 35720
rect 5451 35671 5493 35680
rect 12843 35720 12885 35729
rect 12843 35680 12844 35720
rect 12884 35680 12885 35720
rect 12843 35671 12885 35680
rect 14859 35720 14901 35729
rect 14859 35680 14860 35720
rect 14900 35680 14901 35720
rect 14859 35671 14901 35680
rect 16491 35720 16533 35729
rect 16491 35680 16492 35720
rect 16532 35680 16533 35720
rect 16491 35671 16533 35680
rect 1152 35552 20452 35576
rect 1152 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20452 35552
rect 1152 35488 20452 35512
rect 11115 35384 11157 35393
rect 11115 35344 11116 35384
rect 11156 35344 11157 35384
rect 11115 35335 11157 35344
rect 3723 35300 3765 35309
rect 3723 35260 3724 35300
rect 3764 35260 3765 35300
rect 3723 35251 3765 35260
rect 6027 35300 6069 35309
rect 6027 35260 6028 35300
rect 6068 35260 6069 35300
rect 6027 35251 6069 35260
rect 13995 35300 14037 35309
rect 13995 35260 13996 35300
rect 14036 35260 14037 35300
rect 13995 35251 14037 35260
rect 1995 35216 2037 35225
rect 1995 35176 1996 35216
rect 2036 35176 2037 35216
rect 1995 35167 2037 35176
rect 2091 35216 2133 35225
rect 2091 35176 2092 35216
rect 2132 35176 2133 35216
rect 2091 35167 2133 35176
rect 2571 35216 2613 35225
rect 2571 35176 2572 35216
rect 2612 35176 2613 35216
rect 2571 35167 2613 35176
rect 3043 35216 3101 35217
rect 3043 35176 3052 35216
rect 3092 35176 3101 35216
rect 5259 35216 5301 35225
rect 3043 35175 3101 35176
rect 3531 35202 3573 35211
rect 3531 35162 3532 35202
rect 3572 35162 3573 35202
rect 5259 35176 5260 35216
rect 5300 35176 5301 35216
rect 5259 35167 5301 35176
rect 5355 35216 5397 35225
rect 5355 35176 5356 35216
rect 5396 35176 5397 35216
rect 5355 35167 5397 35176
rect 5451 35216 5493 35225
rect 5451 35176 5452 35216
rect 5492 35176 5493 35216
rect 5451 35167 5493 35176
rect 5547 35216 5589 35225
rect 5547 35176 5548 35216
rect 5588 35176 5589 35216
rect 5547 35167 5589 35176
rect 5739 35216 5781 35225
rect 5739 35176 5740 35216
rect 5780 35176 5781 35216
rect 5739 35167 5781 35176
rect 5835 35216 5877 35225
rect 5835 35176 5836 35216
rect 5876 35176 5877 35216
rect 5835 35167 5877 35176
rect 5931 35216 5973 35225
rect 5931 35176 5932 35216
rect 5972 35176 5973 35216
rect 5931 35167 5973 35176
rect 6307 35216 6365 35217
rect 6307 35176 6316 35216
rect 6356 35176 6365 35216
rect 6307 35175 6365 35176
rect 6603 35216 6645 35225
rect 6603 35176 6604 35216
rect 6644 35176 6645 35216
rect 6603 35167 6645 35176
rect 6699 35216 6741 35225
rect 6699 35176 6700 35216
rect 6740 35176 6741 35216
rect 6699 35167 6741 35176
rect 7171 35216 7229 35217
rect 7171 35176 7180 35216
rect 7220 35176 7229 35216
rect 7171 35175 7229 35176
rect 9667 35216 9725 35217
rect 9667 35176 9676 35216
rect 9716 35176 9725 35216
rect 9667 35175 9725 35176
rect 10915 35216 10973 35217
rect 10915 35176 10924 35216
rect 10964 35176 10973 35216
rect 10915 35175 10973 35176
rect 12267 35216 12309 35225
rect 12267 35176 12268 35216
rect 12308 35176 12309 35216
rect 12267 35167 12309 35176
rect 12363 35216 12405 35225
rect 12363 35176 12364 35216
rect 12404 35176 12405 35216
rect 12363 35167 12405 35176
rect 13315 35216 13373 35217
rect 13315 35176 13324 35216
rect 13364 35176 13373 35216
rect 15619 35216 15677 35217
rect 13315 35175 13373 35176
rect 13803 35202 13845 35211
rect 3531 35153 3573 35162
rect 13803 35162 13804 35202
rect 13844 35162 13845 35202
rect 15619 35176 15628 35216
rect 15668 35176 15677 35216
rect 15619 35175 15677 35176
rect 16867 35216 16925 35217
rect 16867 35176 16876 35216
rect 16916 35176 16925 35216
rect 16867 35175 16925 35176
rect 17251 35216 17309 35217
rect 17251 35176 17260 35216
rect 17300 35176 17309 35216
rect 17251 35175 17309 35176
rect 18499 35216 18557 35217
rect 18499 35176 18508 35216
rect 18548 35176 18557 35216
rect 18499 35175 18557 35176
rect 13803 35153 13845 35162
rect 2475 35132 2517 35141
rect 2475 35092 2476 35132
rect 2516 35092 2517 35132
rect 2475 35083 2517 35092
rect 12747 35132 12789 35141
rect 12747 35092 12748 35132
rect 12788 35092 12789 35132
rect 12747 35083 12789 35092
rect 12843 35132 12885 35141
rect 12843 35092 12844 35132
rect 12884 35092 12885 35132
rect 12843 35083 12885 35092
rect 6979 35048 7037 35049
rect 6979 35008 6988 35048
rect 7028 35008 7037 35048
rect 6979 35007 7037 35008
rect 7275 34964 7317 34973
rect 7275 34924 7276 34964
rect 7316 34924 7317 34964
rect 7275 34915 7317 34924
rect 17067 34964 17109 34973
rect 17067 34924 17068 34964
rect 17108 34924 17109 34964
rect 17067 34915 17109 34924
rect 18699 34964 18741 34973
rect 18699 34924 18700 34964
rect 18740 34924 18741 34964
rect 18699 34915 18741 34924
rect 1152 34796 20352 34820
rect 1152 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 20352 34796
rect 1152 34732 20352 34756
rect 3243 34628 3285 34637
rect 3243 34588 3244 34628
rect 3284 34588 3285 34628
rect 3243 34579 3285 34588
rect 13803 34628 13845 34637
rect 13803 34588 13804 34628
rect 13844 34588 13845 34628
rect 13803 34579 13845 34588
rect 5451 34544 5493 34553
rect 5451 34504 5452 34544
rect 5492 34504 5493 34544
rect 5451 34495 5493 34504
rect 1795 34376 1853 34377
rect 1795 34336 1804 34376
rect 1844 34336 1853 34376
rect 1795 34335 1853 34336
rect 3043 34376 3101 34377
rect 3043 34336 3052 34376
rect 3092 34336 3101 34376
rect 3043 34335 3101 34336
rect 4003 34376 4061 34377
rect 4003 34336 4012 34376
rect 4052 34336 4061 34376
rect 4003 34335 4061 34336
rect 5251 34376 5309 34377
rect 5251 34336 5260 34376
rect 5300 34336 5309 34376
rect 5251 34335 5309 34336
rect 5731 34376 5789 34377
rect 5731 34336 5740 34376
rect 5780 34336 5789 34376
rect 5731 34335 5789 34336
rect 5835 34376 5877 34385
rect 5835 34336 5836 34376
rect 5876 34336 5877 34376
rect 5835 34327 5877 34336
rect 6123 34376 6165 34385
rect 6123 34336 6124 34376
rect 6164 34336 6165 34376
rect 6123 34327 6165 34336
rect 6219 34376 6261 34385
rect 6219 34336 6220 34376
rect 6260 34336 6261 34376
rect 6219 34327 6261 34336
rect 6315 34376 6357 34385
rect 6315 34336 6316 34376
rect 6356 34336 6357 34376
rect 6315 34327 6357 34336
rect 6499 34376 6557 34377
rect 6499 34336 6508 34376
rect 6548 34336 6557 34376
rect 6499 34335 6557 34336
rect 6603 34376 6645 34385
rect 6603 34336 6604 34376
rect 6644 34336 6645 34376
rect 6603 34327 6645 34336
rect 6795 34376 6837 34385
rect 6795 34336 6796 34376
rect 6836 34336 6837 34376
rect 6795 34327 6837 34336
rect 6987 34376 7029 34385
rect 6987 34336 6988 34376
rect 7028 34336 7029 34376
rect 6987 34327 7029 34336
rect 7083 34376 7125 34385
rect 7083 34336 7084 34376
rect 7124 34336 7125 34376
rect 7083 34327 7125 34336
rect 7179 34376 7221 34385
rect 7179 34336 7180 34376
rect 7220 34336 7221 34376
rect 7179 34327 7221 34336
rect 7275 34376 7317 34385
rect 7275 34336 7276 34376
rect 7316 34336 7317 34376
rect 7275 34327 7317 34336
rect 7555 34376 7613 34377
rect 7555 34336 7564 34376
rect 7604 34336 7613 34376
rect 7555 34335 7613 34336
rect 8803 34376 8861 34377
rect 8803 34336 8812 34376
rect 8852 34336 8861 34376
rect 9387 34376 9429 34385
rect 8803 34335 8861 34336
rect 9291 34356 9333 34365
rect 9291 34316 9292 34356
rect 9332 34316 9333 34356
rect 9387 34336 9388 34376
rect 9428 34336 9429 34376
rect 9387 34327 9429 34336
rect 9771 34376 9813 34385
rect 9771 34336 9772 34376
rect 9812 34336 9813 34376
rect 9771 34327 9813 34336
rect 9867 34376 9909 34385
rect 10827 34381 10869 34390
rect 9867 34336 9868 34376
rect 9908 34336 9909 34376
rect 9867 34327 9909 34336
rect 10339 34376 10397 34377
rect 10339 34336 10348 34376
rect 10388 34336 10397 34376
rect 10339 34335 10397 34336
rect 10827 34341 10828 34381
rect 10868 34341 10869 34381
rect 10827 34332 10869 34341
rect 12355 34376 12413 34377
rect 12355 34336 12364 34376
rect 12404 34336 12413 34376
rect 12355 34335 12413 34336
rect 13603 34376 13661 34377
rect 13603 34336 13612 34376
rect 13652 34336 13661 34376
rect 13603 34335 13661 34336
rect 14179 34376 14237 34377
rect 14179 34336 14188 34376
rect 14228 34336 14237 34376
rect 14179 34335 14237 34336
rect 15427 34376 15485 34377
rect 15427 34336 15436 34376
rect 15476 34336 15485 34376
rect 15427 34335 15485 34336
rect 15811 34376 15869 34377
rect 15811 34336 15820 34376
rect 15860 34336 15869 34376
rect 15811 34335 15869 34336
rect 17059 34376 17117 34377
rect 17059 34336 17068 34376
rect 17108 34336 17117 34376
rect 17059 34335 17117 34336
rect 17835 34376 17877 34385
rect 17835 34336 17836 34376
rect 17876 34336 17877 34376
rect 17835 34327 17877 34336
rect 17931 34376 17973 34385
rect 17931 34336 17932 34376
rect 17972 34336 17973 34376
rect 17931 34327 17973 34336
rect 18315 34376 18357 34385
rect 18315 34336 18316 34376
rect 18356 34336 18357 34376
rect 18315 34327 18357 34336
rect 18411 34376 18453 34385
rect 19371 34381 19413 34390
rect 18411 34336 18412 34376
rect 18452 34336 18453 34376
rect 18411 34327 18453 34336
rect 18883 34376 18941 34377
rect 18883 34336 18892 34376
rect 18932 34336 18941 34376
rect 18883 34335 18941 34336
rect 19371 34341 19372 34381
rect 19412 34341 19413 34381
rect 19371 34332 19413 34341
rect 9291 34307 9333 34316
rect 6699 34292 6741 34301
rect 6699 34252 6700 34292
rect 6740 34252 6741 34292
rect 6699 34243 6741 34252
rect 11019 34292 11061 34301
rect 11019 34252 11020 34292
rect 11060 34252 11061 34292
rect 11019 34243 11061 34252
rect 19563 34292 19605 34301
rect 19563 34252 19564 34292
rect 19604 34252 19605 34292
rect 19563 34243 19605 34252
rect 6019 34208 6077 34209
rect 6019 34168 6028 34208
rect 6068 34168 6077 34208
rect 6019 34167 6077 34168
rect 9003 34208 9045 34217
rect 9003 34168 9004 34208
rect 9044 34168 9045 34208
rect 9003 34159 9045 34168
rect 13995 34208 14037 34217
rect 13995 34168 13996 34208
rect 14036 34168 14037 34208
rect 13995 34159 14037 34168
rect 15627 34208 15669 34217
rect 15627 34168 15628 34208
rect 15668 34168 15669 34208
rect 15627 34159 15669 34168
rect 1152 34040 20452 34064
rect 1152 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20452 34040
rect 1152 33976 20452 34000
rect 4011 33872 4053 33881
rect 4011 33832 4012 33872
rect 4052 33832 4053 33872
rect 4011 33823 4053 33832
rect 7363 33872 7421 33873
rect 7363 33832 7372 33872
rect 7412 33832 7421 33872
rect 7363 33831 7421 33832
rect 8995 33872 9053 33873
rect 8995 33832 9004 33872
rect 9044 33832 9053 33872
rect 8995 33831 9053 33832
rect 10635 33872 10677 33881
rect 10635 33832 10636 33872
rect 10676 33832 10677 33872
rect 10635 33823 10677 33832
rect 12651 33872 12693 33881
rect 12651 33832 12652 33872
rect 12692 33832 12693 33872
rect 12651 33823 12693 33832
rect 16395 33872 16437 33881
rect 16395 33832 16396 33872
rect 16436 33832 16437 33872
rect 16395 33823 16437 33832
rect 18027 33872 18069 33881
rect 18027 33832 18028 33872
rect 18068 33832 18069 33872
rect 18027 33823 18069 33832
rect 20235 33872 20277 33881
rect 20235 33832 20236 33872
rect 20276 33832 20277 33872
rect 20235 33823 20277 33832
rect 5739 33788 5781 33797
rect 5739 33748 5740 33788
rect 5780 33748 5781 33788
rect 5739 33739 5781 33748
rect 2283 33704 2325 33713
rect 2283 33664 2284 33704
rect 2324 33664 2325 33704
rect 2283 33655 2325 33664
rect 2379 33704 2421 33713
rect 2379 33664 2380 33704
rect 2420 33664 2421 33704
rect 2379 33655 2421 33664
rect 3331 33704 3389 33705
rect 3331 33664 3340 33704
rect 3380 33664 3389 33704
rect 4291 33704 4349 33705
rect 3331 33663 3389 33664
rect 3819 33690 3861 33699
rect 3819 33650 3820 33690
rect 3860 33650 3861 33690
rect 4291 33664 4300 33704
rect 4340 33664 4349 33704
rect 4291 33663 4349 33664
rect 5539 33704 5597 33705
rect 5539 33664 5548 33704
rect 5588 33664 5597 33704
rect 5539 33663 5597 33664
rect 5923 33704 5981 33705
rect 5923 33664 5932 33704
rect 5972 33664 5981 33704
rect 5923 33663 5981 33664
rect 6027 33704 6069 33713
rect 6027 33664 6028 33704
rect 6068 33664 6069 33704
rect 6027 33655 6069 33664
rect 6307 33704 6365 33705
rect 6307 33664 6316 33704
rect 6356 33664 6365 33704
rect 6307 33663 6365 33664
rect 6603 33704 6645 33713
rect 6603 33664 6604 33704
rect 6644 33664 6645 33704
rect 6603 33655 6645 33664
rect 6699 33704 6741 33713
rect 6699 33664 6700 33704
rect 6740 33664 6741 33704
rect 6699 33655 6741 33664
rect 7171 33704 7229 33705
rect 7171 33664 7180 33704
rect 7220 33664 7229 33704
rect 7171 33663 7229 33664
rect 7275 33704 7317 33713
rect 7275 33664 7276 33704
rect 7316 33664 7317 33704
rect 7275 33655 7317 33664
rect 7467 33704 7509 33713
rect 7467 33664 7468 33704
rect 7508 33664 7509 33704
rect 7467 33655 7509 33664
rect 7659 33704 7701 33713
rect 7659 33664 7660 33704
rect 7700 33664 7701 33704
rect 7659 33655 7701 33664
rect 7851 33704 7893 33713
rect 7851 33664 7852 33704
rect 7892 33664 7893 33704
rect 7851 33655 7893 33664
rect 7939 33704 7997 33705
rect 7939 33664 7948 33704
rect 7988 33664 7997 33704
rect 7939 33663 7997 33664
rect 8235 33704 8277 33713
rect 8235 33664 8236 33704
rect 8276 33664 8277 33704
rect 8235 33655 8277 33664
rect 8427 33704 8469 33713
rect 8427 33664 8428 33704
rect 8468 33664 8469 33704
rect 8427 33655 8469 33664
rect 8523 33704 8565 33713
rect 8523 33664 8524 33704
rect 8564 33664 8565 33704
rect 8523 33655 8565 33664
rect 8715 33704 8757 33713
rect 8715 33664 8716 33704
rect 8756 33664 8757 33704
rect 8715 33655 8757 33664
rect 8811 33704 8853 33713
rect 8811 33664 8812 33704
rect 8852 33664 8853 33704
rect 8811 33655 8853 33664
rect 9187 33704 9245 33705
rect 9187 33664 9196 33704
rect 9236 33664 9245 33704
rect 9187 33663 9245 33664
rect 10435 33704 10493 33705
rect 10435 33664 10444 33704
rect 10484 33664 10493 33704
rect 10435 33663 10493 33664
rect 10923 33704 10965 33713
rect 10923 33664 10924 33704
rect 10964 33664 10965 33704
rect 10923 33655 10965 33664
rect 11019 33704 11061 33713
rect 11019 33664 11020 33704
rect 11060 33664 11061 33704
rect 11019 33655 11061 33664
rect 11403 33704 11445 33713
rect 11403 33664 11404 33704
rect 11444 33664 11445 33704
rect 11403 33655 11445 33664
rect 11971 33704 12029 33705
rect 11971 33664 11980 33704
rect 12020 33664 12029 33704
rect 12931 33704 12989 33705
rect 11971 33663 12029 33664
rect 12459 33690 12501 33699
rect 3819 33641 3861 33650
rect 12459 33650 12460 33690
rect 12500 33650 12501 33690
rect 12931 33664 12940 33704
rect 12980 33664 12989 33704
rect 12931 33663 12989 33664
rect 14179 33704 14237 33705
rect 14179 33664 14188 33704
rect 14228 33664 14237 33704
rect 14179 33663 14237 33664
rect 14667 33704 14709 33713
rect 14667 33664 14668 33704
rect 14708 33664 14709 33704
rect 14667 33655 14709 33664
rect 14763 33704 14805 33713
rect 14763 33664 14764 33704
rect 14804 33664 14805 33704
rect 14763 33655 14805 33664
rect 15715 33704 15773 33705
rect 15715 33664 15724 33704
rect 15764 33664 15773 33704
rect 15715 33663 15773 33664
rect 16203 33699 16245 33708
rect 16203 33659 16204 33699
rect 16244 33659 16245 33699
rect 16579 33704 16637 33705
rect 16579 33664 16588 33704
rect 16628 33664 16637 33704
rect 16579 33663 16637 33664
rect 17827 33704 17885 33705
rect 17827 33664 17836 33704
rect 17876 33664 17885 33704
rect 17827 33663 17885 33664
rect 18507 33704 18549 33713
rect 18507 33664 18508 33704
rect 18548 33664 18549 33704
rect 16203 33650 16245 33659
rect 18507 33655 18549 33664
rect 18603 33704 18645 33713
rect 18603 33664 18604 33704
rect 18644 33664 18645 33704
rect 18603 33655 18645 33664
rect 19555 33704 19613 33705
rect 19555 33664 19564 33704
rect 19604 33664 19613 33704
rect 19555 33663 19613 33664
rect 20043 33690 20085 33699
rect 20043 33650 20044 33690
rect 20084 33650 20085 33690
rect 12459 33641 12501 33650
rect 20043 33641 20085 33650
rect 2763 33620 2805 33629
rect 2763 33580 2764 33620
rect 2804 33580 2805 33620
rect 2763 33571 2805 33580
rect 2859 33620 2901 33629
rect 2859 33580 2860 33620
rect 2900 33580 2901 33620
rect 2859 33571 2901 33580
rect 11499 33620 11541 33629
rect 11499 33580 11500 33620
rect 11540 33580 11541 33620
rect 11499 33571 11541 33580
rect 15147 33620 15189 33629
rect 15147 33580 15148 33620
rect 15188 33580 15189 33620
rect 15147 33571 15189 33580
rect 15243 33620 15285 33629
rect 15243 33580 15244 33620
rect 15284 33580 15285 33620
rect 15243 33571 15285 33580
rect 18987 33620 19029 33629
rect 18987 33580 18988 33620
rect 19028 33580 19029 33620
rect 18987 33571 19029 33580
rect 19083 33620 19125 33629
rect 19083 33580 19084 33620
rect 19124 33580 19125 33620
rect 19083 33571 19125 33580
rect 6979 33536 7037 33537
rect 6979 33496 6988 33536
rect 7028 33496 7037 33536
rect 6979 33495 7037 33496
rect 7659 33536 7701 33545
rect 7659 33496 7660 33536
rect 7700 33496 7701 33536
rect 7659 33487 7701 33496
rect 8515 33536 8573 33537
rect 8515 33496 8524 33536
rect 8564 33496 8573 33536
rect 8515 33495 8573 33496
rect 14379 33452 14421 33461
rect 14379 33412 14380 33452
rect 14420 33412 14421 33452
rect 14379 33403 14421 33412
rect 1152 33284 20352 33308
rect 1152 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 20352 33284
rect 1152 33220 20352 33244
rect 2667 33116 2709 33125
rect 2667 33076 2668 33116
rect 2708 33076 2709 33116
rect 2667 33067 2709 33076
rect 5643 33116 5685 33125
rect 5643 33076 5644 33116
rect 5684 33076 5685 33116
rect 5643 33067 5685 33076
rect 6979 33116 7037 33117
rect 6979 33076 6988 33116
rect 7028 33076 7037 33116
rect 6979 33075 7037 33076
rect 12459 33116 12501 33125
rect 12459 33076 12460 33116
rect 12500 33076 12501 33116
rect 12459 33067 12501 33076
rect 19371 33116 19413 33125
rect 19371 33076 19372 33116
rect 19412 33076 19413 33116
rect 19371 33067 19413 33076
rect 9195 33032 9237 33041
rect 9195 32992 9196 33032
rect 9236 32992 9237 33032
rect 9195 32983 9237 32992
rect 10827 33032 10869 33041
rect 10827 32992 10828 33032
rect 10868 32992 10869 33032
rect 10827 32983 10869 32992
rect 5931 32948 5973 32957
rect 5931 32908 5932 32948
rect 5972 32908 5973 32948
rect 5931 32899 5973 32908
rect 16347 32873 16389 32882
rect 1219 32864 1277 32865
rect 1219 32824 1228 32864
rect 1268 32824 1277 32864
rect 1219 32823 1277 32824
rect 2467 32864 2525 32865
rect 2467 32824 2476 32864
rect 2516 32824 2525 32864
rect 2467 32823 2525 32824
rect 4195 32864 4253 32865
rect 4195 32824 4204 32864
rect 4244 32824 4253 32864
rect 4195 32823 4253 32824
rect 5443 32864 5501 32865
rect 5443 32824 5452 32864
rect 5492 32824 5501 32864
rect 5443 32823 5501 32824
rect 5835 32864 5877 32873
rect 5835 32824 5836 32864
rect 5876 32824 5877 32864
rect 5835 32815 5877 32824
rect 6027 32864 6069 32873
rect 6027 32824 6028 32864
rect 6068 32824 6069 32864
rect 6027 32815 6069 32824
rect 6307 32864 6365 32865
rect 6307 32824 6316 32864
rect 6356 32824 6365 32864
rect 6307 32823 6365 32824
rect 6603 32864 6645 32873
rect 6603 32824 6604 32864
rect 6644 32824 6645 32864
rect 6603 32815 6645 32824
rect 7179 32864 7221 32873
rect 7179 32824 7180 32864
rect 7220 32824 7221 32864
rect 7179 32815 7221 32824
rect 7275 32864 7317 32873
rect 7275 32824 7276 32864
rect 7316 32824 7317 32864
rect 7275 32815 7317 32824
rect 7371 32864 7413 32873
rect 7371 32824 7372 32864
rect 7412 32824 7413 32864
rect 7371 32815 7413 32824
rect 7467 32864 7509 32873
rect 7467 32824 7468 32864
rect 7508 32824 7509 32864
rect 7467 32815 7509 32824
rect 7747 32864 7805 32865
rect 7747 32824 7756 32864
rect 7796 32824 7805 32864
rect 7747 32823 7805 32824
rect 8995 32864 9053 32865
rect 8995 32824 9004 32864
rect 9044 32824 9053 32864
rect 8995 32823 9053 32824
rect 9379 32864 9437 32865
rect 9379 32824 9388 32864
rect 9428 32824 9437 32864
rect 9379 32823 9437 32824
rect 10627 32864 10685 32865
rect 10627 32824 10636 32864
rect 10676 32824 10685 32864
rect 10627 32823 10685 32824
rect 12259 32864 12317 32865
rect 12259 32824 12268 32864
rect 12308 32824 12317 32864
rect 12259 32823 12317 32824
rect 14763 32864 14805 32873
rect 14763 32824 14764 32864
rect 14804 32824 14805 32864
rect 11011 32822 11069 32823
rect 6699 32780 6741 32789
rect 11011 32782 11020 32822
rect 11060 32782 11069 32822
rect 14763 32815 14805 32824
rect 14859 32864 14901 32873
rect 14859 32824 14860 32864
rect 14900 32824 14901 32864
rect 14859 32815 14901 32824
rect 15243 32864 15285 32873
rect 15243 32824 15244 32864
rect 15284 32824 15285 32864
rect 15243 32815 15285 32824
rect 15339 32864 15381 32873
rect 15339 32824 15340 32864
rect 15380 32824 15381 32864
rect 15339 32815 15381 32824
rect 15811 32864 15869 32865
rect 15811 32824 15820 32864
rect 15860 32824 15869 32864
rect 16347 32833 16348 32873
rect 16388 32833 16389 32873
rect 16347 32824 16389 32833
rect 17923 32864 17981 32865
rect 17923 32824 17932 32864
rect 17972 32824 17981 32864
rect 15811 32823 15869 32824
rect 17923 32823 17981 32824
rect 19171 32864 19229 32865
rect 19171 32824 19180 32864
rect 19220 32824 19229 32864
rect 19171 32823 19229 32824
rect 11011 32781 11069 32782
rect 6699 32740 6700 32780
rect 6740 32740 6741 32780
rect 6699 32731 6741 32740
rect 16491 32780 16533 32789
rect 16491 32740 16492 32780
rect 16532 32740 16533 32780
rect 16491 32731 16533 32740
rect 1152 32528 20452 32552
rect 1152 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20452 32528
rect 1152 32464 20452 32488
rect 5451 32360 5493 32369
rect 5451 32320 5452 32360
rect 5492 32320 5493 32360
rect 5451 32311 5493 32320
rect 9099 32360 9141 32369
rect 9099 32320 9100 32360
rect 9140 32320 9141 32360
rect 9099 32311 9141 32320
rect 9475 32360 9533 32361
rect 9475 32320 9484 32360
rect 9524 32320 9533 32360
rect 9475 32319 9533 32320
rect 16491 32360 16533 32369
rect 16491 32320 16492 32360
rect 16532 32320 16533 32360
rect 16491 32311 16533 32320
rect 3723 32276 3765 32285
rect 3723 32236 3724 32276
rect 3764 32236 3765 32276
rect 3723 32227 3765 32236
rect 12171 32276 12213 32285
rect 12171 32236 12172 32276
rect 12212 32236 12213 32276
rect 12171 32227 12213 32236
rect 14187 32276 14229 32285
rect 14187 32236 14188 32276
rect 14228 32236 14229 32276
rect 14187 32227 14229 32236
rect 19467 32276 19509 32285
rect 19467 32236 19468 32276
rect 19508 32236 19509 32276
rect 19467 32227 19509 32236
rect 1995 32192 2037 32201
rect 1995 32152 1996 32192
rect 2036 32152 2037 32192
rect 1995 32143 2037 32152
rect 2091 32192 2133 32201
rect 2091 32152 2092 32192
rect 2132 32152 2133 32192
rect 2091 32143 2133 32152
rect 2571 32192 2613 32201
rect 2571 32152 2572 32192
rect 2612 32152 2613 32192
rect 2571 32143 2613 32152
rect 3043 32192 3101 32193
rect 3043 32152 3052 32192
rect 3092 32152 3101 32192
rect 5731 32192 5789 32193
rect 3043 32151 3101 32152
rect 3531 32178 3573 32187
rect 3531 32138 3532 32178
rect 3572 32138 3573 32178
rect 5731 32152 5740 32192
rect 5780 32152 5789 32192
rect 5731 32151 5789 32152
rect 6979 32192 7037 32193
rect 6979 32152 6988 32192
rect 7028 32152 7037 32192
rect 6979 32151 7037 32152
rect 7651 32192 7709 32193
rect 7651 32152 7660 32192
rect 7700 32152 7709 32192
rect 7651 32151 7709 32152
rect 8899 32192 8957 32193
rect 8899 32152 8908 32192
rect 8948 32152 8957 32192
rect 8899 32151 8957 32152
rect 9283 32192 9341 32193
rect 9283 32152 9292 32192
rect 9332 32152 9341 32192
rect 9283 32151 9341 32152
rect 9379 32192 9437 32193
rect 9379 32152 9388 32192
rect 9428 32152 9437 32192
rect 9379 32151 9437 32152
rect 9579 32192 9621 32201
rect 9579 32152 9580 32192
rect 9620 32152 9621 32192
rect 9579 32143 9621 32152
rect 9675 32192 9717 32201
rect 9675 32152 9676 32192
rect 9716 32152 9717 32192
rect 9675 32143 9717 32152
rect 9768 32192 9826 32193
rect 9768 32152 9777 32192
rect 9817 32152 9826 32192
rect 9768 32151 9826 32152
rect 10051 32192 10109 32193
rect 10051 32152 10060 32192
rect 10100 32152 10109 32192
rect 10051 32151 10109 32152
rect 10155 32192 10197 32201
rect 10155 32152 10156 32192
rect 10196 32152 10197 32192
rect 10155 32143 10197 32152
rect 10723 32192 10781 32193
rect 10723 32152 10732 32192
rect 10772 32152 10781 32192
rect 10723 32151 10781 32152
rect 11971 32192 12029 32193
rect 11971 32152 11980 32192
rect 12020 32152 12029 32192
rect 11971 32151 12029 32152
rect 12459 32192 12501 32201
rect 12459 32152 12460 32192
rect 12500 32152 12501 32192
rect 12459 32143 12501 32152
rect 12555 32192 12597 32201
rect 12555 32152 12556 32192
rect 12596 32152 12597 32192
rect 12555 32143 12597 32152
rect 13507 32192 13565 32193
rect 13507 32152 13516 32192
rect 13556 32152 13565 32192
rect 15043 32192 15101 32193
rect 13507 32151 13565 32152
rect 13995 32178 14037 32187
rect 3531 32129 3573 32138
rect 13995 32138 13996 32178
rect 14036 32138 14037 32178
rect 15043 32152 15052 32192
rect 15092 32152 15101 32192
rect 15043 32151 15101 32152
rect 16291 32192 16349 32193
rect 16291 32152 16300 32192
rect 16340 32152 16349 32192
rect 16291 32151 16349 32152
rect 17739 32192 17781 32201
rect 17739 32152 17740 32192
rect 17780 32152 17781 32192
rect 17739 32143 17781 32152
rect 17835 32192 17877 32201
rect 17835 32152 17836 32192
rect 17876 32152 17877 32192
rect 17835 32143 17877 32152
rect 18219 32192 18261 32201
rect 18219 32152 18220 32192
rect 18260 32152 18261 32192
rect 18219 32143 18261 32152
rect 18787 32192 18845 32193
rect 18787 32152 18796 32192
rect 18836 32152 18845 32192
rect 18787 32151 18845 32152
rect 19275 32178 19317 32187
rect 13995 32129 14037 32138
rect 19275 32138 19276 32178
rect 19316 32138 19317 32178
rect 19275 32129 19317 32138
rect 2475 32108 2517 32117
rect 2475 32068 2476 32108
rect 2516 32068 2517 32108
rect 2475 32059 2517 32068
rect 12939 32108 12981 32117
rect 12939 32068 12940 32108
rect 12980 32068 12981 32108
rect 12939 32059 12981 32068
rect 13035 32108 13077 32117
rect 13035 32068 13036 32108
rect 13076 32068 13077 32108
rect 13035 32059 13077 32068
rect 18315 32108 18357 32117
rect 18315 32068 18316 32108
rect 18356 32068 18357 32108
rect 18315 32059 18357 32068
rect 7179 31940 7221 31949
rect 7179 31900 7180 31940
rect 7220 31900 7221 31940
rect 7179 31891 7221 31900
rect 9291 31940 9333 31949
rect 9291 31900 9292 31940
rect 9332 31900 9333 31940
rect 9291 31891 9333 31900
rect 1152 31772 20352 31796
rect 1152 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 20352 31772
rect 1152 31708 20352 31732
rect 14091 31604 14133 31613
rect 14091 31564 14092 31604
rect 14132 31564 14133 31604
rect 14091 31555 14133 31564
rect 18123 31604 18165 31613
rect 18123 31564 18124 31604
rect 18164 31564 18165 31604
rect 18123 31555 18165 31564
rect 3051 31520 3093 31529
rect 3051 31480 3052 31520
rect 3092 31480 3093 31520
rect 3051 31471 3093 31480
rect 8043 31436 8085 31445
rect 8043 31396 8044 31436
rect 8084 31396 8085 31436
rect 8043 31387 8085 31396
rect 10059 31436 10101 31445
rect 10059 31396 10060 31436
rect 10100 31396 10101 31436
rect 10059 31387 10101 31396
rect 10155 31436 10197 31445
rect 10155 31396 10156 31436
rect 10196 31396 10197 31436
rect 10155 31387 10197 31396
rect 15339 31436 15381 31445
rect 15339 31396 15340 31436
rect 15380 31396 15381 31436
rect 15339 31387 15381 31396
rect 18987 31436 19029 31445
rect 18987 31396 18988 31436
rect 19028 31396 19029 31436
rect 18987 31387 19029 31396
rect 7083 31366 7125 31375
rect 1603 31352 1661 31353
rect 1603 31312 1612 31352
rect 1652 31312 1661 31352
rect 1603 31311 1661 31312
rect 2851 31352 2909 31353
rect 2851 31312 2860 31352
rect 2900 31312 2909 31352
rect 2851 31311 2909 31312
rect 3339 31352 3381 31361
rect 3339 31312 3340 31352
rect 3380 31312 3381 31352
rect 3339 31303 3381 31312
rect 3435 31352 3477 31361
rect 3435 31312 3436 31352
rect 3476 31312 3477 31352
rect 3435 31303 3477 31312
rect 3819 31352 3861 31361
rect 3819 31312 3820 31352
rect 3860 31312 3861 31352
rect 3819 31303 3861 31312
rect 3915 31352 3957 31361
rect 4875 31357 4917 31366
rect 3915 31312 3916 31352
rect 3956 31312 3957 31352
rect 3915 31303 3957 31312
rect 4387 31352 4445 31353
rect 4387 31312 4396 31352
rect 4436 31312 4445 31352
rect 4387 31311 4445 31312
rect 4875 31317 4876 31357
rect 4916 31317 4917 31357
rect 4875 31308 4917 31317
rect 5547 31352 5589 31361
rect 5547 31312 5548 31352
rect 5588 31312 5589 31352
rect 5547 31303 5589 31312
rect 5643 31352 5685 31361
rect 5643 31312 5644 31352
rect 5684 31312 5685 31352
rect 5643 31303 5685 31312
rect 6027 31352 6069 31361
rect 6027 31312 6028 31352
rect 6068 31312 6069 31352
rect 6027 31303 6069 31312
rect 6123 31352 6165 31361
rect 6123 31312 6124 31352
rect 6164 31312 6165 31352
rect 6123 31303 6165 31312
rect 6595 31352 6653 31353
rect 6595 31312 6604 31352
rect 6644 31312 6653 31352
rect 7083 31326 7084 31366
rect 7124 31326 7125 31366
rect 7083 31317 7125 31326
rect 7563 31352 7605 31361
rect 6595 31311 6653 31312
rect 7563 31312 7564 31352
rect 7604 31312 7605 31352
rect 7563 31303 7605 31312
rect 7659 31352 7701 31361
rect 7659 31312 7660 31352
rect 7700 31312 7701 31352
rect 7659 31303 7701 31312
rect 8139 31352 8181 31361
rect 9099 31357 9141 31366
rect 11163 31361 11205 31370
rect 8139 31312 8140 31352
rect 8180 31312 8181 31352
rect 8139 31303 8181 31312
rect 8611 31352 8669 31353
rect 8611 31312 8620 31352
rect 8660 31312 8669 31352
rect 8611 31311 8669 31312
rect 9099 31317 9100 31357
rect 9140 31317 9141 31357
rect 9099 31308 9141 31317
rect 9579 31352 9621 31361
rect 9579 31312 9580 31352
rect 9620 31312 9621 31352
rect 9579 31303 9621 31312
rect 9675 31352 9717 31361
rect 9675 31312 9676 31352
rect 9716 31312 9717 31352
rect 9675 31303 9717 31312
rect 10627 31352 10685 31353
rect 10627 31312 10636 31352
rect 10676 31312 10685 31352
rect 11163 31321 11164 31361
rect 11204 31321 11205 31361
rect 11163 31312 11205 31321
rect 12643 31352 12701 31353
rect 12643 31312 12652 31352
rect 12692 31312 12701 31352
rect 10627 31311 10685 31312
rect 12643 31311 12701 31312
rect 13891 31352 13949 31353
rect 13891 31312 13900 31352
rect 13940 31312 13949 31352
rect 13891 31311 13949 31312
rect 14371 31352 14429 31353
rect 14371 31312 14380 31352
rect 14420 31312 14429 31352
rect 14371 31311 14429 31312
rect 14763 31352 14805 31361
rect 14763 31312 14764 31352
rect 14804 31312 14805 31352
rect 14763 31303 14805 31312
rect 14859 31352 14901 31361
rect 14859 31312 14860 31352
rect 14900 31312 14901 31352
rect 14859 31303 14901 31312
rect 15243 31352 15285 31361
rect 16299 31357 16341 31366
rect 15243 31312 15244 31352
rect 15284 31312 15285 31352
rect 15243 31303 15285 31312
rect 15811 31352 15869 31353
rect 15811 31312 15820 31352
rect 15860 31312 15869 31352
rect 15811 31311 15869 31312
rect 16299 31317 16300 31357
rect 16340 31317 16341 31357
rect 16299 31308 16341 31317
rect 16675 31352 16733 31353
rect 16675 31312 16684 31352
rect 16724 31312 16733 31352
rect 16675 31311 16733 31312
rect 17923 31352 17981 31353
rect 17923 31312 17932 31352
rect 17972 31312 17981 31352
rect 17923 31311 17981 31312
rect 18411 31352 18453 31361
rect 18411 31312 18412 31352
rect 18452 31312 18453 31352
rect 18411 31303 18453 31312
rect 18507 31352 18549 31361
rect 18507 31312 18508 31352
rect 18548 31312 18549 31352
rect 18507 31303 18549 31312
rect 18891 31352 18933 31361
rect 19947 31357 19989 31366
rect 18891 31312 18892 31352
rect 18932 31312 18933 31352
rect 18891 31303 18933 31312
rect 19459 31352 19517 31353
rect 19459 31312 19468 31352
rect 19508 31312 19517 31352
rect 19459 31311 19517 31312
rect 19947 31317 19948 31357
rect 19988 31317 19989 31357
rect 19947 31308 19989 31317
rect 5067 31268 5109 31277
rect 5067 31228 5068 31268
rect 5108 31228 5109 31268
rect 5067 31219 5109 31228
rect 7275 31268 7317 31277
rect 7275 31228 7276 31268
rect 7316 31228 7317 31268
rect 7275 31219 7317 31228
rect 9291 31184 9333 31193
rect 9291 31144 9292 31184
rect 9332 31144 9333 31184
rect 9291 31135 9333 31144
rect 11307 31184 11349 31193
rect 11307 31144 11308 31184
rect 11348 31144 11349 31184
rect 11307 31135 11349 31144
rect 14283 31184 14325 31193
rect 14283 31144 14284 31184
rect 14324 31144 14325 31184
rect 14283 31135 14325 31144
rect 16491 31184 16533 31193
rect 16491 31144 16492 31184
rect 16532 31144 16533 31184
rect 16491 31135 16533 31144
rect 20139 31184 20181 31193
rect 20139 31144 20140 31184
rect 20180 31144 20181 31184
rect 20139 31135 20181 31144
rect 1152 31016 20452 31040
rect 1152 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20452 31016
rect 1152 30952 20452 30976
rect 2667 30848 2709 30857
rect 2667 30808 2668 30848
rect 2708 30808 2709 30848
rect 2667 30799 2709 30808
rect 5259 30848 5301 30857
rect 5259 30808 5260 30848
rect 5300 30808 5301 30848
rect 5259 30799 5301 30808
rect 5451 30848 5493 30857
rect 5451 30808 5452 30848
rect 5492 30808 5493 30848
rect 5451 30799 5493 30808
rect 7467 30848 7509 30857
rect 7467 30808 7468 30848
rect 7508 30808 7509 30848
rect 7467 30799 7509 30808
rect 9675 30848 9717 30857
rect 9675 30808 9676 30848
rect 9716 30808 9717 30848
rect 9675 30799 9717 30808
rect 11307 30848 11349 30857
rect 11307 30808 11308 30848
rect 11348 30808 11349 30848
rect 11307 30799 11349 30808
rect 15051 30848 15093 30857
rect 15051 30808 15052 30848
rect 15092 30808 15093 30848
rect 15051 30799 15093 30808
rect 16683 30848 16725 30857
rect 16683 30808 16684 30848
rect 16724 30808 16725 30848
rect 16683 30799 16725 30808
rect 18315 30848 18357 30857
rect 18315 30808 18316 30848
rect 18356 30808 18357 30848
rect 18315 30799 18357 30808
rect 20235 30848 20277 30857
rect 20235 30808 20236 30848
rect 20276 30808 20277 30848
rect 20235 30799 20277 30808
rect 1219 30680 1277 30681
rect 1219 30640 1228 30680
rect 1268 30640 1277 30680
rect 1219 30639 1277 30640
rect 2467 30680 2525 30681
rect 2467 30640 2476 30680
rect 2516 30640 2525 30680
rect 2467 30639 2525 30640
rect 3811 30680 3869 30681
rect 3811 30640 3820 30680
rect 3860 30640 3869 30680
rect 3811 30639 3869 30640
rect 5059 30680 5117 30681
rect 5059 30640 5068 30680
rect 5108 30640 5117 30680
rect 5059 30639 5117 30640
rect 6019 30680 6077 30681
rect 6019 30640 6028 30680
rect 6068 30640 6077 30680
rect 6019 30639 6077 30640
rect 7267 30680 7325 30681
rect 7267 30640 7276 30680
rect 7316 30640 7325 30680
rect 7267 30639 7325 30640
rect 8227 30680 8285 30681
rect 8227 30640 8236 30680
rect 8276 30640 8285 30680
rect 8227 30639 8285 30640
rect 9475 30680 9533 30681
rect 9475 30640 9484 30680
rect 9524 30640 9533 30680
rect 9475 30639 9533 30640
rect 9859 30680 9917 30681
rect 9859 30640 9868 30680
rect 9908 30640 9917 30680
rect 9859 30639 9917 30640
rect 11107 30680 11165 30681
rect 11107 30640 11116 30680
rect 11156 30640 11165 30680
rect 11107 30639 11165 30640
rect 11491 30680 11549 30681
rect 11491 30640 11500 30680
rect 11540 30640 11549 30680
rect 11491 30639 11549 30640
rect 12739 30680 12797 30681
rect 12739 30640 12748 30680
rect 12788 30640 12797 30680
rect 12739 30639 12797 30640
rect 13131 30680 13173 30689
rect 13131 30640 13132 30680
rect 13172 30640 13173 30680
rect 13131 30631 13173 30640
rect 13227 30680 13269 30689
rect 13227 30640 13228 30680
rect 13268 30640 13269 30680
rect 13227 30631 13269 30640
rect 13323 30680 13365 30689
rect 13323 30640 13324 30680
rect 13364 30640 13365 30680
rect 13323 30631 13365 30640
rect 13419 30680 13461 30689
rect 13419 30640 13420 30680
rect 13460 30640 13461 30680
rect 13419 30631 13461 30640
rect 13603 30680 13661 30681
rect 13603 30640 13612 30680
rect 13652 30640 13661 30680
rect 13603 30639 13661 30640
rect 14851 30680 14909 30681
rect 14851 30640 14860 30680
rect 14900 30640 14909 30680
rect 14851 30639 14909 30640
rect 15235 30680 15293 30681
rect 15235 30640 15244 30680
rect 15284 30640 15293 30680
rect 15235 30639 15293 30640
rect 16483 30680 16541 30681
rect 16483 30640 16492 30680
rect 16532 30640 16541 30680
rect 16483 30639 16541 30640
rect 16867 30680 16925 30681
rect 16867 30640 16876 30680
rect 16916 30640 16925 30680
rect 16867 30639 16925 30640
rect 18115 30680 18173 30681
rect 18115 30640 18124 30680
rect 18164 30640 18173 30680
rect 18115 30639 18173 30640
rect 18787 30680 18845 30681
rect 18787 30640 18796 30680
rect 18836 30640 18845 30680
rect 18787 30639 18845 30640
rect 20035 30680 20093 30681
rect 20035 30640 20044 30680
rect 20084 30640 20093 30680
rect 20035 30639 20093 30640
rect 12939 30428 12981 30437
rect 12939 30388 12940 30428
rect 12980 30388 12981 30428
rect 12939 30379 12981 30388
rect 1152 30260 20352 30284
rect 1152 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 20352 30260
rect 1152 30196 20352 30220
rect 5739 30092 5781 30101
rect 5739 30052 5740 30092
rect 5780 30052 5781 30092
rect 5739 30043 5781 30052
rect 9003 30092 9045 30101
rect 9003 30052 9004 30092
rect 9044 30052 9045 30092
rect 9003 30043 9045 30052
rect 17451 30092 17493 30101
rect 17451 30052 17452 30092
rect 17492 30052 17493 30092
rect 17451 30043 17493 30052
rect 14083 30008 14141 30009
rect 14083 29968 14092 30008
rect 14132 29968 14141 30008
rect 14083 29967 14141 29968
rect 2955 29924 2997 29933
rect 2955 29884 2956 29924
rect 2996 29884 2997 29924
rect 2955 29875 2997 29884
rect 12835 29882 12893 29883
rect 3963 29849 4005 29858
rect 2379 29840 2421 29849
rect 2379 29800 2380 29840
rect 2420 29800 2421 29840
rect 2379 29791 2421 29800
rect 2475 29840 2517 29849
rect 2475 29800 2476 29840
rect 2516 29800 2517 29840
rect 2475 29791 2517 29800
rect 2859 29840 2901 29849
rect 2859 29800 2860 29840
rect 2900 29800 2901 29840
rect 2859 29791 2901 29800
rect 3427 29840 3485 29841
rect 3427 29800 3436 29840
rect 3476 29800 3485 29840
rect 3963 29809 3964 29849
rect 4004 29809 4005 29849
rect 3963 29800 4005 29809
rect 4291 29840 4349 29841
rect 4291 29800 4300 29840
rect 4340 29800 4349 29840
rect 3427 29799 3485 29800
rect 4291 29799 4349 29800
rect 5539 29840 5597 29841
rect 5539 29800 5548 29840
rect 5588 29800 5597 29840
rect 5539 29799 5597 29800
rect 6315 29840 6357 29849
rect 6315 29800 6316 29840
rect 6356 29800 6357 29840
rect 6315 29791 6357 29800
rect 6411 29840 6453 29849
rect 6411 29800 6412 29840
rect 6452 29800 6453 29840
rect 6411 29791 6453 29800
rect 6507 29840 6549 29849
rect 12835 29842 12844 29882
rect 12884 29842 12893 29882
rect 12835 29841 12893 29842
rect 6507 29800 6508 29840
rect 6548 29800 6549 29840
rect 6507 29791 6549 29800
rect 6691 29840 6749 29841
rect 6691 29800 6700 29840
rect 6740 29800 6749 29840
rect 6691 29799 6749 29800
rect 7555 29840 7613 29841
rect 7555 29800 7564 29840
rect 7604 29800 7613 29840
rect 7555 29799 7613 29800
rect 8803 29840 8861 29841
rect 8803 29800 8812 29840
rect 8852 29800 8861 29840
rect 8803 29799 8861 29800
rect 11395 29840 11453 29841
rect 11395 29800 11404 29840
rect 11444 29800 11453 29840
rect 11395 29799 11453 29800
rect 11587 29840 11645 29841
rect 11587 29800 11596 29840
rect 11636 29800 11645 29840
rect 11587 29799 11645 29800
rect 13411 29840 13469 29841
rect 13411 29800 13420 29840
rect 13460 29800 13469 29840
rect 13411 29799 13469 29800
rect 13707 29840 13749 29849
rect 13707 29800 13708 29840
rect 13748 29800 13749 29840
rect 13707 29791 13749 29800
rect 13803 29840 13845 29849
rect 13803 29800 13804 29840
rect 13844 29800 13845 29840
rect 13803 29791 13845 29800
rect 14371 29840 14429 29841
rect 14371 29800 14380 29840
rect 14420 29800 14429 29840
rect 14371 29799 14429 29800
rect 15619 29840 15677 29841
rect 15619 29800 15628 29840
rect 15668 29800 15677 29840
rect 15619 29799 15677 29800
rect 16003 29840 16061 29841
rect 16003 29800 16012 29840
rect 16052 29800 16061 29840
rect 16003 29799 16061 29800
rect 17251 29840 17309 29841
rect 17251 29800 17260 29840
rect 17300 29800 17309 29840
rect 17251 29799 17309 29800
rect 17739 29840 17781 29849
rect 17739 29800 17740 29840
rect 17780 29800 17781 29840
rect 17739 29791 17781 29800
rect 17835 29840 17877 29849
rect 17835 29800 17836 29840
rect 17876 29800 17877 29840
rect 17835 29791 17877 29800
rect 18219 29840 18261 29849
rect 18219 29800 18220 29840
rect 18260 29800 18261 29840
rect 18219 29791 18261 29800
rect 18315 29840 18357 29849
rect 19275 29845 19317 29854
rect 18315 29800 18316 29840
rect 18356 29800 18357 29840
rect 18315 29791 18357 29800
rect 18787 29840 18845 29841
rect 18787 29800 18796 29840
rect 18836 29800 18845 29840
rect 18787 29799 18845 29800
rect 19275 29805 19276 29845
rect 19316 29805 19317 29845
rect 19275 29796 19317 29805
rect 13035 29756 13077 29765
rect 13035 29716 13036 29756
rect 13076 29716 13077 29756
rect 13035 29707 13077 29716
rect 19467 29756 19509 29765
rect 19467 29716 19468 29756
rect 19508 29716 19509 29756
rect 19467 29707 19509 29716
rect 4107 29672 4149 29681
rect 4107 29632 4108 29672
rect 4148 29632 4149 29672
rect 4107 29623 4149 29632
rect 6211 29672 6269 29673
rect 6211 29632 6220 29672
rect 6260 29632 6269 29672
rect 6211 29631 6269 29632
rect 6795 29672 6837 29681
rect 6795 29632 6796 29672
rect 6836 29632 6837 29672
rect 6795 29623 6837 29632
rect 11307 29672 11349 29681
rect 11307 29632 11308 29672
rect 11348 29632 11349 29672
rect 11307 29623 11349 29632
rect 15819 29672 15861 29681
rect 15819 29632 15820 29672
rect 15860 29632 15861 29672
rect 15819 29623 15861 29632
rect 1152 29504 20452 29528
rect 1152 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20452 29504
rect 1152 29440 20452 29464
rect 3147 29336 3189 29345
rect 3147 29296 3148 29336
rect 3188 29296 3189 29336
rect 3147 29287 3189 29296
rect 4299 29336 4341 29345
rect 4299 29296 4300 29336
rect 4340 29296 4341 29336
rect 4299 29287 4341 29296
rect 9003 29336 9045 29345
rect 9003 29296 9004 29336
rect 9044 29296 9045 29336
rect 9003 29287 9045 29296
rect 12747 29336 12789 29345
rect 12747 29296 12748 29336
rect 12788 29296 12789 29336
rect 12747 29287 12789 29296
rect 17451 29336 17493 29345
rect 17451 29296 17452 29336
rect 17492 29296 17493 29336
rect 17451 29287 17493 29296
rect 19659 29336 19701 29345
rect 19659 29296 19660 29336
rect 19700 29296 19701 29336
rect 19659 29287 19701 29296
rect 6603 29252 6645 29261
rect 6603 29212 6604 29252
rect 6644 29212 6645 29252
rect 6603 29203 6645 29212
rect 11019 29252 11061 29261
rect 11019 29212 11020 29252
rect 11060 29212 11061 29252
rect 11019 29203 11061 29212
rect 14283 29189 14325 29198
rect 12939 29179 12981 29188
rect 1699 29168 1757 29169
rect 1699 29128 1708 29168
rect 1748 29128 1757 29168
rect 1699 29127 1757 29128
rect 2947 29168 3005 29169
rect 2947 29128 2956 29168
rect 2996 29128 3005 29168
rect 2947 29127 3005 29128
rect 4483 29168 4541 29169
rect 4483 29128 4492 29168
rect 4532 29128 4541 29168
rect 4483 29127 4541 29128
rect 5731 29168 5789 29169
rect 5731 29128 5740 29168
rect 5780 29128 5789 29168
rect 5731 29127 5789 29128
rect 6027 29168 6069 29177
rect 6027 29128 6028 29168
rect 6068 29128 6069 29168
rect 6027 29119 6069 29128
rect 6115 29168 6173 29169
rect 6115 29128 6124 29168
rect 6164 29128 6173 29168
rect 6115 29127 6173 29128
rect 6699 29168 6741 29177
rect 6699 29128 6700 29168
rect 6740 29128 6741 29168
rect 7267 29168 7325 29169
rect 6699 29119 6741 29128
rect 6979 29151 7037 29152
rect 6979 29111 6988 29151
rect 7028 29111 7037 29151
rect 7267 29128 7276 29168
rect 7316 29128 7325 29168
rect 7267 29127 7325 29128
rect 7555 29168 7613 29169
rect 7555 29128 7564 29168
rect 7604 29128 7613 29168
rect 7555 29127 7613 29128
rect 8803 29168 8861 29169
rect 8803 29128 8812 29168
rect 8852 29128 8861 29168
rect 8803 29127 8861 29128
rect 9291 29168 9333 29177
rect 9291 29128 9292 29168
rect 9332 29128 9333 29168
rect 9291 29119 9333 29128
rect 9387 29168 9429 29177
rect 9387 29128 9388 29168
rect 9428 29128 9429 29168
rect 9387 29119 9429 29128
rect 9867 29168 9909 29177
rect 9867 29128 9868 29168
rect 9908 29128 9909 29168
rect 9867 29119 9909 29128
rect 10339 29168 10397 29169
rect 10339 29128 10348 29168
rect 10388 29128 10397 29168
rect 11299 29168 11357 29169
rect 10339 29127 10397 29128
rect 10827 29154 10869 29163
rect 6979 29110 7037 29111
rect 10827 29114 10828 29154
rect 10868 29114 10869 29154
rect 11299 29128 11308 29168
rect 11348 29128 11357 29168
rect 11299 29127 11357 29128
rect 12547 29168 12605 29169
rect 12547 29128 12556 29168
rect 12596 29128 12605 29168
rect 12939 29139 12940 29179
rect 12980 29139 12981 29179
rect 12939 29130 12981 29139
rect 13131 29168 13173 29177
rect 12547 29127 12605 29128
rect 13131 29128 13132 29168
rect 13172 29128 13173 29168
rect 13131 29119 13173 29128
rect 13411 29168 13469 29169
rect 13411 29128 13420 29168
rect 13460 29128 13469 29168
rect 13411 29127 13469 29128
rect 13707 29168 13749 29177
rect 13707 29128 13708 29168
rect 13748 29128 13749 29168
rect 13707 29119 13749 29128
rect 13803 29168 13845 29177
rect 13803 29128 13804 29168
rect 13844 29128 13845 29168
rect 14283 29149 14284 29189
rect 14324 29149 14325 29189
rect 14475 29189 14517 29198
rect 14283 29140 14325 29149
rect 14379 29168 14421 29177
rect 13803 29119 13845 29128
rect 14379 29128 14380 29168
rect 14420 29128 14421 29168
rect 14475 29149 14476 29189
rect 14516 29149 14517 29189
rect 14475 29140 14517 29149
rect 14571 29168 14613 29177
rect 14379 29119 14421 29128
rect 14571 29128 14572 29168
rect 14612 29128 14613 29168
rect 14571 29119 14613 29128
rect 14763 29168 14805 29177
rect 14763 29128 14764 29168
rect 14804 29128 14805 29168
rect 14763 29119 14805 29128
rect 14859 29168 14901 29177
rect 14859 29128 14860 29168
rect 14900 29128 14901 29168
rect 14859 29119 14901 29128
rect 14955 29168 14997 29177
rect 14955 29128 14956 29168
rect 14996 29128 14997 29168
rect 14955 29119 14997 29128
rect 15051 29168 15093 29177
rect 15051 29128 15052 29168
rect 15092 29128 15093 29168
rect 15051 29119 15093 29128
rect 15243 29168 15285 29177
rect 15243 29128 15244 29168
rect 15284 29128 15285 29168
rect 15243 29119 15285 29128
rect 15435 29168 15477 29177
rect 15435 29128 15436 29168
rect 15476 29128 15477 29168
rect 15435 29119 15477 29128
rect 15523 29168 15581 29169
rect 15523 29128 15532 29168
rect 15572 29128 15581 29168
rect 15523 29127 15581 29128
rect 16003 29168 16061 29169
rect 16003 29128 16012 29168
rect 16052 29128 16061 29168
rect 16003 29127 16061 29128
rect 17251 29168 17309 29169
rect 17251 29128 17260 29168
rect 17300 29128 17309 29168
rect 17251 29127 17309 29128
rect 17931 29168 17973 29177
rect 17931 29128 17932 29168
rect 17972 29128 17973 29168
rect 17931 29119 17973 29128
rect 18027 29168 18069 29177
rect 18027 29128 18028 29168
rect 18068 29128 18069 29168
rect 18027 29119 18069 29128
rect 18507 29168 18549 29177
rect 18507 29128 18508 29168
rect 18548 29128 18549 29168
rect 18507 29119 18549 29128
rect 18979 29168 19037 29169
rect 18979 29128 18988 29168
rect 19028 29128 19037 29168
rect 18979 29127 19037 29128
rect 19515 29158 19557 29167
rect 10827 29105 10869 29114
rect 19515 29118 19516 29158
rect 19556 29118 19557 29158
rect 19515 29109 19557 29118
rect 9771 29084 9813 29093
rect 9771 29044 9772 29084
rect 9812 29044 9813 29084
rect 9771 29035 9813 29044
rect 18411 29084 18453 29093
rect 18411 29044 18412 29084
rect 18452 29044 18453 29084
rect 18411 29035 18453 29044
rect 14083 29000 14141 29001
rect 14083 28960 14092 29000
rect 14132 28960 14141 29000
rect 14083 28959 14141 28960
rect 6307 28916 6365 28917
rect 6307 28876 6316 28916
rect 6356 28876 6365 28916
rect 6307 28875 6365 28876
rect 7371 28916 7413 28925
rect 7371 28876 7372 28916
rect 7412 28876 7413 28916
rect 7371 28867 7413 28876
rect 12939 28916 12981 28925
rect 12939 28876 12940 28916
rect 12980 28876 12981 28916
rect 12939 28867 12981 28876
rect 15243 28916 15285 28925
rect 15243 28876 15244 28916
rect 15284 28876 15285 28916
rect 15243 28867 15285 28876
rect 1152 28748 20352 28772
rect 1152 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 20352 28748
rect 1152 28684 20352 28708
rect 7075 28580 7133 28581
rect 7075 28540 7084 28580
rect 7124 28540 7133 28580
rect 7075 28539 7133 28540
rect 10827 28580 10869 28589
rect 10827 28540 10828 28580
rect 10868 28540 10869 28580
rect 10827 28531 10869 28540
rect 12363 28580 12405 28589
rect 12363 28540 12364 28580
rect 12404 28540 12405 28580
rect 12363 28531 12405 28540
rect 18219 28580 18261 28589
rect 18219 28540 18220 28580
rect 18260 28540 18261 28580
rect 18219 28531 18261 28540
rect 16443 28337 16485 28346
rect 2659 28328 2717 28329
rect 2659 28288 2668 28328
rect 2708 28288 2717 28328
rect 2659 28287 2717 28288
rect 3907 28328 3965 28329
rect 3907 28288 3916 28328
rect 3956 28288 3965 28328
rect 3907 28287 3965 28288
rect 4291 28328 4349 28329
rect 4291 28288 4300 28328
rect 4340 28288 4349 28328
rect 4291 28287 4349 28288
rect 5539 28328 5597 28329
rect 5539 28288 5548 28328
rect 5588 28288 5597 28328
rect 5539 28287 5597 28288
rect 6403 28328 6461 28329
rect 6403 28288 6412 28328
rect 6452 28288 6461 28328
rect 6403 28287 6461 28288
rect 6699 28328 6741 28337
rect 6699 28288 6700 28328
rect 6740 28288 6741 28328
rect 6699 28279 6741 28288
rect 7275 28328 7317 28337
rect 7275 28288 7276 28328
rect 7316 28288 7317 28328
rect 7275 28279 7317 28288
rect 7467 28328 7509 28337
rect 7467 28288 7468 28328
rect 7508 28288 7509 28328
rect 7467 28279 7509 28288
rect 7555 28328 7613 28329
rect 7555 28288 7564 28328
rect 7604 28288 7613 28328
rect 7555 28287 7613 28288
rect 7755 28328 7797 28337
rect 7755 28288 7756 28328
rect 7796 28288 7797 28328
rect 7755 28279 7797 28288
rect 7851 28328 7893 28337
rect 7851 28288 7852 28328
rect 7892 28288 7893 28328
rect 7851 28279 7893 28288
rect 7947 28328 7989 28337
rect 7947 28288 7948 28328
rect 7988 28288 7989 28328
rect 7947 28279 7989 28288
rect 9379 28328 9437 28329
rect 9379 28288 9388 28328
rect 9428 28288 9437 28328
rect 9379 28287 9437 28288
rect 10627 28328 10685 28329
rect 10627 28288 10636 28328
rect 10676 28288 10685 28328
rect 10627 28287 10685 28288
rect 12451 28328 12509 28329
rect 12451 28288 12460 28328
rect 12500 28288 12509 28328
rect 12451 28287 12509 28288
rect 12747 28328 12789 28337
rect 12747 28288 12748 28328
rect 12788 28288 12789 28328
rect 12747 28279 12789 28288
rect 12843 28328 12885 28337
rect 12843 28288 12844 28328
rect 12884 28288 12885 28328
rect 12843 28279 12885 28288
rect 12939 28328 12981 28337
rect 12939 28288 12940 28328
rect 12980 28288 12981 28328
rect 12939 28279 12981 28288
rect 13123 28328 13181 28329
rect 13123 28288 13132 28328
rect 13172 28288 13181 28328
rect 13123 28287 13181 28288
rect 14371 28328 14429 28329
rect 14371 28288 14380 28328
rect 14420 28288 14429 28328
rect 14371 28287 14429 28288
rect 14859 28328 14901 28337
rect 14859 28288 14860 28328
rect 14900 28288 14901 28328
rect 14859 28279 14901 28288
rect 14955 28328 14997 28337
rect 14955 28288 14956 28328
rect 14996 28288 14997 28328
rect 14955 28279 14997 28288
rect 15339 28328 15381 28337
rect 15339 28288 15340 28328
rect 15380 28288 15381 28328
rect 15339 28279 15381 28288
rect 15435 28328 15477 28337
rect 15435 28288 15436 28328
rect 15476 28288 15477 28328
rect 15435 28279 15477 28288
rect 15907 28328 15965 28329
rect 15907 28288 15916 28328
rect 15956 28288 15965 28328
rect 16443 28297 16444 28337
rect 16484 28297 16485 28337
rect 16443 28288 16485 28297
rect 16771 28328 16829 28329
rect 16771 28288 16780 28328
rect 16820 28288 16829 28328
rect 15907 28287 15965 28288
rect 16771 28287 16829 28288
rect 18019 28328 18077 28329
rect 18019 28288 18028 28328
rect 18068 28288 18077 28328
rect 18019 28287 18077 28288
rect 18507 28328 18549 28337
rect 18507 28288 18508 28328
rect 18548 28288 18549 28328
rect 18507 28279 18549 28288
rect 18603 28328 18645 28337
rect 18603 28288 18604 28328
rect 18644 28288 18645 28328
rect 18603 28279 18645 28288
rect 18987 28328 19029 28337
rect 18987 28288 18988 28328
rect 19028 28288 19029 28328
rect 18987 28279 19029 28288
rect 19083 28328 19125 28337
rect 20043 28333 20085 28342
rect 19083 28288 19084 28328
rect 19124 28288 19125 28328
rect 19083 28279 19125 28288
rect 19555 28328 19613 28329
rect 19555 28288 19564 28328
rect 19604 28288 19613 28328
rect 19555 28287 19613 28288
rect 20043 28293 20044 28333
rect 20084 28293 20085 28333
rect 20043 28284 20085 28293
rect 4107 28244 4149 28253
rect 4107 28204 4108 28244
rect 4148 28204 4149 28244
rect 4107 28195 4149 28204
rect 6795 28244 6837 28253
rect 6795 28204 6796 28244
rect 6836 28204 6837 28244
rect 6795 28195 6837 28204
rect 14571 28244 14613 28253
rect 14571 28204 14572 28244
rect 14612 28204 14613 28244
rect 14571 28195 14613 28204
rect 20235 28244 20277 28253
rect 20235 28204 20236 28244
rect 20276 28204 20277 28244
rect 20235 28195 20277 28204
rect 5739 28160 5781 28169
rect 5739 28120 5740 28160
rect 5780 28120 5781 28160
rect 5739 28111 5781 28120
rect 7363 28160 7421 28161
rect 7363 28120 7372 28160
rect 7412 28120 7421 28160
rect 7363 28119 7421 28120
rect 8035 28160 8093 28161
rect 8035 28120 8044 28160
rect 8084 28120 8093 28160
rect 8035 28119 8093 28120
rect 12643 28160 12701 28161
rect 12643 28120 12652 28160
rect 12692 28120 12701 28160
rect 12643 28119 12701 28120
rect 16587 28160 16629 28169
rect 16587 28120 16588 28160
rect 16628 28120 16629 28160
rect 16587 28111 16629 28120
rect 1152 27992 20452 28016
rect 1152 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20452 27992
rect 1152 27928 20452 27952
rect 11971 27824 12029 27825
rect 11971 27784 11980 27824
rect 12020 27784 12029 27824
rect 11971 27783 12029 27784
rect 12835 27824 12893 27825
rect 12835 27784 12844 27824
rect 12884 27784 12893 27824
rect 12835 27783 12893 27784
rect 14467 27824 14525 27825
rect 14467 27784 14476 27824
rect 14516 27784 14525 27824
rect 14467 27783 14525 27784
rect 16587 27824 16629 27833
rect 16587 27784 16588 27824
rect 16628 27784 16629 27824
rect 16587 27775 16629 27784
rect 18219 27824 18261 27833
rect 18219 27784 18220 27824
rect 18260 27784 18261 27824
rect 18219 27775 18261 27784
rect 4587 27740 4629 27749
rect 4587 27700 4588 27740
rect 4628 27700 4629 27740
rect 4587 27691 4629 27700
rect 8907 27740 8949 27749
rect 8907 27700 8908 27740
rect 8948 27700 8949 27740
rect 8907 27691 8949 27700
rect 10923 27740 10965 27749
rect 10923 27700 10924 27740
rect 10964 27700 10965 27740
rect 10923 27691 10965 27700
rect 20235 27740 20277 27749
rect 20235 27700 20236 27740
rect 20276 27700 20277 27740
rect 18787 27698 18845 27699
rect 2859 27656 2901 27665
rect 2859 27616 2860 27656
rect 2900 27616 2901 27656
rect 2859 27607 2901 27616
rect 2955 27656 2997 27665
rect 2955 27616 2956 27656
rect 2996 27616 2997 27656
rect 2955 27607 2997 27616
rect 3435 27656 3477 27665
rect 3435 27616 3436 27656
rect 3476 27616 3477 27656
rect 3435 27607 3477 27616
rect 3907 27656 3965 27657
rect 3907 27616 3916 27656
rect 3956 27616 3965 27656
rect 4867 27656 4925 27657
rect 3907 27615 3965 27616
rect 4395 27642 4437 27651
rect 4395 27602 4396 27642
rect 4436 27602 4437 27642
rect 4867 27616 4876 27656
rect 4916 27616 4925 27656
rect 4867 27615 4925 27616
rect 6115 27656 6173 27657
rect 6115 27616 6124 27656
rect 6164 27616 6173 27656
rect 6115 27615 6173 27616
rect 6507 27656 6549 27665
rect 6507 27616 6508 27656
rect 6548 27616 6549 27656
rect 6507 27607 6549 27616
rect 6699 27656 6741 27665
rect 6699 27616 6700 27656
rect 6740 27616 6741 27656
rect 6699 27607 6741 27616
rect 6883 27656 6941 27657
rect 6883 27616 6892 27656
rect 6932 27616 6941 27656
rect 6883 27615 6941 27616
rect 6987 27656 7029 27665
rect 6987 27616 6988 27656
rect 7028 27616 7029 27656
rect 6987 27607 7029 27616
rect 7179 27656 7221 27665
rect 7179 27616 7180 27656
rect 7220 27616 7221 27656
rect 7179 27607 7221 27616
rect 7459 27656 7517 27657
rect 7459 27616 7468 27656
rect 7508 27616 7517 27656
rect 7459 27615 7517 27616
rect 8707 27656 8765 27657
rect 8707 27616 8716 27656
rect 8756 27616 8765 27656
rect 8707 27615 8765 27616
rect 9195 27656 9237 27665
rect 9195 27616 9196 27656
rect 9236 27616 9237 27656
rect 9195 27607 9237 27616
rect 9291 27656 9333 27665
rect 9291 27616 9292 27656
rect 9332 27616 9333 27656
rect 9291 27607 9333 27616
rect 9771 27656 9813 27665
rect 9771 27616 9772 27656
rect 9812 27616 9813 27656
rect 9771 27607 9813 27616
rect 10243 27656 10301 27657
rect 10243 27616 10252 27656
rect 10292 27616 10301 27656
rect 11491 27656 11549 27657
rect 10243 27615 10301 27616
rect 10731 27642 10773 27651
rect 4395 27593 4437 27602
rect 10731 27602 10732 27642
rect 10772 27602 10773 27642
rect 11491 27616 11500 27656
rect 11540 27616 11549 27656
rect 11491 27615 11549 27616
rect 11595 27656 11637 27665
rect 11595 27616 11596 27656
rect 11636 27616 11637 27656
rect 11979 27656 12021 27665
rect 11595 27607 11637 27616
rect 11821 27641 11863 27650
rect 10731 27593 10773 27602
rect 11821 27601 11822 27641
rect 11862 27601 11863 27641
rect 11979 27616 11980 27656
rect 12020 27616 12021 27656
rect 11979 27607 12021 27616
rect 12075 27656 12117 27665
rect 12075 27616 12076 27656
rect 12116 27616 12117 27656
rect 12075 27607 12117 27616
rect 12259 27656 12317 27657
rect 12259 27616 12268 27656
rect 12308 27616 12317 27656
rect 12259 27615 12317 27616
rect 12355 27656 12413 27657
rect 12355 27616 12364 27656
rect 12404 27616 12413 27656
rect 12355 27615 12413 27616
rect 12555 27656 12597 27665
rect 12555 27616 12556 27656
rect 12596 27616 12597 27656
rect 12555 27607 12597 27616
rect 12651 27656 12693 27665
rect 12651 27616 12652 27656
rect 12692 27616 12693 27656
rect 12651 27607 12693 27616
rect 13219 27656 13277 27657
rect 13219 27616 13228 27656
rect 13268 27616 13277 27656
rect 13219 27615 13277 27616
rect 13323 27656 13365 27665
rect 13323 27616 13324 27656
rect 13364 27616 13365 27656
rect 13323 27607 13365 27616
rect 13515 27656 13557 27665
rect 13515 27616 13516 27656
rect 13556 27616 13557 27656
rect 13515 27607 13557 27616
rect 13707 27656 13749 27665
rect 13707 27616 13708 27656
rect 13748 27616 13749 27656
rect 13707 27607 13749 27616
rect 13899 27656 13941 27665
rect 13899 27616 13900 27656
rect 13940 27616 13941 27656
rect 13899 27607 13941 27616
rect 13987 27656 14045 27657
rect 13987 27616 13996 27656
rect 14036 27616 14045 27656
rect 13987 27615 14045 27616
rect 14462 27656 14520 27657
rect 14462 27616 14471 27656
rect 14511 27616 14520 27656
rect 14462 27615 14520 27616
rect 14571 27656 14613 27665
rect 14571 27616 14572 27656
rect 14612 27616 14613 27656
rect 14571 27607 14613 27616
rect 14667 27656 14709 27665
rect 18787 27658 18796 27698
rect 18836 27658 18845 27698
rect 20235 27691 20277 27700
rect 18787 27657 18845 27658
rect 14667 27616 14668 27656
rect 14708 27616 14709 27656
rect 14667 27607 14709 27616
rect 14851 27656 14909 27657
rect 14851 27616 14860 27656
rect 14900 27616 14909 27656
rect 14851 27615 14909 27616
rect 14947 27656 15005 27657
rect 14947 27616 14956 27656
rect 14996 27616 15005 27656
rect 14947 27615 15005 27616
rect 15139 27656 15197 27657
rect 15139 27616 15148 27656
rect 15188 27616 15197 27656
rect 15139 27615 15197 27616
rect 16387 27656 16445 27657
rect 16387 27616 16396 27656
rect 16436 27616 16445 27656
rect 16387 27615 16445 27616
rect 16771 27656 16829 27657
rect 16771 27616 16780 27656
rect 16820 27616 16829 27656
rect 16771 27615 16829 27616
rect 18019 27656 18077 27657
rect 18019 27616 18028 27656
rect 18068 27616 18077 27656
rect 18019 27615 18077 27616
rect 20035 27656 20093 27657
rect 20035 27616 20044 27656
rect 20084 27616 20093 27656
rect 20035 27615 20093 27616
rect 11821 27592 11863 27601
rect 3339 27572 3381 27581
rect 3339 27532 3340 27572
rect 3380 27532 3381 27572
rect 3339 27523 3381 27532
rect 9675 27572 9717 27581
rect 9675 27532 9676 27572
rect 9716 27532 9717 27572
rect 9675 27523 9717 27532
rect 13707 27488 13749 27497
rect 13707 27448 13708 27488
rect 13748 27448 13749 27488
rect 13707 27439 13749 27448
rect 6315 27404 6357 27413
rect 6315 27364 6316 27404
rect 6356 27364 6357 27404
rect 6315 27355 6357 27364
rect 6507 27404 6549 27413
rect 6507 27364 6508 27404
rect 6548 27364 6549 27404
rect 6507 27355 6549 27364
rect 7179 27404 7221 27413
rect 7179 27364 7180 27404
rect 7220 27364 7221 27404
rect 7179 27355 7221 27364
rect 12363 27404 12405 27413
rect 12363 27364 12364 27404
rect 12404 27364 12405 27404
rect 12363 27355 12405 27364
rect 13515 27404 13557 27413
rect 13515 27364 13516 27404
rect 13556 27364 13557 27404
rect 13515 27355 13557 27364
rect 14955 27404 14997 27413
rect 14955 27364 14956 27404
rect 14996 27364 14997 27404
rect 14955 27355 14997 27364
rect 1152 27236 20352 27260
rect 1152 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 20352 27236
rect 1152 27172 20352 27196
rect 6219 27068 6261 27077
rect 6219 27028 6220 27068
rect 6260 27028 6261 27068
rect 6219 27019 6261 27028
rect 10443 27068 10485 27077
rect 10443 27028 10444 27068
rect 10484 27028 10485 27068
rect 10443 27019 10485 27028
rect 14763 27068 14805 27077
rect 14763 27028 14764 27068
rect 14804 27028 14805 27068
rect 14763 27019 14805 27028
rect 4299 26984 4341 26993
rect 4299 26944 4300 26984
rect 4340 26944 4341 26984
rect 4299 26935 4341 26944
rect 7467 26984 7509 26993
rect 7467 26944 7468 26984
rect 7508 26944 7509 26984
rect 7467 26935 7509 26944
rect 12459 26984 12501 26993
rect 12459 26944 12460 26984
rect 12500 26944 12501 26984
rect 12459 26935 12501 26944
rect 15043 26984 15101 26985
rect 15043 26944 15052 26984
rect 15092 26944 15101 26984
rect 15043 26943 15101 26944
rect 16971 26984 17013 26993
rect 16971 26944 16972 26984
rect 17012 26944 17013 26984
rect 16971 26935 17013 26944
rect 2955 26900 2997 26909
rect 2955 26860 2956 26900
rect 2996 26860 2997 26900
rect 17739 26900 17781 26909
rect 2955 26851 2997 26860
rect 3963 26858 4005 26867
rect 2379 26816 2421 26825
rect 2379 26776 2380 26816
rect 2420 26776 2421 26816
rect 2379 26767 2421 26776
rect 2475 26816 2517 26825
rect 2475 26776 2476 26816
rect 2516 26776 2517 26816
rect 2475 26767 2517 26776
rect 2859 26816 2901 26825
rect 3963 26818 3964 26858
rect 4004 26818 4005 26858
rect 17739 26860 17740 26900
rect 17780 26860 17781 26900
rect 17739 26851 17781 26860
rect 2859 26776 2860 26816
rect 2900 26776 2901 26816
rect 2859 26767 2901 26776
rect 3427 26816 3485 26817
rect 3427 26776 3436 26816
rect 3476 26776 3485 26816
rect 3963 26809 4005 26818
rect 4483 26816 4541 26817
rect 3427 26775 3485 26776
rect 4483 26776 4492 26816
rect 4532 26776 4541 26816
rect 4483 26775 4541 26776
rect 5731 26816 5789 26817
rect 5731 26776 5740 26816
rect 5780 26776 5789 26816
rect 5731 26775 5789 26776
rect 5923 26816 5981 26817
rect 5923 26776 5932 26816
rect 5972 26776 5981 26816
rect 5923 26775 5981 26776
rect 6027 26816 6069 26825
rect 6027 26776 6028 26816
rect 6068 26776 6069 26816
rect 6027 26767 6069 26776
rect 6219 26816 6261 26825
rect 6219 26776 6220 26816
rect 6260 26776 6261 26816
rect 6219 26767 6261 26776
rect 6507 26816 6549 26825
rect 6507 26776 6508 26816
rect 6548 26776 6549 26816
rect 6507 26767 6549 26776
rect 6603 26816 6645 26825
rect 6603 26776 6604 26816
rect 6644 26776 6645 26816
rect 6603 26767 6645 26776
rect 6699 26816 6741 26825
rect 6699 26776 6700 26816
rect 6740 26776 6741 26816
rect 6699 26767 6741 26776
rect 6795 26816 6837 26825
rect 6795 26776 6796 26816
rect 6836 26776 6837 26816
rect 6795 26767 6837 26776
rect 6979 26816 7037 26817
rect 6979 26776 6988 26816
rect 7028 26776 7037 26816
rect 6979 26775 7037 26776
rect 7083 26816 7125 26825
rect 7083 26776 7084 26816
rect 7124 26776 7125 26816
rect 7083 26767 7125 26776
rect 7275 26816 7317 26825
rect 7275 26776 7276 26816
rect 7316 26776 7317 26816
rect 7275 26767 7317 26776
rect 7467 26816 7509 26825
rect 7467 26776 7468 26816
rect 7508 26776 7509 26816
rect 7467 26767 7509 26776
rect 7755 26816 7797 26825
rect 7755 26776 7756 26816
rect 7796 26776 7797 26816
rect 7755 26767 7797 26776
rect 8523 26816 8565 26825
rect 8523 26776 8524 26816
rect 8564 26776 8565 26816
rect 8523 26767 8565 26776
rect 8715 26816 8757 26825
rect 8715 26776 8716 26816
rect 8756 26776 8757 26816
rect 8715 26767 8757 26776
rect 8803 26816 8861 26817
rect 8803 26776 8812 26816
rect 8852 26776 8861 26816
rect 8803 26775 8861 26776
rect 8995 26816 9053 26817
rect 8995 26776 9004 26816
rect 9044 26776 9053 26816
rect 8995 26775 9053 26776
rect 10243 26816 10301 26817
rect 10243 26776 10252 26816
rect 10292 26776 10301 26816
rect 10243 26775 10301 26776
rect 10627 26816 10685 26817
rect 10627 26776 10636 26816
rect 10676 26776 10685 26816
rect 10627 26775 10685 26776
rect 11875 26816 11933 26817
rect 11875 26776 11884 26816
rect 11924 26776 11933 26816
rect 11875 26775 11933 26776
rect 12267 26816 12309 26825
rect 12267 26776 12268 26816
rect 12308 26776 12309 26816
rect 12267 26767 12309 26776
rect 12363 26816 12405 26825
rect 12363 26776 12364 26816
rect 12404 26776 12405 26816
rect 12363 26767 12405 26776
rect 12555 26816 12597 26825
rect 12555 26776 12556 26816
rect 12596 26776 12597 26816
rect 12555 26767 12597 26776
rect 13315 26816 13373 26817
rect 13315 26776 13324 26816
rect 13364 26776 13373 26816
rect 13315 26775 13373 26776
rect 14563 26816 14621 26817
rect 14563 26776 14572 26816
rect 14612 26776 14621 26816
rect 14563 26775 14621 26776
rect 14955 26816 14997 26825
rect 14955 26776 14956 26816
rect 14996 26776 14997 26816
rect 14955 26767 14997 26776
rect 15051 26816 15093 26825
rect 15051 26776 15052 26816
rect 15092 26776 15093 26816
rect 15051 26767 15093 26776
rect 15243 26816 15285 26825
rect 15243 26776 15244 26816
rect 15284 26776 15285 26816
rect 15243 26767 15285 26776
rect 15523 26816 15581 26817
rect 15523 26776 15532 26816
rect 15572 26776 15581 26816
rect 15523 26775 15581 26776
rect 16771 26816 16829 26817
rect 16771 26776 16780 26816
rect 16820 26776 16829 26816
rect 16771 26775 16829 26776
rect 17259 26816 17301 26825
rect 17259 26776 17260 26816
rect 17300 26776 17301 26816
rect 17259 26767 17301 26776
rect 17355 26816 17397 26825
rect 17355 26776 17356 26816
rect 17396 26776 17397 26816
rect 17355 26767 17397 26776
rect 17835 26816 17877 26825
rect 18795 26821 18837 26830
rect 17835 26776 17836 26816
rect 17876 26776 17877 26816
rect 17835 26767 17877 26776
rect 18307 26816 18365 26817
rect 18307 26776 18316 26816
rect 18356 26776 18365 26816
rect 18307 26775 18365 26776
rect 18795 26781 18796 26821
rect 18836 26781 18837 26821
rect 18795 26772 18837 26781
rect 18987 26732 19029 26741
rect 18987 26692 18988 26732
rect 19028 26692 19029 26732
rect 18987 26683 19029 26692
rect 4107 26648 4149 26657
rect 4107 26608 4108 26648
rect 4148 26608 4149 26648
rect 4107 26599 4149 26608
rect 7171 26648 7229 26649
rect 7171 26608 7180 26648
rect 7220 26608 7229 26648
rect 7171 26607 7229 26608
rect 8611 26648 8669 26649
rect 8611 26608 8620 26648
rect 8660 26608 8669 26648
rect 8611 26607 8669 26608
rect 12075 26648 12117 26657
rect 12075 26608 12076 26648
rect 12116 26608 12117 26648
rect 12075 26599 12117 26608
rect 1152 26480 20452 26504
rect 1152 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20452 26480
rect 1152 26416 20452 26440
rect 2667 26312 2709 26321
rect 2667 26272 2668 26312
rect 2708 26272 2709 26312
rect 2667 26263 2709 26272
rect 4491 26312 4533 26321
rect 4491 26272 4492 26312
rect 4532 26272 4533 26312
rect 4491 26263 4533 26272
rect 7563 26312 7605 26321
rect 7563 26272 7564 26312
rect 7604 26272 7605 26312
rect 7563 26263 7605 26272
rect 9963 26312 10005 26321
rect 9963 26272 9964 26312
rect 10004 26272 10005 26312
rect 9963 26263 10005 26272
rect 12075 26312 12117 26321
rect 12075 26272 12076 26312
rect 12116 26272 12117 26312
rect 12075 26263 12117 26272
rect 15051 26312 15093 26321
rect 15051 26272 15052 26312
rect 15092 26272 15093 26312
rect 15051 26263 15093 26272
rect 15523 26312 15581 26313
rect 15523 26272 15532 26312
rect 15572 26272 15581 26312
rect 15523 26271 15581 26272
rect 15723 26312 15765 26321
rect 15723 26272 15724 26312
rect 15764 26272 15765 26312
rect 15723 26263 15765 26272
rect 17931 26312 17973 26321
rect 17931 26272 17932 26312
rect 17972 26272 17973 26312
rect 17931 26263 17973 26272
rect 19947 26312 19989 26321
rect 19947 26272 19948 26312
rect 19988 26272 19989 26312
rect 19947 26263 19989 26272
rect 6123 26228 6165 26237
rect 6123 26188 6124 26228
rect 6164 26188 6165 26228
rect 6123 26179 6165 26188
rect 9291 26228 9333 26237
rect 9291 26188 9292 26228
rect 9332 26188 9333 26228
rect 9291 26179 9333 26188
rect 10443 26228 10485 26237
rect 10443 26188 10444 26228
rect 10484 26188 10485 26228
rect 10443 26179 10485 26188
rect 16107 26228 16149 26237
rect 16107 26188 16108 26228
rect 16148 26188 16149 26228
rect 16107 26179 16149 26188
rect 1219 26144 1277 26145
rect 1219 26104 1228 26144
rect 1268 26104 1277 26144
rect 1219 26103 1277 26104
rect 2467 26144 2525 26145
rect 2467 26104 2476 26144
rect 2516 26104 2525 26144
rect 2467 26103 2525 26104
rect 3043 26144 3101 26145
rect 3043 26104 3052 26144
rect 3092 26104 3101 26144
rect 3043 26103 3101 26104
rect 4291 26144 4349 26145
rect 4291 26104 4300 26144
rect 4340 26104 4349 26144
rect 4291 26103 4349 26104
rect 4675 26144 4733 26145
rect 4675 26104 4684 26144
rect 4724 26104 4733 26144
rect 4675 26103 4733 26104
rect 5923 26144 5981 26145
rect 5923 26104 5932 26144
rect 5972 26104 5981 26144
rect 5923 26103 5981 26104
rect 6411 26144 6453 26153
rect 6411 26104 6412 26144
rect 6452 26104 6453 26144
rect 7371 26144 7413 26153
rect 6411 26095 6453 26104
rect 6603 26129 6645 26138
rect 6499 26102 6557 26103
rect 6499 26062 6508 26102
rect 6548 26062 6557 26102
rect 6603 26089 6604 26129
rect 6644 26089 6645 26129
rect 7371 26104 7372 26144
rect 7412 26104 7413 26144
rect 7371 26095 7413 26104
rect 7659 26144 7701 26153
rect 7659 26104 7660 26144
rect 7700 26104 7701 26144
rect 7659 26095 7701 26104
rect 7843 26144 7901 26145
rect 7843 26104 7852 26144
rect 7892 26104 7901 26144
rect 7843 26103 7901 26104
rect 9091 26144 9149 26145
rect 9091 26104 9100 26144
rect 9140 26104 9149 26144
rect 9091 26103 9149 26104
rect 9579 26144 9621 26153
rect 9579 26104 9580 26144
rect 9620 26104 9621 26144
rect 9579 26095 9621 26104
rect 9675 26144 9717 26153
rect 9675 26104 9676 26144
rect 9716 26104 9717 26144
rect 9675 26095 9717 26104
rect 9771 26144 9813 26153
rect 9771 26104 9772 26144
rect 9812 26104 9813 26144
rect 9771 26095 9813 26104
rect 10155 26144 10197 26153
rect 10155 26104 10156 26144
rect 10196 26104 10197 26144
rect 10155 26095 10197 26104
rect 10251 26144 10293 26153
rect 10251 26104 10252 26144
rect 10292 26104 10293 26144
rect 10251 26095 10293 26104
rect 10347 26144 10389 26153
rect 10347 26104 10348 26144
rect 10388 26104 10389 26144
rect 10347 26095 10389 26104
rect 10627 26144 10685 26145
rect 10627 26104 10636 26144
rect 10676 26104 10685 26144
rect 10627 26103 10685 26104
rect 11875 26144 11933 26145
rect 11875 26104 11884 26144
rect 11924 26104 11933 26144
rect 11875 26103 11933 26104
rect 13603 26144 13661 26145
rect 13603 26104 13612 26144
rect 13652 26104 13661 26144
rect 13603 26103 13661 26104
rect 14851 26144 14909 26145
rect 14851 26104 14860 26144
rect 14900 26104 14909 26144
rect 14851 26103 14909 26104
rect 15243 26144 15285 26153
rect 15243 26104 15244 26144
rect 15284 26104 15285 26144
rect 15811 26144 15869 26145
rect 15243 26095 15285 26104
rect 15336 26134 15394 26135
rect 15336 26094 15345 26134
rect 15385 26094 15394 26134
rect 15811 26104 15820 26144
rect 15860 26104 15869 26144
rect 15811 26103 15869 26104
rect 16011 26144 16053 26153
rect 16011 26104 16012 26144
rect 16052 26104 16053 26144
rect 16011 26095 16053 26104
rect 16203 26144 16245 26153
rect 16203 26104 16204 26144
rect 16244 26104 16245 26144
rect 16203 26095 16245 26104
rect 16291 26144 16349 26145
rect 16291 26104 16300 26144
rect 16340 26104 16349 26144
rect 16291 26103 16349 26104
rect 16483 26144 16541 26145
rect 16483 26104 16492 26144
rect 16532 26104 16541 26144
rect 16483 26103 16541 26104
rect 17731 26144 17789 26145
rect 17731 26104 17740 26144
rect 17780 26104 17789 26144
rect 17731 26103 17789 26104
rect 18219 26144 18261 26153
rect 18219 26104 18220 26144
rect 18260 26104 18261 26144
rect 18219 26095 18261 26104
rect 18315 26144 18357 26153
rect 18315 26104 18316 26144
rect 18356 26104 18357 26144
rect 18315 26095 18357 26104
rect 18699 26144 18741 26153
rect 18699 26104 18700 26144
rect 18740 26104 18741 26144
rect 18699 26095 18741 26104
rect 18795 26144 18837 26153
rect 18795 26104 18796 26144
rect 18836 26104 18837 26144
rect 18795 26095 18837 26104
rect 19267 26144 19325 26145
rect 19267 26104 19276 26144
rect 19316 26104 19325 26144
rect 19267 26103 19325 26104
rect 19803 26134 19845 26143
rect 15336 26093 15394 26094
rect 19803 26094 19804 26134
rect 19844 26094 19845 26134
rect 6603 26080 6645 26089
rect 19803 26085 19845 26094
rect 6499 26061 6557 26062
rect 6787 25892 6845 25893
rect 6787 25852 6796 25892
rect 6836 25852 6845 25892
rect 6787 25851 6845 25852
rect 1152 25724 20352 25748
rect 1152 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 20352 25724
rect 1152 25660 20352 25684
rect 2667 25556 2709 25565
rect 2667 25516 2668 25556
rect 2708 25516 2709 25556
rect 2667 25507 2709 25516
rect 2859 25556 2901 25565
rect 2859 25516 2860 25556
rect 2900 25516 2901 25556
rect 2859 25507 2901 25516
rect 5931 25556 5973 25565
rect 5931 25516 5932 25556
rect 5972 25516 5973 25556
rect 5931 25507 5973 25516
rect 8523 25556 8565 25565
rect 8523 25516 8524 25556
rect 8564 25516 8565 25556
rect 8523 25507 8565 25516
rect 18123 25556 18165 25565
rect 18123 25516 18124 25556
rect 18164 25516 18165 25556
rect 18123 25507 18165 25516
rect 19755 25556 19797 25565
rect 19755 25516 19756 25556
rect 19796 25516 19797 25556
rect 19755 25507 19797 25516
rect 13035 25388 13077 25397
rect 13035 25348 13036 25388
rect 13076 25348 13077 25388
rect 13035 25339 13077 25348
rect 14139 25313 14181 25322
rect 1219 25304 1277 25305
rect 1219 25264 1228 25304
rect 1268 25264 1277 25304
rect 1219 25263 1277 25264
rect 2467 25304 2525 25305
rect 2467 25264 2476 25304
rect 2516 25264 2525 25304
rect 2467 25263 2525 25264
rect 3043 25304 3101 25305
rect 3043 25264 3052 25304
rect 3092 25264 3101 25304
rect 3043 25263 3101 25264
rect 4291 25304 4349 25305
rect 4291 25264 4300 25304
rect 4340 25264 4349 25304
rect 4291 25263 4349 25264
rect 4483 25304 4541 25305
rect 4483 25264 4492 25304
rect 4532 25264 4541 25304
rect 4483 25263 4541 25264
rect 5731 25304 5789 25305
rect 5731 25264 5740 25304
rect 5780 25264 5789 25304
rect 5731 25263 5789 25264
rect 6123 25304 6165 25313
rect 6123 25264 6124 25304
rect 6164 25264 6165 25304
rect 6123 25255 6165 25264
rect 6219 25304 6261 25313
rect 6219 25264 6220 25304
rect 6260 25264 6261 25304
rect 6219 25255 6261 25264
rect 6315 25304 6357 25313
rect 6315 25264 6316 25304
rect 6356 25264 6357 25304
rect 6315 25255 6357 25264
rect 6411 25304 6453 25313
rect 6411 25264 6412 25304
rect 6452 25264 6453 25304
rect 6411 25255 6453 25264
rect 6603 25304 6645 25313
rect 6603 25264 6604 25304
rect 6644 25264 6645 25304
rect 6603 25255 6645 25264
rect 6699 25304 6741 25313
rect 6699 25264 6700 25304
rect 6740 25264 6741 25304
rect 6699 25255 6741 25264
rect 6795 25304 6837 25313
rect 6795 25264 6796 25304
rect 6836 25264 6837 25304
rect 6795 25255 6837 25264
rect 7075 25304 7133 25305
rect 7075 25264 7084 25304
rect 7124 25264 7133 25304
rect 7075 25263 7133 25264
rect 8323 25304 8381 25305
rect 8323 25264 8332 25304
rect 8372 25264 8381 25304
rect 8323 25263 8381 25264
rect 8899 25304 8957 25305
rect 8899 25264 8908 25304
rect 8948 25264 8957 25304
rect 8899 25263 8957 25264
rect 10147 25304 10205 25305
rect 10147 25264 10156 25304
rect 10196 25264 10205 25304
rect 10147 25263 10205 25264
rect 10819 25304 10877 25305
rect 10819 25264 10828 25304
rect 10868 25264 10877 25304
rect 10819 25263 10877 25264
rect 12067 25304 12125 25305
rect 12067 25264 12076 25304
rect 12116 25264 12125 25304
rect 12067 25263 12125 25264
rect 12555 25304 12597 25313
rect 12555 25264 12556 25304
rect 12596 25264 12597 25304
rect 12555 25255 12597 25264
rect 12651 25304 12693 25313
rect 12651 25264 12652 25304
rect 12692 25264 12693 25304
rect 12651 25255 12693 25264
rect 13131 25304 13173 25313
rect 13131 25264 13132 25304
rect 13172 25264 13173 25304
rect 13131 25255 13173 25264
rect 13603 25304 13661 25305
rect 13603 25264 13612 25304
rect 13652 25264 13661 25304
rect 14139 25273 14140 25313
rect 14180 25273 14181 25313
rect 14139 25264 14181 25273
rect 15147 25304 15189 25313
rect 15147 25264 15148 25304
rect 15188 25264 15189 25304
rect 13603 25263 13661 25264
rect 15147 25255 15189 25264
rect 15339 25304 15381 25313
rect 15339 25264 15340 25304
rect 15380 25264 15381 25304
rect 15339 25255 15381 25264
rect 15531 25304 15573 25313
rect 15531 25264 15532 25304
rect 15572 25264 15573 25304
rect 15531 25255 15573 25264
rect 15627 25304 15669 25313
rect 15627 25264 15628 25304
rect 15668 25264 15669 25304
rect 15627 25255 15669 25264
rect 15723 25304 15765 25313
rect 15723 25264 15724 25304
rect 15764 25264 15765 25304
rect 15723 25255 15765 25264
rect 15819 25304 15861 25313
rect 15819 25264 15820 25304
rect 15860 25264 15861 25304
rect 15819 25255 15861 25264
rect 16011 25304 16053 25313
rect 16011 25264 16012 25304
rect 16052 25264 16053 25304
rect 16011 25255 16053 25264
rect 16107 25304 16149 25313
rect 16107 25264 16108 25304
rect 16148 25264 16149 25304
rect 16107 25255 16149 25264
rect 16203 25304 16245 25313
rect 16203 25264 16204 25304
rect 16244 25264 16245 25304
rect 16203 25255 16245 25264
rect 16299 25304 16341 25313
rect 16299 25264 16300 25304
rect 16340 25264 16341 25304
rect 16299 25255 16341 25264
rect 16675 25304 16733 25305
rect 16675 25264 16684 25304
rect 16724 25264 16733 25304
rect 16675 25263 16733 25264
rect 17923 25304 17981 25305
rect 17923 25264 17932 25304
rect 17972 25264 17981 25304
rect 17923 25263 17981 25264
rect 18307 25304 18365 25305
rect 18307 25264 18316 25304
rect 18356 25264 18365 25304
rect 18307 25263 18365 25264
rect 19555 25304 19613 25305
rect 19555 25264 19564 25304
rect 19604 25264 19613 25304
rect 19555 25263 19613 25264
rect 8715 25220 8757 25229
rect 8715 25180 8716 25220
rect 8756 25180 8757 25220
rect 8715 25171 8757 25180
rect 12267 25220 12309 25229
rect 12267 25180 12268 25220
rect 12308 25180 12309 25220
rect 12267 25171 12309 25180
rect 15243 25220 15285 25229
rect 15243 25180 15244 25220
rect 15284 25180 15285 25220
rect 15243 25171 15285 25180
rect 6883 25136 6941 25137
rect 6883 25096 6892 25136
rect 6932 25096 6941 25136
rect 6883 25095 6941 25096
rect 14283 25136 14325 25145
rect 14283 25096 14284 25136
rect 14324 25096 14325 25136
rect 14283 25087 14325 25096
rect 1152 24968 20452 24992
rect 1152 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20452 24968
rect 1152 24904 20452 24928
rect 3915 24800 3957 24809
rect 3915 24760 3916 24800
rect 3956 24760 3957 24800
rect 3915 24751 3957 24760
rect 11883 24800 11925 24809
rect 11883 24760 11884 24800
rect 11924 24760 11925 24800
rect 11883 24751 11925 24760
rect 14187 24800 14229 24809
rect 14187 24760 14188 24800
rect 14228 24760 14229 24800
rect 14187 24751 14229 24760
rect 16387 24800 16445 24801
rect 16387 24760 16396 24800
rect 16436 24760 16445 24800
rect 16387 24759 16445 24760
rect 7563 24716 7605 24725
rect 7563 24676 7564 24716
rect 7604 24676 7605 24716
rect 7563 24667 7605 24676
rect 9579 24716 9621 24725
rect 9579 24676 9580 24716
rect 9620 24676 9621 24716
rect 9579 24667 9621 24676
rect 18219 24716 18261 24725
rect 18219 24676 18220 24716
rect 18260 24676 18261 24716
rect 18219 24667 18261 24676
rect 20235 24716 20277 24725
rect 20235 24676 20236 24716
rect 20276 24676 20277 24716
rect 20235 24667 20277 24676
rect 12267 24644 12309 24653
rect 1611 24632 1653 24641
rect 1611 24592 1612 24632
rect 1652 24592 1653 24632
rect 1611 24583 1653 24592
rect 1899 24632 1941 24641
rect 1899 24592 1900 24632
rect 1940 24592 1941 24632
rect 1899 24583 1941 24592
rect 2187 24632 2229 24641
rect 2187 24592 2188 24632
rect 2228 24592 2229 24632
rect 2187 24583 2229 24592
rect 2283 24632 2325 24641
rect 2283 24592 2284 24632
rect 2324 24592 2325 24632
rect 2283 24583 2325 24592
rect 2763 24632 2805 24641
rect 2763 24592 2764 24632
rect 2804 24592 2805 24632
rect 2763 24583 2805 24592
rect 3235 24632 3293 24633
rect 3235 24592 3244 24632
rect 3284 24592 3293 24632
rect 4291 24632 4349 24633
rect 3235 24591 3293 24592
rect 3723 24618 3765 24627
rect 3723 24578 3724 24618
rect 3764 24578 3765 24618
rect 4291 24592 4300 24632
rect 4340 24592 4349 24632
rect 4291 24591 4349 24592
rect 5539 24632 5597 24633
rect 5539 24592 5548 24632
rect 5588 24592 5597 24632
rect 5539 24591 5597 24592
rect 6115 24632 6173 24633
rect 6115 24592 6124 24632
rect 6164 24592 6173 24632
rect 6115 24591 6173 24592
rect 7363 24632 7421 24633
rect 7363 24592 7372 24632
rect 7412 24592 7421 24632
rect 7363 24591 7421 24592
rect 7851 24632 7893 24641
rect 7851 24592 7852 24632
rect 7892 24592 7893 24632
rect 7851 24583 7893 24592
rect 7947 24632 7989 24641
rect 7947 24592 7948 24632
rect 7988 24592 7989 24632
rect 7947 24583 7989 24592
rect 8331 24632 8373 24641
rect 8331 24592 8332 24632
rect 8372 24592 8373 24632
rect 8331 24583 8373 24592
rect 8427 24632 8469 24641
rect 8427 24592 8428 24632
rect 8468 24592 8469 24632
rect 8427 24583 8469 24592
rect 8899 24632 8957 24633
rect 8899 24592 8908 24632
rect 8948 24592 8957 24632
rect 8899 24591 8957 24592
rect 9387 24627 9429 24636
rect 9387 24587 9388 24627
rect 9428 24587 9429 24627
rect 9387 24578 9429 24587
rect 9963 24632 10005 24641
rect 9963 24592 9964 24632
rect 10004 24592 10005 24632
rect 9963 24583 10005 24592
rect 10251 24632 10293 24641
rect 10251 24592 10252 24632
rect 10292 24592 10293 24632
rect 10251 24583 10293 24592
rect 10435 24632 10493 24633
rect 10435 24592 10444 24632
rect 10484 24592 10493 24632
rect 10435 24591 10493 24592
rect 11683 24632 11741 24633
rect 11683 24592 11692 24632
rect 11732 24592 11741 24632
rect 12267 24604 12268 24644
rect 12308 24604 12309 24644
rect 12267 24595 12309 24604
rect 12363 24632 12405 24641
rect 11683 24591 11741 24592
rect 12363 24592 12364 24632
rect 12404 24592 12405 24632
rect 12363 24583 12405 24592
rect 12459 24632 12501 24641
rect 12459 24592 12460 24632
rect 12500 24592 12501 24632
rect 12459 24583 12501 24592
rect 12739 24632 12797 24633
rect 12739 24592 12748 24632
rect 12788 24592 12797 24632
rect 12739 24591 12797 24592
rect 13987 24632 14045 24633
rect 13987 24592 13996 24632
rect 14036 24592 14045 24632
rect 13987 24591 14045 24592
rect 14659 24632 14717 24633
rect 14659 24592 14668 24632
rect 14708 24592 14717 24632
rect 14659 24591 14717 24592
rect 15907 24632 15965 24633
rect 15907 24592 15916 24632
rect 15956 24592 15965 24632
rect 15907 24591 15965 24592
rect 16299 24632 16341 24641
rect 16299 24592 16300 24632
rect 16340 24592 16341 24632
rect 16299 24583 16341 24592
rect 16491 24632 16533 24641
rect 16491 24592 16492 24632
rect 16532 24592 16533 24632
rect 16491 24583 16533 24592
rect 16579 24632 16637 24633
rect 16579 24592 16588 24632
rect 16628 24592 16637 24632
rect 16579 24591 16637 24592
rect 16771 24632 16829 24633
rect 16771 24592 16780 24632
rect 16820 24592 16829 24632
rect 16771 24591 16829 24592
rect 18019 24632 18077 24633
rect 18019 24592 18028 24632
rect 18068 24592 18077 24632
rect 18019 24591 18077 24592
rect 18507 24632 18549 24641
rect 18507 24592 18508 24632
rect 18548 24592 18549 24632
rect 18507 24583 18549 24592
rect 18603 24632 18645 24641
rect 18603 24592 18604 24632
rect 18644 24592 18645 24632
rect 18603 24583 18645 24592
rect 18987 24632 19029 24641
rect 18987 24592 18988 24632
rect 19028 24592 19029 24632
rect 18987 24583 19029 24592
rect 19555 24632 19613 24633
rect 19555 24592 19564 24632
rect 19604 24592 19613 24632
rect 19555 24591 19613 24592
rect 20043 24618 20085 24627
rect 20043 24578 20044 24618
rect 20084 24578 20085 24618
rect 3723 24569 3765 24578
rect 20043 24569 20085 24578
rect 2667 24548 2709 24557
rect 2667 24508 2668 24548
rect 2708 24508 2709 24548
rect 2667 24499 2709 24508
rect 19083 24548 19125 24557
rect 19083 24508 19084 24548
rect 19124 24508 19125 24548
rect 19083 24499 19125 24508
rect 1899 24380 1941 24389
rect 1899 24340 1900 24380
rect 1940 24340 1941 24380
rect 1899 24331 1941 24340
rect 5739 24380 5781 24389
rect 5739 24340 5740 24380
rect 5780 24340 5781 24380
rect 5739 24331 5781 24340
rect 10251 24380 10293 24389
rect 10251 24340 10252 24380
rect 10292 24340 10293 24380
rect 10251 24331 10293 24340
rect 11883 24380 11925 24389
rect 11883 24340 11884 24380
rect 11924 24340 11925 24380
rect 11883 24331 11925 24340
rect 12067 24380 12125 24381
rect 12067 24340 12076 24380
rect 12116 24340 12125 24380
rect 12067 24339 12125 24340
rect 16107 24380 16149 24389
rect 16107 24340 16108 24380
rect 16148 24340 16149 24380
rect 16107 24331 16149 24340
rect 1152 24212 20352 24236
rect 1152 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 20352 24212
rect 1152 24148 20352 24172
rect 16003 24044 16061 24045
rect 16003 24004 16012 24044
rect 16052 24004 16061 24044
rect 16003 24003 16061 24004
rect 5643 23960 5685 23969
rect 5643 23920 5644 23960
rect 5684 23920 5685 23960
rect 5643 23911 5685 23920
rect 15811 23960 15869 23961
rect 15811 23920 15820 23960
rect 15860 23920 15869 23960
rect 15811 23919 15869 23920
rect 18603 23960 18645 23969
rect 18603 23920 18604 23960
rect 18644 23920 18645 23960
rect 18603 23911 18645 23920
rect 20235 23960 20277 23969
rect 20235 23920 20236 23960
rect 20276 23920 20277 23960
rect 20235 23911 20277 23920
rect 2763 23876 2805 23885
rect 2763 23836 2764 23876
rect 2804 23836 2805 23876
rect 2763 23827 2805 23836
rect 13227 23876 13269 23885
rect 13227 23836 13228 23876
rect 13268 23836 13269 23876
rect 5923 23834 5981 23835
rect 3867 23801 3909 23810
rect 2283 23792 2325 23801
rect 2283 23752 2284 23792
rect 2324 23752 2325 23792
rect 2283 23743 2325 23752
rect 2379 23792 2421 23801
rect 2379 23752 2380 23792
rect 2420 23752 2421 23792
rect 2379 23743 2421 23752
rect 2859 23792 2901 23801
rect 2859 23752 2860 23792
rect 2900 23752 2901 23792
rect 2859 23743 2901 23752
rect 3331 23792 3389 23793
rect 3331 23752 3340 23792
rect 3380 23752 3389 23792
rect 3867 23761 3868 23801
rect 3908 23761 3909 23801
rect 5923 23794 5932 23834
rect 5972 23794 5981 23834
rect 13227 23827 13269 23836
rect 5923 23793 5981 23794
rect 3867 23752 3909 23761
rect 4195 23792 4253 23793
rect 4195 23752 4204 23792
rect 4244 23752 4253 23792
rect 3331 23751 3389 23752
rect 4195 23751 4253 23752
rect 5443 23792 5501 23793
rect 5443 23752 5452 23792
rect 5492 23752 5501 23792
rect 5443 23751 5501 23752
rect 6027 23792 6069 23801
rect 6027 23752 6028 23792
rect 6068 23752 6069 23792
rect 6027 23743 6069 23752
rect 6123 23792 6165 23801
rect 6123 23752 6124 23792
rect 6164 23752 6165 23792
rect 6123 23743 6165 23752
rect 6499 23792 6557 23793
rect 6499 23752 6508 23792
rect 6548 23752 6557 23792
rect 6499 23751 6557 23752
rect 7747 23792 7805 23793
rect 7747 23752 7756 23792
rect 7796 23752 7805 23792
rect 7747 23751 7805 23752
rect 8331 23792 8373 23801
rect 8331 23752 8332 23792
rect 8372 23752 8373 23792
rect 8331 23743 8373 23752
rect 8427 23792 8469 23801
rect 8427 23752 8428 23792
rect 8468 23752 8469 23792
rect 8427 23743 8469 23752
rect 8811 23792 8853 23801
rect 8811 23752 8812 23792
rect 8852 23752 8853 23792
rect 8811 23743 8853 23752
rect 8907 23792 8949 23801
rect 9867 23797 9909 23806
rect 14235 23801 14277 23810
rect 8907 23752 8908 23792
rect 8948 23752 8949 23792
rect 8907 23743 8949 23752
rect 9379 23792 9437 23793
rect 9379 23752 9388 23792
rect 9428 23752 9437 23792
rect 9379 23751 9437 23752
rect 9867 23757 9868 23797
rect 9908 23757 9909 23797
rect 9867 23748 9909 23757
rect 10443 23792 10485 23801
rect 10443 23752 10444 23792
rect 10484 23752 10485 23792
rect 10443 23743 10485 23752
rect 10635 23792 10677 23801
rect 10635 23752 10636 23792
rect 10676 23752 10677 23792
rect 10635 23743 10677 23752
rect 10723 23792 10781 23793
rect 10723 23752 10732 23792
rect 10772 23752 10781 23792
rect 10723 23751 10781 23752
rect 10915 23792 10973 23793
rect 10915 23752 10924 23792
rect 10964 23752 10973 23792
rect 10915 23751 10973 23752
rect 12163 23792 12221 23793
rect 12163 23752 12172 23792
rect 12212 23752 12221 23792
rect 12163 23751 12221 23752
rect 12651 23792 12693 23801
rect 12651 23752 12652 23792
rect 12692 23752 12693 23792
rect 12651 23743 12693 23752
rect 12747 23792 12789 23801
rect 12747 23752 12748 23792
rect 12788 23752 12789 23792
rect 12747 23743 12789 23752
rect 13131 23792 13173 23801
rect 13131 23752 13132 23792
rect 13172 23752 13173 23792
rect 13131 23743 13173 23752
rect 13699 23792 13757 23793
rect 13699 23752 13708 23792
rect 13748 23752 13757 23792
rect 14235 23761 14236 23801
rect 14276 23761 14277 23801
rect 14235 23752 14277 23761
rect 14571 23792 14613 23801
rect 14571 23752 14572 23792
rect 14612 23752 14613 23792
rect 15139 23792 15197 23793
rect 13699 23751 13757 23752
rect 14571 23743 14613 23752
rect 14667 23771 14709 23780
rect 14667 23731 14668 23771
rect 14708 23731 14709 23771
rect 14667 23722 14709 23731
rect 14763 23771 14805 23780
rect 14763 23731 14764 23771
rect 14804 23731 14805 23771
rect 15139 23752 15148 23792
rect 15188 23752 15197 23792
rect 15139 23751 15197 23752
rect 15435 23792 15477 23801
rect 15435 23752 15436 23792
rect 15476 23752 15477 23792
rect 15435 23743 15477 23752
rect 16299 23792 16341 23801
rect 16299 23752 16300 23792
rect 16340 23752 16341 23792
rect 16299 23743 16341 23752
rect 16395 23792 16437 23801
rect 16395 23752 16396 23792
rect 16436 23752 16437 23792
rect 16395 23743 16437 23752
rect 16675 23792 16733 23793
rect 16675 23752 16684 23792
rect 16724 23752 16733 23792
rect 16675 23751 16733 23752
rect 17155 23792 17213 23793
rect 17155 23752 17164 23792
rect 17204 23752 17213 23792
rect 17155 23751 17213 23752
rect 18403 23792 18461 23793
rect 18403 23752 18412 23792
rect 18452 23752 18461 23792
rect 18403 23751 18461 23752
rect 18787 23792 18845 23793
rect 18787 23752 18796 23792
rect 18836 23752 18845 23792
rect 18787 23751 18845 23752
rect 20035 23792 20093 23793
rect 20035 23752 20044 23792
rect 20084 23752 20093 23792
rect 20035 23751 20093 23752
rect 14763 23722 14805 23731
rect 7947 23708 7989 23717
rect 7947 23668 7948 23708
rect 7988 23668 7989 23708
rect 7947 23659 7989 23668
rect 10059 23708 10101 23717
rect 10059 23668 10060 23708
rect 10100 23668 10101 23708
rect 10059 23659 10101 23668
rect 12363 23708 12405 23717
rect 12363 23668 12364 23708
rect 12404 23668 12405 23708
rect 12363 23659 12405 23668
rect 14379 23708 14421 23717
rect 14379 23668 14380 23708
rect 14420 23668 14421 23708
rect 14379 23659 14421 23668
rect 15531 23708 15573 23717
rect 15531 23668 15532 23708
rect 15572 23668 15573 23708
rect 15531 23659 15573 23668
rect 4011 23624 4053 23633
rect 4011 23584 4012 23624
rect 4052 23584 4053 23624
rect 4011 23575 4053 23584
rect 6315 23624 6357 23633
rect 6315 23584 6316 23624
rect 6356 23584 6357 23624
rect 6315 23575 6357 23584
rect 10531 23624 10589 23625
rect 10531 23584 10540 23624
rect 10580 23584 10589 23624
rect 10531 23583 10589 23584
rect 14851 23624 14909 23625
rect 14851 23584 14860 23624
rect 14900 23584 14909 23624
rect 14851 23583 14909 23584
rect 1152 23456 20452 23480
rect 1152 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20452 23456
rect 1152 23392 20452 23416
rect 2667 23288 2709 23297
rect 2667 23248 2668 23288
rect 2708 23248 2709 23288
rect 2667 23239 2709 23248
rect 5443 23288 5501 23289
rect 5443 23248 5452 23288
rect 5492 23248 5501 23288
rect 5443 23247 5501 23248
rect 6115 23288 6173 23289
rect 6115 23248 6124 23288
rect 6164 23248 6173 23288
rect 6115 23247 6173 23248
rect 9867 23288 9909 23297
rect 9867 23248 9868 23288
rect 9908 23248 9909 23288
rect 9867 23239 9909 23248
rect 11499 23288 11541 23297
rect 11499 23248 11500 23288
rect 11540 23248 11541 23288
rect 11499 23239 11541 23248
rect 12067 23288 12125 23289
rect 12067 23248 12076 23288
rect 12116 23248 12125 23288
rect 12067 23247 12125 23248
rect 14379 23288 14421 23297
rect 14379 23248 14380 23288
rect 14420 23248 14421 23288
rect 14379 23239 14421 23248
rect 14859 23288 14901 23297
rect 14859 23248 14860 23288
rect 14900 23248 14901 23288
rect 14859 23239 14901 23248
rect 15051 23288 15093 23297
rect 15051 23248 15052 23288
rect 15092 23248 15093 23288
rect 15051 23239 15093 23248
rect 16771 23288 16829 23289
rect 16771 23248 16780 23288
rect 16820 23248 16829 23288
rect 16771 23247 16829 23248
rect 17443 23288 17501 23289
rect 17443 23248 17452 23288
rect 17492 23248 17501 23288
rect 17443 23247 17501 23248
rect 17739 23288 17781 23297
rect 17739 23248 17740 23288
rect 17780 23248 17781 23288
rect 17739 23239 17781 23248
rect 20139 23288 20181 23297
rect 20139 23248 20140 23288
rect 20180 23248 20181 23288
rect 20139 23239 20181 23248
rect 18027 23204 18069 23213
rect 18027 23164 18028 23204
rect 18068 23164 18069 23204
rect 18027 23155 18069 23164
rect 1219 23120 1277 23121
rect 1219 23080 1228 23120
rect 1268 23080 1277 23120
rect 1219 23079 1277 23080
rect 2467 23120 2525 23121
rect 2467 23080 2476 23120
rect 2516 23080 2525 23120
rect 2467 23079 2525 23080
rect 3715 23120 3773 23121
rect 3715 23080 3724 23120
rect 3764 23080 3773 23120
rect 3715 23079 3773 23080
rect 4963 23120 5021 23121
rect 4963 23080 4972 23120
rect 5012 23080 5021 23120
rect 4963 23079 5021 23080
rect 5355 23120 5397 23129
rect 5355 23080 5356 23120
rect 5396 23080 5397 23120
rect 5355 23071 5397 23080
rect 5547 23120 5589 23129
rect 5547 23080 5548 23120
rect 5588 23080 5589 23120
rect 5547 23071 5589 23080
rect 5635 23120 5693 23121
rect 5635 23080 5644 23120
rect 5684 23080 5693 23120
rect 5635 23079 5693 23080
rect 5835 23120 5877 23129
rect 5835 23080 5836 23120
rect 5876 23080 5877 23120
rect 5835 23071 5877 23080
rect 5931 23120 5973 23129
rect 5931 23080 5932 23120
rect 5972 23080 5973 23120
rect 5931 23071 5973 23080
rect 6027 23120 6069 23129
rect 6027 23080 6028 23120
rect 6068 23080 6069 23120
rect 6027 23071 6069 23080
rect 6307 23120 6365 23121
rect 6307 23080 6316 23120
rect 6356 23080 6365 23120
rect 6307 23079 6365 23080
rect 7555 23120 7613 23121
rect 7555 23080 7564 23120
rect 7604 23080 7613 23120
rect 7555 23079 7613 23080
rect 8419 23120 8477 23121
rect 8419 23080 8428 23120
rect 8468 23080 8477 23120
rect 8419 23079 8477 23080
rect 9667 23120 9725 23121
rect 9667 23080 9676 23120
rect 9716 23080 9725 23120
rect 9667 23079 9725 23080
rect 10051 23120 10109 23121
rect 10051 23080 10060 23120
rect 10100 23080 10109 23120
rect 10051 23079 10109 23080
rect 11299 23120 11357 23121
rect 11299 23080 11308 23120
rect 11348 23080 11357 23120
rect 11299 23079 11357 23080
rect 11787 23120 11829 23129
rect 11787 23080 11788 23120
rect 11828 23080 11829 23120
rect 11787 23071 11829 23080
rect 11883 23120 11925 23129
rect 11883 23080 11884 23120
rect 11924 23080 11925 23120
rect 11883 23071 11925 23080
rect 11979 23120 12021 23129
rect 11979 23080 11980 23120
rect 12020 23080 12021 23120
rect 11979 23071 12021 23080
rect 12931 23120 12989 23121
rect 12931 23080 12940 23120
rect 12980 23080 12989 23120
rect 12931 23079 12989 23080
rect 14179 23120 14237 23121
rect 14179 23080 14188 23120
rect 14228 23080 14237 23120
rect 14179 23079 14237 23080
rect 14755 23120 14813 23121
rect 14755 23080 14764 23120
rect 14804 23080 14813 23120
rect 14755 23079 14813 23080
rect 15235 23120 15293 23121
rect 15235 23080 15244 23120
rect 15284 23080 15293 23120
rect 15235 23079 15293 23080
rect 16683 23120 16725 23129
rect 16683 23080 16684 23120
rect 16724 23080 16725 23120
rect 16483 23078 16541 23079
rect 16483 23038 16492 23078
rect 16532 23038 16541 23078
rect 16683 23071 16725 23080
rect 16875 23120 16917 23129
rect 16875 23080 16876 23120
rect 16916 23080 16917 23120
rect 16875 23071 16917 23080
rect 16963 23120 17021 23121
rect 16963 23080 16972 23120
rect 17012 23080 17021 23120
rect 16963 23079 17021 23080
rect 17163 23120 17205 23129
rect 17163 23080 17164 23120
rect 17204 23080 17205 23120
rect 17163 23071 17205 23080
rect 17259 23120 17301 23129
rect 17259 23080 17260 23120
rect 17300 23080 17301 23120
rect 17259 23071 17301 23080
rect 17355 23120 17397 23129
rect 17355 23080 17356 23120
rect 17396 23080 17397 23120
rect 17355 23071 17397 23080
rect 17635 23120 17693 23121
rect 17635 23080 17644 23120
rect 17684 23080 17693 23120
rect 17635 23079 17693 23080
rect 17923 23120 17981 23121
rect 17923 23080 17932 23120
rect 17972 23080 17981 23120
rect 17923 23079 17981 23080
rect 18691 23120 18749 23121
rect 18691 23080 18700 23120
rect 18740 23080 18749 23120
rect 18691 23079 18749 23080
rect 19939 23120 19997 23121
rect 19939 23080 19948 23120
rect 19988 23080 19997 23120
rect 19939 23079 19997 23080
rect 16483 23037 16541 23038
rect 5163 22868 5205 22877
rect 5163 22828 5164 22868
rect 5204 22828 5205 22868
rect 5163 22819 5205 22828
rect 7755 22868 7797 22877
rect 7755 22828 7756 22868
rect 7796 22828 7797 22868
rect 7755 22819 7797 22828
rect 1152 22700 20352 22724
rect 1152 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 20352 22700
rect 1152 22636 20352 22660
rect 2667 22532 2709 22541
rect 2667 22492 2668 22532
rect 2708 22492 2709 22532
rect 2667 22483 2709 22492
rect 4299 22532 4341 22541
rect 4299 22492 4300 22532
rect 4340 22492 4341 22532
rect 4299 22483 4341 22492
rect 15147 22532 15189 22541
rect 15147 22492 15148 22532
rect 15188 22492 15189 22532
rect 15147 22483 15189 22492
rect 18219 22448 18261 22457
rect 18219 22408 18220 22448
rect 18260 22408 18261 22448
rect 18219 22399 18261 22408
rect 5259 22364 5301 22373
rect 5259 22324 5260 22364
rect 5300 22324 5301 22364
rect 5259 22315 5301 22324
rect 5355 22364 5397 22373
rect 5355 22324 5356 22364
rect 5396 22324 5397 22364
rect 5355 22315 5397 22324
rect 8331 22364 8373 22373
rect 8331 22324 8332 22364
rect 8372 22324 8373 22364
rect 8331 22315 8373 22324
rect 12843 22364 12885 22373
rect 12843 22324 12844 22364
rect 12884 22324 12885 22364
rect 12843 22315 12885 22324
rect 18987 22364 19029 22373
rect 18987 22324 18988 22364
rect 19028 22324 19029 22364
rect 18987 22315 19029 22324
rect 19083 22364 19125 22373
rect 19083 22324 19084 22364
rect 19124 22324 19125 22364
rect 19083 22315 19125 22324
rect 4779 22299 4821 22308
rect 1219 22280 1277 22281
rect 1219 22240 1228 22280
rect 1268 22240 1277 22280
rect 1219 22239 1277 22240
rect 2467 22280 2525 22281
rect 2467 22240 2476 22280
rect 2516 22240 2525 22280
rect 2467 22239 2525 22240
rect 2851 22280 2909 22281
rect 2851 22240 2860 22280
rect 2900 22240 2909 22280
rect 2851 22239 2909 22240
rect 4099 22280 4157 22281
rect 4099 22240 4108 22280
rect 4148 22240 4157 22280
rect 4779 22259 4780 22299
rect 4820 22259 4821 22299
rect 4779 22250 4821 22259
rect 4875 22280 4917 22289
rect 6315 22285 6357 22294
rect 4099 22239 4157 22240
rect 4875 22240 4876 22280
rect 4916 22240 4917 22280
rect 4875 22231 4917 22240
rect 5827 22280 5885 22281
rect 5827 22240 5836 22280
rect 5876 22240 5885 22280
rect 5827 22239 5885 22240
rect 6315 22245 6316 22285
rect 6356 22245 6357 22285
rect 6315 22236 6357 22245
rect 7755 22280 7797 22289
rect 7755 22240 7756 22280
rect 7796 22240 7797 22280
rect 7755 22231 7797 22240
rect 7851 22280 7893 22289
rect 7851 22240 7852 22280
rect 7892 22240 7893 22280
rect 7851 22231 7893 22240
rect 8235 22280 8277 22289
rect 9291 22285 9333 22294
rect 8235 22240 8236 22280
rect 8276 22240 8277 22280
rect 8235 22231 8277 22240
rect 8803 22280 8861 22281
rect 8803 22240 8812 22280
rect 8852 22240 8861 22280
rect 8803 22239 8861 22240
rect 9291 22245 9292 22285
rect 9332 22245 9333 22285
rect 9291 22236 9333 22245
rect 10531 22280 10589 22281
rect 10531 22240 10540 22280
rect 10580 22240 10589 22280
rect 10531 22239 10589 22240
rect 11779 22280 11837 22281
rect 11779 22240 11788 22280
rect 11828 22240 11837 22280
rect 11779 22239 11837 22240
rect 12267 22280 12309 22289
rect 12267 22240 12268 22280
rect 12308 22240 12309 22280
rect 12267 22231 12309 22240
rect 12363 22280 12405 22289
rect 12363 22240 12364 22280
rect 12404 22240 12405 22280
rect 12363 22231 12405 22240
rect 12747 22280 12789 22289
rect 13803 22285 13845 22294
rect 12747 22240 12748 22280
rect 12788 22240 12789 22280
rect 12747 22231 12789 22240
rect 13315 22280 13373 22281
rect 13315 22240 13324 22280
rect 13364 22240 13373 22280
rect 13315 22239 13373 22240
rect 13803 22245 13804 22285
rect 13844 22245 13845 22285
rect 14366 22293 14424 22294
rect 14366 22253 14375 22293
rect 14415 22253 14424 22293
rect 14366 22252 14424 22253
rect 14667 22280 14709 22289
rect 13803 22236 13845 22245
rect 14667 22240 14668 22280
rect 14708 22240 14709 22280
rect 14667 22231 14709 22240
rect 14859 22280 14901 22289
rect 14859 22240 14860 22280
rect 14900 22240 14901 22280
rect 14859 22231 14901 22240
rect 14955 22280 14997 22289
rect 14955 22240 14956 22280
rect 14996 22240 14997 22280
rect 14955 22231 14997 22240
rect 15331 22280 15389 22281
rect 15331 22240 15340 22280
rect 15380 22240 15389 22280
rect 15331 22239 15389 22240
rect 16579 22280 16637 22281
rect 16579 22240 16588 22280
rect 16628 22240 16637 22280
rect 16579 22239 16637 22240
rect 16771 22280 16829 22281
rect 16771 22240 16780 22280
rect 16820 22240 16829 22280
rect 16771 22239 16829 22240
rect 18019 22280 18077 22281
rect 18019 22240 18028 22280
rect 18068 22240 18077 22280
rect 18019 22239 18077 22240
rect 18507 22280 18549 22289
rect 18507 22240 18508 22280
rect 18548 22240 18549 22280
rect 18507 22231 18549 22240
rect 18603 22280 18645 22289
rect 20043 22285 20085 22294
rect 18603 22240 18604 22280
rect 18644 22240 18645 22280
rect 18603 22231 18645 22240
rect 19555 22280 19613 22281
rect 19555 22240 19564 22280
rect 19604 22240 19613 22280
rect 19555 22239 19613 22240
rect 20043 22245 20044 22285
rect 20084 22245 20085 22285
rect 20043 22236 20085 22245
rect 11979 22196 12021 22205
rect 11979 22156 11980 22196
rect 12020 22156 12021 22196
rect 11979 22147 12021 22156
rect 20235 22196 20277 22205
rect 20235 22156 20236 22196
rect 20276 22156 20277 22196
rect 20235 22147 20277 22156
rect 6507 22112 6549 22121
rect 6507 22072 6508 22112
rect 6548 22072 6549 22112
rect 6507 22063 6549 22072
rect 9483 22112 9525 22121
rect 9483 22072 9484 22112
rect 9524 22072 9525 22112
rect 9483 22063 9525 22072
rect 13995 22112 14037 22121
rect 13995 22072 13996 22112
rect 14036 22072 14037 22112
rect 13995 22063 14037 22072
rect 14475 22112 14517 22121
rect 14475 22072 14476 22112
rect 14516 22072 14517 22112
rect 14475 22063 14517 22072
rect 14763 22112 14805 22121
rect 14763 22072 14764 22112
rect 14804 22072 14805 22112
rect 14763 22063 14805 22072
rect 1152 21944 20452 21968
rect 1152 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20452 21944
rect 1152 21880 20452 21904
rect 9291 21776 9333 21785
rect 9291 21736 9292 21776
rect 9332 21736 9333 21776
rect 9291 21727 9333 21736
rect 13707 21776 13749 21785
rect 13707 21736 13708 21776
rect 13748 21736 13749 21776
rect 13707 21727 13749 21736
rect 15339 21776 15381 21785
rect 15339 21736 15340 21776
rect 15380 21736 15381 21776
rect 15339 21727 15381 21736
rect 15715 21776 15773 21777
rect 15715 21736 15724 21776
rect 15764 21736 15773 21776
rect 15715 21735 15773 21736
rect 20139 21776 20181 21785
rect 20139 21736 20140 21776
rect 20180 21736 20181 21776
rect 20139 21727 20181 21736
rect 2475 21692 2517 21701
rect 2475 21652 2476 21692
rect 2516 21652 2517 21692
rect 2475 21643 2517 21652
rect 6219 21692 6261 21701
rect 6219 21652 6220 21692
rect 6260 21652 6261 21692
rect 6219 21643 6261 21652
rect 18123 21692 18165 21701
rect 18123 21652 18124 21692
rect 18164 21652 18165 21692
rect 18123 21643 18165 21652
rect 3139 21608 3197 21609
rect 2667 21594 2709 21603
rect 2667 21554 2668 21594
rect 2708 21554 2709 21594
rect 3139 21568 3148 21608
rect 3188 21568 3197 21608
rect 3139 21567 3197 21568
rect 4107 21608 4149 21617
rect 4107 21568 4108 21608
rect 4148 21568 4149 21608
rect 4107 21559 4149 21568
rect 4203 21608 4245 21617
rect 4203 21568 4204 21608
rect 4244 21568 4245 21608
rect 4203 21559 4245 21568
rect 4771 21608 4829 21609
rect 4771 21568 4780 21608
rect 4820 21568 4829 21608
rect 4771 21567 4829 21568
rect 6019 21608 6077 21609
rect 6019 21568 6028 21608
rect 6068 21568 6077 21608
rect 6019 21567 6077 21568
rect 7843 21608 7901 21609
rect 7843 21568 7852 21608
rect 7892 21568 7901 21608
rect 7843 21567 7901 21568
rect 9091 21608 9149 21609
rect 9091 21568 9100 21608
rect 9140 21568 9149 21608
rect 9091 21567 9149 21568
rect 9475 21608 9533 21609
rect 9475 21568 9484 21608
rect 9524 21568 9533 21608
rect 9475 21567 9533 21568
rect 10723 21608 10781 21609
rect 10723 21568 10732 21608
rect 10772 21568 10781 21608
rect 10723 21567 10781 21568
rect 12259 21608 12317 21609
rect 12259 21568 12268 21608
rect 12308 21568 12317 21608
rect 12259 21567 12317 21568
rect 13507 21608 13565 21609
rect 13507 21568 13516 21608
rect 13556 21568 13565 21608
rect 13507 21567 13565 21568
rect 13891 21608 13949 21609
rect 13891 21568 13900 21608
rect 13940 21568 13949 21608
rect 13891 21567 13949 21568
rect 15139 21608 15197 21609
rect 15139 21568 15148 21608
rect 15188 21568 15197 21608
rect 15139 21567 15197 21568
rect 15523 21608 15581 21609
rect 15523 21568 15532 21608
rect 15572 21568 15581 21608
rect 15523 21567 15581 21568
rect 15619 21608 15677 21609
rect 15619 21568 15628 21608
rect 15668 21568 15677 21608
rect 15619 21567 15677 21568
rect 15819 21608 15861 21617
rect 15819 21568 15820 21608
rect 15860 21568 15861 21608
rect 15819 21559 15861 21568
rect 15915 21608 15957 21617
rect 15915 21568 15916 21608
rect 15956 21568 15957 21608
rect 15915 21559 15957 21568
rect 16008 21608 16066 21609
rect 16008 21568 16017 21608
rect 16057 21568 16066 21608
rect 16008 21567 16066 21568
rect 16675 21608 16733 21609
rect 16675 21568 16684 21608
rect 16724 21568 16733 21608
rect 16675 21567 16733 21568
rect 17923 21608 17981 21609
rect 17923 21568 17932 21608
rect 17972 21568 17981 21608
rect 17923 21567 17981 21568
rect 18411 21608 18453 21617
rect 18411 21568 18412 21608
rect 18452 21568 18453 21608
rect 18411 21559 18453 21568
rect 18507 21608 18549 21617
rect 18507 21568 18508 21608
rect 18548 21568 18549 21608
rect 18507 21559 18549 21568
rect 18891 21608 18933 21617
rect 18891 21568 18892 21608
rect 18932 21568 18933 21608
rect 18891 21559 18933 21568
rect 18987 21608 19029 21617
rect 18987 21568 18988 21608
rect 19028 21568 19029 21608
rect 18987 21559 19029 21568
rect 19459 21608 19517 21609
rect 19459 21568 19468 21608
rect 19508 21568 19517 21608
rect 19459 21567 19517 21568
rect 19947 21594 19989 21603
rect 2667 21545 2709 21554
rect 19947 21554 19948 21594
rect 19988 21554 19989 21594
rect 19947 21545 19989 21554
rect 2083 21524 2141 21525
rect 2083 21484 2092 21524
rect 2132 21484 2141 21524
rect 2083 21483 2141 21484
rect 3627 21524 3669 21533
rect 3627 21484 3628 21524
rect 3668 21484 3669 21524
rect 3627 21475 3669 21484
rect 3723 21524 3765 21533
rect 3723 21484 3724 21524
rect 3764 21484 3765 21524
rect 3723 21475 3765 21484
rect 1899 21356 1941 21365
rect 1899 21316 1900 21356
rect 1940 21316 1941 21356
rect 1899 21307 1941 21316
rect 10923 21356 10965 21365
rect 10923 21316 10924 21356
rect 10964 21316 10965 21356
rect 10923 21307 10965 21316
rect 1152 21188 20352 21212
rect 1152 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 20352 21188
rect 1152 21124 20352 21148
rect 15147 21020 15189 21029
rect 15147 20980 15148 21020
rect 15188 20980 15189 21020
rect 15147 20971 15189 20980
rect 6315 20852 6357 20861
rect 6315 20812 6316 20852
rect 6356 20812 6357 20852
rect 6315 20803 6357 20812
rect 9099 20852 9141 20861
rect 9099 20812 9100 20852
rect 9140 20812 9141 20852
rect 9099 20803 9141 20812
rect 11115 20852 11157 20861
rect 11115 20812 11116 20852
rect 11156 20812 11157 20852
rect 11115 20803 11157 20812
rect 1219 20768 1277 20769
rect 1219 20728 1228 20768
rect 1268 20728 1277 20768
rect 1219 20727 1277 20728
rect 2467 20768 2525 20769
rect 2467 20728 2476 20768
rect 2516 20728 2525 20768
rect 2467 20727 2525 20728
rect 4003 20768 4061 20769
rect 4003 20728 4012 20768
rect 4052 20728 4061 20768
rect 4003 20727 4061 20728
rect 5251 20768 5309 20769
rect 5251 20728 5260 20768
rect 5300 20728 5309 20768
rect 5251 20727 5309 20728
rect 5739 20768 5781 20777
rect 5739 20728 5740 20768
rect 5780 20728 5781 20768
rect 5739 20719 5781 20728
rect 5835 20768 5877 20777
rect 5835 20728 5836 20768
rect 5876 20728 5877 20768
rect 5835 20719 5877 20728
rect 6219 20768 6261 20777
rect 7275 20773 7317 20782
rect 10107 20777 10149 20786
rect 12123 20777 12165 20786
rect 6219 20728 6220 20768
rect 6260 20728 6261 20768
rect 6219 20719 6261 20728
rect 6787 20768 6845 20769
rect 6787 20728 6796 20768
rect 6836 20728 6845 20768
rect 6787 20727 6845 20728
rect 7275 20733 7276 20773
rect 7316 20733 7317 20773
rect 7275 20724 7317 20733
rect 8523 20768 8565 20777
rect 8523 20728 8524 20768
rect 8564 20728 8565 20768
rect 8523 20719 8565 20728
rect 8619 20768 8661 20777
rect 8619 20728 8620 20768
rect 8660 20728 8661 20768
rect 8619 20719 8661 20728
rect 9003 20768 9045 20777
rect 9003 20728 9004 20768
rect 9044 20728 9045 20768
rect 9003 20719 9045 20728
rect 9571 20768 9629 20769
rect 9571 20728 9580 20768
rect 9620 20728 9629 20768
rect 10107 20737 10108 20777
rect 10148 20737 10149 20777
rect 10107 20728 10149 20737
rect 10539 20768 10581 20777
rect 10539 20728 10540 20768
rect 10580 20728 10581 20768
rect 9571 20727 9629 20728
rect 10539 20719 10581 20728
rect 10635 20768 10677 20777
rect 10635 20728 10636 20768
rect 10676 20728 10677 20768
rect 10635 20719 10677 20728
rect 11019 20768 11061 20777
rect 11019 20728 11020 20768
rect 11060 20728 11061 20768
rect 11019 20719 11061 20728
rect 11587 20768 11645 20769
rect 11587 20728 11596 20768
rect 11636 20728 11645 20768
rect 12123 20737 12124 20777
rect 12164 20737 12165 20777
rect 12123 20728 12165 20737
rect 13699 20768 13757 20769
rect 13699 20728 13708 20768
rect 13748 20728 13757 20768
rect 11587 20727 11645 20728
rect 13699 20727 13757 20728
rect 14947 20768 15005 20769
rect 14947 20728 14956 20768
rect 14996 20728 15005 20768
rect 14947 20727 15005 20728
rect 15339 20768 15381 20777
rect 15339 20728 15340 20768
rect 15380 20728 15381 20768
rect 15339 20719 15381 20728
rect 15435 20768 15477 20777
rect 15435 20728 15436 20768
rect 15476 20728 15477 20768
rect 15435 20719 15477 20728
rect 16099 20768 16157 20769
rect 16099 20728 16108 20768
rect 16148 20728 16157 20768
rect 16099 20727 16157 20728
rect 16299 20768 16341 20777
rect 16299 20728 16300 20768
rect 16340 20728 16341 20768
rect 16299 20719 16341 20728
rect 16395 20768 16437 20777
rect 16395 20728 16396 20768
rect 16436 20728 16437 20768
rect 16395 20719 16437 20728
rect 16491 20768 16533 20777
rect 16491 20728 16492 20768
rect 16532 20728 16533 20768
rect 16491 20719 16533 20728
rect 16771 20768 16829 20769
rect 16771 20728 16780 20768
rect 16820 20728 16829 20768
rect 16771 20727 16829 20728
rect 16875 20768 16917 20777
rect 16875 20728 16876 20768
rect 16916 20728 16917 20768
rect 16875 20719 16917 20728
rect 17067 20768 17109 20777
rect 17067 20728 17068 20768
rect 17108 20728 17109 20768
rect 17067 20719 17109 20728
rect 18499 20768 18557 20769
rect 18499 20728 18508 20768
rect 18548 20728 18557 20768
rect 18499 20727 18557 20728
rect 19747 20768 19805 20769
rect 19747 20728 19756 20768
rect 19796 20728 19805 20768
rect 19747 20727 19805 20728
rect 2667 20684 2709 20693
rect 2667 20644 2668 20684
rect 2708 20644 2709 20684
rect 2667 20635 2709 20644
rect 5451 20684 5493 20693
rect 5451 20644 5452 20684
rect 5492 20644 5493 20684
rect 5451 20635 5493 20644
rect 10251 20684 10293 20693
rect 10251 20644 10252 20684
rect 10292 20644 10293 20684
rect 10251 20635 10293 20644
rect 7467 20600 7509 20609
rect 7467 20560 7468 20600
rect 7508 20560 7509 20600
rect 7467 20551 7509 20560
rect 12267 20600 12309 20609
rect 12267 20560 12268 20600
rect 12308 20560 12309 20600
rect 12267 20551 12309 20560
rect 15619 20600 15677 20601
rect 15619 20560 15628 20600
rect 15668 20560 15677 20600
rect 15619 20559 15677 20560
rect 16011 20600 16053 20609
rect 16011 20560 16012 20600
rect 16052 20560 16053 20600
rect 16011 20551 16053 20560
rect 16579 20600 16637 20601
rect 16579 20560 16588 20600
rect 16628 20560 16637 20600
rect 16579 20559 16637 20560
rect 16963 20600 17021 20601
rect 16963 20560 16972 20600
rect 17012 20560 17021 20600
rect 16963 20559 17021 20560
rect 19947 20600 19989 20609
rect 19947 20560 19948 20600
rect 19988 20560 19989 20600
rect 19947 20551 19989 20560
rect 1152 20432 20452 20456
rect 1152 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20452 20432
rect 1152 20368 20452 20392
rect 2667 20264 2709 20273
rect 2667 20224 2668 20264
rect 2708 20224 2709 20264
rect 2667 20215 2709 20224
rect 6795 20264 6837 20273
rect 6795 20224 6796 20264
rect 6836 20224 6837 20264
rect 6795 20215 6837 20224
rect 8427 20264 8469 20273
rect 8427 20224 8428 20264
rect 8468 20224 8469 20264
rect 8427 20215 8469 20224
rect 10155 20264 10197 20273
rect 10155 20224 10156 20264
rect 10196 20224 10197 20264
rect 10155 20215 10197 20224
rect 12267 20264 12309 20273
rect 12267 20224 12268 20264
rect 12308 20224 12309 20264
rect 12267 20215 12309 20224
rect 16971 20180 17013 20189
rect 16971 20140 16972 20180
rect 17012 20140 17013 20180
rect 16971 20131 17013 20140
rect 20235 20180 20277 20189
rect 20235 20140 20236 20180
rect 20276 20140 20277 20180
rect 20235 20131 20277 20140
rect 1219 20096 1277 20097
rect 1219 20056 1228 20096
rect 1268 20056 1277 20096
rect 1219 20055 1277 20056
rect 2467 20096 2525 20097
rect 2467 20056 2476 20096
rect 2516 20056 2525 20096
rect 2467 20055 2525 20056
rect 3715 20096 3773 20097
rect 3715 20056 3724 20096
rect 3764 20056 3773 20096
rect 3715 20055 3773 20056
rect 4963 20096 5021 20097
rect 4963 20056 4972 20096
rect 5012 20056 5021 20096
rect 4963 20055 5021 20056
rect 5347 20096 5405 20097
rect 5347 20056 5356 20096
rect 5396 20056 5405 20096
rect 5347 20055 5405 20056
rect 6595 20096 6653 20097
rect 6595 20056 6604 20096
rect 6644 20056 6653 20096
rect 6595 20055 6653 20056
rect 6979 20096 7037 20097
rect 6979 20056 6988 20096
rect 7028 20056 7037 20096
rect 6979 20055 7037 20056
rect 8227 20096 8285 20097
rect 8227 20056 8236 20096
rect 8276 20056 8285 20096
rect 8227 20055 8285 20056
rect 8707 20096 8765 20097
rect 8707 20056 8716 20096
rect 8756 20056 8765 20096
rect 8707 20055 8765 20056
rect 9955 20096 10013 20097
rect 9955 20056 9964 20096
rect 10004 20056 10013 20096
rect 9955 20055 10013 20056
rect 10819 20096 10877 20097
rect 10819 20056 10828 20096
rect 10868 20056 10877 20096
rect 10819 20055 10877 20056
rect 12067 20096 12125 20097
rect 12067 20056 12076 20096
rect 12116 20056 12125 20096
rect 12067 20055 12125 20056
rect 12835 20096 12893 20097
rect 12835 20056 12844 20096
rect 12884 20056 12893 20096
rect 12835 20055 12893 20056
rect 14083 20096 14141 20097
rect 14083 20056 14092 20096
rect 14132 20056 14141 20096
rect 14083 20055 14141 20056
rect 14851 20096 14909 20097
rect 14851 20056 14860 20096
rect 14900 20056 14909 20096
rect 14851 20055 14909 20056
rect 16099 20096 16157 20097
rect 16099 20056 16108 20096
rect 16148 20056 16157 20096
rect 16099 20055 16157 20056
rect 16579 20096 16637 20097
rect 16579 20056 16588 20096
rect 16628 20056 16637 20096
rect 16579 20055 16637 20056
rect 16875 20096 16917 20105
rect 16875 20056 16876 20096
rect 16916 20056 16917 20096
rect 16875 20047 16917 20056
rect 17451 20096 17493 20105
rect 17451 20056 17452 20096
rect 17492 20056 17493 20096
rect 17451 20047 17493 20056
rect 17643 20096 17685 20105
rect 17643 20056 17644 20096
rect 17684 20056 17685 20096
rect 17643 20047 17685 20056
rect 17731 20096 17789 20097
rect 17731 20056 17740 20096
rect 17780 20056 17789 20096
rect 17731 20055 17789 20056
rect 17923 20096 17981 20097
rect 17923 20056 17932 20096
rect 17972 20056 17981 20096
rect 17923 20055 17981 20056
rect 18507 20096 18549 20105
rect 18507 20056 18508 20096
rect 18548 20056 18549 20096
rect 18507 20047 18549 20056
rect 18603 20096 18645 20105
rect 18603 20056 18604 20096
rect 18644 20056 18645 20096
rect 18603 20047 18645 20056
rect 18987 20096 19029 20105
rect 18987 20056 18988 20096
rect 19028 20056 19029 20096
rect 18987 20047 19029 20056
rect 19555 20096 19613 20097
rect 19555 20056 19564 20096
rect 19604 20056 19613 20096
rect 19555 20055 19613 20056
rect 20043 20082 20085 20091
rect 20043 20042 20044 20082
rect 20084 20042 20085 20082
rect 20043 20033 20085 20042
rect 19083 20012 19125 20021
rect 19083 19972 19084 20012
rect 19124 19972 19125 20012
rect 19083 19963 19125 19972
rect 17251 19928 17309 19929
rect 17251 19888 17260 19928
rect 17300 19888 17309 19928
rect 17251 19887 17309 19888
rect 5163 19844 5205 19853
rect 5163 19804 5164 19844
rect 5204 19804 5205 19844
rect 5163 19795 5205 19804
rect 14283 19844 14325 19853
rect 14283 19804 14284 19844
rect 14324 19804 14325 19844
rect 14283 19795 14325 19804
rect 16299 19844 16341 19853
rect 16299 19804 16300 19844
rect 16340 19804 16341 19844
rect 16299 19795 16341 19804
rect 17451 19844 17493 19853
rect 17451 19804 17452 19844
rect 17492 19804 17493 19844
rect 17451 19795 17493 19804
rect 18027 19844 18069 19853
rect 18027 19804 18028 19844
rect 18068 19804 18069 19844
rect 18027 19795 18069 19804
rect 1152 19676 20352 19700
rect 1152 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 20352 19676
rect 1152 19612 20352 19636
rect 2667 19508 2709 19517
rect 2667 19468 2668 19508
rect 2708 19468 2709 19508
rect 2667 19459 2709 19468
rect 16771 19508 16829 19509
rect 16771 19468 16780 19508
rect 16820 19468 16829 19508
rect 16771 19467 16829 19468
rect 18411 19508 18453 19517
rect 18411 19468 18412 19508
rect 18452 19468 18453 19508
rect 18411 19459 18453 19468
rect 20043 19508 20085 19517
rect 20043 19468 20044 19508
rect 20084 19468 20085 19508
rect 20043 19459 20085 19468
rect 4491 19270 4533 19279
rect 1219 19256 1277 19257
rect 1219 19216 1228 19256
rect 1268 19216 1277 19256
rect 1219 19215 1277 19216
rect 2467 19256 2525 19257
rect 2467 19216 2476 19256
rect 2516 19216 2525 19256
rect 2467 19215 2525 19216
rect 2955 19256 2997 19265
rect 2955 19216 2956 19256
rect 2996 19216 2997 19256
rect 2955 19207 2997 19216
rect 3051 19256 3093 19265
rect 3051 19216 3052 19256
rect 3092 19216 3093 19256
rect 3051 19207 3093 19216
rect 3435 19256 3477 19265
rect 3435 19216 3436 19256
rect 3476 19216 3477 19256
rect 3435 19207 3477 19216
rect 3531 19256 3573 19265
rect 3531 19216 3532 19256
rect 3572 19216 3573 19256
rect 3531 19207 3573 19216
rect 4003 19256 4061 19257
rect 4003 19216 4012 19256
rect 4052 19216 4061 19256
rect 4491 19230 4492 19270
rect 4532 19230 4533 19270
rect 4491 19221 4533 19230
rect 5347 19256 5405 19257
rect 4003 19215 4061 19216
rect 5347 19216 5356 19256
rect 5396 19216 5405 19256
rect 5347 19215 5405 19216
rect 6595 19256 6653 19257
rect 6595 19216 6604 19256
rect 6644 19216 6653 19256
rect 6595 19215 6653 19216
rect 6979 19256 7037 19257
rect 6979 19216 6988 19256
rect 7028 19216 7037 19256
rect 6979 19215 7037 19216
rect 8227 19256 8285 19257
rect 8227 19216 8236 19256
rect 8276 19216 8285 19256
rect 8227 19215 8285 19216
rect 8715 19256 8757 19265
rect 8715 19216 8716 19256
rect 8756 19216 8757 19256
rect 8715 19207 8757 19216
rect 8811 19256 8853 19265
rect 8811 19216 8812 19256
rect 8852 19216 8853 19256
rect 8811 19207 8853 19216
rect 9195 19256 9237 19265
rect 9195 19216 9196 19256
rect 9236 19216 9237 19256
rect 9195 19207 9237 19216
rect 9291 19256 9333 19265
rect 10251 19261 10293 19270
rect 14139 19265 14181 19274
rect 9291 19216 9292 19256
rect 9332 19216 9333 19256
rect 9291 19207 9333 19216
rect 9763 19256 9821 19257
rect 9763 19216 9772 19256
rect 9812 19216 9821 19256
rect 9763 19215 9821 19216
rect 10251 19221 10252 19261
rect 10292 19221 10293 19261
rect 10251 19212 10293 19221
rect 10819 19256 10877 19257
rect 10819 19216 10828 19256
rect 10868 19216 10877 19256
rect 10819 19215 10877 19216
rect 12067 19256 12125 19257
rect 12067 19216 12076 19256
rect 12116 19216 12125 19256
rect 12067 19215 12125 19216
rect 12555 19256 12597 19265
rect 12555 19216 12556 19256
rect 12596 19216 12597 19256
rect 12555 19207 12597 19216
rect 12651 19256 12693 19265
rect 12651 19216 12652 19256
rect 12692 19216 12693 19256
rect 12651 19207 12693 19216
rect 13035 19256 13077 19265
rect 13035 19216 13036 19256
rect 13076 19216 13077 19256
rect 13035 19207 13077 19216
rect 13131 19256 13173 19265
rect 13131 19216 13132 19256
rect 13172 19216 13173 19256
rect 13131 19207 13173 19216
rect 13603 19256 13661 19257
rect 13603 19216 13612 19256
rect 13652 19216 13661 19256
rect 14139 19225 14140 19265
rect 14180 19225 14181 19265
rect 14139 19216 14181 19225
rect 14667 19256 14709 19265
rect 14667 19216 14668 19256
rect 14708 19216 14709 19256
rect 13603 19215 13661 19216
rect 14667 19207 14709 19216
rect 14859 19256 14901 19265
rect 14859 19216 14860 19256
rect 14900 19216 14901 19256
rect 14859 19207 14901 19216
rect 15043 19256 15101 19257
rect 15043 19216 15052 19256
rect 15092 19216 15101 19256
rect 15043 19215 15101 19216
rect 15147 19256 15189 19265
rect 15147 19216 15148 19256
rect 15188 19216 15189 19256
rect 15147 19207 15189 19216
rect 15339 19256 15381 19265
rect 15339 19216 15340 19256
rect 15380 19216 15381 19256
rect 15339 19207 15381 19216
rect 15627 19256 15669 19265
rect 15627 19216 15628 19256
rect 15668 19216 15669 19256
rect 15627 19207 15669 19216
rect 15723 19256 15765 19265
rect 15723 19216 15724 19256
rect 15764 19216 15765 19256
rect 15723 19207 15765 19216
rect 15819 19256 15861 19265
rect 15819 19216 15820 19256
rect 15860 19216 15861 19256
rect 15819 19207 15861 19216
rect 16099 19256 16157 19257
rect 16099 19216 16108 19256
rect 16148 19216 16157 19256
rect 16099 19215 16157 19216
rect 16395 19256 16437 19265
rect 16395 19216 16396 19256
rect 16436 19216 16437 19256
rect 16395 19207 16437 19216
rect 16491 19256 16533 19265
rect 16491 19216 16492 19256
rect 16532 19216 16533 19256
rect 16491 19207 16533 19216
rect 16963 19256 17021 19257
rect 16963 19216 16972 19256
rect 17012 19216 17021 19256
rect 16963 19215 17021 19216
rect 18211 19256 18269 19257
rect 18211 19216 18220 19256
rect 18260 19216 18269 19256
rect 18211 19215 18269 19216
rect 18595 19256 18653 19257
rect 18595 19216 18604 19256
rect 18644 19216 18653 19256
rect 18595 19215 18653 19216
rect 19843 19256 19901 19257
rect 19843 19216 19852 19256
rect 19892 19216 19901 19256
rect 19843 19215 19901 19216
rect 8427 19172 8469 19181
rect 8427 19132 8428 19172
rect 8468 19132 8469 19172
rect 8427 19123 8469 19132
rect 12267 19172 12309 19181
rect 12267 19132 12268 19172
rect 12308 19132 12309 19172
rect 12267 19123 12309 19132
rect 4683 19088 4725 19097
rect 4683 19048 4684 19088
rect 4724 19048 4725 19088
rect 4683 19039 4725 19048
rect 6795 19088 6837 19097
rect 6795 19048 6796 19088
rect 6836 19048 6837 19088
rect 14283 19088 14325 19097
rect 6795 19039 6837 19048
rect 10443 19046 10485 19055
rect 10443 19006 10444 19046
rect 10484 19006 10485 19046
rect 14283 19048 14284 19088
rect 14324 19048 14325 19088
rect 14283 19039 14325 19048
rect 14763 19088 14805 19097
rect 14763 19048 14764 19088
rect 14804 19048 14805 19088
rect 14763 19039 14805 19048
rect 15235 19088 15293 19089
rect 15235 19048 15244 19088
rect 15284 19048 15293 19088
rect 15235 19047 15293 19048
rect 15523 19088 15581 19089
rect 15523 19048 15532 19088
rect 15572 19048 15581 19088
rect 15523 19047 15581 19048
rect 10443 18997 10485 19006
rect 1152 18920 20452 18944
rect 1152 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20452 18920
rect 1152 18856 20452 18880
rect 10539 18752 10581 18761
rect 10539 18712 10540 18752
rect 10580 18712 10581 18752
rect 10539 18703 10581 18712
rect 16491 18752 16533 18761
rect 16491 18712 16492 18752
rect 16532 18712 16533 18752
rect 16491 18703 16533 18712
rect 17443 18752 17501 18753
rect 17443 18712 17452 18752
rect 17492 18712 17501 18752
rect 17443 18711 17501 18712
rect 17739 18752 17781 18761
rect 17739 18712 17740 18752
rect 17780 18712 17781 18752
rect 17739 18703 17781 18712
rect 20235 18752 20277 18761
rect 20235 18712 20236 18752
rect 20276 18712 20277 18752
rect 20235 18703 20277 18712
rect 2475 18668 2517 18677
rect 2475 18628 2476 18668
rect 2516 18628 2517 18668
rect 2475 18619 2517 18628
rect 7371 18668 7413 18677
rect 7371 18628 7372 18668
rect 7412 18628 7413 18668
rect 7371 18619 7413 18628
rect 12459 18668 12501 18677
rect 12459 18628 12460 18668
rect 12500 18628 12501 18668
rect 12459 18619 12501 18628
rect 14475 18668 14517 18677
rect 14475 18628 14476 18668
rect 14516 18628 14517 18668
rect 14475 18619 14517 18628
rect 17163 18605 17205 18614
rect 3139 18584 3197 18585
rect 2667 18570 2709 18579
rect 2667 18530 2668 18570
rect 2708 18530 2709 18570
rect 3139 18544 3148 18584
rect 3188 18544 3197 18584
rect 3139 18543 3197 18544
rect 3627 18584 3669 18593
rect 3627 18544 3628 18584
rect 3668 18544 3669 18584
rect 3627 18535 3669 18544
rect 4107 18584 4149 18593
rect 4107 18544 4108 18584
rect 4148 18544 4149 18584
rect 4107 18535 4149 18544
rect 4203 18584 4245 18593
rect 4203 18544 4204 18584
rect 4244 18544 4245 18584
rect 4203 18535 4245 18544
rect 5643 18584 5685 18593
rect 5643 18544 5644 18584
rect 5684 18544 5685 18584
rect 5643 18535 5685 18544
rect 5739 18584 5781 18593
rect 5739 18544 5740 18584
rect 5780 18544 5781 18584
rect 5739 18535 5781 18544
rect 6691 18584 6749 18585
rect 6691 18544 6700 18584
rect 6740 18544 6749 18584
rect 6691 18543 6749 18544
rect 7179 18579 7221 18588
rect 7179 18539 7180 18579
rect 7220 18539 7221 18579
rect 9091 18584 9149 18585
rect 9091 18544 9100 18584
rect 9140 18544 9149 18584
rect 9091 18543 9149 18544
rect 10339 18584 10397 18585
rect 10339 18544 10348 18584
rect 10388 18544 10397 18584
rect 10339 18543 10397 18544
rect 11011 18584 11069 18585
rect 11011 18544 11020 18584
rect 11060 18544 11069 18584
rect 11011 18543 11069 18544
rect 12259 18584 12317 18585
rect 12259 18544 12268 18584
rect 12308 18544 12317 18584
rect 12259 18543 12317 18544
rect 12747 18584 12789 18593
rect 12747 18544 12748 18584
rect 12788 18544 12789 18584
rect 7179 18530 7221 18539
rect 12747 18535 12789 18544
rect 12843 18584 12885 18593
rect 12843 18544 12844 18584
rect 12884 18544 12885 18584
rect 12843 18535 12885 18544
rect 13795 18584 13853 18585
rect 13795 18544 13804 18584
rect 13844 18544 13853 18584
rect 15043 18584 15101 18585
rect 13795 18543 13853 18544
rect 14283 18570 14325 18579
rect 14283 18530 14284 18570
rect 14324 18530 14325 18570
rect 15043 18544 15052 18584
rect 15092 18544 15101 18584
rect 15043 18543 15101 18544
rect 16291 18584 16349 18585
rect 16291 18544 16300 18584
rect 16340 18544 16349 18584
rect 16291 18543 16349 18544
rect 16683 18584 16725 18593
rect 16683 18544 16684 18584
rect 16724 18544 16725 18584
rect 16683 18535 16725 18544
rect 16779 18584 16821 18593
rect 16779 18544 16780 18584
rect 16820 18544 16821 18584
rect 16779 18535 16821 18544
rect 16875 18584 16917 18593
rect 16875 18544 16876 18584
rect 16916 18544 16917 18584
rect 16875 18535 16917 18544
rect 16971 18584 17013 18593
rect 16971 18544 16972 18584
rect 17012 18544 17013 18584
rect 17163 18565 17164 18605
rect 17204 18565 17205 18605
rect 17163 18556 17205 18565
rect 17259 18584 17301 18593
rect 16971 18535 17013 18544
rect 17259 18544 17260 18584
rect 17300 18544 17301 18584
rect 17259 18535 17301 18544
rect 17355 18584 17397 18593
rect 17355 18544 17356 18584
rect 17396 18544 17397 18584
rect 17355 18535 17397 18544
rect 17635 18584 17693 18585
rect 17635 18544 17644 18584
rect 17684 18544 17693 18584
rect 17635 18543 17693 18544
rect 18411 18584 18453 18593
rect 18411 18544 18412 18584
rect 18452 18544 18453 18584
rect 18411 18535 18453 18544
rect 18603 18584 18645 18593
rect 18603 18544 18604 18584
rect 18644 18544 18645 18584
rect 18603 18535 18645 18544
rect 18787 18584 18845 18585
rect 18787 18544 18796 18584
rect 18836 18544 18845 18584
rect 18787 18543 18845 18544
rect 20035 18584 20093 18585
rect 20035 18544 20044 18584
rect 20084 18544 20093 18584
rect 20035 18543 20093 18544
rect 2667 18521 2709 18530
rect 14283 18521 14325 18530
rect 3723 18500 3765 18509
rect 3723 18460 3724 18500
rect 3764 18460 3765 18500
rect 3723 18451 3765 18460
rect 6123 18500 6165 18509
rect 6123 18460 6124 18500
rect 6164 18460 6165 18500
rect 6123 18451 6165 18460
rect 6219 18500 6261 18509
rect 6219 18460 6220 18500
rect 6260 18460 6261 18500
rect 6219 18451 6261 18460
rect 13227 18500 13269 18509
rect 13227 18460 13228 18500
rect 13268 18460 13269 18500
rect 13227 18451 13269 18460
rect 13323 18500 13365 18509
rect 13323 18460 13324 18500
rect 13364 18460 13365 18500
rect 13323 18451 13365 18460
rect 18507 18500 18549 18509
rect 18507 18460 18508 18500
rect 18548 18460 18549 18500
rect 18507 18451 18549 18460
rect 1152 18164 20352 18188
rect 1152 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 20352 18164
rect 1152 18100 20352 18124
rect 2667 17996 2709 18005
rect 2667 17956 2668 17996
rect 2708 17956 2709 17996
rect 2667 17947 2709 17956
rect 5835 17996 5877 18005
rect 5835 17956 5836 17996
rect 5876 17956 5877 17996
rect 5835 17947 5877 17956
rect 14859 17996 14901 18005
rect 14859 17956 14860 17996
rect 14900 17956 14901 17996
rect 14859 17947 14901 17956
rect 16875 17996 16917 18005
rect 16875 17956 16876 17996
rect 16916 17956 16917 17996
rect 16875 17947 16917 17956
rect 17643 17996 17685 18005
rect 17643 17956 17644 17996
rect 17684 17956 17685 17996
rect 17643 17947 17685 17956
rect 10395 17753 10437 17762
rect 1219 17744 1277 17745
rect 1219 17704 1228 17744
rect 1268 17704 1277 17744
rect 1219 17703 1277 17704
rect 2467 17744 2525 17745
rect 2467 17704 2476 17744
rect 2516 17704 2525 17744
rect 2467 17703 2525 17704
rect 4387 17744 4445 17745
rect 4387 17704 4396 17744
rect 4436 17704 4445 17744
rect 4387 17703 4445 17704
rect 5635 17744 5693 17745
rect 5635 17704 5644 17744
rect 5684 17704 5693 17744
rect 5635 17703 5693 17704
rect 7075 17744 7133 17745
rect 7075 17704 7084 17744
rect 7124 17704 7133 17744
rect 7075 17703 7133 17704
rect 8323 17744 8381 17745
rect 8323 17704 8332 17744
rect 8372 17704 8381 17744
rect 8323 17703 8381 17704
rect 8811 17744 8853 17753
rect 8811 17704 8812 17744
rect 8852 17704 8853 17744
rect 8811 17695 8853 17704
rect 8907 17744 8949 17753
rect 8907 17704 8908 17744
rect 8948 17704 8949 17744
rect 8907 17695 8949 17704
rect 9291 17744 9333 17753
rect 9291 17704 9292 17744
rect 9332 17704 9333 17744
rect 9291 17695 9333 17704
rect 9387 17744 9429 17753
rect 9387 17704 9388 17744
rect 9428 17704 9429 17744
rect 9387 17695 9429 17704
rect 9859 17744 9917 17745
rect 9859 17704 9868 17744
rect 9908 17704 9917 17744
rect 10395 17713 10396 17753
rect 10436 17713 10437 17753
rect 10395 17704 10437 17713
rect 13411 17744 13469 17745
rect 13411 17704 13420 17744
rect 13460 17704 13469 17744
rect 9859 17703 9917 17704
rect 13411 17703 13469 17704
rect 14659 17744 14717 17745
rect 14659 17704 14668 17744
rect 14708 17704 14717 17744
rect 14659 17703 14717 17704
rect 15427 17744 15485 17745
rect 15427 17704 15436 17744
rect 15476 17704 15485 17744
rect 15427 17703 15485 17704
rect 16675 17744 16733 17745
rect 16675 17704 16684 17744
rect 16724 17704 16733 17744
rect 16675 17703 16733 17704
rect 17731 17744 17789 17745
rect 17731 17704 17740 17744
rect 17780 17704 17789 17744
rect 17731 17703 17789 17704
rect 17923 17744 17981 17745
rect 17923 17704 17932 17744
rect 17972 17704 17981 17744
rect 17923 17703 17981 17704
rect 19171 17744 19229 17745
rect 19171 17704 19180 17744
rect 19220 17704 19229 17744
rect 19171 17703 19229 17704
rect 19563 17744 19605 17753
rect 19563 17704 19564 17744
rect 19604 17704 19605 17744
rect 19563 17695 19605 17704
rect 19659 17744 19701 17753
rect 19659 17704 19660 17744
rect 19700 17704 19701 17744
rect 19659 17695 19701 17704
rect 19755 17744 19797 17753
rect 19755 17704 19756 17744
rect 19796 17704 19797 17744
rect 19755 17695 19797 17704
rect 20043 17744 20085 17753
rect 20043 17704 20044 17744
rect 20084 17704 20085 17744
rect 20043 17695 20085 17704
rect 20131 17744 20189 17745
rect 20131 17704 20140 17744
rect 20180 17704 20189 17744
rect 20131 17703 20189 17704
rect 8523 17660 8565 17669
rect 8523 17620 8524 17660
rect 8564 17620 8565 17660
rect 8523 17611 8565 17620
rect 19371 17660 19413 17669
rect 19371 17620 19372 17660
rect 19412 17620 19413 17660
rect 19371 17611 19413 17620
rect 10539 17576 10581 17585
rect 10539 17536 10540 17576
rect 10580 17536 10581 17576
rect 10539 17527 10581 17536
rect 19843 17576 19901 17577
rect 19843 17536 19852 17576
rect 19892 17536 19901 17576
rect 19843 17535 19901 17536
rect 1152 17408 20452 17432
rect 1152 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20452 17408
rect 1152 17344 20452 17368
rect 10635 17240 10677 17249
rect 10635 17200 10636 17240
rect 10676 17200 10677 17240
rect 10635 17191 10677 17200
rect 18795 17240 18837 17249
rect 18795 17200 18796 17240
rect 18836 17200 18837 17240
rect 18795 17191 18837 17200
rect 20227 17240 20285 17241
rect 20227 17200 20236 17240
rect 20276 17200 20285 17240
rect 20227 17199 20285 17200
rect 2187 17156 2229 17165
rect 2187 17116 2188 17156
rect 2228 17116 2229 17156
rect 2187 17107 2229 17116
rect 6987 17156 7029 17165
rect 6987 17116 6988 17156
rect 7028 17116 7029 17156
rect 6987 17107 7029 17116
rect 19467 17156 19509 17165
rect 19467 17116 19468 17156
rect 19508 17116 19509 17156
rect 19467 17107 19509 17116
rect 2851 17072 2909 17073
rect 2379 17058 2421 17067
rect 2379 17018 2380 17058
rect 2420 17018 2421 17058
rect 2851 17032 2860 17072
rect 2900 17032 2909 17072
rect 3435 17072 3477 17081
rect 2851 17031 2909 17032
rect 2379 17009 2421 17018
rect 3339 17030 3381 17039
rect 3339 16990 3340 17030
rect 3380 16990 3381 17030
rect 3435 17032 3436 17072
rect 3476 17032 3477 17072
rect 3435 17023 3477 17032
rect 3819 17072 3861 17081
rect 3819 17032 3820 17072
rect 3860 17032 3861 17072
rect 3819 17023 3861 17032
rect 3915 17072 3957 17081
rect 3915 17032 3916 17072
rect 3956 17032 3957 17072
rect 3915 17023 3957 17032
rect 5259 17072 5301 17081
rect 5259 17032 5260 17072
rect 5300 17032 5301 17072
rect 5259 17023 5301 17032
rect 5355 17072 5397 17081
rect 5355 17032 5356 17072
rect 5396 17032 5397 17072
rect 5355 17023 5397 17032
rect 6307 17072 6365 17073
rect 6307 17032 6316 17072
rect 6356 17032 6365 17072
rect 7363 17072 7421 17073
rect 6307 17031 6365 17032
rect 6795 17058 6837 17067
rect 6795 17018 6796 17058
rect 6836 17018 6837 17058
rect 7363 17032 7372 17072
rect 7412 17032 7421 17072
rect 7363 17031 7421 17032
rect 8611 17072 8669 17073
rect 8611 17032 8620 17072
rect 8660 17032 8669 17072
rect 8611 17031 8669 17032
rect 9187 17072 9245 17073
rect 9187 17032 9196 17072
rect 9236 17032 9245 17072
rect 9187 17031 9245 17032
rect 10435 17072 10493 17073
rect 10435 17032 10444 17072
rect 10484 17032 10493 17072
rect 10435 17031 10493 17032
rect 11299 17072 11357 17073
rect 11299 17032 11308 17072
rect 11348 17032 11357 17072
rect 11299 17031 11357 17032
rect 12547 17072 12605 17073
rect 12547 17032 12556 17072
rect 12596 17032 12605 17072
rect 12547 17031 12605 17032
rect 13315 17072 13373 17073
rect 13315 17032 13324 17072
rect 13364 17032 13373 17072
rect 13315 17031 13373 17032
rect 14563 17072 14621 17073
rect 14563 17032 14572 17072
rect 14612 17032 14621 17072
rect 14563 17031 14621 17032
rect 15715 17072 15773 17073
rect 15715 17032 15724 17072
rect 15764 17032 15773 17072
rect 15715 17031 15773 17032
rect 16963 17072 17021 17073
rect 16963 17032 16972 17072
rect 17012 17032 17021 17072
rect 16963 17031 17021 17032
rect 17347 17072 17405 17073
rect 17347 17032 17356 17072
rect 17396 17032 17405 17072
rect 17347 17031 17405 17032
rect 18595 17072 18653 17073
rect 18595 17032 18604 17072
rect 18644 17032 18653 17072
rect 18595 17031 18653 17032
rect 19075 17072 19133 17073
rect 19075 17032 19084 17072
rect 19124 17032 19133 17072
rect 19075 17031 19133 17032
rect 19371 17072 19413 17081
rect 19371 17032 19372 17072
rect 19412 17032 19413 17072
rect 19371 17023 19413 17032
rect 19947 17072 19989 17081
rect 19947 17032 19948 17072
rect 19988 17032 19989 17072
rect 19947 17023 19989 17032
rect 20043 17072 20085 17081
rect 20043 17032 20044 17072
rect 20084 17032 20085 17072
rect 20043 17023 20085 17032
rect 20131 17030 20189 17031
rect 6795 17009 6837 17018
rect 3339 16981 3381 16990
rect 5739 16988 5781 16997
rect 5739 16948 5740 16988
rect 5780 16948 5781 16988
rect 5739 16939 5781 16948
rect 5835 16988 5877 16997
rect 20131 16990 20140 17030
rect 20180 16990 20189 17030
rect 20131 16989 20189 16990
rect 5835 16948 5836 16988
rect 5876 16948 5877 16988
rect 5835 16939 5877 16948
rect 7179 16820 7221 16829
rect 7179 16780 7180 16820
rect 7220 16780 7221 16820
rect 7179 16771 7221 16780
rect 12747 16820 12789 16829
rect 12747 16780 12748 16820
rect 12788 16780 12789 16820
rect 12747 16771 12789 16780
rect 14763 16820 14805 16829
rect 14763 16780 14764 16820
rect 14804 16780 14805 16820
rect 14763 16771 14805 16780
rect 17163 16820 17205 16829
rect 17163 16780 17164 16820
rect 17204 16780 17205 16820
rect 17163 16771 17205 16780
rect 19747 16820 19805 16821
rect 19747 16780 19756 16820
rect 19796 16780 19805 16820
rect 19747 16779 19805 16780
rect 1152 16652 20352 16676
rect 1152 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 20352 16652
rect 1152 16588 20352 16612
rect 19555 16400 19613 16401
rect 19555 16360 19564 16400
rect 19604 16360 19613 16400
rect 19555 16359 19613 16360
rect 1411 16316 1469 16317
rect 1411 16276 1420 16316
rect 1460 16276 1469 16316
rect 1411 16275 1469 16276
rect 3243 16316 3285 16325
rect 3243 16276 3244 16316
rect 3284 16276 3285 16316
rect 3243 16267 3285 16276
rect 6123 16316 6165 16325
rect 6123 16276 6124 16316
rect 6164 16276 6165 16316
rect 6123 16267 6165 16276
rect 6219 16316 6261 16325
rect 6219 16276 6220 16316
rect 6260 16276 6261 16316
rect 6219 16267 6261 16276
rect 10827 16316 10869 16325
rect 10827 16276 10828 16316
rect 10868 16276 10869 16316
rect 10827 16267 10869 16276
rect 17635 16316 17693 16317
rect 17635 16276 17644 16316
rect 17684 16276 17693 16316
rect 17635 16275 17693 16276
rect 4251 16241 4293 16250
rect 7227 16241 7269 16250
rect 9819 16241 9861 16250
rect 11835 16241 11877 16250
rect 14283 16246 14325 16255
rect 2667 16232 2709 16241
rect 2667 16192 2668 16232
rect 2708 16192 2709 16232
rect 2667 16183 2709 16192
rect 2763 16232 2805 16241
rect 2763 16192 2764 16232
rect 2804 16192 2805 16232
rect 2763 16183 2805 16192
rect 3147 16232 3189 16241
rect 3147 16192 3148 16232
rect 3188 16192 3189 16232
rect 3147 16183 3189 16192
rect 3715 16232 3773 16233
rect 3715 16192 3724 16232
rect 3764 16192 3773 16232
rect 4251 16201 4252 16241
rect 4292 16201 4293 16241
rect 4251 16192 4293 16201
rect 5643 16232 5685 16241
rect 5643 16192 5644 16232
rect 5684 16192 5685 16232
rect 3715 16191 3773 16192
rect 5643 16183 5685 16192
rect 5739 16232 5781 16241
rect 5739 16192 5740 16232
rect 5780 16192 5781 16232
rect 5739 16183 5781 16192
rect 6691 16232 6749 16233
rect 6691 16192 6700 16232
rect 6740 16192 6749 16232
rect 7227 16201 7228 16241
rect 7268 16201 7269 16241
rect 7227 16192 7269 16201
rect 8235 16232 8277 16241
rect 8235 16192 8236 16232
rect 8276 16192 8277 16232
rect 6691 16191 6749 16192
rect 8235 16183 8277 16192
rect 8331 16232 8373 16241
rect 8331 16192 8332 16232
rect 8372 16192 8373 16232
rect 8331 16183 8373 16192
rect 8715 16232 8757 16241
rect 8715 16192 8716 16232
rect 8756 16192 8757 16232
rect 8715 16183 8757 16192
rect 8811 16232 8853 16241
rect 8811 16192 8812 16232
rect 8852 16192 8853 16232
rect 8811 16183 8853 16192
rect 9283 16232 9341 16233
rect 9283 16192 9292 16232
rect 9332 16192 9341 16232
rect 9819 16201 9820 16241
rect 9860 16201 9861 16241
rect 9819 16192 9861 16201
rect 10251 16232 10293 16241
rect 10251 16192 10252 16232
rect 10292 16192 10293 16232
rect 9283 16191 9341 16192
rect 10251 16183 10293 16192
rect 10347 16232 10389 16241
rect 10347 16192 10348 16232
rect 10388 16192 10389 16232
rect 10347 16183 10389 16192
rect 10731 16232 10773 16241
rect 10731 16192 10732 16232
rect 10772 16192 10773 16232
rect 10731 16183 10773 16192
rect 11299 16232 11357 16233
rect 11299 16192 11308 16232
rect 11348 16192 11357 16232
rect 11835 16201 11836 16241
rect 11876 16201 11877 16241
rect 11835 16192 11877 16201
rect 12747 16232 12789 16241
rect 12747 16192 12748 16232
rect 12788 16192 12789 16232
rect 11299 16191 11357 16192
rect 12747 16183 12789 16192
rect 12843 16232 12885 16241
rect 12843 16192 12844 16232
rect 12884 16192 12885 16232
rect 12843 16183 12885 16192
rect 13227 16232 13269 16241
rect 13227 16192 13228 16232
rect 13268 16192 13269 16232
rect 13227 16183 13269 16192
rect 13323 16232 13365 16241
rect 13323 16192 13324 16232
rect 13364 16192 13365 16232
rect 13323 16183 13365 16192
rect 13795 16232 13853 16233
rect 13795 16192 13804 16232
rect 13844 16192 13853 16232
rect 14283 16206 14284 16246
rect 14324 16206 14325 16246
rect 17067 16246 17109 16255
rect 14283 16197 14325 16206
rect 15531 16232 15573 16241
rect 13795 16191 13853 16192
rect 15531 16192 15532 16232
rect 15572 16192 15573 16232
rect 15531 16183 15573 16192
rect 15627 16232 15669 16241
rect 15627 16192 15628 16232
rect 15668 16192 15669 16232
rect 15627 16183 15669 16192
rect 16011 16232 16053 16241
rect 16011 16192 16012 16232
rect 16052 16192 16053 16232
rect 16011 16183 16053 16192
rect 16107 16232 16149 16241
rect 16107 16192 16108 16232
rect 16148 16192 16149 16232
rect 16107 16183 16149 16192
rect 16579 16232 16637 16233
rect 16579 16192 16588 16232
rect 16628 16192 16637 16232
rect 17067 16206 17068 16246
rect 17108 16206 17109 16246
rect 17067 16197 17109 16206
rect 17827 16232 17885 16233
rect 16579 16191 16637 16192
rect 17827 16192 17836 16232
rect 17876 16192 17885 16232
rect 17827 16191 17885 16192
rect 17931 16232 17973 16241
rect 17931 16192 17932 16232
rect 17972 16192 17973 16232
rect 17931 16183 17973 16192
rect 18123 16232 18165 16241
rect 18123 16192 18124 16232
rect 18164 16192 18165 16232
rect 18123 16183 18165 16192
rect 18315 16232 18357 16241
rect 18315 16192 18316 16232
rect 18356 16192 18357 16232
rect 18315 16183 18357 16192
rect 18411 16232 18453 16241
rect 18411 16192 18412 16232
rect 18452 16192 18453 16232
rect 18411 16183 18453 16192
rect 18507 16232 18549 16241
rect 18507 16192 18508 16232
rect 18548 16192 18549 16232
rect 18507 16183 18549 16192
rect 18603 16232 18645 16241
rect 18603 16192 18604 16232
rect 18644 16192 18645 16232
rect 18603 16183 18645 16192
rect 18883 16232 18941 16233
rect 18883 16192 18892 16232
rect 18932 16192 18941 16232
rect 18883 16191 18941 16192
rect 19179 16232 19221 16241
rect 19179 16192 19180 16232
rect 19220 16192 19221 16232
rect 19179 16183 19221 16192
rect 19755 16232 19797 16241
rect 19755 16192 19756 16232
rect 19796 16192 19797 16232
rect 19755 16183 19797 16192
rect 19851 16232 19893 16241
rect 19851 16192 19852 16232
rect 19892 16192 19893 16232
rect 19851 16183 19893 16192
rect 19947 16232 19989 16241
rect 19947 16192 19948 16232
rect 19988 16192 19989 16232
rect 19947 16183 19989 16192
rect 9963 16148 10005 16157
rect 9963 16108 9964 16148
rect 10004 16108 10005 16148
rect 9963 16099 10005 16108
rect 17259 16148 17301 16157
rect 17259 16108 17260 16148
rect 17300 16108 17301 16148
rect 17259 16099 17301 16108
rect 19275 16148 19317 16157
rect 19275 16108 19276 16148
rect 19316 16108 19317 16148
rect 19275 16099 19317 16108
rect 1227 16064 1269 16073
rect 1227 16024 1228 16064
rect 1268 16024 1269 16064
rect 1227 16015 1269 16024
rect 4395 16064 4437 16073
rect 4395 16024 4396 16064
rect 4436 16024 4437 16064
rect 4395 16015 4437 16024
rect 7371 16064 7413 16073
rect 7371 16024 7372 16064
rect 7412 16024 7413 16064
rect 7371 16015 7413 16024
rect 11979 16064 12021 16073
rect 11979 16024 11980 16064
rect 12020 16024 12021 16064
rect 11979 16015 12021 16024
rect 14475 16064 14517 16073
rect 14475 16024 14476 16064
rect 14516 16024 14517 16064
rect 14475 16015 14517 16024
rect 17451 16064 17493 16073
rect 17451 16024 17452 16064
rect 17492 16024 17493 16064
rect 17451 16015 17493 16024
rect 18019 16064 18077 16065
rect 18019 16024 18028 16064
rect 18068 16024 18077 16064
rect 18019 16023 18077 16024
rect 20035 16064 20093 16065
rect 20035 16024 20044 16064
rect 20084 16024 20093 16064
rect 20035 16023 20093 16024
rect 1152 15896 20452 15920
rect 1152 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20452 15896
rect 1152 15832 20452 15856
rect 2667 15728 2709 15737
rect 2667 15688 2668 15728
rect 2708 15688 2709 15728
rect 2667 15679 2709 15688
rect 5163 15728 5205 15737
rect 5163 15688 5164 15728
rect 5204 15688 5205 15728
rect 5163 15679 5205 15688
rect 6795 15728 6837 15737
rect 6795 15688 6796 15728
rect 6836 15688 6837 15728
rect 6795 15679 6837 15688
rect 8427 15728 8469 15737
rect 8427 15688 8428 15728
rect 8468 15688 8469 15728
rect 8427 15679 8469 15688
rect 10251 15728 10293 15737
rect 10251 15688 10252 15728
rect 10292 15688 10293 15728
rect 10251 15679 10293 15688
rect 12459 15644 12501 15653
rect 12459 15604 12460 15644
rect 12500 15604 12501 15644
rect 12459 15595 12501 15604
rect 14475 15644 14517 15653
rect 14475 15604 14476 15644
rect 14516 15604 14517 15644
rect 14475 15595 14517 15604
rect 16107 15644 16149 15653
rect 16107 15604 16108 15644
rect 16148 15604 16149 15644
rect 16107 15595 16149 15604
rect 19563 15644 19605 15653
rect 19563 15604 19564 15644
rect 19604 15604 19605 15644
rect 19563 15595 19605 15604
rect 1219 15560 1277 15561
rect 1219 15520 1228 15560
rect 1268 15520 1277 15560
rect 1219 15519 1277 15520
rect 2467 15560 2525 15561
rect 2467 15520 2476 15560
rect 2516 15520 2525 15560
rect 2467 15519 2525 15520
rect 3715 15560 3773 15561
rect 3715 15520 3724 15560
rect 3764 15520 3773 15560
rect 3715 15519 3773 15520
rect 4963 15560 5021 15561
rect 4963 15520 4972 15560
rect 5012 15520 5021 15560
rect 4963 15519 5021 15520
rect 5347 15560 5405 15561
rect 5347 15520 5356 15560
rect 5396 15520 5405 15560
rect 5347 15519 5405 15520
rect 6595 15560 6653 15561
rect 6595 15520 6604 15560
rect 6644 15520 6653 15560
rect 6595 15519 6653 15520
rect 8227 15560 8285 15561
rect 8227 15520 8236 15560
rect 8276 15520 8285 15560
rect 8227 15519 8285 15520
rect 8803 15560 8861 15561
rect 8803 15520 8812 15560
rect 8852 15520 8861 15560
rect 8803 15519 8861 15520
rect 10051 15560 10109 15561
rect 10051 15520 10060 15560
rect 10100 15520 10109 15560
rect 10051 15519 10109 15520
rect 11011 15560 11069 15561
rect 11011 15520 11020 15560
rect 11060 15520 11069 15560
rect 11011 15519 11069 15520
rect 12259 15560 12317 15561
rect 12259 15520 12268 15560
rect 12308 15520 12317 15560
rect 12259 15519 12317 15520
rect 12747 15560 12789 15569
rect 12747 15520 12748 15560
rect 12788 15520 12789 15560
rect 6979 15518 7037 15519
rect 6979 15478 6988 15518
rect 7028 15478 7037 15518
rect 12747 15511 12789 15520
rect 12843 15560 12885 15569
rect 12843 15520 12844 15560
rect 12884 15520 12885 15560
rect 12843 15511 12885 15520
rect 13227 15560 13269 15569
rect 13227 15520 13228 15560
rect 13268 15520 13269 15560
rect 13227 15511 13269 15520
rect 13795 15560 13853 15561
rect 13795 15520 13804 15560
rect 13844 15520 13853 15560
rect 14659 15560 14717 15561
rect 13795 15519 13853 15520
rect 14331 15550 14373 15559
rect 14331 15510 14332 15550
rect 14372 15510 14373 15550
rect 14659 15520 14668 15560
rect 14708 15520 14717 15560
rect 14659 15519 14717 15520
rect 15907 15560 15965 15561
rect 15907 15520 15916 15560
rect 15956 15520 15965 15560
rect 15907 15519 15965 15520
rect 16483 15560 16541 15561
rect 16483 15520 16492 15560
rect 16532 15520 16541 15560
rect 16483 15519 16541 15520
rect 17731 15560 17789 15561
rect 17731 15520 17740 15560
rect 17780 15520 17789 15560
rect 17731 15519 17789 15520
rect 18115 15560 18173 15561
rect 18115 15520 18124 15560
rect 18164 15520 18173 15560
rect 18115 15519 18173 15520
rect 19363 15560 19421 15561
rect 19363 15520 19372 15560
rect 19412 15520 19421 15560
rect 19363 15519 19421 15520
rect 19747 15560 19805 15561
rect 19747 15520 19756 15560
rect 19796 15520 19805 15560
rect 19747 15519 19805 15520
rect 19851 15560 19893 15569
rect 19851 15520 19852 15560
rect 19892 15520 19893 15560
rect 19851 15511 19893 15520
rect 20043 15560 20085 15569
rect 20043 15520 20044 15560
rect 20084 15520 20085 15560
rect 20043 15511 20085 15520
rect 14331 15501 14373 15510
rect 6979 15477 7037 15478
rect 3043 15476 3101 15477
rect 3043 15436 3052 15476
rect 3092 15436 3101 15476
rect 3043 15435 3101 15436
rect 13323 15476 13365 15485
rect 13323 15436 13324 15476
rect 13364 15436 13365 15476
rect 13323 15427 13365 15436
rect 2859 15392 2901 15401
rect 2859 15352 2860 15392
rect 2900 15352 2901 15392
rect 2859 15343 2901 15352
rect 20043 15392 20085 15401
rect 20043 15352 20044 15392
rect 20084 15352 20085 15392
rect 20043 15343 20085 15352
rect 16299 15308 16341 15317
rect 16299 15268 16300 15308
rect 16340 15268 16341 15308
rect 16299 15259 16341 15268
rect 1152 15140 20352 15164
rect 1152 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 20352 15140
rect 1152 15076 20352 15100
rect 3435 14972 3477 14981
rect 3435 14932 3436 14972
rect 3476 14932 3477 14972
rect 3435 14923 3477 14932
rect 5643 14972 5685 14981
rect 5643 14932 5644 14972
rect 5684 14932 5685 14972
rect 5643 14923 5685 14932
rect 7467 14972 7509 14981
rect 7467 14932 7468 14972
rect 7508 14932 7509 14972
rect 7467 14923 7509 14932
rect 9867 14972 9909 14981
rect 9867 14932 9868 14972
rect 9908 14932 9909 14972
rect 9867 14923 9909 14932
rect 11979 14972 12021 14981
rect 11979 14932 11980 14972
rect 12020 14932 12021 14972
rect 11979 14923 12021 14932
rect 14571 14972 14613 14981
rect 14571 14932 14572 14972
rect 14612 14932 14613 14972
rect 14571 14923 14613 14932
rect 19179 14972 19221 14981
rect 19179 14932 19180 14972
rect 19220 14932 19221 14972
rect 19179 14923 19221 14932
rect 19659 14972 19701 14981
rect 19659 14932 19660 14972
rect 19700 14932 19701 14972
rect 19659 14923 19701 14932
rect 1699 14804 1757 14805
rect 1699 14764 1708 14804
rect 1748 14764 1757 14804
rect 1699 14763 1757 14764
rect 3811 14804 3869 14805
rect 3811 14764 3820 14804
rect 3860 14764 3869 14804
rect 3811 14763 3869 14764
rect 15627 14804 15669 14813
rect 15627 14764 15628 14804
rect 15668 14764 15669 14804
rect 15627 14755 15669 14764
rect 15723 14804 15765 14813
rect 15723 14764 15724 14804
rect 15764 14764 15765 14804
rect 15723 14755 15765 14764
rect 17251 14804 17309 14805
rect 17251 14764 17260 14804
rect 17300 14764 17309 14804
rect 17251 14763 17309 14764
rect 16683 14734 16725 14743
rect 1987 14720 2045 14721
rect 1987 14680 1996 14720
rect 2036 14680 2045 14720
rect 1987 14679 2045 14680
rect 3235 14720 3293 14721
rect 3235 14680 3244 14720
rect 3284 14680 3293 14720
rect 3235 14679 3293 14680
rect 4195 14720 4253 14721
rect 4195 14680 4204 14720
rect 4244 14680 4253 14720
rect 4195 14679 4253 14680
rect 5443 14720 5501 14721
rect 5443 14680 5452 14720
rect 5492 14680 5501 14720
rect 5443 14679 5501 14680
rect 6019 14720 6077 14721
rect 6019 14680 6028 14720
rect 6068 14680 6077 14720
rect 6019 14679 6077 14680
rect 7267 14720 7325 14721
rect 7267 14680 7276 14720
rect 7316 14680 7325 14720
rect 7267 14679 7325 14680
rect 8419 14720 8477 14721
rect 8419 14680 8428 14720
rect 8468 14680 8477 14720
rect 8419 14679 8477 14680
rect 9667 14720 9725 14721
rect 9667 14680 9676 14720
rect 9716 14680 9725 14720
rect 9667 14679 9725 14680
rect 10531 14720 10589 14721
rect 10531 14680 10540 14720
rect 10580 14680 10589 14720
rect 10531 14679 10589 14680
rect 11779 14720 11837 14721
rect 11779 14680 11788 14720
rect 11828 14680 11837 14720
rect 11779 14679 11837 14680
rect 13123 14720 13181 14721
rect 13123 14680 13132 14720
rect 13172 14680 13181 14720
rect 13123 14679 13181 14680
rect 14371 14720 14429 14721
rect 14371 14680 14380 14720
rect 14420 14680 14429 14720
rect 14371 14679 14429 14680
rect 15147 14720 15189 14729
rect 15147 14680 15148 14720
rect 15188 14680 15189 14720
rect 15147 14671 15189 14680
rect 15243 14720 15285 14729
rect 15243 14680 15244 14720
rect 15284 14680 15285 14720
rect 15243 14671 15285 14680
rect 16195 14720 16253 14721
rect 16195 14680 16204 14720
rect 16244 14680 16253 14720
rect 16683 14694 16684 14734
rect 16724 14694 16725 14734
rect 16683 14685 16725 14694
rect 17539 14720 17597 14721
rect 16195 14679 16253 14680
rect 17539 14680 17548 14720
rect 17588 14680 17597 14720
rect 17539 14679 17597 14680
rect 18787 14720 18845 14721
rect 18787 14680 18796 14720
rect 18836 14680 18845 14720
rect 18787 14679 18845 14680
rect 19179 14720 19221 14729
rect 19179 14680 19180 14720
rect 19220 14680 19221 14720
rect 19179 14671 19221 14680
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19371 14671 19413 14680
rect 19459 14720 19517 14721
rect 19459 14680 19468 14720
rect 19508 14680 19517 14720
rect 19459 14679 19517 14680
rect 19747 14720 19805 14721
rect 19747 14680 19756 14720
rect 19796 14680 19805 14720
rect 19747 14679 19805 14680
rect 16875 14636 16917 14645
rect 16875 14596 16876 14636
rect 16916 14596 16917 14636
rect 16875 14587 16917 14596
rect 1515 14552 1557 14561
rect 1515 14512 1516 14552
rect 1556 14512 1557 14552
rect 1515 14503 1557 14512
rect 3627 14552 3669 14561
rect 3627 14512 3628 14552
rect 3668 14512 3669 14552
rect 3627 14503 3669 14512
rect 17067 14552 17109 14561
rect 17067 14512 17068 14552
rect 17108 14512 17109 14552
rect 17067 14503 17109 14512
rect 18987 14552 19029 14561
rect 18987 14512 18988 14552
rect 19028 14512 19029 14552
rect 18987 14503 19029 14512
rect 1152 14384 20452 14408
rect 1152 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20452 14384
rect 1152 14320 20452 14344
rect 2667 14216 2709 14225
rect 2667 14176 2668 14216
rect 2708 14176 2709 14216
rect 2667 14167 2709 14176
rect 7947 14216 7989 14225
rect 7947 14176 7948 14216
rect 7988 14176 7989 14216
rect 7947 14167 7989 14176
rect 15147 14216 15189 14225
rect 15147 14176 15148 14216
rect 15188 14176 15189 14216
rect 15147 14167 15189 14176
rect 20139 14216 20181 14225
rect 20139 14176 20140 14216
rect 20180 14176 20181 14216
rect 20139 14167 20181 14176
rect 4683 14132 4725 14141
rect 4683 14092 4684 14132
rect 4724 14092 4725 14132
rect 4683 14083 4725 14092
rect 10347 14132 10389 14141
rect 10347 14092 10348 14132
rect 10388 14092 10389 14132
rect 10347 14083 10389 14092
rect 12939 14132 12981 14141
rect 12939 14092 12940 14132
rect 12980 14092 12981 14132
rect 12939 14083 12981 14092
rect 14955 14132 14997 14141
rect 14955 14092 14956 14132
rect 14996 14092 14997 14132
rect 14955 14083 14997 14092
rect 1219 14048 1277 14049
rect 1219 14008 1228 14048
rect 1268 14008 1277 14048
rect 1219 14007 1277 14008
rect 2467 14048 2525 14049
rect 2467 14008 2476 14048
rect 2516 14008 2525 14048
rect 2467 14007 2525 14008
rect 2955 14048 2997 14057
rect 2955 14008 2956 14048
rect 2996 14008 2997 14048
rect 2955 13999 2997 14008
rect 3051 14048 3093 14057
rect 3051 14008 3052 14048
rect 3092 14008 3093 14048
rect 3051 13999 3093 14008
rect 3435 14048 3477 14057
rect 3435 14008 3436 14048
rect 3476 14008 3477 14048
rect 3435 13999 3477 14008
rect 3531 14048 3573 14057
rect 3531 14008 3532 14048
rect 3572 14008 3573 14048
rect 3531 13999 3573 14008
rect 4003 14048 4061 14049
rect 4003 14008 4012 14048
rect 4052 14008 4061 14048
rect 6219 14048 6261 14057
rect 4003 14007 4061 14008
rect 4491 14034 4533 14043
rect 4491 13994 4492 14034
rect 4532 13994 4533 14034
rect 6219 14008 6220 14048
rect 6260 14008 6261 14048
rect 6219 13999 6261 14008
rect 6315 14048 6357 14057
rect 6315 14008 6316 14048
rect 6356 14008 6357 14048
rect 6315 13999 6357 14008
rect 6699 14048 6741 14057
rect 6699 14008 6700 14048
rect 6740 14008 6741 14048
rect 6699 13999 6741 14008
rect 6795 14048 6837 14057
rect 6795 14008 6796 14048
rect 6836 14008 6837 14048
rect 6795 13999 6837 14008
rect 7267 14048 7325 14049
rect 7267 14008 7276 14048
rect 7316 14008 7325 14048
rect 8619 14048 8661 14057
rect 7267 14007 7325 14008
rect 7755 14034 7797 14043
rect 4491 13985 4533 13994
rect 7755 13994 7756 14034
rect 7796 13994 7797 14034
rect 8619 14008 8620 14048
rect 8660 14008 8661 14048
rect 8619 13999 8661 14008
rect 8715 14048 8757 14057
rect 8715 14008 8716 14048
rect 8756 14008 8757 14048
rect 8715 13999 8757 14008
rect 9099 14048 9141 14057
rect 9099 14008 9100 14048
rect 9140 14008 9141 14048
rect 9099 13999 9141 14008
rect 9195 14048 9237 14057
rect 9195 14008 9196 14048
rect 9236 14008 9237 14048
rect 9195 13999 9237 14008
rect 9667 14048 9725 14049
rect 9667 14008 9676 14048
rect 9716 14008 9725 14048
rect 11211 14048 11253 14057
rect 9667 14007 9725 14008
rect 10155 14034 10197 14043
rect 7755 13985 7797 13994
rect 10155 13994 10156 14034
rect 10196 13994 10197 14034
rect 11211 14008 11212 14048
rect 11252 14008 11253 14048
rect 11211 13999 11253 14008
rect 11307 14048 11349 14057
rect 11307 14008 11308 14048
rect 11348 14008 11349 14048
rect 11307 13999 11349 14008
rect 11787 14048 11829 14057
rect 11787 14008 11788 14048
rect 11828 14008 11829 14048
rect 11787 13999 11829 14008
rect 12259 14048 12317 14049
rect 12259 14008 12268 14048
rect 12308 14008 12317 14048
rect 13227 14048 13269 14057
rect 12259 14007 12317 14008
rect 12747 14034 12789 14043
rect 10155 13985 10197 13994
rect 12747 13994 12748 14034
rect 12788 13994 12789 14034
rect 13227 14008 13228 14048
rect 13268 14008 13269 14048
rect 13227 13999 13269 14008
rect 13323 14048 13365 14057
rect 13323 14008 13324 14048
rect 13364 14008 13365 14048
rect 13323 13999 13365 14008
rect 14275 14048 14333 14049
rect 14275 14008 14284 14048
rect 14324 14008 14333 14048
rect 15331 14048 15389 14049
rect 14275 14007 14333 14008
rect 14763 14034 14805 14043
rect 12747 13985 12789 13994
rect 14763 13994 14764 14034
rect 14804 13994 14805 14034
rect 15331 14008 15340 14048
rect 15380 14008 15389 14048
rect 15331 14007 15389 14008
rect 16579 14048 16637 14049
rect 16579 14008 16588 14048
rect 16628 14008 16637 14048
rect 16579 14007 16637 14008
rect 18411 14048 18453 14057
rect 18411 14008 18412 14048
rect 18452 14008 18453 14048
rect 18411 13999 18453 14008
rect 18507 14048 18549 14057
rect 18507 14008 18508 14048
rect 18548 14008 18549 14048
rect 18507 13999 18549 14008
rect 18987 14048 19029 14057
rect 18987 14008 18988 14048
rect 19028 14008 19029 14048
rect 18987 13999 19029 14008
rect 19459 14048 19517 14049
rect 19459 14008 19468 14048
rect 19508 14008 19517 14048
rect 19459 14007 19517 14008
rect 19995 14038 20037 14047
rect 14763 13985 14805 13994
rect 19995 13998 19996 14038
rect 20036 13998 20037 14038
rect 19995 13989 20037 13998
rect 11691 13964 11733 13973
rect 11691 13924 11692 13964
rect 11732 13924 11733 13964
rect 11691 13915 11733 13924
rect 13707 13964 13749 13973
rect 13707 13924 13708 13964
rect 13748 13924 13749 13964
rect 13707 13915 13749 13924
rect 13803 13964 13845 13973
rect 13803 13924 13804 13964
rect 13844 13924 13845 13964
rect 13803 13915 13845 13924
rect 18891 13964 18933 13973
rect 18891 13924 18892 13964
rect 18932 13924 18933 13964
rect 18891 13915 18933 13924
rect 1152 13628 20352 13652
rect 1152 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 20352 13628
rect 1152 13564 20352 13588
rect 1803 13460 1845 13469
rect 1803 13420 1804 13460
rect 1844 13420 1845 13460
rect 1803 13411 1845 13420
rect 4395 13460 4437 13469
rect 4395 13420 4396 13460
rect 4436 13420 4437 13460
rect 4395 13411 4437 13420
rect 8907 13460 8949 13469
rect 8907 13420 8908 13460
rect 8948 13420 8949 13460
rect 8907 13411 8949 13420
rect 10923 13460 10965 13469
rect 10923 13420 10924 13460
rect 10964 13420 10965 13460
rect 10923 13411 10965 13420
rect 12555 13460 12597 13469
rect 12555 13420 12556 13460
rect 12596 13420 12597 13460
rect 12555 13411 12597 13420
rect 14571 13460 14613 13469
rect 14571 13420 14572 13460
rect 14612 13420 14613 13460
rect 14571 13411 14613 13420
rect 20235 13460 20277 13469
rect 20235 13420 20236 13460
rect 20276 13420 20277 13460
rect 20235 13411 20277 13420
rect 1603 13292 1661 13293
rect 1603 13252 1612 13292
rect 1652 13252 1661 13292
rect 1603 13251 1661 13252
rect 1987 13292 2045 13293
rect 1987 13252 1996 13292
rect 2036 13252 2045 13292
rect 1987 13251 2045 13252
rect 2763 13292 2805 13301
rect 2763 13252 2764 13292
rect 2804 13252 2805 13292
rect 2763 13243 2805 13252
rect 4195 13292 4253 13293
rect 4195 13252 4204 13292
rect 4244 13252 4253 13292
rect 4195 13251 4253 13252
rect 5931 13292 5973 13301
rect 5931 13252 5932 13292
rect 5972 13252 5973 13292
rect 5931 13243 5973 13252
rect 16491 13292 16533 13301
rect 16491 13252 16492 13292
rect 16532 13252 16533 13292
rect 16491 13243 16533 13252
rect 16587 13292 16629 13301
rect 16587 13252 16588 13292
rect 16628 13252 16629 13292
rect 16587 13243 16629 13252
rect 18115 13292 18173 13293
rect 18115 13252 18124 13292
rect 18164 13252 18173 13292
rect 18115 13251 18173 13252
rect 2283 13208 2325 13217
rect 2283 13168 2284 13208
rect 2324 13168 2325 13208
rect 2283 13159 2325 13168
rect 2379 13208 2421 13217
rect 2379 13168 2380 13208
rect 2420 13168 2421 13208
rect 2379 13159 2421 13168
rect 2859 13208 2901 13217
rect 3819 13213 3861 13222
rect 7035 13217 7077 13226
rect 17595 13217 17637 13226
rect 2859 13168 2860 13208
rect 2900 13168 2901 13208
rect 2859 13159 2901 13168
rect 3331 13208 3389 13209
rect 3331 13168 3340 13208
rect 3380 13168 3389 13208
rect 3331 13167 3389 13168
rect 3819 13173 3820 13213
rect 3860 13173 3861 13213
rect 3819 13164 3861 13173
rect 5451 13208 5493 13217
rect 5451 13168 5452 13208
rect 5492 13168 5493 13208
rect 5451 13159 5493 13168
rect 5547 13208 5589 13217
rect 5547 13168 5548 13208
rect 5588 13168 5589 13208
rect 5547 13159 5589 13168
rect 6027 13208 6069 13217
rect 6027 13168 6028 13208
rect 6068 13168 6069 13208
rect 6027 13159 6069 13168
rect 6499 13208 6557 13209
rect 6499 13168 6508 13208
rect 6548 13168 6557 13208
rect 7035 13177 7036 13217
rect 7076 13177 7077 13217
rect 7035 13168 7077 13177
rect 7459 13208 7517 13209
rect 7459 13168 7468 13208
rect 7508 13168 7517 13208
rect 6499 13167 6557 13168
rect 7459 13167 7517 13168
rect 8707 13208 8765 13209
rect 8707 13168 8716 13208
rect 8756 13168 8765 13208
rect 8707 13167 8765 13168
rect 9475 13208 9533 13209
rect 9475 13168 9484 13208
rect 9524 13168 9533 13208
rect 9475 13167 9533 13168
rect 10723 13208 10781 13209
rect 10723 13168 10732 13208
rect 10772 13168 10781 13208
rect 10723 13167 10781 13168
rect 11107 13208 11165 13209
rect 11107 13168 11116 13208
rect 11156 13168 11165 13208
rect 11107 13167 11165 13168
rect 12355 13208 12413 13209
rect 12355 13168 12364 13208
rect 12404 13168 12413 13208
rect 12355 13167 12413 13168
rect 13123 13208 13181 13209
rect 13123 13168 13132 13208
rect 13172 13168 13181 13208
rect 13123 13167 13181 13168
rect 14371 13208 14429 13209
rect 14371 13168 14380 13208
rect 14420 13168 14429 13208
rect 14371 13167 14429 13168
rect 16011 13208 16053 13217
rect 16011 13168 16012 13208
rect 16052 13168 16053 13208
rect 16011 13159 16053 13168
rect 16107 13208 16149 13217
rect 16107 13168 16108 13208
rect 16148 13168 16149 13208
rect 16107 13159 16149 13168
rect 17059 13208 17117 13209
rect 17059 13168 17068 13208
rect 17108 13168 17117 13208
rect 17595 13177 17596 13217
rect 17636 13177 17637 13217
rect 17595 13168 17637 13177
rect 18787 13208 18845 13209
rect 18787 13168 18796 13208
rect 18836 13168 18845 13208
rect 17059 13167 17117 13168
rect 18787 13167 18845 13168
rect 20035 13208 20093 13209
rect 20035 13168 20044 13208
rect 20084 13168 20093 13208
rect 20035 13167 20093 13168
rect 7179 13124 7221 13133
rect 7179 13084 7180 13124
rect 7220 13084 7221 13124
rect 7179 13075 7221 13084
rect 17739 13124 17781 13133
rect 17739 13084 17740 13124
rect 17780 13084 17781 13124
rect 17739 13075 17781 13084
rect 1419 13040 1461 13049
rect 1419 13000 1420 13040
rect 1460 13000 1461 13040
rect 1419 12991 1461 13000
rect 4011 13040 4053 13049
rect 4011 13000 4012 13040
rect 4052 13000 4053 13040
rect 4011 12991 4053 13000
rect 17931 13040 17973 13049
rect 17931 13000 17932 13040
rect 17972 13000 17973 13040
rect 17931 12991 17973 13000
rect 1152 12872 20452 12896
rect 1152 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20452 12872
rect 1152 12808 20452 12832
rect 10251 12704 10293 12713
rect 10251 12664 10252 12704
rect 10292 12664 10293 12704
rect 10251 12655 10293 12664
rect 10443 12704 10485 12713
rect 10443 12664 10444 12704
rect 10484 12664 10485 12704
rect 10443 12655 10485 12664
rect 16011 12704 16053 12713
rect 16011 12664 16012 12704
rect 16052 12664 16053 12704
rect 16011 12655 16053 12664
rect 4203 12620 4245 12629
rect 4203 12580 4204 12620
rect 4244 12580 4245 12620
rect 4203 12571 4245 12580
rect 6123 12620 6165 12629
rect 6123 12580 6124 12620
rect 6164 12580 6165 12620
rect 6123 12571 6165 12580
rect 8235 12620 8277 12629
rect 8235 12580 8236 12620
rect 8276 12580 8277 12620
rect 8235 12571 8277 12580
rect 12939 12620 12981 12629
rect 12939 12580 12940 12620
rect 12980 12580 12981 12620
rect 12939 12571 12981 12580
rect 17739 12620 17781 12629
rect 17739 12580 17740 12620
rect 17780 12580 17781 12620
rect 17739 12571 17781 12580
rect 20043 12620 20085 12629
rect 20043 12580 20044 12620
rect 20084 12580 20085 12620
rect 20043 12571 20085 12580
rect 2755 12536 2813 12537
rect 2755 12496 2764 12536
rect 2804 12496 2813 12536
rect 2755 12495 2813 12496
rect 4003 12536 4061 12537
rect 4003 12496 4012 12536
rect 4052 12496 4061 12536
rect 4003 12495 4061 12496
rect 4675 12536 4733 12537
rect 4675 12496 4684 12536
rect 4724 12496 4733 12536
rect 4675 12495 4733 12496
rect 5923 12536 5981 12537
rect 5923 12496 5932 12536
rect 5972 12496 5981 12536
rect 5923 12495 5981 12496
rect 6787 12536 6845 12537
rect 6787 12496 6796 12536
rect 6836 12496 6845 12536
rect 6787 12495 6845 12496
rect 8035 12536 8093 12537
rect 8035 12496 8044 12536
rect 8084 12496 8093 12536
rect 8035 12495 8093 12496
rect 8803 12536 8861 12537
rect 8803 12496 8812 12536
rect 8852 12496 8861 12536
rect 8803 12495 8861 12496
rect 10051 12536 10109 12537
rect 10051 12496 10060 12536
rect 10100 12496 10109 12536
rect 10051 12495 10109 12496
rect 11491 12536 11549 12537
rect 11491 12496 11500 12536
rect 11540 12496 11549 12536
rect 11491 12495 11549 12496
rect 12739 12536 12797 12537
rect 12739 12496 12748 12536
rect 12788 12496 12797 12536
rect 12739 12495 12797 12496
rect 14563 12536 14621 12537
rect 14563 12496 14572 12536
rect 14612 12496 14621 12536
rect 14563 12495 14621 12496
rect 15811 12536 15869 12537
rect 15811 12496 15820 12536
rect 15860 12496 15869 12536
rect 15811 12495 15869 12496
rect 16291 12536 16349 12537
rect 16291 12496 16300 12536
rect 16340 12496 16349 12536
rect 16291 12495 16349 12496
rect 17539 12536 17597 12537
rect 17539 12496 17548 12536
rect 17588 12496 17597 12536
rect 17539 12495 17597 12496
rect 18315 12536 18357 12545
rect 18315 12496 18316 12536
rect 18356 12496 18357 12536
rect 18315 12487 18357 12496
rect 18411 12536 18453 12545
rect 18411 12496 18412 12536
rect 18452 12496 18453 12536
rect 18411 12487 18453 12496
rect 18795 12536 18837 12545
rect 18795 12496 18796 12536
rect 18836 12496 18837 12536
rect 18795 12487 18837 12496
rect 18891 12536 18933 12545
rect 18891 12496 18892 12536
rect 18932 12496 18933 12536
rect 18891 12487 18933 12496
rect 19363 12536 19421 12537
rect 19363 12496 19372 12536
rect 19412 12496 19421 12536
rect 19363 12495 19421 12496
rect 19899 12494 19941 12503
rect 19899 12454 19900 12494
rect 19940 12454 19941 12494
rect 1699 12452 1757 12453
rect 1699 12412 1708 12452
rect 1748 12412 1757 12452
rect 1699 12411 1757 12412
rect 2083 12452 2141 12453
rect 2083 12412 2092 12452
rect 2132 12412 2141 12452
rect 2083 12411 2141 12412
rect 2467 12452 2525 12453
rect 2467 12412 2476 12452
rect 2516 12412 2525 12452
rect 2467 12411 2525 12412
rect 10627 12452 10685 12453
rect 10627 12412 10636 12452
rect 10676 12412 10685 12452
rect 10627 12411 10685 12412
rect 11299 12452 11357 12453
rect 11299 12412 11308 12452
rect 11348 12412 11357 12452
rect 11299 12411 11357 12412
rect 14179 12452 14237 12453
rect 14179 12412 14188 12452
rect 14228 12412 14237 12452
rect 19899 12445 19941 12454
rect 14179 12411 14237 12412
rect 11115 12368 11157 12377
rect 11115 12328 11116 12368
rect 11156 12328 11157 12368
rect 11115 12319 11157 12328
rect 13995 12368 14037 12377
rect 13995 12328 13996 12368
rect 14036 12328 14037 12368
rect 13995 12319 14037 12328
rect 1515 12284 1557 12293
rect 1515 12244 1516 12284
rect 1556 12244 1557 12284
rect 1515 12235 1557 12244
rect 1899 12284 1941 12293
rect 1899 12244 1900 12284
rect 1940 12244 1941 12284
rect 1899 12235 1941 12244
rect 2283 12284 2325 12293
rect 2283 12244 2284 12284
rect 2324 12244 2325 12284
rect 2283 12235 2325 12244
rect 1152 12116 20352 12140
rect 1152 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 20352 12116
rect 1152 12052 20352 12076
rect 2667 11948 2709 11957
rect 2667 11908 2668 11948
rect 2708 11908 2709 11948
rect 2667 11899 2709 11908
rect 5547 11948 5589 11957
rect 5547 11908 5548 11948
rect 5588 11908 5589 11948
rect 5547 11899 5589 11908
rect 12171 11948 12213 11957
rect 12171 11908 12172 11948
rect 12212 11908 12213 11948
rect 12171 11899 12213 11908
rect 18699 11948 18741 11957
rect 18699 11908 18700 11948
rect 18740 11908 18741 11948
rect 18699 11899 18741 11908
rect 3243 11864 3285 11873
rect 3243 11824 3244 11864
rect 3284 11824 3285 11864
rect 3243 11815 3285 11824
rect 3043 11780 3101 11781
rect 3043 11740 3052 11780
rect 3092 11740 3101 11780
rect 3043 11739 3101 11740
rect 3427 11780 3485 11781
rect 3427 11740 3436 11780
rect 3476 11740 3485 11780
rect 3427 11739 3485 11740
rect 3811 11780 3869 11781
rect 3811 11740 3820 11780
rect 3860 11740 3869 11780
rect 3811 11739 3869 11740
rect 6411 11780 6453 11789
rect 6411 11740 6412 11780
rect 6452 11740 6453 11780
rect 6411 11731 6453 11740
rect 9003 11780 9045 11789
rect 9003 11740 9004 11780
rect 9044 11740 9045 11780
rect 9003 11731 9045 11740
rect 9099 11780 9141 11789
rect 9099 11740 9100 11780
rect 9140 11740 9141 11780
rect 9099 11731 9141 11740
rect 12355 11780 12413 11781
rect 12355 11740 12364 11780
rect 12404 11740 12413 11780
rect 12355 11739 12413 11740
rect 15051 11780 15093 11789
rect 15051 11740 15052 11780
rect 15092 11740 15093 11780
rect 15051 11731 15093 11740
rect 1219 11696 1277 11697
rect 1219 11656 1228 11696
rect 1268 11656 1277 11696
rect 1219 11655 1277 11656
rect 2467 11696 2525 11697
rect 2467 11656 2476 11696
rect 2516 11656 2525 11696
rect 2467 11655 2525 11656
rect 4099 11696 4157 11697
rect 4099 11656 4108 11696
rect 4148 11656 4157 11696
rect 4099 11655 4157 11656
rect 5347 11696 5405 11697
rect 5347 11656 5356 11696
rect 5396 11656 5405 11696
rect 5347 11655 5405 11656
rect 5835 11696 5877 11705
rect 5835 11656 5836 11696
rect 5876 11656 5877 11696
rect 5835 11647 5877 11656
rect 5931 11696 5973 11705
rect 5931 11656 5932 11696
rect 5972 11656 5973 11696
rect 5931 11647 5973 11656
rect 6315 11696 6357 11705
rect 7371 11701 7413 11710
rect 6315 11656 6316 11696
rect 6356 11656 6357 11696
rect 6315 11647 6357 11656
rect 6883 11696 6941 11697
rect 6883 11656 6892 11696
rect 6932 11656 6941 11696
rect 6883 11655 6941 11656
rect 7371 11661 7372 11701
rect 7412 11661 7413 11701
rect 7371 11652 7413 11661
rect 8523 11696 8565 11705
rect 8523 11656 8524 11696
rect 8564 11656 8565 11696
rect 8523 11647 8565 11656
rect 8619 11696 8661 11705
rect 10059 11701 10101 11710
rect 8619 11656 8620 11696
rect 8660 11656 8661 11696
rect 8619 11647 8661 11656
rect 9571 11696 9629 11697
rect 9571 11656 9580 11696
rect 9620 11656 9629 11696
rect 9571 11655 9629 11656
rect 10059 11661 10060 11701
rect 10100 11661 10101 11701
rect 10059 11652 10101 11661
rect 10531 11696 10589 11697
rect 10531 11656 10540 11696
rect 10580 11656 10589 11696
rect 10531 11655 10589 11656
rect 11779 11696 11837 11697
rect 11779 11656 11788 11696
rect 11828 11656 11837 11696
rect 11779 11655 11837 11656
rect 12643 11696 12701 11697
rect 12643 11656 12652 11696
rect 12692 11656 12701 11696
rect 12643 11655 12701 11656
rect 13891 11696 13949 11697
rect 13891 11656 13900 11696
rect 13940 11656 13949 11696
rect 13891 11655 13949 11656
rect 14571 11696 14613 11705
rect 14571 11656 14572 11696
rect 14612 11656 14613 11696
rect 14571 11647 14613 11656
rect 14667 11696 14709 11705
rect 14667 11656 14668 11696
rect 14708 11656 14709 11696
rect 14667 11647 14709 11656
rect 15147 11696 15189 11705
rect 16107 11701 16149 11710
rect 15147 11656 15148 11696
rect 15188 11656 15189 11696
rect 15147 11647 15189 11656
rect 15619 11696 15677 11697
rect 15619 11656 15628 11696
rect 15668 11656 15677 11696
rect 15619 11655 15677 11656
rect 16107 11661 16108 11701
rect 16148 11661 16149 11701
rect 16107 11652 16149 11661
rect 17251 11696 17309 11697
rect 17251 11656 17260 11696
rect 17300 11656 17309 11696
rect 17251 11655 17309 11656
rect 18499 11696 18557 11697
rect 18499 11656 18508 11696
rect 18548 11656 18557 11696
rect 18499 11655 18557 11656
rect 7563 11612 7605 11621
rect 7563 11572 7564 11612
rect 7604 11572 7605 11612
rect 7563 11563 7605 11572
rect 10251 11612 10293 11621
rect 10251 11572 10252 11612
rect 10292 11572 10293 11612
rect 10251 11563 10293 11572
rect 16299 11612 16341 11621
rect 16299 11572 16300 11612
rect 16340 11572 16341 11612
rect 16299 11563 16341 11572
rect 2859 11528 2901 11537
rect 2859 11488 2860 11528
rect 2900 11488 2901 11528
rect 2859 11479 2901 11488
rect 3627 11528 3669 11537
rect 3627 11488 3628 11528
rect 3668 11488 3669 11528
rect 3627 11479 3669 11488
rect 11979 11528 12021 11537
rect 11979 11488 11980 11528
rect 12020 11488 12021 11528
rect 11979 11479 12021 11488
rect 14091 11528 14133 11537
rect 14091 11488 14092 11528
rect 14132 11488 14133 11528
rect 14091 11479 14133 11488
rect 1152 11360 20452 11384
rect 1152 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20452 11360
rect 1152 11296 20452 11320
rect 1899 11192 1941 11201
rect 1899 11152 1900 11192
rect 1940 11152 1941 11192
rect 1899 11143 1941 11152
rect 9963 11192 10005 11201
rect 9963 11152 9964 11192
rect 10004 11152 10005 11192
rect 9963 11143 10005 11152
rect 11979 11192 12021 11201
rect 11979 11152 11980 11192
rect 12020 11152 12021 11192
rect 11979 11143 12021 11152
rect 14283 11192 14325 11201
rect 14283 11152 14284 11192
rect 14324 11152 14325 11192
rect 14283 11143 14325 11152
rect 20139 11192 20181 11201
rect 20139 11152 20140 11192
rect 20180 11152 20181 11192
rect 20139 11143 20181 11152
rect 4299 11108 4341 11117
rect 4299 11068 4300 11108
rect 4340 11068 4341 11108
rect 4299 11059 4341 11068
rect 7179 11108 7221 11117
rect 7179 11068 7180 11108
rect 7220 11068 7221 11108
rect 7179 11059 7221 11068
rect 17451 11108 17493 11117
rect 17451 11068 17452 11108
rect 17492 11068 17493 11108
rect 17451 11059 17493 11068
rect 2571 11024 2613 11033
rect 2571 10984 2572 11024
rect 2612 10984 2613 11024
rect 2571 10975 2613 10984
rect 2667 11024 2709 11033
rect 2667 10984 2668 11024
rect 2708 10984 2709 11024
rect 2667 10975 2709 10984
rect 3619 11024 3677 11025
rect 3619 10984 3628 11024
rect 3668 10984 3677 11024
rect 5451 11024 5493 11033
rect 3619 10983 3677 10984
rect 4107 11010 4149 11019
rect 4107 10970 4108 11010
rect 4148 10970 4149 11010
rect 5451 10984 5452 11024
rect 5492 10984 5493 11024
rect 5451 10975 5493 10984
rect 5547 11024 5589 11033
rect 5547 10984 5548 11024
rect 5588 10984 5589 11024
rect 5547 10975 5589 10984
rect 5931 11024 5973 11033
rect 5931 10984 5932 11024
rect 5972 10984 5973 11024
rect 5931 10975 5973 10984
rect 6027 11024 6069 11033
rect 6027 10984 6028 11024
rect 6068 10984 6069 11024
rect 6027 10975 6069 10984
rect 6499 11024 6557 11025
rect 6499 10984 6508 11024
rect 6548 10984 6557 11024
rect 8515 11024 8573 11025
rect 6499 10983 6557 10984
rect 6987 11010 7029 11019
rect 4107 10961 4149 10970
rect 6987 10970 6988 11010
rect 7028 10970 7029 11010
rect 8515 10984 8524 11024
rect 8564 10984 8573 11024
rect 8515 10983 8573 10984
rect 9763 11024 9821 11025
rect 9763 10984 9772 11024
rect 9812 10984 9821 11024
rect 9763 10983 9821 10984
rect 10251 11024 10293 11033
rect 10251 10984 10252 11024
rect 10292 10984 10293 11024
rect 10251 10975 10293 10984
rect 10347 11024 10389 11033
rect 10347 10984 10348 11024
rect 10388 10984 10389 11024
rect 10347 10975 10389 10984
rect 10731 11024 10773 11033
rect 10731 10984 10732 11024
rect 10772 10984 10773 11024
rect 10731 10975 10773 10984
rect 11299 11024 11357 11025
rect 11299 10984 11308 11024
rect 11348 10984 11357 11024
rect 12555 11024 12597 11033
rect 11299 10983 11357 10984
rect 11835 11014 11877 11023
rect 6987 10961 7029 10970
rect 11835 10974 11836 11014
rect 11876 10974 11877 11014
rect 12555 10984 12556 11024
rect 12596 10984 12597 11024
rect 12555 10975 12597 10984
rect 12651 11024 12693 11033
rect 12651 10984 12652 11024
rect 12692 10984 12693 11024
rect 12651 10975 12693 10984
rect 13131 11024 13173 11033
rect 13131 10984 13132 11024
rect 13172 10984 13173 11024
rect 13131 10975 13173 10984
rect 13603 11024 13661 11025
rect 13603 10984 13612 11024
rect 13652 10984 13661 11024
rect 13603 10983 13661 10984
rect 14091 11019 14133 11028
rect 14091 10979 14092 11019
rect 14132 10979 14133 11019
rect 11835 10965 11877 10974
rect 14091 10970 14133 10979
rect 15723 11024 15765 11033
rect 15723 10984 15724 11024
rect 15764 10984 15765 11024
rect 15723 10975 15765 10984
rect 15819 11024 15861 11033
rect 15819 10984 15820 11024
rect 15860 10984 15861 11024
rect 15819 10975 15861 10984
rect 16299 11024 16341 11033
rect 16299 10984 16300 11024
rect 16340 10984 16341 11024
rect 16299 10975 16341 10984
rect 16771 11024 16829 11025
rect 16771 10984 16780 11024
rect 16820 10984 16829 11024
rect 18691 11024 18749 11025
rect 16771 10983 16829 10984
rect 17259 11010 17301 11019
rect 17259 10970 17260 11010
rect 17300 10970 17301 11010
rect 18691 10984 18700 11024
rect 18740 10984 18749 11024
rect 18691 10983 18749 10984
rect 19939 11024 19997 11025
rect 19939 10984 19948 11024
rect 19988 10984 19997 11024
rect 19939 10983 19997 10984
rect 17259 10961 17301 10970
rect 1699 10940 1757 10941
rect 1699 10900 1708 10940
rect 1748 10900 1757 10940
rect 1699 10899 1757 10900
rect 2083 10940 2141 10941
rect 2083 10900 2092 10940
rect 2132 10900 2141 10940
rect 2083 10899 2141 10900
rect 3051 10940 3093 10949
rect 3051 10900 3052 10940
rect 3092 10900 3093 10940
rect 3051 10891 3093 10900
rect 3147 10940 3189 10949
rect 3147 10900 3148 10940
rect 3188 10900 3189 10940
rect 3147 10891 3189 10900
rect 4675 10940 4733 10941
rect 4675 10900 4684 10940
rect 4724 10900 4733 10940
rect 4675 10899 4733 10900
rect 4867 10940 4925 10941
rect 4867 10900 4876 10940
rect 4916 10900 4925 10940
rect 4867 10899 4925 10900
rect 10827 10940 10869 10949
rect 10827 10900 10828 10940
rect 10868 10900 10869 10940
rect 10827 10891 10869 10900
rect 13035 10940 13077 10949
rect 13035 10900 13036 10940
rect 13076 10900 13077 10940
rect 13035 10891 13077 10900
rect 14659 10940 14717 10941
rect 14659 10900 14668 10940
rect 14708 10900 14717 10940
rect 14659 10899 14717 10900
rect 16203 10940 16245 10949
rect 16203 10900 16204 10940
rect 16244 10900 16245 10940
rect 16203 10891 16245 10900
rect 14475 10856 14517 10865
rect 14475 10816 14476 10856
rect 14516 10816 14517 10856
rect 14475 10807 14517 10816
rect 1515 10772 1557 10781
rect 1515 10732 1516 10772
rect 1556 10732 1557 10772
rect 1515 10723 1557 10732
rect 4491 10772 4533 10781
rect 4491 10732 4492 10772
rect 4532 10732 4533 10772
rect 4491 10723 4533 10732
rect 5067 10772 5109 10781
rect 5067 10732 5068 10772
rect 5108 10732 5109 10772
rect 5067 10723 5109 10732
rect 1152 10604 20352 10628
rect 1152 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 20352 10604
rect 1152 10540 20352 10564
rect 2667 10436 2709 10445
rect 2667 10396 2668 10436
rect 2708 10396 2709 10436
rect 2667 10387 2709 10396
rect 4971 10436 5013 10445
rect 4971 10396 4972 10436
rect 5012 10396 5013 10436
rect 4971 10387 5013 10396
rect 5163 10436 5205 10445
rect 5163 10396 5164 10436
rect 5204 10396 5205 10436
rect 5163 10387 5205 10396
rect 7083 10436 7125 10445
rect 7083 10396 7084 10436
rect 7124 10396 7125 10436
rect 7083 10387 7125 10396
rect 10155 10436 10197 10445
rect 10155 10396 10156 10436
rect 10196 10396 10197 10436
rect 10155 10387 10197 10396
rect 12747 10436 12789 10445
rect 12747 10396 12748 10436
rect 12788 10396 12789 10436
rect 12747 10387 12789 10396
rect 14475 10436 14517 10445
rect 14475 10396 14476 10436
rect 14516 10396 14517 10436
rect 14475 10387 14517 10396
rect 16203 10436 16245 10445
rect 16203 10396 16204 10436
rect 16244 10396 16245 10436
rect 16203 10387 16245 10396
rect 17835 10436 17877 10445
rect 17835 10396 17836 10436
rect 17876 10396 17877 10436
rect 17835 10387 17877 10396
rect 2859 10352 2901 10361
rect 2859 10312 2860 10352
rect 2900 10312 2901 10352
rect 2859 10303 2901 10312
rect 3043 10268 3101 10269
rect 3043 10228 3052 10268
rect 3092 10228 3101 10268
rect 3043 10227 3101 10228
rect 5347 10268 5405 10269
rect 5347 10228 5356 10268
rect 5396 10228 5405 10268
rect 5347 10227 5405 10228
rect 7459 10268 7517 10269
rect 7459 10228 7468 10268
rect 7508 10228 7517 10268
rect 7459 10227 7517 10228
rect 18699 10268 18741 10277
rect 18699 10228 18700 10268
rect 18740 10228 18741 10268
rect 18699 10219 18741 10228
rect 18795 10268 18837 10277
rect 18795 10228 18796 10268
rect 18836 10228 18837 10268
rect 18795 10219 18837 10228
rect 19803 10193 19845 10202
rect 1219 10184 1277 10185
rect 1219 10144 1228 10184
rect 1268 10144 1277 10184
rect 1219 10143 1277 10144
rect 2467 10184 2525 10185
rect 2467 10144 2476 10184
rect 2516 10144 2525 10184
rect 2467 10143 2525 10144
rect 4771 10184 4829 10185
rect 4771 10144 4780 10184
rect 4820 10144 4829 10184
rect 4771 10143 4829 10144
rect 5635 10184 5693 10185
rect 5635 10144 5644 10184
rect 5684 10144 5693 10184
rect 5635 10143 5693 10144
rect 6883 10184 6941 10185
rect 6883 10144 6892 10184
rect 6932 10144 6941 10184
rect 6883 10143 6941 10144
rect 8707 10184 8765 10185
rect 8707 10144 8716 10184
rect 8756 10144 8765 10184
rect 8707 10143 8765 10144
rect 9955 10184 10013 10185
rect 9955 10144 9964 10184
rect 10004 10144 10013 10184
rect 9955 10143 10013 10144
rect 11299 10184 11357 10185
rect 11299 10144 11308 10184
rect 11348 10144 11357 10184
rect 11299 10143 11357 10144
rect 12547 10184 12605 10185
rect 12547 10144 12556 10184
rect 12596 10144 12605 10184
rect 12547 10143 12605 10144
rect 13027 10184 13085 10185
rect 13027 10144 13036 10184
rect 13076 10144 13085 10184
rect 13027 10143 13085 10144
rect 14275 10184 14333 10185
rect 14275 10144 14284 10184
rect 14324 10144 14333 10184
rect 14275 10143 14333 10144
rect 14755 10184 14813 10185
rect 14755 10144 14764 10184
rect 14804 10144 14813 10184
rect 14755 10143 14813 10144
rect 16003 10184 16061 10185
rect 16003 10144 16012 10184
rect 16052 10144 16061 10184
rect 16003 10143 16061 10144
rect 16387 10184 16445 10185
rect 16387 10144 16396 10184
rect 16436 10144 16445 10184
rect 16387 10143 16445 10144
rect 17635 10184 17693 10185
rect 17635 10144 17644 10184
rect 17684 10144 17693 10184
rect 17635 10143 17693 10144
rect 18219 10184 18261 10193
rect 18219 10144 18220 10184
rect 18260 10144 18261 10184
rect 3523 10142 3581 10143
rect 3523 10102 3532 10142
rect 3572 10102 3581 10142
rect 18219 10135 18261 10144
rect 18315 10184 18357 10193
rect 18315 10144 18316 10184
rect 18356 10144 18357 10184
rect 18315 10135 18357 10144
rect 19267 10184 19325 10185
rect 19267 10144 19276 10184
rect 19316 10144 19325 10184
rect 19803 10153 19804 10193
rect 19844 10153 19845 10193
rect 19803 10144 19845 10153
rect 19267 10143 19325 10144
rect 3523 10101 3581 10102
rect 19947 10100 19989 10109
rect 19947 10060 19948 10100
rect 19988 10060 19989 10100
rect 19947 10051 19989 10060
rect 7275 10016 7317 10025
rect 7275 9976 7276 10016
rect 7316 9976 7317 10016
rect 7275 9967 7317 9976
rect 1152 9848 20452 9872
rect 1152 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20452 9848
rect 1152 9784 20452 9808
rect 19947 9722 19989 9731
rect 1419 9680 1461 9689
rect 1419 9640 1420 9680
rect 1460 9640 1461 9680
rect 1419 9631 1461 9640
rect 2187 9680 2229 9689
rect 2187 9640 2188 9680
rect 2228 9640 2229 9680
rect 2187 9631 2229 9640
rect 4395 9680 4437 9689
rect 4395 9640 4396 9680
rect 4436 9640 4437 9680
rect 4395 9631 4437 9640
rect 7083 9680 7125 9689
rect 7083 9640 7084 9680
rect 7124 9640 7125 9680
rect 7083 9631 7125 9640
rect 8715 9680 8757 9689
rect 8715 9640 8716 9680
rect 8756 9640 8757 9680
rect 8715 9631 8757 9640
rect 13515 9680 13557 9689
rect 13515 9640 13516 9680
rect 13556 9640 13557 9680
rect 13515 9631 13557 9640
rect 15819 9680 15861 9689
rect 15819 9640 15820 9680
rect 15860 9640 15861 9680
rect 15819 9631 15861 9640
rect 17931 9680 17973 9689
rect 17931 9640 17932 9680
rect 17972 9640 17973 9680
rect 19947 9682 19948 9722
rect 19988 9682 19989 9722
rect 19947 9673 19989 9682
rect 17931 9631 17973 9640
rect 11691 9596 11733 9605
rect 11691 9556 11692 9596
rect 11732 9556 11733 9596
rect 11691 9547 11733 9556
rect 11883 9596 11925 9605
rect 11883 9556 11884 9596
rect 11924 9556 11925 9596
rect 11883 9547 11925 9556
rect 2667 9512 2709 9521
rect 2667 9472 2668 9512
rect 2708 9472 2709 9512
rect 2667 9463 2709 9472
rect 2763 9512 2805 9521
rect 2763 9472 2764 9512
rect 2804 9472 2805 9512
rect 2763 9463 2805 9472
rect 3147 9512 3189 9521
rect 3147 9472 3148 9512
rect 3188 9472 3189 9512
rect 3147 9463 3189 9472
rect 3243 9512 3285 9521
rect 3243 9472 3244 9512
rect 3284 9472 3285 9512
rect 3243 9463 3285 9472
rect 3715 9512 3773 9513
rect 3715 9472 3724 9512
rect 3764 9472 3773 9512
rect 3715 9471 3773 9472
rect 4203 9507 4245 9516
rect 4203 9467 4204 9507
rect 4244 9467 4245 9507
rect 5635 9512 5693 9513
rect 5635 9472 5644 9512
rect 5684 9472 5693 9512
rect 5635 9471 5693 9472
rect 6883 9512 6941 9513
rect 6883 9472 6892 9512
rect 6932 9472 6941 9512
rect 6883 9471 6941 9472
rect 7267 9512 7325 9513
rect 7267 9472 7276 9512
rect 7316 9472 7325 9512
rect 7267 9471 7325 9472
rect 8515 9512 8573 9513
rect 8515 9472 8524 9512
rect 8564 9472 8573 9512
rect 8515 9471 8573 9472
rect 9963 9512 10005 9521
rect 9963 9472 9964 9512
rect 10004 9472 10005 9512
rect 4203 9458 4245 9467
rect 9963 9463 10005 9472
rect 10059 9512 10101 9521
rect 10059 9472 10060 9512
rect 10100 9472 10101 9512
rect 10059 9463 10101 9472
rect 10539 9512 10581 9521
rect 10539 9472 10540 9512
rect 10580 9472 10581 9512
rect 10539 9463 10581 9472
rect 11011 9512 11069 9513
rect 11011 9472 11020 9512
rect 11060 9472 11069 9512
rect 11011 9471 11069 9472
rect 11499 9507 11541 9516
rect 11499 9467 11500 9507
rect 11540 9467 11541 9507
rect 12067 9512 12125 9513
rect 12067 9472 12076 9512
rect 12116 9472 12125 9512
rect 12067 9471 12125 9472
rect 13315 9512 13373 9513
rect 13315 9472 13324 9512
rect 13364 9472 13373 9512
rect 13315 9471 13373 9472
rect 14371 9512 14429 9513
rect 14371 9472 14380 9512
rect 14420 9472 14429 9512
rect 14371 9471 14429 9472
rect 15619 9512 15677 9513
rect 15619 9472 15628 9512
rect 15668 9472 15677 9512
rect 15619 9471 15677 9472
rect 16483 9512 16541 9513
rect 16483 9472 16492 9512
rect 16532 9472 16541 9512
rect 16483 9471 16541 9472
rect 17731 9512 17789 9513
rect 17731 9472 17740 9512
rect 17780 9472 17789 9512
rect 17731 9471 17789 9472
rect 18219 9512 18261 9521
rect 18219 9472 18220 9512
rect 18260 9472 18261 9512
rect 11499 9458 11541 9467
rect 18219 9463 18261 9472
rect 18315 9512 18357 9521
rect 18315 9472 18316 9512
rect 18356 9472 18357 9512
rect 18315 9463 18357 9472
rect 18699 9512 18741 9521
rect 18699 9472 18700 9512
rect 18740 9472 18741 9512
rect 18699 9463 18741 9472
rect 18795 9512 18837 9521
rect 18795 9472 18796 9512
rect 18836 9472 18837 9512
rect 18795 9463 18837 9472
rect 19267 9512 19325 9513
rect 19267 9472 19276 9512
rect 19316 9472 19325 9512
rect 19267 9471 19325 9472
rect 19803 9470 19845 9479
rect 1603 9428 1661 9429
rect 1603 9388 1612 9428
rect 1652 9388 1661 9428
rect 1603 9387 1661 9388
rect 1987 9428 2045 9429
rect 1987 9388 1996 9428
rect 2036 9388 2045 9428
rect 1987 9387 2045 9388
rect 2371 9428 2429 9429
rect 2371 9388 2380 9428
rect 2420 9388 2429 9428
rect 2371 9387 2429 9388
rect 4771 9428 4829 9429
rect 4771 9388 4780 9428
rect 4820 9388 4829 9428
rect 4771 9387 4829 9388
rect 5155 9428 5213 9429
rect 5155 9388 5164 9428
rect 5204 9388 5213 9428
rect 5155 9387 5213 9388
rect 10443 9428 10485 9437
rect 19803 9430 19804 9470
rect 19844 9430 19845 9470
rect 10443 9388 10444 9428
rect 10484 9388 10485 9428
rect 10443 9379 10485 9388
rect 13699 9428 13757 9429
rect 13699 9388 13708 9428
rect 13748 9388 13757 9428
rect 19803 9421 19845 9430
rect 13699 9387 13757 9388
rect 1803 9260 1845 9269
rect 1803 9220 1804 9260
rect 1844 9220 1845 9260
rect 1803 9211 1845 9220
rect 4587 9260 4629 9269
rect 4587 9220 4588 9260
rect 4628 9220 4629 9260
rect 4587 9211 4629 9220
rect 4971 9260 5013 9269
rect 4971 9220 4972 9260
rect 5012 9220 5013 9260
rect 4971 9211 5013 9220
rect 1152 9092 20352 9116
rect 1152 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 20352 9092
rect 1152 9028 20352 9052
rect 18315 8924 18357 8933
rect 18315 8884 18316 8924
rect 18356 8884 18357 8924
rect 18315 8875 18357 8884
rect 20139 8924 20181 8933
rect 20139 8884 20140 8924
rect 20180 8884 20181 8924
rect 20139 8875 20181 8884
rect 2667 8840 2709 8849
rect 2667 8800 2668 8840
rect 2708 8800 2709 8840
rect 2667 8791 2709 8800
rect 4299 8840 4341 8849
rect 4299 8800 4300 8840
rect 4340 8800 4341 8840
rect 4299 8791 4341 8800
rect 4675 8756 4733 8757
rect 4675 8716 4684 8756
rect 4724 8716 4733 8756
rect 4675 8715 4733 8716
rect 5643 8756 5685 8765
rect 5643 8716 5644 8756
rect 5684 8716 5685 8756
rect 5643 8707 5685 8716
rect 5739 8756 5781 8765
rect 5739 8716 5740 8756
rect 5780 8716 5781 8756
rect 5739 8707 5781 8716
rect 7851 8756 7893 8765
rect 7851 8716 7852 8756
rect 7892 8716 7893 8756
rect 7851 8707 7893 8716
rect 7947 8756 7989 8765
rect 7947 8716 7948 8756
rect 7988 8716 7989 8756
rect 7947 8707 7989 8716
rect 16107 8756 16149 8765
rect 16107 8716 16108 8756
rect 16148 8716 16149 8756
rect 16107 8707 16149 8716
rect 1219 8672 1277 8673
rect 1219 8632 1228 8672
rect 1268 8632 1277 8672
rect 1219 8631 1277 8632
rect 2467 8672 2525 8673
rect 2467 8632 2476 8672
rect 2516 8632 2525 8672
rect 2467 8631 2525 8632
rect 2851 8672 2909 8673
rect 2851 8632 2860 8672
rect 2900 8632 2909 8672
rect 2851 8631 2909 8632
rect 4099 8672 4157 8673
rect 4099 8632 4108 8672
rect 4148 8632 4157 8672
rect 4099 8631 4157 8632
rect 5163 8672 5205 8681
rect 5163 8632 5164 8672
rect 5204 8632 5205 8672
rect 5163 8623 5205 8632
rect 5259 8672 5301 8681
rect 6699 8677 6741 8686
rect 8955 8681 8997 8690
rect 5259 8632 5260 8672
rect 5300 8632 5301 8672
rect 5259 8623 5301 8632
rect 6211 8672 6269 8673
rect 6211 8632 6220 8672
rect 6260 8632 6269 8672
rect 6211 8631 6269 8632
rect 6699 8637 6700 8677
rect 6740 8637 6741 8677
rect 6699 8628 6741 8637
rect 7371 8672 7413 8681
rect 7371 8632 7372 8672
rect 7412 8632 7413 8672
rect 7371 8623 7413 8632
rect 7467 8672 7509 8681
rect 7467 8632 7468 8672
rect 7508 8632 7509 8672
rect 7467 8623 7509 8632
rect 8419 8672 8477 8673
rect 8419 8632 8428 8672
rect 8468 8632 8477 8672
rect 8955 8641 8956 8681
rect 8996 8641 8997 8681
rect 8955 8632 8997 8641
rect 10627 8672 10685 8673
rect 10627 8632 10636 8672
rect 10676 8632 10685 8672
rect 8419 8631 8477 8632
rect 10627 8631 10685 8632
rect 11875 8672 11933 8673
rect 11875 8632 11884 8672
rect 11924 8632 11933 8672
rect 11875 8631 11933 8632
rect 12363 8672 12405 8681
rect 12363 8632 12364 8672
rect 12404 8632 12405 8672
rect 12363 8623 12405 8632
rect 12459 8672 12501 8681
rect 12459 8632 12460 8672
rect 12500 8632 12501 8672
rect 12459 8623 12501 8632
rect 12843 8672 12885 8681
rect 12843 8632 12844 8672
rect 12884 8632 12885 8672
rect 12843 8623 12885 8632
rect 12939 8672 12981 8681
rect 13899 8677 13941 8686
rect 12939 8632 12940 8672
rect 12980 8632 12981 8672
rect 12939 8623 12981 8632
rect 13411 8672 13469 8673
rect 13411 8632 13420 8672
rect 13460 8632 13469 8672
rect 13411 8631 13469 8632
rect 13899 8637 13900 8677
rect 13940 8637 13941 8677
rect 13899 8628 13941 8637
rect 15051 8677 15093 8686
rect 15051 8637 15052 8677
rect 15092 8637 15093 8677
rect 15051 8628 15093 8637
rect 15523 8672 15581 8673
rect 15523 8632 15532 8672
rect 15572 8632 15581 8672
rect 15523 8631 15581 8632
rect 16011 8672 16053 8681
rect 16011 8632 16012 8672
rect 16052 8632 16053 8672
rect 16011 8623 16053 8632
rect 16491 8672 16533 8681
rect 16491 8632 16492 8672
rect 16532 8632 16533 8672
rect 16491 8623 16533 8632
rect 16587 8672 16629 8681
rect 16587 8632 16588 8672
rect 16628 8632 16629 8672
rect 16587 8623 16629 8632
rect 16867 8672 16925 8673
rect 16867 8632 16876 8672
rect 16916 8632 16925 8672
rect 16867 8631 16925 8632
rect 18115 8672 18173 8673
rect 18115 8632 18124 8672
rect 18164 8632 18173 8672
rect 18115 8631 18173 8632
rect 18691 8672 18749 8673
rect 18691 8632 18700 8672
rect 18740 8632 18749 8672
rect 18691 8631 18749 8632
rect 19939 8672 19997 8673
rect 19939 8632 19948 8672
rect 19988 8632 19997 8672
rect 19939 8631 19997 8632
rect 12075 8588 12117 8597
rect 12075 8548 12076 8588
rect 12116 8548 12117 8588
rect 12075 8539 12117 8548
rect 14091 8588 14133 8597
rect 14091 8548 14092 8588
rect 14132 8548 14133 8588
rect 14091 8539 14133 8548
rect 4875 8504 4917 8513
rect 4875 8464 4876 8504
rect 4916 8464 4917 8504
rect 4875 8455 4917 8464
rect 6891 8504 6933 8513
rect 6891 8464 6892 8504
rect 6932 8464 6933 8504
rect 6891 8455 6933 8464
rect 9099 8504 9141 8513
rect 9099 8464 9100 8504
rect 9140 8464 9141 8504
rect 9099 8455 9141 8464
rect 14859 8504 14901 8513
rect 14859 8464 14860 8504
rect 14900 8464 14901 8504
rect 14859 8455 14901 8464
rect 1152 8336 20452 8360
rect 1152 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20452 8336
rect 1152 8272 20452 8296
rect 2667 8168 2709 8177
rect 2667 8128 2668 8168
rect 2708 8128 2709 8168
rect 2667 8119 2709 8128
rect 2859 8168 2901 8177
rect 2859 8128 2860 8168
rect 2900 8128 2901 8168
rect 2859 8119 2901 8128
rect 3243 8168 3285 8177
rect 3243 8128 3244 8168
rect 3284 8128 3285 8168
rect 3243 8119 3285 8128
rect 5643 8168 5685 8177
rect 5643 8128 5644 8168
rect 5684 8128 5685 8168
rect 5643 8119 5685 8128
rect 7275 8168 7317 8177
rect 7275 8128 7276 8168
rect 7316 8128 7317 8168
rect 7275 8119 7317 8128
rect 9675 8168 9717 8177
rect 9675 8128 9676 8168
rect 9716 8128 9717 8168
rect 9675 8119 9717 8128
rect 9867 8168 9909 8177
rect 9867 8128 9868 8168
rect 9908 8128 9909 8168
rect 9867 8119 9909 8128
rect 13899 8168 13941 8177
rect 13899 8128 13900 8168
rect 13940 8128 13941 8168
rect 13899 8119 13941 8128
rect 15531 8168 15573 8177
rect 15531 8128 15532 8168
rect 15572 8128 15573 8168
rect 15531 8119 15573 8128
rect 15723 8168 15765 8177
rect 15723 8128 15724 8168
rect 15764 8128 15765 8168
rect 15723 8119 15765 8128
rect 19659 8168 19701 8177
rect 19659 8128 19660 8168
rect 19700 8128 19701 8168
rect 19659 8119 19701 8128
rect 1219 8000 1277 8001
rect 1219 7960 1228 8000
rect 1268 7960 1277 8000
rect 1219 7959 1277 7960
rect 2467 8000 2525 8001
rect 2467 7960 2476 8000
rect 2516 7960 2525 8000
rect 2467 7959 2525 7960
rect 4195 8000 4253 8001
rect 4195 7960 4204 8000
rect 4244 7960 4253 8000
rect 4195 7959 4253 7960
rect 5443 8000 5501 8001
rect 5443 7960 5452 8000
rect 5492 7960 5501 8000
rect 5443 7959 5501 7960
rect 5827 8000 5885 8001
rect 5827 7960 5836 8000
rect 5876 7960 5885 8000
rect 5827 7959 5885 7960
rect 7075 8000 7133 8001
rect 7075 7960 7084 8000
rect 7124 7960 7133 8000
rect 7075 7959 7133 7960
rect 8227 8000 8285 8001
rect 8227 7960 8236 8000
rect 8276 7960 8285 8000
rect 8227 7959 8285 7960
rect 9475 8000 9533 8001
rect 9475 7960 9484 8000
rect 9524 7960 9533 8000
rect 9475 7959 9533 7960
rect 10059 7995 10101 8004
rect 10059 7955 10060 7995
rect 10100 7955 10101 7995
rect 10531 8000 10589 8001
rect 10531 7960 10540 8000
rect 10580 7960 10589 8000
rect 10531 7959 10589 7960
rect 11019 8000 11061 8009
rect 11019 7960 11020 8000
rect 11060 7960 11061 8000
rect 10059 7946 10101 7955
rect 11019 7951 11061 7960
rect 11499 8000 11541 8009
rect 11499 7960 11500 8000
rect 11540 7960 11541 8000
rect 11499 7951 11541 7960
rect 11595 8000 11637 8009
rect 11595 7960 11596 8000
rect 11636 7960 11637 8000
rect 11595 7951 11637 7960
rect 12451 8000 12509 8001
rect 12451 7960 12460 8000
rect 12500 7960 12509 8000
rect 12451 7959 12509 7960
rect 13699 8000 13757 8001
rect 13699 7960 13708 8000
rect 13748 7960 13757 8000
rect 13699 7959 13757 7960
rect 14083 8000 14141 8001
rect 14083 7960 14092 8000
rect 14132 7960 14141 8000
rect 14083 7959 14141 7960
rect 15331 8000 15389 8001
rect 15331 7960 15340 8000
rect 15380 7960 15389 8000
rect 15331 7959 15389 7960
rect 15907 8000 15965 8001
rect 15907 7960 15916 8000
rect 15956 7960 15965 8000
rect 15907 7959 15965 7960
rect 17155 8000 17213 8001
rect 17155 7960 17164 8000
rect 17204 7960 17213 8000
rect 17155 7959 17213 7960
rect 17931 8000 17973 8009
rect 17931 7960 17932 8000
rect 17972 7960 17973 8000
rect 17931 7951 17973 7960
rect 18027 8000 18069 8009
rect 18027 7960 18028 8000
rect 18068 7960 18069 8000
rect 18027 7951 18069 7960
rect 18411 8000 18453 8009
rect 18411 7960 18412 8000
rect 18452 7960 18453 8000
rect 18411 7951 18453 7960
rect 18507 8000 18549 8009
rect 18507 7960 18508 8000
rect 18548 7960 18549 8000
rect 18507 7951 18549 7960
rect 18979 8000 19037 8001
rect 18979 7960 18988 8000
rect 19028 7960 19037 8000
rect 18979 7959 19037 7960
rect 19467 7986 19509 7995
rect 19467 7946 19468 7986
rect 19508 7946 19509 7986
rect 19467 7937 19509 7946
rect 3043 7916 3101 7917
rect 3043 7876 3052 7916
rect 3092 7876 3101 7916
rect 3043 7875 3101 7876
rect 3427 7916 3485 7917
rect 3427 7876 3436 7916
rect 3476 7876 3485 7916
rect 3427 7875 3485 7876
rect 3811 7916 3869 7917
rect 3811 7876 3820 7916
rect 3860 7876 3869 7916
rect 3811 7875 3869 7876
rect 7651 7916 7709 7917
rect 7651 7876 7660 7916
rect 7700 7876 7709 7916
rect 7651 7875 7709 7876
rect 8035 7916 8093 7917
rect 8035 7876 8044 7916
rect 8084 7876 8093 7916
rect 8035 7875 8093 7876
rect 11115 7916 11157 7925
rect 11115 7876 11116 7916
rect 11156 7876 11157 7916
rect 11115 7867 11157 7876
rect 4011 7832 4053 7841
rect 4011 7792 4012 7832
rect 4052 7792 4053 7832
rect 4011 7783 4053 7792
rect 7467 7748 7509 7757
rect 7467 7708 7468 7748
rect 7508 7708 7509 7748
rect 7467 7699 7509 7708
rect 7851 7748 7893 7757
rect 7851 7708 7852 7748
rect 7892 7708 7893 7748
rect 7851 7699 7893 7708
rect 1152 7580 20352 7604
rect 1152 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 20352 7580
rect 1152 7516 20352 7540
rect 2955 7412 2997 7421
rect 2955 7372 2956 7412
rect 2996 7372 2997 7412
rect 2955 7363 2997 7372
rect 9579 7412 9621 7421
rect 9579 7372 9580 7412
rect 9620 7372 9621 7412
rect 9579 7363 9621 7372
rect 11691 7412 11733 7421
rect 11691 7372 11692 7412
rect 11732 7372 11733 7412
rect 11691 7363 11733 7372
rect 20043 7412 20085 7421
rect 20043 7372 20044 7412
rect 20084 7372 20085 7412
rect 20043 7363 20085 7372
rect 18027 7328 18069 7337
rect 18027 7288 18028 7328
rect 18068 7288 18069 7328
rect 18027 7279 18069 7288
rect 3723 7244 3765 7253
rect 3723 7204 3724 7244
rect 3764 7204 3765 7244
rect 3723 7195 3765 7204
rect 3819 7244 3861 7253
rect 3819 7204 3820 7244
rect 3860 7204 3861 7244
rect 3819 7195 3861 7204
rect 8803 7244 8861 7245
rect 8803 7204 8812 7244
rect 8852 7204 8861 7244
rect 8803 7203 8861 7204
rect 9379 7244 9437 7245
rect 9379 7204 9388 7244
rect 9428 7204 9437 7244
rect 9379 7203 9437 7204
rect 9763 7244 9821 7245
rect 9763 7204 9772 7244
rect 9812 7204 9821 7244
rect 9763 7203 9821 7204
rect 15051 7244 15093 7253
rect 15051 7204 15052 7244
rect 15092 7204 15093 7244
rect 15051 7195 15093 7204
rect 1507 7160 1565 7161
rect 1507 7120 1516 7160
rect 1556 7120 1565 7160
rect 1507 7119 1565 7120
rect 2755 7160 2813 7161
rect 2755 7120 2764 7160
rect 2804 7120 2813 7160
rect 2755 7119 2813 7120
rect 3243 7160 3285 7169
rect 3243 7120 3244 7160
rect 3284 7120 3285 7160
rect 3243 7111 3285 7120
rect 3339 7160 3381 7169
rect 4779 7165 4821 7174
rect 3339 7120 3340 7160
rect 3380 7120 3381 7160
rect 3339 7111 3381 7120
rect 4291 7160 4349 7161
rect 4291 7120 4300 7160
rect 4340 7120 4349 7160
rect 4291 7119 4349 7120
rect 4779 7125 4780 7165
rect 4820 7125 4821 7165
rect 6987 7165 7029 7174
rect 16155 7169 16197 7178
rect 4779 7116 4821 7125
rect 5155 7160 5213 7161
rect 5155 7120 5164 7160
rect 5204 7120 5213 7160
rect 5155 7119 5213 7120
rect 6403 7160 6461 7161
rect 6403 7120 6412 7160
rect 6452 7120 6461 7160
rect 6403 7119 6461 7120
rect 6987 7125 6988 7165
rect 7028 7125 7029 7165
rect 6987 7116 7029 7125
rect 7459 7160 7517 7161
rect 7459 7120 7468 7160
rect 7508 7120 7517 7160
rect 7459 7119 7517 7120
rect 7947 7160 7989 7169
rect 7947 7120 7948 7160
rect 7988 7120 7989 7160
rect 7947 7111 7989 7120
rect 8043 7160 8085 7169
rect 8043 7120 8044 7160
rect 8084 7120 8085 7160
rect 8043 7111 8085 7120
rect 8427 7160 8469 7169
rect 8427 7120 8428 7160
rect 8468 7120 8469 7160
rect 8427 7111 8469 7120
rect 8523 7160 8565 7169
rect 8523 7120 8524 7160
rect 8564 7120 8565 7160
rect 8523 7111 8565 7120
rect 10243 7160 10301 7161
rect 10243 7120 10252 7160
rect 10292 7120 10301 7160
rect 10243 7119 10301 7120
rect 11491 7160 11549 7161
rect 11491 7120 11500 7160
rect 11540 7120 11549 7160
rect 11491 7119 11549 7120
rect 12835 7160 12893 7161
rect 12835 7120 12844 7160
rect 12884 7120 12893 7160
rect 12835 7119 12893 7120
rect 14083 7160 14141 7161
rect 14083 7120 14092 7160
rect 14132 7120 14141 7160
rect 14083 7119 14141 7120
rect 14571 7160 14613 7169
rect 14571 7120 14572 7160
rect 14612 7120 14613 7160
rect 14571 7111 14613 7120
rect 14667 7160 14709 7169
rect 14667 7120 14668 7160
rect 14708 7120 14709 7160
rect 14667 7111 14709 7120
rect 15147 7160 15189 7169
rect 15147 7120 15148 7160
rect 15188 7120 15189 7160
rect 15147 7111 15189 7120
rect 15619 7160 15677 7161
rect 15619 7120 15628 7160
rect 15668 7120 15677 7160
rect 16155 7129 16156 7169
rect 16196 7129 16197 7169
rect 16155 7120 16197 7129
rect 16579 7160 16637 7161
rect 16579 7120 16588 7160
rect 16628 7120 16637 7160
rect 15619 7119 15677 7120
rect 16579 7119 16637 7120
rect 17827 7160 17885 7161
rect 17827 7120 17836 7160
rect 17876 7120 17885 7160
rect 17827 7119 17885 7120
rect 18595 7160 18653 7161
rect 18595 7120 18604 7160
rect 18644 7120 18653 7160
rect 18595 7119 18653 7120
rect 19843 7160 19901 7161
rect 19843 7120 19852 7160
rect 19892 7120 19901 7160
rect 19843 7119 19901 7120
rect 4971 7076 5013 7085
rect 4971 7036 4972 7076
rect 5012 7036 5013 7076
rect 4971 7027 5013 7036
rect 14283 7076 14325 7085
rect 14283 7036 14284 7076
rect 14324 7036 14325 7076
rect 14283 7027 14325 7036
rect 6603 6992 6645 7001
rect 6603 6952 6604 6992
rect 6644 6952 6645 6992
rect 6603 6943 6645 6952
rect 6795 6992 6837 7001
rect 6795 6952 6796 6992
rect 6836 6952 6837 6992
rect 6795 6943 6837 6952
rect 9003 6992 9045 7001
rect 9003 6952 9004 6992
rect 9044 6952 9045 6992
rect 9003 6943 9045 6952
rect 9195 6992 9237 7001
rect 9195 6952 9196 6992
rect 9236 6952 9237 6992
rect 9195 6943 9237 6952
rect 16299 6992 16341 7001
rect 16299 6952 16300 6992
rect 16340 6952 16341 6992
rect 16299 6943 16341 6952
rect 1152 6824 20452 6848
rect 1152 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20452 6824
rect 1152 6760 20452 6784
rect 2667 6656 2709 6665
rect 2667 6616 2668 6656
rect 2708 6616 2709 6656
rect 2667 6607 2709 6616
rect 7467 6656 7509 6665
rect 7467 6616 7468 6656
rect 7508 6616 7509 6656
rect 7467 6607 7509 6616
rect 9099 6656 9141 6665
rect 9099 6616 9100 6656
rect 9140 6616 9141 6656
rect 9099 6607 9141 6616
rect 10731 6656 10773 6665
rect 10731 6616 10732 6656
rect 10772 6616 10773 6656
rect 10731 6607 10773 6616
rect 13803 6656 13845 6665
rect 13803 6616 13804 6656
rect 13844 6616 13845 6656
rect 13803 6607 13845 6616
rect 16299 6656 16341 6665
rect 16299 6616 16300 6656
rect 16340 6616 16341 6656
rect 16299 6607 16341 6616
rect 19947 6656 19989 6665
rect 19947 6616 19948 6656
rect 19988 6616 19989 6656
rect 19947 6607 19989 6616
rect 4779 6572 4821 6581
rect 4779 6532 4780 6572
rect 4820 6532 4821 6572
rect 4779 6523 4821 6532
rect 1219 6488 1277 6489
rect 1219 6448 1228 6488
rect 1268 6448 1277 6488
rect 1219 6447 1277 6448
rect 2467 6488 2525 6489
rect 2467 6448 2476 6488
rect 2516 6448 2525 6488
rect 2467 6447 2525 6448
rect 3051 6488 3093 6497
rect 3051 6448 3052 6488
rect 3092 6448 3093 6488
rect 3051 6439 3093 6448
rect 3147 6488 3189 6497
rect 3147 6448 3148 6488
rect 3188 6448 3189 6488
rect 3147 6439 3189 6448
rect 3531 6488 3573 6497
rect 3531 6448 3532 6488
rect 3572 6448 3573 6488
rect 3531 6439 3573 6448
rect 3627 6488 3669 6497
rect 3627 6448 3628 6488
rect 3668 6448 3669 6488
rect 3627 6439 3669 6448
rect 4099 6488 4157 6489
rect 4099 6448 4108 6488
rect 4148 6448 4157 6488
rect 6019 6488 6077 6489
rect 4099 6447 4157 6448
rect 4587 6474 4629 6483
rect 4587 6434 4588 6474
rect 4628 6434 4629 6474
rect 6019 6448 6028 6488
rect 6068 6448 6077 6488
rect 6019 6447 6077 6448
rect 7267 6488 7325 6489
rect 7267 6448 7276 6488
rect 7316 6448 7325 6488
rect 7267 6447 7325 6448
rect 7651 6488 7709 6489
rect 7651 6448 7660 6488
rect 7700 6448 7709 6488
rect 7651 6447 7709 6448
rect 8899 6488 8957 6489
rect 8899 6448 8908 6488
rect 8948 6448 8957 6488
rect 8899 6447 8957 6448
rect 9283 6488 9341 6489
rect 9283 6448 9292 6488
rect 9332 6448 9341 6488
rect 9283 6447 9341 6448
rect 10531 6488 10589 6489
rect 10531 6448 10540 6488
rect 10580 6448 10589 6488
rect 10531 6447 10589 6448
rect 12075 6488 12117 6497
rect 12075 6448 12076 6488
rect 12116 6448 12117 6488
rect 12075 6439 12117 6448
rect 12171 6488 12213 6497
rect 12171 6448 12172 6488
rect 12212 6448 12213 6488
rect 12171 6439 12213 6448
rect 12555 6488 12597 6497
rect 12555 6448 12556 6488
rect 12596 6448 12597 6488
rect 12555 6439 12597 6448
rect 12651 6488 12693 6497
rect 12651 6448 12652 6488
rect 12692 6448 12693 6488
rect 12651 6439 12693 6448
rect 13123 6488 13181 6489
rect 13123 6448 13132 6488
rect 13172 6448 13181 6488
rect 14851 6488 14909 6489
rect 13123 6447 13181 6448
rect 13611 6474 13653 6483
rect 4587 6425 4629 6434
rect 13611 6434 13612 6474
rect 13652 6434 13653 6474
rect 14851 6448 14860 6488
rect 14900 6448 14909 6488
rect 14851 6447 14909 6448
rect 16099 6488 16157 6489
rect 16099 6448 16108 6488
rect 16148 6448 16157 6488
rect 16099 6447 16157 6448
rect 16483 6488 16541 6489
rect 16483 6448 16492 6488
rect 16532 6448 16541 6488
rect 16483 6447 16541 6448
rect 17731 6488 17789 6489
rect 17731 6448 17740 6488
rect 17780 6448 17789 6488
rect 17731 6447 17789 6448
rect 18499 6488 18557 6489
rect 18499 6448 18508 6488
rect 18548 6448 18557 6488
rect 18499 6447 18557 6448
rect 19747 6488 19805 6489
rect 19747 6448 19756 6488
rect 19796 6448 19805 6488
rect 19747 6447 19805 6448
rect 13611 6425 13653 6434
rect 5155 6404 5213 6405
rect 5155 6364 5164 6404
rect 5204 6364 5213 6404
rect 5155 6363 5213 6364
rect 5347 6404 5405 6405
rect 5347 6364 5356 6404
rect 5396 6364 5405 6404
rect 5347 6363 5405 6364
rect 11107 6404 11165 6405
rect 11107 6364 11116 6404
rect 11156 6364 11165 6404
rect 11107 6363 11165 6364
rect 4971 6320 5013 6329
rect 4971 6280 4972 6320
rect 5012 6280 5013 6320
rect 4971 6271 5013 6280
rect 5547 6320 5589 6329
rect 5547 6280 5548 6320
rect 5588 6280 5589 6320
rect 5547 6271 5589 6280
rect 10923 6320 10965 6329
rect 10923 6280 10924 6320
rect 10964 6280 10965 6320
rect 10923 6271 10965 6280
rect 17931 6236 17973 6245
rect 17931 6196 17932 6236
rect 17972 6196 17973 6236
rect 17931 6187 17973 6196
rect 1152 6068 20352 6092
rect 1152 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 20352 6068
rect 1152 6004 20352 6028
rect 1515 5900 1557 5909
rect 1515 5860 1516 5900
rect 1556 5860 1557 5900
rect 1515 5851 1557 5860
rect 1899 5900 1941 5909
rect 1899 5860 1900 5900
rect 1940 5860 1941 5900
rect 1899 5851 1941 5860
rect 3819 5900 3861 5909
rect 3819 5860 3820 5900
rect 3860 5860 3861 5900
rect 3819 5851 3861 5860
rect 4395 5900 4437 5909
rect 4395 5860 4396 5900
rect 4436 5860 4437 5900
rect 4395 5851 4437 5860
rect 6507 5900 6549 5909
rect 6507 5860 6508 5900
rect 6548 5860 6549 5900
rect 6507 5851 6549 5860
rect 11595 5900 11637 5909
rect 11595 5860 11596 5900
rect 11636 5860 11637 5900
rect 11595 5851 11637 5860
rect 13707 5900 13749 5909
rect 13707 5860 13708 5900
rect 13748 5860 13749 5900
rect 13707 5851 13749 5860
rect 4203 5816 4245 5825
rect 4203 5776 4204 5816
rect 4244 5776 4245 5816
rect 4203 5767 4245 5776
rect 9291 5816 9333 5825
rect 9291 5776 9292 5816
rect 9332 5776 9333 5816
rect 9291 5767 9333 5776
rect 11779 5743 11837 5744
rect 1699 5732 1757 5733
rect 1699 5692 1708 5732
rect 1748 5692 1757 5732
rect 1699 5691 1757 5692
rect 2083 5732 2141 5733
rect 2083 5692 2092 5732
rect 2132 5692 2141 5732
rect 2083 5691 2141 5692
rect 4003 5732 4061 5733
rect 4003 5692 4012 5732
rect 4052 5692 4061 5732
rect 4003 5691 4061 5692
rect 4579 5732 4637 5733
rect 4579 5692 4588 5732
rect 4628 5692 4637 5732
rect 4579 5691 4637 5692
rect 4875 5732 4917 5741
rect 4875 5692 4876 5732
rect 4916 5692 4917 5732
rect 4875 5683 4917 5692
rect 7275 5732 7317 5741
rect 7275 5692 7276 5732
rect 7316 5692 7317 5732
rect 7275 5683 7317 5692
rect 7371 5732 7413 5741
rect 7371 5692 7372 5732
rect 7412 5692 7413 5732
rect 7371 5683 7413 5692
rect 8899 5732 8957 5733
rect 8899 5692 8908 5732
rect 8948 5692 8957 5732
rect 8899 5691 8957 5692
rect 10251 5732 10293 5741
rect 10251 5692 10252 5732
rect 10292 5692 10293 5732
rect 11779 5703 11788 5743
rect 11828 5703 11837 5743
rect 11779 5702 11837 5703
rect 14475 5732 14517 5741
rect 10251 5683 10293 5692
rect 14475 5692 14476 5732
rect 14516 5692 14517 5732
rect 14475 5683 14517 5692
rect 14571 5732 14613 5741
rect 14571 5692 14572 5732
rect 14612 5692 14613 5732
rect 14571 5683 14613 5692
rect 17259 5732 17301 5741
rect 17259 5692 17260 5732
rect 17300 5692 17301 5732
rect 17259 5683 17301 5692
rect 17355 5732 17397 5741
rect 17355 5692 17356 5732
rect 17396 5692 17397 5732
rect 17355 5683 17397 5692
rect 2371 5648 2429 5649
rect 2371 5608 2380 5648
rect 2420 5608 2429 5648
rect 2371 5607 2429 5608
rect 3619 5648 3677 5649
rect 3619 5608 3628 5648
rect 3668 5608 3677 5648
rect 3619 5607 3677 5608
rect 5059 5648 5117 5649
rect 5059 5608 5068 5648
rect 5108 5608 5117 5648
rect 5059 5607 5117 5608
rect 6307 5648 6365 5649
rect 6307 5608 6316 5648
rect 6356 5608 6365 5648
rect 6307 5607 6365 5608
rect 6795 5648 6837 5657
rect 6795 5608 6796 5648
rect 6836 5608 6837 5648
rect 6795 5599 6837 5608
rect 6891 5648 6933 5657
rect 8331 5653 8373 5662
rect 6891 5608 6892 5648
rect 6932 5608 6933 5648
rect 6891 5599 6933 5608
rect 7843 5648 7901 5649
rect 7843 5608 7852 5648
rect 7892 5608 7901 5648
rect 7843 5607 7901 5608
rect 8331 5613 8332 5653
rect 8372 5613 8373 5653
rect 8331 5604 8373 5613
rect 9675 5648 9717 5657
rect 9675 5608 9676 5648
rect 9716 5608 9717 5648
rect 9675 5599 9717 5608
rect 9771 5648 9813 5657
rect 9771 5608 9772 5648
rect 9812 5608 9813 5648
rect 9771 5599 9813 5608
rect 10155 5648 10197 5657
rect 11211 5653 11253 5662
rect 15579 5657 15621 5666
rect 18315 5662 18357 5671
rect 10155 5608 10156 5648
rect 10196 5608 10197 5648
rect 10155 5599 10197 5608
rect 10723 5648 10781 5649
rect 10723 5608 10732 5648
rect 10772 5608 10781 5648
rect 10723 5607 10781 5608
rect 11211 5613 11212 5653
rect 11252 5613 11253 5653
rect 11211 5604 11253 5613
rect 12259 5648 12317 5649
rect 12259 5608 12268 5648
rect 12308 5608 12317 5648
rect 12259 5607 12317 5608
rect 13507 5648 13565 5649
rect 13507 5608 13516 5648
rect 13556 5608 13565 5648
rect 13507 5607 13565 5608
rect 13995 5648 14037 5657
rect 13995 5608 13996 5648
rect 14036 5608 14037 5648
rect 13995 5599 14037 5608
rect 14091 5648 14133 5657
rect 14091 5608 14092 5648
rect 14132 5608 14133 5648
rect 14091 5599 14133 5608
rect 15043 5648 15101 5649
rect 15043 5608 15052 5648
rect 15092 5608 15101 5648
rect 15579 5617 15580 5657
rect 15620 5617 15621 5657
rect 15579 5608 15621 5617
rect 16779 5648 16821 5657
rect 16779 5608 16780 5648
rect 16820 5608 16821 5648
rect 15043 5607 15101 5608
rect 16779 5599 16821 5608
rect 16875 5648 16917 5657
rect 16875 5608 16876 5648
rect 16916 5608 16917 5648
rect 16875 5599 16917 5608
rect 17827 5648 17885 5649
rect 17827 5608 17836 5648
rect 17876 5608 17885 5648
rect 18315 5622 18316 5662
rect 18356 5622 18357 5662
rect 18315 5613 18357 5622
rect 18691 5648 18749 5649
rect 17827 5607 17885 5608
rect 18691 5608 18700 5648
rect 18740 5608 18749 5648
rect 18691 5607 18749 5608
rect 19939 5648 19997 5649
rect 19939 5608 19948 5648
rect 19988 5608 19997 5648
rect 19939 5607 19997 5608
rect 8523 5564 8565 5573
rect 8523 5524 8524 5564
rect 8564 5524 8565 5564
rect 8523 5515 8565 5524
rect 11403 5564 11445 5573
rect 11403 5524 11404 5564
rect 11444 5524 11445 5564
rect 11403 5515 11445 5524
rect 18507 5564 18549 5573
rect 18507 5524 18508 5564
rect 18548 5524 18549 5564
rect 18507 5515 18549 5524
rect 9099 5480 9141 5489
rect 9099 5440 9100 5480
rect 9140 5440 9141 5480
rect 9099 5431 9141 5440
rect 11971 5480 12029 5481
rect 11971 5440 11980 5480
rect 12020 5440 12029 5480
rect 11971 5439 12029 5440
rect 15723 5480 15765 5489
rect 15723 5440 15724 5480
rect 15764 5440 15765 5480
rect 15723 5431 15765 5440
rect 20139 5480 20181 5489
rect 20139 5440 20140 5480
rect 20180 5440 20181 5480
rect 20139 5431 20181 5440
rect 1152 5312 20452 5336
rect 1152 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20452 5312
rect 1152 5248 20452 5272
rect 4779 5144 4821 5153
rect 4779 5104 4780 5144
rect 4820 5104 4821 5144
rect 4779 5095 4821 5104
rect 7179 5144 7221 5153
rect 7179 5104 7180 5144
rect 7220 5104 7221 5144
rect 7179 5095 7221 5104
rect 9003 5144 9045 5153
rect 9003 5104 9004 5144
rect 9044 5104 9045 5144
rect 9003 5095 9045 5104
rect 13995 5144 14037 5153
rect 13995 5104 13996 5144
rect 14036 5104 14037 5144
rect 13995 5095 14037 5104
rect 15723 5144 15765 5153
rect 15723 5104 15724 5144
rect 15764 5104 15765 5144
rect 15723 5095 15765 5104
rect 17355 5144 17397 5153
rect 17355 5104 17356 5144
rect 17396 5104 17397 5144
rect 17355 5095 17397 5104
rect 2667 5060 2709 5069
rect 2667 5020 2668 5060
rect 2708 5020 2709 5060
rect 2667 5011 2709 5020
rect 4299 5060 4341 5069
rect 4299 5020 4300 5060
rect 4340 5020 4341 5060
rect 4299 5011 4341 5020
rect 12267 5060 12309 5069
rect 12267 5020 12268 5060
rect 12308 5020 12309 5060
rect 12267 5011 12309 5020
rect 18315 5060 18357 5069
rect 18315 5020 18316 5060
rect 18356 5020 18357 5060
rect 18315 5011 18357 5020
rect 1219 4976 1277 4977
rect 1219 4936 1228 4976
rect 1268 4936 1277 4976
rect 1219 4935 1277 4936
rect 2467 4976 2525 4977
rect 2467 4936 2476 4976
rect 2516 4936 2525 4976
rect 2467 4935 2525 4936
rect 2851 4976 2909 4977
rect 2851 4936 2860 4976
rect 2900 4936 2909 4976
rect 2851 4935 2909 4936
rect 4099 4976 4157 4977
rect 4099 4936 4108 4976
rect 4148 4936 4157 4976
rect 5443 4976 5501 4977
rect 4099 4935 4157 4936
rect 4923 4934 4965 4943
rect 5443 4936 5452 4976
rect 5492 4936 5501 4976
rect 6507 4976 6549 4985
rect 5443 4935 5501 4936
rect 6411 4957 6453 4966
rect 4923 4894 4924 4934
rect 4964 4894 4965 4934
rect 6411 4917 6412 4957
rect 6452 4917 6453 4957
rect 6507 4936 6508 4976
rect 6548 4936 6549 4976
rect 6507 4927 6549 4936
rect 7555 4976 7613 4977
rect 7555 4936 7564 4976
rect 7604 4936 7613 4976
rect 7555 4935 7613 4936
rect 8803 4976 8861 4977
rect 8803 4936 8812 4976
rect 8852 4936 8861 4976
rect 8803 4935 8861 4936
rect 9187 4976 9245 4977
rect 9187 4936 9196 4976
rect 9236 4936 9245 4976
rect 9187 4935 9245 4936
rect 10435 4976 10493 4977
rect 10435 4936 10444 4976
rect 10484 4936 10493 4976
rect 10435 4935 10493 4936
rect 10819 4976 10877 4977
rect 10819 4936 10828 4976
rect 10868 4936 10877 4976
rect 10819 4935 10877 4936
rect 12067 4976 12125 4977
rect 12067 4936 12076 4976
rect 12116 4936 12125 4976
rect 12067 4935 12125 4936
rect 12547 4976 12605 4977
rect 12547 4936 12556 4976
rect 12596 4936 12605 4976
rect 12547 4935 12605 4936
rect 13795 4976 13853 4977
rect 13795 4936 13804 4976
rect 13844 4936 13853 4976
rect 13795 4935 13853 4936
rect 14275 4976 14333 4977
rect 14275 4936 14284 4976
rect 14324 4936 14333 4976
rect 14275 4935 14333 4936
rect 15523 4976 15581 4977
rect 15523 4936 15532 4976
rect 15572 4936 15581 4976
rect 15523 4935 15581 4936
rect 15907 4976 15965 4977
rect 15907 4936 15916 4976
rect 15956 4936 15965 4976
rect 15907 4935 15965 4936
rect 17155 4976 17213 4977
rect 17155 4936 17164 4976
rect 17204 4936 17213 4976
rect 18979 4976 19037 4977
rect 17155 4935 17213 4936
rect 18507 4962 18549 4971
rect 6411 4908 6453 4917
rect 18507 4922 18508 4962
rect 18548 4922 18549 4962
rect 18979 4936 18988 4976
rect 19028 4936 19037 4976
rect 18979 4935 19037 4936
rect 19467 4976 19509 4985
rect 19467 4936 19468 4976
rect 19508 4936 19509 4976
rect 19467 4927 19509 4936
rect 19563 4976 19605 4985
rect 19563 4936 19564 4976
rect 19604 4936 19605 4976
rect 19563 4927 19605 4936
rect 19947 4976 19989 4985
rect 19947 4936 19948 4976
rect 19988 4936 19989 4976
rect 19947 4927 19989 4936
rect 20043 4976 20085 4985
rect 20043 4936 20044 4976
rect 20084 4936 20085 4976
rect 20043 4927 20085 4936
rect 18507 4913 18549 4922
rect 4923 4885 4965 4894
rect 5931 4892 5973 4901
rect 5931 4852 5932 4892
rect 5972 4852 5973 4892
rect 5931 4843 5973 4852
rect 6027 4892 6069 4901
rect 6027 4852 6028 4892
rect 6068 4852 6069 4892
rect 6027 4843 6069 4852
rect 6979 4892 7037 4893
rect 6979 4852 6988 4892
rect 7028 4852 7037 4892
rect 6979 4851 7037 4852
rect 7363 4892 7421 4893
rect 7363 4852 7372 4892
rect 7412 4852 7421 4892
rect 7363 4851 7421 4852
rect 4587 4808 4629 4817
rect 4587 4768 4588 4808
rect 4628 4768 4629 4808
rect 4587 4759 4629 4768
rect 6795 4808 6837 4817
rect 6795 4768 6796 4808
rect 6836 4768 6837 4808
rect 6795 4759 6837 4768
rect 10635 4724 10677 4733
rect 10635 4684 10636 4724
rect 10676 4684 10677 4724
rect 10635 4675 10677 4684
rect 1152 4556 20352 4580
rect 1152 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 20352 4556
rect 1152 4492 20352 4516
rect 2667 4388 2709 4397
rect 2667 4348 2668 4388
rect 2708 4348 2709 4388
rect 2667 4339 2709 4348
rect 4587 4388 4629 4397
rect 4587 4348 4588 4388
rect 4628 4348 4629 4388
rect 4587 4339 4629 4348
rect 6795 4388 6837 4397
rect 6795 4348 6796 4388
rect 6836 4348 6837 4388
rect 6795 4339 6837 4348
rect 2859 4304 2901 4313
rect 2859 4264 2860 4304
rect 2900 4264 2901 4304
rect 2859 4255 2901 4264
rect 4963 4220 5021 4221
rect 4963 4180 4972 4220
rect 5012 4180 5021 4220
rect 4963 4179 5021 4180
rect 9771 4220 9813 4229
rect 9771 4180 9772 4220
rect 9812 4180 9813 4220
rect 9771 4171 9813 4180
rect 9867 4220 9909 4229
rect 9867 4180 9868 4220
rect 9908 4180 9909 4220
rect 9867 4171 9909 4180
rect 10819 4220 10877 4221
rect 10819 4180 10828 4220
rect 10868 4180 10877 4220
rect 10819 4179 10877 4180
rect 11203 4220 11261 4221
rect 11203 4180 11212 4220
rect 11252 4180 11261 4220
rect 11203 4179 11261 4180
rect 11587 4220 11645 4221
rect 11587 4180 11596 4220
rect 11636 4180 11645 4220
rect 11587 4179 11645 4180
rect 18315 4220 18357 4229
rect 18315 4180 18316 4220
rect 18356 4180 18357 4220
rect 18315 4171 18357 4180
rect 18411 4220 18453 4229
rect 18411 4180 18412 4220
rect 18452 4180 18453 4220
rect 18411 4171 18453 4180
rect 8763 4145 8805 4154
rect 19419 4145 19461 4154
rect 1219 4136 1277 4137
rect 1219 4096 1228 4136
rect 1268 4096 1277 4136
rect 1219 4095 1277 4096
rect 2467 4136 2525 4137
rect 2467 4096 2476 4136
rect 2516 4096 2525 4136
rect 2467 4095 2525 4096
rect 3139 4136 3197 4137
rect 3139 4096 3148 4136
rect 3188 4096 3197 4136
rect 3139 4095 3197 4096
rect 4387 4136 4445 4137
rect 4387 4096 4396 4136
rect 4436 4096 4445 4136
rect 4387 4095 4445 4096
rect 5347 4136 5405 4137
rect 5347 4096 5356 4136
rect 5396 4096 5405 4136
rect 5347 4095 5405 4096
rect 6595 4136 6653 4137
rect 6595 4096 6604 4136
rect 6644 4096 6653 4136
rect 6595 4095 6653 4096
rect 6979 4136 7037 4137
rect 6979 4096 6988 4136
rect 7028 4096 7037 4136
rect 6979 4095 7037 4096
rect 8227 4136 8285 4137
rect 8227 4096 8236 4136
rect 8276 4096 8285 4136
rect 8763 4105 8764 4145
rect 8804 4105 8805 4145
rect 8763 4096 8805 4105
rect 9283 4136 9341 4137
rect 9283 4096 9292 4136
rect 9332 4096 9341 4136
rect 8227 4095 8285 4096
rect 9283 4095 9341 4096
rect 10251 4136 10293 4145
rect 10251 4096 10252 4136
rect 10292 4096 10293 4136
rect 11875 4136 11933 4137
rect 10251 4087 10293 4096
rect 10347 4116 10389 4125
rect 10347 4076 10348 4116
rect 10388 4076 10389 4116
rect 11875 4096 11884 4136
rect 11924 4096 11933 4136
rect 11875 4095 11933 4096
rect 13123 4136 13181 4137
rect 13123 4096 13132 4136
rect 13172 4096 13181 4136
rect 13123 4095 13181 4096
rect 13699 4136 13757 4137
rect 13699 4096 13708 4136
rect 13748 4096 13757 4136
rect 13699 4095 13757 4096
rect 14947 4136 15005 4137
rect 14947 4096 14956 4136
rect 14996 4096 15005 4136
rect 14947 4095 15005 4096
rect 15331 4136 15389 4137
rect 15331 4096 15340 4136
rect 15380 4096 15389 4136
rect 15331 4095 15389 4096
rect 16579 4136 16637 4137
rect 16579 4096 16588 4136
rect 16628 4096 16637 4136
rect 16579 4095 16637 4096
rect 17835 4136 17877 4145
rect 17835 4096 17836 4136
rect 17876 4096 17877 4136
rect 17835 4087 17877 4096
rect 17931 4136 17973 4145
rect 17931 4096 17932 4136
rect 17972 4096 17973 4136
rect 17931 4087 17973 4096
rect 18883 4136 18941 4137
rect 18883 4096 18892 4136
rect 18932 4096 18941 4136
rect 19419 4105 19420 4145
rect 19460 4105 19461 4145
rect 19419 4096 19461 4105
rect 18883 4095 18941 4096
rect 10347 4067 10389 4076
rect 8427 4052 8469 4061
rect 8427 4012 8428 4052
rect 8468 4012 8469 4052
rect 8427 4003 8469 4012
rect 5163 3968 5205 3977
rect 5163 3928 5164 3968
rect 5204 3928 5205 3968
rect 5163 3919 5205 3928
rect 8619 3968 8661 3977
rect 8619 3928 8620 3968
rect 8660 3928 8661 3968
rect 8619 3919 8661 3928
rect 10635 3968 10677 3977
rect 10635 3928 10636 3968
rect 10676 3928 10677 3968
rect 10635 3919 10677 3928
rect 11019 3968 11061 3977
rect 11019 3928 11020 3968
rect 11060 3928 11061 3968
rect 11019 3919 11061 3928
rect 11403 3968 11445 3977
rect 11403 3928 11404 3968
rect 11444 3928 11445 3968
rect 11403 3919 11445 3928
rect 13323 3968 13365 3977
rect 13323 3928 13324 3968
rect 13364 3928 13365 3968
rect 13323 3919 13365 3928
rect 15147 3968 15189 3977
rect 15147 3928 15148 3968
rect 15188 3928 15189 3968
rect 15147 3919 15189 3928
rect 16779 3968 16821 3977
rect 16779 3928 16780 3968
rect 16820 3928 16821 3968
rect 16779 3919 16821 3928
rect 19563 3968 19605 3977
rect 19563 3928 19564 3968
rect 19604 3928 19605 3968
rect 19563 3919 19605 3928
rect 1152 3800 20452 3824
rect 1152 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20452 3800
rect 1152 3736 20452 3760
rect 1515 3632 1557 3641
rect 1515 3592 1516 3632
rect 1556 3592 1557 3632
rect 1515 3583 1557 3592
rect 2091 3632 2133 3641
rect 2091 3592 2092 3632
rect 2132 3592 2133 3632
rect 2091 3583 2133 3592
rect 3723 3632 3765 3641
rect 3723 3592 3724 3632
rect 3764 3592 3765 3632
rect 3723 3583 3765 3592
rect 5835 3632 5877 3641
rect 5835 3592 5836 3632
rect 5876 3592 5877 3632
rect 5835 3583 5877 3592
rect 10347 3632 10389 3641
rect 10347 3592 10348 3632
rect 10388 3592 10389 3632
rect 10347 3583 10389 3592
rect 13515 3632 13557 3641
rect 13515 3592 13516 3632
rect 13556 3592 13557 3632
rect 13515 3583 13557 3592
rect 16203 3632 16245 3641
rect 16203 3592 16204 3632
rect 16244 3592 16245 3632
rect 16203 3583 16245 3592
rect 19659 3632 19701 3641
rect 19659 3592 19660 3632
rect 19700 3592 19701 3632
rect 19659 3583 19701 3592
rect 1323 3548 1365 3557
rect 1323 3508 1324 3548
rect 1364 3508 1365 3548
rect 1323 3499 1365 3508
rect 2275 3464 2333 3465
rect 2275 3424 2284 3464
rect 2324 3424 2333 3464
rect 2275 3423 2333 3424
rect 3523 3464 3581 3465
rect 3523 3424 3532 3464
rect 3572 3424 3581 3464
rect 3523 3423 3581 3424
rect 4107 3464 4149 3473
rect 4107 3424 4108 3464
rect 4148 3424 4149 3464
rect 4107 3415 4149 3424
rect 4203 3464 4245 3473
rect 4203 3424 4204 3464
rect 4244 3424 4245 3464
rect 4203 3415 4245 3424
rect 5155 3464 5213 3465
rect 5155 3424 5164 3464
rect 5204 3424 5213 3464
rect 6211 3464 6269 3465
rect 5155 3423 5213 3424
rect 5643 3450 5685 3459
rect 5643 3410 5644 3450
rect 5684 3410 5685 3450
rect 6211 3424 6220 3464
rect 6260 3424 6269 3464
rect 6211 3423 6269 3424
rect 7459 3464 7517 3465
rect 7459 3424 7468 3464
rect 7508 3424 7517 3464
rect 7459 3423 7517 3424
rect 8619 3464 8661 3473
rect 8619 3424 8620 3464
rect 8660 3424 8661 3464
rect 8619 3415 8661 3424
rect 8715 3464 8757 3473
rect 8715 3424 8716 3464
rect 8756 3424 8757 3464
rect 8715 3415 8757 3424
rect 9099 3464 9141 3473
rect 9099 3424 9100 3464
rect 9140 3424 9141 3464
rect 9099 3415 9141 3424
rect 9667 3464 9725 3465
rect 9667 3424 9676 3464
rect 9716 3424 9725 3464
rect 11787 3464 11829 3473
rect 9667 3423 9725 3424
rect 10203 3422 10245 3431
rect 5643 3401 5685 3410
rect 1699 3380 1757 3381
rect 1699 3340 1708 3380
rect 1748 3340 1757 3380
rect 1699 3339 1757 3340
rect 1891 3380 1949 3381
rect 1891 3340 1900 3380
rect 1940 3340 1949 3380
rect 1891 3339 1949 3340
rect 4587 3380 4629 3389
rect 4587 3340 4588 3380
rect 4628 3340 4629 3380
rect 4587 3331 4629 3340
rect 4683 3380 4725 3389
rect 4683 3340 4684 3380
rect 4724 3340 4725 3380
rect 4683 3331 4725 3340
rect 7747 3380 7805 3381
rect 7747 3340 7756 3380
rect 7796 3340 7805 3380
rect 7747 3339 7805 3340
rect 8131 3380 8189 3381
rect 8131 3340 8140 3380
rect 8180 3340 8189 3380
rect 8131 3339 8189 3340
rect 9195 3380 9237 3389
rect 9195 3340 9196 3380
rect 9236 3340 9237 3380
rect 10203 3382 10204 3422
rect 10244 3382 10245 3422
rect 11787 3424 11788 3464
rect 11828 3424 11829 3464
rect 11787 3415 11829 3424
rect 11883 3464 11925 3473
rect 11883 3424 11884 3464
rect 11924 3424 11925 3464
rect 11883 3415 11925 3424
rect 12363 3464 12405 3473
rect 12363 3424 12364 3464
rect 12404 3424 12405 3464
rect 12363 3415 12405 3424
rect 12835 3464 12893 3465
rect 12835 3424 12844 3464
rect 12884 3424 12893 3464
rect 12835 3423 12893 3424
rect 13323 3459 13365 3468
rect 13323 3419 13324 3459
rect 13364 3419 13365 3459
rect 13323 3410 13365 3419
rect 14475 3464 14517 3473
rect 14475 3424 14476 3464
rect 14516 3424 14517 3464
rect 14475 3415 14517 3424
rect 14571 3464 14613 3473
rect 14571 3424 14572 3464
rect 14612 3424 14613 3464
rect 14571 3415 14613 3424
rect 14955 3464 14997 3473
rect 14955 3424 14956 3464
rect 14996 3424 14997 3464
rect 14955 3415 14997 3424
rect 15051 3464 15093 3473
rect 15051 3424 15052 3464
rect 15092 3424 15093 3464
rect 15051 3415 15093 3424
rect 15523 3464 15581 3465
rect 15523 3424 15532 3464
rect 15572 3424 15581 3464
rect 17931 3464 17973 3473
rect 15523 3423 15581 3424
rect 16059 3422 16101 3431
rect 10203 3373 10245 3382
rect 10531 3380 10589 3381
rect 9195 3331 9237 3340
rect 10531 3340 10540 3380
rect 10580 3340 10589 3380
rect 10531 3339 10589 3340
rect 10915 3380 10973 3381
rect 10915 3340 10924 3380
rect 10964 3340 10973 3380
rect 10915 3339 10973 3340
rect 11491 3380 11549 3381
rect 11491 3340 11500 3380
rect 11540 3340 11549 3380
rect 11491 3339 11549 3340
rect 12267 3380 12309 3389
rect 16059 3382 16060 3422
rect 16100 3382 16101 3422
rect 17931 3424 17932 3464
rect 17972 3424 17973 3464
rect 17931 3415 17973 3424
rect 18027 3464 18069 3473
rect 18027 3424 18028 3464
rect 18068 3424 18069 3464
rect 18027 3415 18069 3424
rect 18507 3464 18549 3473
rect 18507 3424 18508 3464
rect 18548 3424 18549 3464
rect 18507 3415 18549 3424
rect 18979 3464 19037 3465
rect 18979 3424 18988 3464
rect 19028 3424 19037 3464
rect 18979 3423 19037 3424
rect 19515 3422 19557 3431
rect 12267 3340 12268 3380
rect 12308 3340 12309 3380
rect 12267 3331 12309 3340
rect 13699 3380 13757 3381
rect 13699 3340 13708 3380
rect 13748 3340 13757 3380
rect 16059 3373 16101 3382
rect 16579 3380 16637 3381
rect 13699 3339 13757 3340
rect 16579 3340 16588 3380
rect 16628 3340 16637 3380
rect 16579 3339 16637 3340
rect 16963 3380 17021 3381
rect 16963 3340 16972 3380
rect 17012 3340 17021 3380
rect 16963 3339 17021 3340
rect 17347 3380 17405 3381
rect 17347 3340 17356 3380
rect 17396 3340 17405 3380
rect 17347 3339 17405 3340
rect 18411 3380 18453 3389
rect 18411 3340 18412 3380
rect 18452 3340 18453 3380
rect 19515 3382 19516 3422
rect 19556 3382 19557 3422
rect 19515 3373 19557 3382
rect 18411 3331 18453 3340
rect 6027 3212 6069 3221
rect 6027 3172 6028 3212
rect 6068 3172 6069 3212
rect 6027 3163 6069 3172
rect 7947 3212 7989 3221
rect 7947 3172 7948 3212
rect 7988 3172 7989 3212
rect 7947 3163 7989 3172
rect 8331 3212 8373 3221
rect 8331 3172 8332 3212
rect 8372 3172 8373 3212
rect 8331 3163 8373 3172
rect 10731 3212 10773 3221
rect 10731 3172 10732 3212
rect 10772 3172 10773 3212
rect 10731 3163 10773 3172
rect 11115 3212 11157 3221
rect 11115 3172 11116 3212
rect 11156 3172 11157 3212
rect 11115 3163 11157 3172
rect 11307 3212 11349 3221
rect 11307 3172 11308 3212
rect 11348 3172 11349 3212
rect 11307 3163 11349 3172
rect 13899 3212 13941 3221
rect 13899 3172 13900 3212
rect 13940 3172 13941 3212
rect 13899 3163 13941 3172
rect 16395 3212 16437 3221
rect 16395 3172 16396 3212
rect 16436 3172 16437 3212
rect 16395 3163 16437 3172
rect 16779 3212 16821 3221
rect 16779 3172 16780 3212
rect 16820 3172 16821 3212
rect 16779 3163 16821 3172
rect 17163 3212 17205 3221
rect 17163 3172 17164 3212
rect 17204 3172 17205 3212
rect 17163 3163 17205 3172
rect 1152 3044 20352 3068
rect 1152 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 20352 3044
rect 1152 2980 20352 3004
rect 3435 2876 3477 2885
rect 3435 2836 3436 2876
rect 3476 2836 3477 2876
rect 3435 2827 3477 2836
rect 5067 2876 5109 2885
rect 5067 2836 5068 2876
rect 5108 2836 5109 2876
rect 5067 2827 5109 2836
rect 6699 2876 6741 2885
rect 6699 2836 6700 2876
rect 6740 2836 6741 2876
rect 6699 2827 6741 2836
rect 9483 2876 9525 2885
rect 9483 2836 9484 2876
rect 9524 2836 9525 2876
rect 9483 2827 9525 2836
rect 11499 2876 11541 2885
rect 11499 2836 11500 2876
rect 11540 2836 11541 2876
rect 11499 2827 11541 2836
rect 18507 2876 18549 2885
rect 18507 2836 18508 2876
rect 18548 2836 18549 2876
rect 18507 2827 18549 2836
rect 20235 2876 20277 2885
rect 20235 2836 20236 2876
rect 20276 2836 20277 2876
rect 20235 2827 20277 2836
rect 2859 2792 2901 2801
rect 2859 2752 2860 2792
rect 2900 2752 2901 2792
rect 2859 2743 2901 2752
rect 9099 2792 9141 2801
rect 9099 2752 9100 2792
rect 9140 2752 9141 2792
rect 9099 2743 9141 2752
rect 9867 2792 9909 2801
rect 9867 2752 9868 2792
rect 9908 2752 9909 2792
rect 9867 2743 9909 2752
rect 13707 2792 13749 2801
rect 13707 2752 13708 2792
rect 13748 2752 13749 2792
rect 13707 2743 13749 2752
rect 3235 2708 3293 2709
rect 3235 2668 3244 2708
rect 3284 2668 3293 2708
rect 3235 2667 3293 2668
rect 7563 2708 7605 2717
rect 7563 2668 7564 2708
rect 7604 2668 7605 2708
rect 3619 2666 3677 2667
rect 3619 2626 3628 2666
rect 3668 2626 3677 2666
rect 7563 2659 7605 2668
rect 8899 2708 8957 2709
rect 8899 2668 8908 2708
rect 8948 2668 8957 2708
rect 8899 2667 8957 2668
rect 9283 2708 9341 2709
rect 9283 2668 9292 2708
rect 9332 2668 9341 2708
rect 9283 2667 9341 2668
rect 9667 2708 9725 2709
rect 9667 2668 9676 2708
rect 9716 2668 9725 2708
rect 9667 2667 9725 2668
rect 12267 2708 12309 2717
rect 12267 2668 12268 2708
rect 12308 2668 12309 2708
rect 12267 2659 12309 2668
rect 12363 2708 12405 2717
rect 12363 2668 12364 2708
rect 12404 2668 12405 2708
rect 12363 2659 12405 2668
rect 14179 2708 14237 2709
rect 14179 2668 14188 2708
rect 14228 2668 14237 2708
rect 14179 2667 14237 2668
rect 14563 2708 14621 2709
rect 14563 2668 14572 2708
rect 14612 2668 14621 2708
rect 14563 2667 14621 2668
rect 15627 2708 15669 2717
rect 15627 2668 15628 2708
rect 15668 2668 15669 2708
rect 15627 2659 15669 2668
rect 15723 2708 15765 2717
rect 15723 2668 15724 2708
rect 15764 2668 15765 2708
rect 15723 2659 15765 2668
rect 8523 2638 8565 2647
rect 16683 2638 16725 2647
rect 3619 2625 3677 2626
rect 1411 2624 1469 2625
rect 1411 2584 1420 2624
rect 1460 2584 1469 2624
rect 1411 2583 1469 2584
rect 2659 2624 2717 2625
rect 2659 2584 2668 2624
rect 2708 2584 2717 2624
rect 2659 2583 2717 2584
rect 4867 2624 4925 2625
rect 4867 2584 4876 2624
rect 4916 2584 4925 2624
rect 4867 2583 4925 2584
rect 5251 2624 5309 2625
rect 5251 2584 5260 2624
rect 5300 2584 5309 2624
rect 5251 2583 5309 2584
rect 6499 2624 6557 2625
rect 6499 2584 6508 2624
rect 6548 2584 6557 2624
rect 6499 2583 6557 2584
rect 6987 2624 7029 2633
rect 6987 2584 6988 2624
rect 7028 2584 7029 2624
rect 6987 2575 7029 2584
rect 7083 2624 7125 2633
rect 7083 2584 7084 2624
rect 7124 2584 7125 2624
rect 7083 2575 7125 2584
rect 7467 2624 7509 2633
rect 7467 2584 7468 2624
rect 7508 2584 7509 2624
rect 7467 2575 7509 2584
rect 8035 2624 8093 2625
rect 8035 2584 8044 2624
rect 8084 2584 8093 2624
rect 8523 2598 8524 2638
rect 8564 2598 8565 2638
rect 8523 2589 8565 2598
rect 10051 2624 10109 2625
rect 8035 2583 8093 2584
rect 10051 2584 10060 2624
rect 10100 2584 10109 2624
rect 10051 2583 10109 2584
rect 11299 2624 11357 2625
rect 11299 2584 11308 2624
rect 11348 2584 11357 2624
rect 11299 2583 11357 2584
rect 11787 2624 11829 2633
rect 11787 2584 11788 2624
rect 11828 2584 11829 2624
rect 11787 2575 11829 2584
rect 11883 2624 11925 2633
rect 13323 2629 13365 2638
rect 11883 2584 11884 2624
rect 11924 2584 11925 2624
rect 11883 2575 11925 2584
rect 12835 2624 12893 2625
rect 12835 2584 12844 2624
rect 12884 2584 12893 2624
rect 12835 2583 12893 2584
rect 13323 2589 13324 2629
rect 13364 2589 13365 2629
rect 13323 2580 13365 2589
rect 15147 2624 15189 2633
rect 15147 2584 15148 2624
rect 15188 2584 15189 2624
rect 15147 2575 15189 2584
rect 15243 2624 15285 2633
rect 15243 2584 15244 2624
rect 15284 2584 15285 2624
rect 15243 2575 15285 2584
rect 16195 2624 16253 2625
rect 16195 2584 16204 2624
rect 16244 2584 16253 2624
rect 16683 2598 16684 2638
rect 16724 2598 16725 2638
rect 16683 2589 16725 2598
rect 17059 2624 17117 2625
rect 16195 2583 16253 2584
rect 17059 2584 17068 2624
rect 17108 2584 17117 2624
rect 17059 2583 17117 2584
rect 18307 2624 18365 2625
rect 18307 2584 18316 2624
rect 18356 2584 18365 2624
rect 18307 2583 18365 2584
rect 18787 2624 18845 2625
rect 18787 2584 18796 2624
rect 18836 2584 18845 2624
rect 18787 2583 18845 2584
rect 20035 2624 20093 2625
rect 20035 2584 20044 2624
rect 20084 2584 20093 2624
rect 20035 2583 20093 2584
rect 8715 2540 8757 2549
rect 8715 2500 8716 2540
rect 8756 2500 8757 2540
rect 8715 2491 8757 2500
rect 13515 2540 13557 2549
rect 13515 2500 13516 2540
rect 13556 2500 13557 2540
rect 13515 2491 13557 2500
rect 16875 2540 16917 2549
rect 16875 2500 16876 2540
rect 16916 2500 16917 2540
rect 16875 2491 16917 2500
rect 13995 2456 14037 2465
rect 13995 2416 13996 2456
rect 14036 2416 14037 2456
rect 13995 2407 14037 2416
rect 14379 2456 14421 2465
rect 14379 2416 14380 2456
rect 14420 2416 14421 2456
rect 14379 2407 14421 2416
rect 1152 2288 20452 2312
rect 1152 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20452 2288
rect 1152 2224 20452 2248
rect 2667 2120 2709 2129
rect 2667 2080 2668 2120
rect 2708 2080 2709 2120
rect 2667 2071 2709 2080
rect 2859 2120 2901 2129
rect 2859 2080 2860 2120
rect 2900 2080 2901 2120
rect 2859 2071 2901 2080
rect 5067 2120 5109 2129
rect 5067 2080 5068 2120
rect 5108 2080 5109 2120
rect 5067 2071 5109 2080
rect 6699 2120 6741 2129
rect 6699 2080 6700 2120
rect 6740 2080 6741 2120
rect 6699 2071 6741 2080
rect 6979 2120 7037 2121
rect 6979 2080 6988 2120
rect 7028 2080 7037 2120
rect 6979 2079 7037 2080
rect 8619 2120 8661 2129
rect 8619 2080 8620 2120
rect 8660 2080 8661 2120
rect 8619 2071 8661 2080
rect 11307 2120 11349 2129
rect 11307 2080 11308 2120
rect 11348 2080 11349 2120
rect 11307 2071 11349 2080
rect 12939 2120 12981 2129
rect 12939 2080 12940 2120
rect 12980 2080 12981 2120
rect 12939 2071 12981 2080
rect 14571 2120 14613 2129
rect 14571 2080 14572 2120
rect 14612 2080 14613 2120
rect 14571 2071 14613 2080
rect 16203 2120 16245 2129
rect 16203 2080 16204 2120
rect 16244 2080 16245 2120
rect 16203 2071 16245 2080
rect 17931 2120 17973 2129
rect 17931 2080 17932 2120
rect 17972 2080 17973 2120
rect 17931 2071 17973 2080
rect 19851 2120 19893 2129
rect 19851 2080 19852 2120
rect 19892 2080 19893 2120
rect 19851 2071 19893 2080
rect 8811 2036 8853 2045
rect 8811 1996 8812 2036
rect 8852 1996 8853 2036
rect 8811 1987 8853 1996
rect 1219 1952 1277 1953
rect 1219 1912 1228 1952
rect 1268 1912 1277 1952
rect 1219 1911 1277 1912
rect 2467 1952 2525 1953
rect 2467 1912 2476 1952
rect 2516 1912 2525 1952
rect 2467 1911 2525 1912
rect 3339 1952 3381 1961
rect 3339 1912 3340 1952
rect 3380 1912 3381 1952
rect 3339 1903 3381 1912
rect 3435 1952 3477 1961
rect 3435 1912 3436 1952
rect 3476 1912 3477 1952
rect 3435 1903 3477 1912
rect 3915 1952 3957 1961
rect 3915 1912 3916 1952
rect 3956 1912 3957 1952
rect 3915 1903 3957 1912
rect 4387 1952 4445 1953
rect 4387 1912 4396 1952
rect 4436 1912 4445 1952
rect 5251 1952 5309 1953
rect 4387 1911 4445 1912
rect 4875 1938 4917 1947
rect 4875 1898 4876 1938
rect 4916 1898 4917 1938
rect 5251 1912 5260 1952
rect 5300 1912 5309 1952
rect 5251 1911 5309 1912
rect 6499 1952 6557 1953
rect 6499 1912 6508 1952
rect 6548 1912 6557 1952
rect 6499 1911 6557 1912
rect 7171 1952 7229 1953
rect 7171 1912 7180 1952
rect 7220 1912 7229 1952
rect 7171 1911 7229 1912
rect 8419 1952 8477 1953
rect 8419 1912 8428 1952
rect 8468 1912 8477 1952
rect 8419 1911 8477 1912
rect 9859 1952 9917 1953
rect 9859 1912 9868 1952
rect 9908 1912 9917 1952
rect 9859 1911 9917 1912
rect 11107 1952 11165 1953
rect 11107 1912 11116 1952
rect 11156 1912 11165 1952
rect 11107 1911 11165 1912
rect 11491 1952 11549 1953
rect 11491 1912 11500 1952
rect 11540 1912 11549 1952
rect 11491 1911 11549 1912
rect 12739 1952 12797 1953
rect 12739 1912 12748 1952
rect 12788 1912 12797 1952
rect 12739 1911 12797 1912
rect 13123 1952 13181 1953
rect 13123 1912 13132 1952
rect 13172 1912 13181 1952
rect 13123 1911 13181 1912
rect 14371 1952 14429 1953
rect 14371 1912 14380 1952
rect 14420 1912 14429 1952
rect 14371 1911 14429 1912
rect 14755 1952 14813 1953
rect 14755 1912 14764 1952
rect 14804 1912 14813 1952
rect 14755 1911 14813 1912
rect 16003 1952 16061 1953
rect 16003 1912 16012 1952
rect 16052 1912 16061 1952
rect 16003 1911 16061 1912
rect 16483 1952 16541 1953
rect 16483 1912 16492 1952
rect 16532 1912 16541 1952
rect 16483 1911 16541 1912
rect 17731 1952 17789 1953
rect 17731 1912 17740 1952
rect 17780 1912 17789 1952
rect 17731 1911 17789 1912
rect 18403 1952 18461 1953
rect 18403 1912 18412 1952
rect 18452 1912 18461 1952
rect 18403 1911 18461 1912
rect 19651 1952 19709 1953
rect 19651 1912 19660 1952
rect 19700 1912 19709 1952
rect 19651 1911 19709 1912
rect 4875 1889 4917 1898
rect 3043 1868 3101 1869
rect 3043 1828 3052 1868
rect 3092 1828 3101 1868
rect 3043 1827 3101 1828
rect 3819 1868 3861 1877
rect 3819 1828 3820 1868
rect 3860 1828 3861 1868
rect 3819 1819 3861 1828
rect 9091 1868 9149 1869
rect 9091 1828 9100 1868
rect 9140 1828 9149 1868
rect 9091 1827 9149 1828
rect 9475 1868 9533 1869
rect 9475 1828 9484 1868
rect 9524 1828 9533 1868
rect 9475 1827 9533 1828
rect 20227 1868 20285 1869
rect 20227 1828 20236 1868
rect 20276 1828 20285 1868
rect 20227 1827 20285 1828
rect 9291 1700 9333 1709
rect 9291 1660 9292 1700
rect 9332 1660 9333 1700
rect 9291 1651 9333 1660
rect 9675 1700 9717 1709
rect 9675 1660 9676 1700
rect 9716 1660 9717 1700
rect 9675 1651 9717 1660
rect 20043 1700 20085 1709
rect 20043 1660 20044 1700
rect 20084 1660 20085 1700
rect 20043 1651 20085 1660
rect 1152 1532 20352 1556
rect 1152 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 20352 1532
rect 1152 1468 20352 1492
rect 2763 1280 2805 1289
rect 2763 1240 2764 1280
rect 2804 1240 2805 1280
rect 2763 1231 2805 1240
rect 4971 1280 5013 1289
rect 4971 1240 4972 1280
rect 5012 1240 5013 1280
rect 4971 1231 5013 1240
rect 6699 1280 6741 1289
rect 6699 1240 6700 1280
rect 6740 1240 6741 1280
rect 6699 1231 6741 1240
rect 6987 1280 7029 1289
rect 6987 1240 6988 1280
rect 7028 1240 7029 1280
rect 6987 1231 7029 1240
rect 8619 1280 8661 1289
rect 8619 1240 8620 1280
rect 8660 1240 8661 1280
rect 8619 1231 8661 1240
rect 10251 1280 10293 1289
rect 10251 1240 10252 1280
rect 10292 1240 10293 1280
rect 10251 1231 10293 1240
rect 12075 1280 12117 1289
rect 12075 1240 12076 1280
rect 12116 1240 12117 1280
rect 12075 1231 12117 1240
rect 13707 1280 13749 1289
rect 13707 1240 13708 1280
rect 13748 1240 13749 1280
rect 13707 1231 13749 1240
rect 15339 1280 15381 1289
rect 15339 1240 15340 1280
rect 15380 1240 15381 1280
rect 15339 1231 15381 1240
rect 19851 1280 19893 1289
rect 19851 1240 19852 1280
rect 19892 1240 19893 1280
rect 19851 1231 19893 1240
rect 3139 1196 3197 1197
rect 3139 1156 3148 1196
rect 3188 1156 3197 1196
rect 3139 1155 3197 1156
rect 17155 1196 17213 1197
rect 17155 1156 17164 1196
rect 17204 1156 17213 1196
rect 17155 1155 17213 1156
rect 17539 1196 17597 1197
rect 17539 1156 17548 1196
rect 17588 1156 17597 1196
rect 17539 1155 17597 1156
rect 18211 1196 18269 1197
rect 18211 1156 18220 1196
rect 18260 1156 18269 1196
rect 18211 1155 18269 1156
rect 1315 1112 1373 1113
rect 1315 1072 1324 1112
rect 1364 1072 1373 1112
rect 1315 1071 1373 1072
rect 2563 1112 2621 1113
rect 2563 1072 2572 1112
rect 2612 1072 2621 1112
rect 2563 1071 2621 1072
rect 3523 1112 3581 1113
rect 3523 1072 3532 1112
rect 3572 1072 3581 1112
rect 3523 1071 3581 1072
rect 4771 1112 4829 1113
rect 4771 1072 4780 1112
rect 4820 1072 4829 1112
rect 4771 1071 4829 1072
rect 5251 1112 5309 1113
rect 5251 1072 5260 1112
rect 5300 1072 5309 1112
rect 5251 1071 5309 1072
rect 6499 1112 6557 1113
rect 6499 1072 6508 1112
rect 6548 1072 6557 1112
rect 6499 1071 6557 1072
rect 7171 1112 7229 1113
rect 7171 1072 7180 1112
rect 7220 1072 7229 1112
rect 7171 1071 7229 1072
rect 8419 1112 8477 1113
rect 8419 1072 8428 1112
rect 8468 1072 8477 1112
rect 8419 1071 8477 1072
rect 8803 1112 8861 1113
rect 8803 1072 8812 1112
rect 8852 1072 8861 1112
rect 8803 1071 8861 1072
rect 10051 1112 10109 1113
rect 10051 1072 10060 1112
rect 10100 1072 10109 1112
rect 10051 1071 10109 1072
rect 10627 1112 10685 1113
rect 10627 1072 10636 1112
rect 10676 1072 10685 1112
rect 10627 1071 10685 1072
rect 11875 1112 11933 1113
rect 11875 1072 11884 1112
rect 11924 1072 11933 1112
rect 11875 1071 11933 1072
rect 12259 1112 12317 1113
rect 12259 1072 12268 1112
rect 12308 1072 12317 1112
rect 12259 1071 12317 1072
rect 13507 1112 13565 1113
rect 13507 1072 13516 1112
rect 13556 1072 13565 1112
rect 13507 1071 13565 1072
rect 13891 1112 13949 1113
rect 13891 1072 13900 1112
rect 13940 1072 13949 1112
rect 13891 1071 13949 1072
rect 15139 1112 15197 1113
rect 15139 1072 15148 1112
rect 15188 1072 15197 1112
rect 15139 1071 15197 1072
rect 15523 1112 15581 1113
rect 15523 1072 15532 1112
rect 15572 1072 15581 1112
rect 15523 1071 15581 1072
rect 16771 1112 16829 1113
rect 16771 1072 16780 1112
rect 16820 1072 16829 1112
rect 16771 1071 16829 1072
rect 18403 1112 18461 1113
rect 18403 1072 18412 1112
rect 18452 1072 18461 1112
rect 18403 1071 18461 1072
rect 19651 1112 19709 1113
rect 19651 1072 19660 1112
rect 19700 1072 19709 1112
rect 19651 1071 19709 1072
rect 2955 944 2997 953
rect 2955 904 2956 944
rect 2996 904 2997 944
rect 2955 895 2997 904
rect 10443 944 10485 953
rect 10443 904 10444 944
rect 10484 904 10485 944
rect 10443 895 10485 904
rect 16971 944 17013 953
rect 16971 904 16972 944
rect 17012 904 17013 944
rect 16971 895 17013 904
rect 17355 944 17397 953
rect 17355 904 17356 944
rect 17396 904 17397 944
rect 17355 895 17397 904
rect 18027 944 18069 953
rect 18027 904 18028 944
rect 18068 904 18069 944
rect 18027 895 18069 904
rect 1152 776 20452 800
rect 1152 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20452 776
rect 1152 712 20452 736
<< via1 >>
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 5164 84484 5204 84524
rect 13132 84484 13172 84524
rect 18892 84484 18932 84524
rect 1516 84400 1556 84440
rect 1900 84400 1940 84440
rect 7276 84400 7316 84440
rect 7852 84400 7892 84440
rect 8044 84400 8084 84440
rect 19276 84400 19316 84440
rect 20044 84400 20084 84440
rect 1324 84316 1364 84356
rect 1708 84316 1748 84356
rect 7084 84316 7124 84356
rect 7660 84316 7700 84356
rect 8236 84316 8276 84356
rect 11788 84316 11828 84356
rect 12268 84316 12308 84356
rect 12940 84316 12980 84356
rect 13516 84316 13556 84356
rect 19084 84316 19124 84356
rect 19468 84316 19508 84356
rect 19852 84316 19892 84356
rect 20236 84316 20276 84356
rect 2092 84232 2132 84272
rect 3340 84232 3380 84272
rect 3724 84232 3764 84272
rect 4972 84232 5012 84272
rect 5548 84232 5588 84272
rect 6796 84232 6836 84272
rect 8428 84232 8468 84272
rect 9676 84232 9716 84272
rect 10252 84232 10292 84272
rect 11500 84232 11540 84272
rect 11692 84232 11732 84272
rect 11884 84232 11924 84272
rect 13708 84232 13748 84272
rect 14956 84232 14996 84272
rect 15340 84232 15380 84272
rect 16588 84232 16628 84272
rect 17260 84232 17300 84272
rect 18508 84232 18548 84272
rect 3532 84064 3572 84104
rect 5356 84064 5396 84104
rect 9868 84064 9908 84104
rect 10060 84064 10100 84104
rect 12460 84064 12500 84104
rect 12748 84064 12788 84104
rect 13324 84064 13364 84104
rect 15148 84064 15188 84104
rect 16780 84064 16820 84104
rect 17068 84064 17108 84104
rect 18700 84064 18740 84104
rect 19660 84064 19700 84104
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 1516 83728 1556 83768
rect 6700 83728 6740 83768
rect 7084 83728 7124 83768
rect 9004 83728 9044 83768
rect 18508 83728 18548 83768
rect 19564 83728 19604 83768
rect 19948 83728 19988 83768
rect 11788 83644 11828 83684
rect 1708 83560 1748 83600
rect 2956 83560 2996 83600
rect 3340 83560 3380 83600
rect 4588 83560 4628 83600
rect 4972 83560 5012 83600
rect 6220 83560 6260 83600
rect 7372 83560 7412 83600
rect 8620 83560 8660 83600
rect 10060 83560 10100 83600
rect 19084 83602 19124 83642
rect 10156 83560 10196 83600
rect 11116 83560 11156 83600
rect 11596 83546 11636 83586
rect 13996 83560 14036 83600
rect 15244 83560 15284 83600
rect 16492 83560 16532 83600
rect 17740 83560 17780 83600
rect 19276 83560 19316 83600
rect 19372 83560 19412 83600
rect 1324 83476 1364 83516
rect 9196 83476 9236 83516
rect 10540 83476 10580 83516
rect 10636 83476 10676 83516
rect 12172 83476 12212 83516
rect 12748 83476 12788 83516
rect 13420 83476 13460 83516
rect 13804 83476 13844 83516
rect 15820 83476 15860 83516
rect 16204 83476 16244 83516
rect 18316 83476 18356 83516
rect 18700 83476 18740 83516
rect 19756 83476 19796 83516
rect 20121 83473 20161 83513
rect 6604 83392 6644 83432
rect 7180 83392 7220 83432
rect 9484 83392 9524 83432
rect 9676 83392 9716 83432
rect 12556 83392 12596 83432
rect 12940 83392 12980 83432
rect 19084 83392 19124 83432
rect 3148 83308 3188 83348
rect 4780 83308 4820 83348
rect 6412 83308 6452 83348
rect 8812 83308 8852 83348
rect 12364 83308 12404 83348
rect 13228 83308 13268 83348
rect 13612 83308 13652 83348
rect 15436 83308 15476 83348
rect 15628 83308 15668 83348
rect 16012 83308 16052 83348
rect 17932 83308 17972 83348
rect 18124 83308 18164 83348
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 5644 82972 5684 83012
rect 6028 82972 6068 83012
rect 6412 82972 6452 83012
rect 11788 82972 11828 83012
rect 19084 82972 19124 83012
rect 20044 82972 20084 83012
rect 5164 82888 5204 82928
rect 3052 82804 3092 82844
rect 5452 82804 5492 82844
rect 5836 82804 5876 82844
rect 6220 82804 6260 82844
rect 7180 82804 7220 82844
rect 13612 82804 13652 82844
rect 14476 82804 14516 82844
rect 1324 82720 1364 82760
rect 2572 82720 2612 82760
rect 4684 82720 4724 82760
rect 6700 82720 6740 82760
rect 3436 82678 3476 82718
rect 6796 82720 6836 82760
rect 8284 82762 8324 82802
rect 20236 82804 20276 82844
rect 7276 82720 7316 82760
rect 7756 82720 7796 82760
rect 8716 82720 8756 82760
rect 9964 82720 10004 82760
rect 10348 82720 10388 82760
rect 11596 82720 11636 82760
rect 12460 82720 12500 82760
rect 12556 82720 12596 82760
rect 12652 82720 12692 82760
rect 13900 82720 13940 82760
rect 13996 82720 14036 82760
rect 14380 82720 14420 82760
rect 14956 82720 14996 82760
rect 15436 82734 15476 82774
rect 15820 82720 15860 82760
rect 17068 82720 17108 82760
rect 17452 82720 17492 82760
rect 18700 82720 18740 82760
rect 19468 82720 19508 82760
rect 19756 82720 19796 82760
rect 10156 82636 10196 82676
rect 18892 82636 18932 82676
rect 19372 82636 19412 82676
rect 2764 82552 2804 82592
rect 3244 82552 3284 82592
rect 4876 82552 4916 82592
rect 8428 82552 8468 82592
rect 12172 82552 12212 82592
rect 12748 82552 12788 82592
rect 12940 82552 12980 82592
rect 13420 82552 13460 82592
rect 15628 82552 15668 82592
rect 17260 82552 17300 82592
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 3052 82216 3092 82256
rect 3628 82216 3668 82256
rect 4012 82216 4052 82256
rect 4396 82216 4436 82256
rect 6604 82216 6644 82256
rect 6892 82216 6932 82256
rect 7180 82216 7220 82256
rect 10636 82216 10676 82256
rect 11020 82216 11060 82256
rect 12364 82216 12404 82256
rect 6412 82132 6452 82172
rect 14092 82132 14132 82172
rect 16204 82132 16244 82172
rect 1228 82048 1268 82088
rect 2476 82048 2516 82088
rect 4684 82048 4724 82088
rect 4780 82048 4820 82088
rect 5164 82048 5204 82088
rect 5740 82048 5780 82088
rect 6220 82043 6260 82083
rect 7564 82048 7604 82088
rect 8812 82048 8852 82088
rect 9196 82048 9236 82088
rect 10444 82048 10484 82088
rect 10828 82048 10868 82088
rect 11116 82048 11156 82088
rect 11404 82048 11444 82088
rect 11692 82048 11732 82088
rect 11788 82048 11828 82088
rect 12268 82048 12308 82088
rect 12460 82048 12500 82088
rect 12652 82048 12692 82088
rect 13900 82048 13940 82088
rect 14476 82048 14516 82088
rect 14572 82048 14612 82088
rect 15532 82048 15572 82088
rect 16012 82043 16052 82083
rect 16780 82048 16820 82088
rect 18028 82048 18068 82088
rect 18604 82048 18644 82088
rect 19852 82048 19892 82088
rect 2860 81964 2900 82004
rect 3436 81964 3476 82004
rect 3820 81964 3860 82004
rect 4204 81964 4244 82004
rect 5260 81964 5300 82004
rect 7372 81964 7412 82004
rect 14956 81964 14996 82004
rect 15052 81964 15092 82004
rect 16492 81880 16532 81920
rect 2668 81796 2708 81836
rect 9004 81796 9044 81836
rect 12076 81796 12116 81836
rect 18220 81796 18260 81836
rect 20044 81796 20084 81836
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 5356 81460 5396 81500
rect 11692 81460 11732 81500
rect 13612 81460 13652 81500
rect 15724 81460 15764 81500
rect 16588 81460 16628 81500
rect 3052 81376 3092 81416
rect 18604 81376 18644 81416
rect 4012 81292 4052 81332
rect 5548 81292 5588 81332
rect 15916 81292 15956 81332
rect 16396 81292 16436 81332
rect 1228 81208 1268 81248
rect 2476 81208 2516 81248
rect 3436 81208 3476 81248
rect 3532 81208 3572 81248
rect 3916 81208 3956 81248
rect 4492 81208 4532 81248
rect 4972 81222 5012 81262
rect 5740 81208 5780 81248
rect 6988 81208 7028 81248
rect 8908 81250 8948 81290
rect 7372 81208 7412 81248
rect 7660 81208 7700 81248
rect 9484 81208 9524 81248
rect 10732 81208 10772 81248
rect 11212 81208 11252 81248
rect 11308 81208 11348 81248
rect 11404 81208 11444 81248
rect 11500 81208 11540 81248
rect 11692 81208 11732 81248
rect 11884 81208 11924 81248
rect 11980 81208 12020 81248
rect 12172 81208 12212 81248
rect 13420 81208 13460 81248
rect 13804 81208 13844 81248
rect 15052 81208 15092 81248
rect 16780 81208 16820 81248
rect 18028 81208 18068 81248
rect 18796 81208 18836 81248
rect 20044 81208 20084 81248
rect 5164 81124 5204 81164
rect 2668 81040 2708 81080
rect 3148 81040 3188 81080
rect 7180 81040 7220 81080
rect 9100 81040 9140 81080
rect 9292 81040 9332 81080
rect 15244 81040 15284 81080
rect 15436 81040 15476 81080
rect 16108 81040 16148 81080
rect 18220 81040 18260 81080
rect 18508 81040 18548 81080
rect 20236 81040 20276 81080
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 3340 80704 3380 80744
rect 3724 80704 3764 80744
rect 11884 80704 11924 80744
rect 3052 80620 3092 80660
rect 9196 80620 9236 80660
rect 11500 80620 11540 80660
rect 13516 80620 13556 80660
rect 15532 80620 15572 80660
rect 1324 80536 1364 80576
rect 1420 80536 1460 80576
rect 2380 80536 2420 80576
rect 2860 80531 2900 80571
rect 4396 80536 4436 80576
rect 4972 80536 5012 80576
rect 1804 80452 1844 80492
rect 1900 80452 1940 80492
rect 3868 80494 3908 80534
rect 5356 80536 5396 80576
rect 5452 80536 5492 80576
rect 6028 80536 6068 80576
rect 6220 80536 6260 80576
rect 6604 80536 6644 80576
rect 6892 80536 6932 80576
rect 7468 80536 7508 80576
rect 7564 80536 7604 80576
rect 8524 80536 8564 80576
rect 9004 80531 9044 80571
rect 9772 80536 9812 80576
rect 9868 80536 9908 80576
rect 10828 80536 10868 80576
rect 11356 80526 11396 80566
rect 11788 80536 11828 80576
rect 12076 80536 12116 80576
rect 13324 80536 13364 80576
rect 13804 80536 13844 80576
rect 13900 80536 13940 80576
rect 14380 80536 14420 80576
rect 14860 80536 14900 80576
rect 15340 80531 15380 80571
rect 15820 80536 15860 80576
rect 16012 80536 16052 80576
rect 16204 80536 16244 80576
rect 16492 80536 16532 80576
rect 16876 80536 16916 80576
rect 18124 80536 18164 80576
rect 18892 80536 18932 80576
rect 4876 80452 4916 80492
rect 5740 80452 5780 80492
rect 6796 80452 6836 80492
rect 7084 80452 7124 80492
rect 7948 80452 7988 80492
rect 8044 80452 8084 80492
rect 10252 80452 10292 80492
rect 10348 80452 10388 80492
rect 20140 80494 20180 80534
rect 14284 80452 14324 80492
rect 6028 80368 6068 80408
rect 18508 80368 18548 80408
rect 15820 80284 15860 80324
rect 16204 80284 16244 80324
rect 16684 80284 16724 80324
rect 18700 80284 18740 80324
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 3532 79948 3572 79988
rect 15532 79948 15572 79988
rect 7468 79780 7508 79820
rect 16300 79780 16340 79820
rect 16396 79780 16436 79820
rect 1415 79696 1455 79736
rect 1516 79696 1556 79736
rect 1612 79696 1652 79736
rect 1804 79696 1844 79736
rect 1900 79696 1940 79736
rect 2092 79696 2132 79736
rect 3340 79696 3380 79736
rect 4012 79696 4052 79736
rect 5260 79696 5300 79736
rect 5740 79696 5780 79736
rect 6988 79696 7028 79736
rect 7852 79696 7892 79736
rect 9100 79696 9140 79736
rect 9484 79696 9524 79736
rect 10732 79696 10772 79736
rect 11116 79696 11156 79736
rect 12364 79717 12404 79757
rect 13708 79696 13748 79736
rect 14956 79696 14996 79736
rect 15340 79696 15380 79736
rect 15532 79696 15572 79736
rect 15820 79696 15860 79736
rect 15916 79696 15956 79736
rect 16876 79696 16916 79736
rect 17356 79710 17396 79750
rect 17932 79710 17972 79750
rect 18412 79696 18452 79736
rect 18892 79696 18932 79736
rect 18988 79696 19028 79736
rect 19372 79696 19412 79736
rect 19468 79715 19508 79755
rect 19756 79696 19796 79736
rect 19852 79696 19892 79736
rect 19948 79696 19988 79736
rect 15148 79612 15188 79652
rect 17740 79612 17780 79652
rect 1420 79528 1460 79568
rect 3820 79528 3860 79568
rect 5452 79528 5492 79568
rect 7180 79528 7220 79568
rect 9292 79528 9332 79568
rect 10924 79528 10964 79568
rect 12556 79528 12596 79568
rect 17548 79528 17588 79568
rect 20044 79528 20084 79568
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 3052 79192 3092 79232
rect 7468 79192 7508 79232
rect 17548 79192 17588 79232
rect 18124 79192 18164 79232
rect 10252 79108 10292 79148
rect 12364 79108 12404 79148
rect 20140 79108 20180 79148
rect 1228 79024 1268 79064
rect 2476 79024 2516 79064
rect 3244 79024 3284 79064
rect 4492 79024 4532 79064
rect 4972 79024 5012 79064
rect 6220 79024 6260 79064
rect 6892 79024 6932 79064
rect 6988 79024 7028 79064
rect 7084 79024 7124 79064
rect 7180 79024 7220 79064
rect 7756 79024 7796 79064
rect 7948 79024 7988 79064
rect 8044 79024 8084 79064
rect 8236 79024 8276 79064
rect 8428 79024 8468 79064
rect 8812 79024 8852 79064
rect 10060 79024 10100 79064
rect 10636 79024 10676 79064
rect 10732 79024 10772 79064
rect 11212 79024 11252 79064
rect 11692 79024 11732 79064
rect 12220 79014 12260 79054
rect 12556 79024 12596 79064
rect 13804 79024 13844 79064
rect 14380 79024 14420 79064
rect 15628 79024 15668 79064
rect 15916 79024 15956 79064
rect 17164 79024 17204 79064
rect 17644 79024 17684 79064
rect 17836 79024 17876 79064
rect 17932 79024 17972 79064
rect 18028 79024 18068 79064
rect 18412 79005 18452 79045
rect 18508 79005 18548 79045
rect 19468 79024 19508 79064
rect 19948 79019 19988 79059
rect 2860 78940 2900 78980
rect 11116 78940 11156 78980
rect 18892 78940 18932 78980
rect 18988 78940 19028 78980
rect 7372 78856 7412 78896
rect 7756 78856 7796 78896
rect 8236 78856 8276 78896
rect 2668 78772 2708 78812
rect 4684 78772 4724 78812
rect 6412 78772 6452 78812
rect 13996 78772 14036 78812
rect 14188 78772 14228 78812
rect 17356 78772 17396 78812
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 5356 78436 5396 78476
rect 7084 78436 7124 78476
rect 8044 78436 8084 78476
rect 17644 78436 17684 78476
rect 18508 78436 18548 78476
rect 3532 78268 3572 78308
rect 11116 78268 11156 78308
rect 13804 78268 13844 78308
rect 15820 78268 15860 78308
rect 17452 78268 17492 78308
rect 17836 78268 17876 78308
rect 18028 78268 18068 78308
rect 18316 78268 18356 78308
rect 1228 78184 1268 78224
rect 2476 78184 2516 78224
rect 2956 78184 2996 78224
rect 3052 78184 3092 78224
rect 3436 78184 3476 78224
rect 4012 78184 4052 78224
rect 4492 78198 4532 78238
rect 4876 78184 4916 78224
rect 4972 78184 5012 78224
rect 5452 78184 5492 78224
rect 5644 78184 5684 78224
rect 6892 78184 6932 78224
rect 7372 78184 7412 78224
rect 7660 78184 7700 78224
rect 7756 78184 7796 78224
rect 8428 78184 8468 78224
rect 9676 78184 9716 78224
rect 10540 78184 10580 78224
rect 10636 78184 10676 78224
rect 11020 78184 11060 78224
rect 11596 78184 11636 78224
rect 12076 78189 12116 78229
rect 13324 78184 13364 78224
rect 13420 78184 13460 78224
rect 13900 78184 13940 78224
rect 14380 78184 14420 78224
rect 14860 78198 14900 78238
rect 15340 78184 15380 78224
rect 15436 78184 15476 78224
rect 15916 78184 15956 78224
rect 16396 78184 16436 78224
rect 16876 78198 16916 78238
rect 18700 78184 18740 78224
rect 19948 78184 19988 78224
rect 2668 78100 2708 78140
rect 4684 78100 4724 78140
rect 12268 78100 12308 78140
rect 15052 78100 15092 78140
rect 5164 78016 5204 78056
rect 7084 78016 7124 78056
rect 9868 78016 9908 78056
rect 17068 78016 17108 78056
rect 17260 78016 17300 78056
rect 20140 78016 20180 78056
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 4972 77680 5012 77720
rect 7852 77680 7892 77720
rect 8332 77680 8372 77720
rect 8620 77680 8660 77720
rect 10444 77596 10484 77636
rect 12460 77638 12500 77678
rect 14860 77680 14900 77720
rect 17356 77680 17396 77720
rect 17548 77680 17588 77720
rect 17932 77680 17972 77720
rect 1228 77512 1268 77552
rect 2476 77512 2516 77552
rect 2956 77512 2996 77552
rect 4204 77512 4244 77552
rect 6124 77512 6164 77552
rect 6220 77512 6260 77552
rect 7180 77512 7220 77552
rect 7660 77507 7700 77547
rect 8044 77512 8084 77552
rect 8140 77512 8180 77552
rect 8236 77512 8276 77552
rect 8524 77512 8564 77552
rect 9004 77512 9044 77552
rect 10252 77512 10292 77552
rect 10732 77512 10772 77552
rect 10828 77512 10868 77552
rect 11308 77512 11348 77552
rect 11788 77512 11828 77552
rect 13420 77512 13460 77552
rect 14668 77512 14708 77552
rect 15532 77512 15572 77552
rect 16780 77512 16820 77552
rect 18604 77512 18644 77552
rect 19852 77512 19892 77552
rect 4780 77428 4820 77468
rect 5164 77428 5204 77468
rect 6604 77428 6644 77468
rect 6700 77428 6740 77468
rect 11212 77428 11252 77468
rect 12316 77470 12356 77510
rect 15244 77428 15284 77468
rect 17164 77428 17204 77468
rect 17740 77428 17780 77468
rect 18124 77428 18164 77468
rect 18316 77344 18356 77384
rect 2668 77260 2708 77300
rect 4396 77260 4436 77300
rect 4588 77260 4628 77300
rect 15052 77260 15092 77300
rect 16972 77260 17012 77300
rect 20044 77260 20084 77300
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 2092 76840 2132 76880
rect 4588 76840 4628 76880
rect 12556 76840 12596 76880
rect 17932 76840 17972 76880
rect 1324 76756 1364 76796
rect 1708 76756 1748 76796
rect 3148 76756 3188 76796
rect 4780 76756 4820 76796
rect 8908 76756 8948 76796
rect 2092 76672 2132 76712
rect 2188 76672 2228 76712
rect 2380 76672 2420 76712
rect 2668 76672 2708 76712
rect 2764 76672 2804 76712
rect 3244 76672 3284 76712
rect 3724 76672 3764 76712
rect 4204 76686 4244 76726
rect 6700 76714 6740 76754
rect 18124 76756 18164 76796
rect 18892 76756 18932 76796
rect 18988 76756 19028 76796
rect 5068 76672 5108 76712
rect 6316 76672 6356 76712
rect 7948 76672 7988 76712
rect 8428 76672 8468 76712
rect 8524 76672 8564 76712
rect 9004 76672 9044 76712
rect 9484 76672 9524 76712
rect 9964 76686 10004 76726
rect 11116 76672 11156 76712
rect 12364 76672 12404 76712
rect 14572 76672 14612 76712
rect 15820 76672 15860 76712
rect 16204 76672 16244 76712
rect 17452 76672 17492 76712
rect 18412 76672 18452 76712
rect 18508 76672 18548 76712
rect 19468 76672 19508 76712
rect 19948 76686 19988 76726
rect 4396 76588 4436 76628
rect 8140 76588 8180 76628
rect 1516 76504 1556 76544
rect 1900 76504 1940 76544
rect 6508 76504 6548 76544
rect 10156 76504 10196 76544
rect 16012 76504 16052 76544
rect 17644 76504 17684 76544
rect 20140 76504 20180 76544
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 1420 76168 1460 76208
rect 6700 76168 6740 76208
rect 7372 76168 7412 76208
rect 19660 76168 19700 76208
rect 20044 76168 20084 76208
rect 6412 76084 6452 76124
rect 15436 76084 15476 76124
rect 1612 76000 1652 76040
rect 2860 76000 2900 76040
rect 3436 76000 3476 76040
rect 4684 76000 4724 76040
rect 4972 76000 5012 76040
rect 6220 76000 6260 76040
rect 6638 75985 6678 76025
rect 6796 76000 6836 76040
rect 6892 76000 6932 76040
rect 7084 76000 7124 76040
rect 7180 76000 7220 76040
rect 7564 76000 7604 76040
rect 7660 76000 7700 76040
rect 7852 76000 7892 76040
rect 7948 76000 7988 76040
rect 8044 76000 8084 76040
rect 8140 76000 8180 76040
rect 10156 76000 10196 76040
rect 11404 76000 11444 76040
rect 12172 76000 12212 76040
rect 13420 76000 13460 76040
rect 13996 76000 14036 76040
rect 15244 76000 15284 76040
rect 15628 76000 15668 76040
rect 15724 76000 15764 76040
rect 15916 76000 15956 76040
rect 16204 76000 16244 76040
rect 17452 76000 17492 76040
rect 18028 76000 18068 76040
rect 19276 76000 19316 76040
rect 1228 75916 1268 75956
rect 20236 75916 20276 75956
rect 15724 75832 15764 75872
rect 3052 75748 3092 75788
rect 3244 75748 3284 75788
rect 11596 75748 11636 75788
rect 13612 75748 13652 75788
rect 17644 75748 17684 75788
rect 17836 75748 17876 75788
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 1612 75412 1652 75452
rect 2188 75412 2228 75452
rect 6316 75412 6356 75452
rect 7948 75412 7988 75452
rect 20140 75328 20180 75368
rect 1420 75244 1460 75284
rect 2380 75244 2420 75284
rect 2668 75160 2708 75200
rect 2764 75160 2804 75200
rect 3148 75160 3188 75200
rect 4252 75202 4292 75242
rect 11980 75244 12020 75284
rect 12076 75244 12116 75284
rect 17164 75244 17204 75284
rect 3244 75160 3284 75200
rect 3724 75160 3764 75200
rect 4588 75160 4628 75200
rect 5836 75160 5876 75200
rect 6220 75160 6260 75200
rect 6508 75160 6548 75200
rect 7756 75160 7796 75200
rect 8140 75160 8180 75200
rect 9388 75160 9428 75200
rect 9772 75160 9812 75200
rect 11020 75160 11060 75200
rect 11500 75160 11540 75200
rect 11596 75160 11636 75200
rect 12556 75160 12596 75200
rect 13036 75174 13076 75214
rect 13516 75160 13556 75200
rect 14764 75160 14804 75200
rect 15244 75160 15284 75200
rect 15340 75160 15380 75200
rect 15724 75160 15764 75200
rect 15820 75160 15860 75200
rect 16012 75160 16052 75200
rect 16108 75160 16148 75200
rect 16209 75160 16249 75200
rect 16684 75160 16724 75200
rect 16780 75160 16820 75200
rect 17260 75160 17300 75200
rect 17740 75160 17780 75200
rect 18220 75174 18260 75214
rect 4396 75076 4436 75116
rect 6028 74992 6068 75032
rect 9580 74992 9620 75032
rect 11212 74992 11252 75032
rect 13228 74992 13268 75032
rect 14956 74992 14996 75032
rect 15532 74992 15572 75032
rect 15916 74992 15956 75032
rect 18412 74992 18452 75032
rect 20044 74992 20084 75032
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 9964 74656 10004 74696
rect 11980 74656 12020 74696
rect 12460 74656 12500 74696
rect 7756 74572 7796 74612
rect 15148 74572 15188 74612
rect 15628 74572 15668 74612
rect 20236 74572 20276 74612
rect 1900 74488 1940 74528
rect 3148 74488 3188 74528
rect 4204 74488 4244 74528
rect 5452 74488 5492 74528
rect 6028 74488 6068 74528
rect 6124 74488 6164 74528
rect 6508 74488 6548 74528
rect 6604 74488 6644 74528
rect 7084 74488 7124 74528
rect 7612 74478 7652 74518
rect 9676 74488 9716 74528
rect 9772 74488 9812 74528
rect 10252 74488 10292 74528
rect 10348 74488 10388 74528
rect 10828 74488 10868 74528
rect 11308 74488 11348 74528
rect 11788 74483 11828 74523
rect 12844 74488 12884 74528
rect 12940 74488 12980 74528
rect 13036 74488 13076 74528
rect 13132 74488 13172 74528
rect 13420 74488 13460 74528
rect 13516 74488 13556 74528
rect 13900 74488 13940 74528
rect 13996 74488 14036 74528
rect 14476 74488 14516 74528
rect 14956 74483 14996 74523
rect 16492 74488 16532 74528
rect 16780 74488 16820 74528
rect 18028 74488 18068 74528
rect 18508 74488 18548 74528
rect 18604 74488 18644 74528
rect 18988 74488 19028 74528
rect 19564 74488 19604 74528
rect 20044 74483 20084 74523
rect 10732 74404 10772 74444
rect 12652 74404 12692 74444
rect 19084 74404 19124 74444
rect 3340 74236 3380 74276
rect 4012 74236 4052 74276
rect 18220 74236 18260 74276
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 10060 73900 10100 73940
rect 13900 73900 13940 73940
rect 16108 73900 16148 73940
rect 7084 73816 7124 73856
rect 2092 73732 2132 73772
rect 2188 73732 2228 73772
rect 1612 73648 1652 73688
rect 1708 73648 1748 73688
rect 2668 73648 2708 73688
rect 3148 73662 3188 73702
rect 3532 73648 3572 73688
rect 4780 73648 4820 73688
rect 5356 73648 5396 73688
rect 6604 73648 6644 73688
rect 6796 73648 6836 73688
rect 6988 73648 7028 73688
rect 7084 73648 7124 73688
rect 7276 73648 7316 73688
rect 7372 73648 7412 73688
rect 7564 73648 7604 73688
rect 7660 73648 7700 73688
rect 7815 73648 7855 73688
rect 8044 73648 8084 73688
rect 8140 73648 8180 73688
rect 8428 73648 8468 73688
rect 9676 73648 9716 73688
rect 10060 73648 10100 73688
rect 10156 73663 10196 73703
rect 10348 73648 10388 73688
rect 10444 73677 10484 73717
rect 10545 73648 10585 73688
rect 10828 73648 10868 73688
rect 12076 73648 12116 73688
rect 12460 73648 12500 73688
rect 13708 73648 13748 73688
rect 14284 73648 14324 73688
rect 15532 73648 15572 73688
rect 16012 73648 16052 73688
rect 16876 73648 16916 73688
rect 18124 73648 18164 73688
rect 18508 73648 18548 73688
rect 19756 73648 19796 73688
rect 9868 73564 9908 73604
rect 3340 73438 3380 73478
rect 4972 73480 5012 73520
rect 5164 73480 5204 73520
rect 7660 73480 7700 73520
rect 12268 73480 12308 73520
rect 15724 73480 15764 73520
rect 18316 73480 18356 73520
rect 19948 73480 19988 73520
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 7468 73144 7508 73184
rect 7948 73144 7988 73184
rect 10060 73144 10100 73184
rect 10444 73144 10484 73184
rect 3628 73060 3668 73100
rect 9772 73060 9812 73100
rect 13324 73060 13364 73100
rect 17452 73060 17492 73100
rect 1228 72976 1268 73016
rect 2476 72976 2516 73016
rect 3820 72971 3860 73011
rect 4300 72976 4340 73016
rect 5260 72976 5300 73016
rect 5356 72976 5396 73016
rect 6028 72976 6068 73016
rect 7276 72976 7316 73016
rect 7660 72976 7700 73016
rect 7756 72976 7796 73016
rect 8332 72976 8372 73016
rect 9580 72976 9620 73016
rect 9964 72976 10004 73016
rect 10156 72976 10196 73016
rect 10252 72976 10292 73016
rect 10540 72976 10580 73016
rect 11692 72976 11732 73016
rect 12940 72976 12980 73016
rect 13420 72976 13460 73016
rect 13516 72976 13556 73016
rect 13612 72976 13652 73016
rect 13996 72976 14036 73016
rect 15244 72976 15284 73016
rect 15724 72957 15764 72997
rect 15820 72976 15860 73016
rect 16780 72976 16820 73016
rect 17260 72971 17300 73011
rect 18412 72976 18452 73016
rect 19660 72976 19700 73016
rect 4780 72892 4820 72932
rect 4876 72892 4916 72932
rect 16204 72892 16244 72932
rect 16300 72892 16340 72932
rect 15436 72808 15476 72848
rect 2668 72724 2708 72764
rect 13132 72724 13172 72764
rect 19852 72724 19892 72764
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 7372 72388 7412 72428
rect 13324 72388 13364 72428
rect 13612 72220 13652 72260
rect 16300 72220 16340 72260
rect 19084 72220 19124 72260
rect 1708 72136 1748 72176
rect 2956 72136 2996 72176
rect 4300 72136 4340 72176
rect 5548 72136 5588 72176
rect 5932 72136 5972 72176
rect 7180 72136 7220 72176
rect 7756 72136 7796 72176
rect 9004 72136 9044 72176
rect 9388 72136 9428 72176
rect 10636 72136 10676 72176
rect 11212 72136 11252 72176
rect 11308 72136 11348 72176
rect 11692 72136 11732 72176
rect 11884 72136 11924 72176
rect 13132 72136 13172 72176
rect 13516 72136 13556 72176
rect 13804 72136 13844 72176
rect 13996 72136 14036 72176
rect 15244 72136 15284 72176
rect 15724 72136 15764 72176
rect 15820 72136 15860 72176
rect 16204 72136 16244 72176
rect 16780 72136 16820 72176
rect 17260 72150 17300 72190
rect 18508 72136 18548 72176
rect 18604 72136 18644 72176
rect 18988 72136 19028 72176
rect 19564 72136 19604 72176
rect 20044 72150 20084 72190
rect 3148 71968 3188 72008
rect 5740 71968 5780 72008
rect 9196 71968 9236 72008
rect 10828 71968 10868 72008
rect 11020 71968 11060 72008
rect 11596 71968 11636 72008
rect 13324 71968 13364 72008
rect 15436 71968 15476 72008
rect 17452 71968 17492 72008
rect 20236 71968 20276 72008
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 3244 71632 3284 71672
rect 7660 71632 7700 71672
rect 6028 71548 6068 71588
rect 9676 71548 9716 71588
rect 13996 71548 14036 71588
rect 1516 71464 1556 71504
rect 1612 71464 1652 71504
rect 2092 71464 2132 71504
rect 2572 71464 2612 71504
rect 3052 71459 3092 71499
rect 4300 71464 4340 71504
rect 4396 71464 4436 71504
rect 5356 71464 5396 71504
rect 5836 71459 5876 71499
rect 6220 71464 6260 71504
rect 7468 71464 7508 71504
rect 7948 71464 7988 71504
rect 8044 71464 8084 71504
rect 8524 71464 8564 71504
rect 9004 71464 9044 71504
rect 9484 71459 9524 71499
rect 9868 71464 9908 71504
rect 11116 71464 11156 71504
rect 11500 71464 11540 71504
rect 11596 71464 11636 71504
rect 11788 71464 11828 71504
rect 12268 71464 12308 71504
rect 12364 71464 12404 71504
rect 1996 71380 2036 71420
rect 4780 71380 4820 71420
rect 4876 71380 4916 71420
rect 8428 71380 8468 71420
rect 12748 71422 12788 71462
rect 12844 71464 12884 71504
rect 13324 71464 13364 71504
rect 13804 71459 13844 71499
rect 14188 71464 14228 71504
rect 14380 71464 14420 71504
rect 14572 71464 14612 71504
rect 15820 71464 15860 71504
rect 16204 71464 16244 71504
rect 17452 71464 17492 71504
rect 18316 71464 18356 71504
rect 19564 71464 19604 71504
rect 11500 71296 11540 71336
rect 11308 71212 11348 71252
rect 14380 71212 14420 71252
rect 16012 71212 16052 71252
rect 17644 71212 17684 71252
rect 19756 71212 19796 71252
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 10924 70876 10964 70916
rect 12268 70876 12308 70916
rect 12460 70792 12500 70832
rect 4780 70666 4820 70706
rect 1228 70624 1268 70664
rect 2476 70624 2516 70664
rect 3148 70624 3188 70664
rect 4396 70624 4436 70664
rect 6028 70624 6068 70664
rect 6604 70624 6644 70664
rect 7852 70624 7892 70664
rect 8332 70624 8372 70664
rect 8428 70624 8468 70664
rect 8812 70624 8852 70664
rect 8908 70624 8948 70664
rect 9388 70624 9428 70664
rect 9916 70633 9956 70673
rect 10439 70624 10479 70664
rect 10540 70624 10580 70664
rect 10636 70624 10676 70664
rect 10828 70624 10868 70664
rect 10924 70624 10964 70664
rect 11212 70624 11252 70664
rect 11980 70624 12020 70664
rect 12076 70624 12116 70664
rect 12748 70666 12788 70706
rect 12268 70624 12308 70664
rect 12844 70624 12884 70664
rect 13132 70624 13172 70664
rect 13420 70624 13460 70664
rect 14668 70624 14708 70664
rect 15052 70624 15092 70664
rect 15244 70624 15284 70664
rect 16204 70624 16244 70664
rect 17452 70624 17492 70664
rect 18508 70624 18548 70664
rect 19756 70624 19796 70664
rect 8044 70540 8084 70580
rect 10060 70540 10100 70580
rect 11116 70540 11156 70580
rect 15148 70540 15188 70580
rect 17644 70540 17684 70580
rect 2668 70456 2708 70496
rect 4588 70456 4628 70496
rect 6220 70456 6260 70496
rect 14860 70456 14900 70496
rect 19948 70456 19988 70496
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 5164 70120 5204 70160
rect 10156 70120 10196 70160
rect 7948 70036 7988 70076
rect 12844 70036 12884 70076
rect 14668 70036 14708 70076
rect 16684 70036 16724 70076
rect 19948 70036 19988 70076
rect 1228 69952 1268 69992
rect 2476 69952 2516 69992
rect 3436 69952 3476 69992
rect 3532 69952 3572 69992
rect 3916 69952 3956 69992
rect 4492 69952 4532 69992
rect 4972 69947 5012 69987
rect 6220 69952 6260 69992
rect 6316 69952 6356 69992
rect 6700 69952 6740 69992
rect 6796 69952 6836 69992
rect 7276 69952 7316 69992
rect 7756 69938 7796 69978
rect 9964 69952 10004 69992
rect 11116 69952 11156 69992
rect 8716 69910 8756 69950
rect 11212 69952 11252 69992
rect 11692 69952 11732 69992
rect 12172 69952 12212 69992
rect 12652 69938 12692 69978
rect 13228 69952 13268 69992
rect 14476 69952 14516 69992
rect 14956 69952 14996 69992
rect 15052 69952 15092 69992
rect 16012 69952 16052 69992
rect 16492 69947 16532 69987
rect 18220 69952 18260 69992
rect 18316 69952 18356 69992
rect 18700 69952 18740 69992
rect 18796 69952 18836 69992
rect 19276 69952 19316 69992
rect 19804 69942 19844 69982
rect 4012 69868 4052 69908
rect 11596 69868 11636 69908
rect 15436 69868 15476 69908
rect 15532 69868 15572 69908
rect 2668 69700 2708 69740
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 7660 69364 7700 69404
rect 11020 69364 11060 69404
rect 12652 69364 12692 69404
rect 8524 69196 8564 69236
rect 15532 69196 15572 69236
rect 18892 69196 18932 69236
rect 1228 69112 1268 69152
rect 2476 69112 2516 69152
rect 2860 69112 2900 69152
rect 4108 69112 4148 69152
rect 4684 69112 4724 69152
rect 5932 69112 5972 69152
rect 6220 69112 6260 69152
rect 7468 69112 7508 69152
rect 8428 69112 8468 69152
rect 8620 69112 8660 69152
rect 8812 69112 8852 69152
rect 8908 69112 8948 69152
rect 9004 69112 9044 69152
rect 9580 69112 9620 69152
rect 10828 69112 10868 69152
rect 11212 69112 11252 69152
rect 12460 69112 12500 69152
rect 13228 69112 13268 69152
rect 14476 69112 14516 69152
rect 14956 69112 14996 69152
rect 15052 69112 15092 69152
rect 15436 69112 15476 69152
rect 16012 69112 16052 69152
rect 16492 69126 16532 69166
rect 18316 69112 18356 69152
rect 18412 69112 18452 69152
rect 18796 69112 18836 69152
rect 19372 69112 19412 69152
rect 19852 69126 19892 69166
rect 2668 68944 2708 68984
rect 4300 68944 4340 68984
rect 4492 68944 4532 68984
rect 9100 68944 9140 68984
rect 14668 68944 14708 68984
rect 16684 68944 16724 68984
rect 20044 68944 20084 68984
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 9580 68608 9620 68648
rect 3436 68524 3476 68564
rect 1708 68440 1748 68480
rect 1804 68440 1844 68480
rect 2284 68440 2324 68480
rect 2764 68440 2804 68480
rect 3244 68435 3284 68475
rect 4780 68440 4820 68480
rect 6028 68440 6068 68480
rect 6508 68440 6548 68480
rect 7756 68440 7796 68480
rect 8140 68440 8180 68480
rect 9388 68440 9428 68480
rect 9772 68440 9812 68480
rect 9964 68440 10004 68480
rect 10156 68440 10196 68480
rect 11404 68419 11444 68459
rect 12556 68440 12596 68480
rect 13804 68440 13844 68480
rect 14188 68440 14228 68480
rect 15436 68440 15476 68480
rect 15916 68440 15956 68480
rect 17164 68440 17204 68480
rect 18412 68440 18452 68480
rect 19660 68440 19700 68480
rect 2188 68356 2228 68396
rect 9868 68356 9908 68396
rect 6220 68188 6260 68228
rect 7948 68188 7988 68228
rect 11596 68188 11636 68228
rect 12364 68188 12404 68228
rect 13996 68188 14036 68228
rect 17356 68188 17396 68228
rect 19852 68188 19892 68228
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 10348 67852 10388 67892
rect 5164 67684 5204 67724
rect 8428 67684 8468 67724
rect 11980 67684 12020 67724
rect 18412 67684 18452 67724
rect 1804 67600 1844 67640
rect 3052 67600 3092 67640
rect 4684 67600 4724 67640
rect 4780 67600 4820 67640
rect 5260 67600 5300 67640
rect 5740 67600 5780 67640
rect 6220 67614 6260 67654
rect 7372 67600 7412 67640
rect 7468 67600 7508 67640
rect 7660 67600 7700 67640
rect 7948 67600 7988 67640
rect 8044 67600 8084 67640
rect 8524 67600 8564 67640
rect 9004 67600 9044 67640
rect 9484 67614 9524 67654
rect 9868 67600 9908 67640
rect 9964 67600 10004 67640
rect 10060 67600 10100 67640
rect 10156 67600 10196 67640
rect 10348 67600 10388 67640
rect 10540 67600 10580 67640
rect 10636 67600 10676 67640
rect 11500 67600 11540 67640
rect 11596 67600 11636 67640
rect 12076 67600 12116 67640
rect 12556 67600 12596 67640
rect 13036 67614 13076 67654
rect 13612 67600 13652 67640
rect 14860 67600 14900 67640
rect 15916 67600 15956 67640
rect 17164 67600 17204 67640
rect 17932 67600 17972 67640
rect 18028 67600 18068 67640
rect 18508 67600 18548 67640
rect 18988 67600 19028 67640
rect 19468 67614 19508 67654
rect 9676 67516 9716 67556
rect 3244 67432 3284 67472
rect 6412 67432 6452 67472
rect 13228 67432 13268 67472
rect 13420 67432 13460 67472
rect 17356 67432 17396 67472
rect 19660 67390 19700 67430
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 4204 67096 4244 67136
rect 8620 67096 8660 67136
rect 9292 67012 9332 67052
rect 11212 67012 11252 67052
rect 13228 67012 13268 67052
rect 16108 67012 16148 67052
rect 19660 67012 19700 67052
rect 2476 66928 2516 66968
rect 2572 66928 2612 66968
rect 3052 66928 3092 66968
rect 3532 66928 3572 66968
rect 4060 66918 4100 66958
rect 5164 66928 5204 66968
rect 6412 66928 6452 66968
rect 6879 66931 6919 66971
rect 7180 66928 7220 66968
rect 8428 66928 8468 66968
rect 8908 66928 8948 66968
rect 9196 66928 9236 66968
rect 9772 66928 9812 66968
rect 11020 66928 11060 66968
rect 11500 66928 11540 66968
rect 11596 66928 11636 66968
rect 11980 66928 12020 66968
rect 12556 66928 12596 66968
rect 13084 66918 13124 66958
rect 14380 66928 14420 66968
rect 14476 66928 14516 66968
rect 14860 66928 14900 66968
rect 14956 66928 14996 66968
rect 15436 66928 15476 66968
rect 15916 66923 15956 66963
rect 16684 66928 16724 66968
rect 17932 66928 17972 66968
rect 18028 66928 18068 66968
rect 18412 66928 18452 66968
rect 18508 66928 18548 66968
rect 18988 66928 19028 66968
rect 19468 66923 19508 66963
rect 2956 66844 2996 66884
rect 12076 66844 12116 66884
rect 9580 66760 9620 66800
rect 16972 66760 17012 66800
rect 6604 66676 6644 66716
rect 6988 66676 7028 66716
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 9004 66256 9044 66296
rect 1420 66088 1460 66128
rect 2668 66088 2708 66128
rect 3340 66088 3380 66128
rect 4588 66088 4628 66128
rect 5068 66088 5108 66128
rect 6316 66088 6356 66128
rect 6690 66097 6730 66137
rect 6796 66088 6836 66128
rect 6988 66088 7028 66128
rect 7084 66117 7124 66157
rect 7185 66088 7225 66128
rect 7468 66088 7508 66128
rect 7564 66088 7604 66128
rect 8716 66088 8756 66128
rect 8908 66088 8948 66128
rect 9004 66088 9044 66128
rect 9196 66088 9236 66128
rect 9292 66088 9332 66128
rect 11212 66088 11252 66128
rect 12460 66088 12500 66128
rect 12844 66088 12884 66128
rect 14092 66088 14132 66128
rect 14476 66088 14516 66128
rect 15724 66088 15764 66128
rect 16684 66088 16724 66128
rect 17932 66088 17972 66128
rect 18316 66088 18356 66128
rect 19564 66088 19604 66128
rect 2860 65920 2900 65960
rect 4780 65920 4820 65960
rect 6508 65920 6548 65960
rect 7084 65920 7124 65960
rect 7756 65920 7796 65960
rect 12652 65920 12692 65960
rect 14284 65920 14324 65960
rect 15916 65920 15956 65960
rect 18124 65920 18164 65960
rect 19756 65920 19796 65960
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 5740 65584 5780 65624
rect 9196 65584 9236 65624
rect 4588 65500 4628 65540
rect 10828 65500 10868 65540
rect 12844 65500 12884 65540
rect 16012 65500 16052 65540
rect 19180 65500 19220 65540
rect 2860 65416 2900 65456
rect 2956 65416 2996 65456
rect 3436 65416 3476 65456
rect 3916 65416 3956 65456
rect 4444 65406 4484 65446
rect 5644 65416 5684 65456
rect 5836 65416 5876 65456
rect 5932 65416 5972 65456
rect 6124 65416 6164 65456
rect 7372 65416 7412 65456
rect 7756 65416 7796 65456
rect 9388 65416 9428 65456
rect 10636 65416 10676 65456
rect 11116 65416 11156 65456
rect 9004 65374 9044 65414
rect 11212 65416 11252 65456
rect 11596 65416 11636 65456
rect 11692 65416 11732 65456
rect 12172 65416 12212 65456
rect 12652 65411 12692 65451
rect 14284 65416 14324 65456
rect 14380 65416 14420 65456
rect 14764 65416 14804 65456
rect 14860 65416 14900 65456
rect 15340 65416 15380 65456
rect 15868 65406 15908 65446
rect 17452 65416 17492 65456
rect 17548 65416 17588 65456
rect 18028 65416 18068 65456
rect 18508 65416 18548 65456
rect 18988 65411 19028 65451
rect 3340 65332 3380 65372
rect 16492 65332 16532 65372
rect 17932 65332 17972 65372
rect 16684 65248 16724 65288
rect 7564 65164 7604 65204
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 9292 64828 9332 64868
rect 2668 64660 2708 64700
rect 6220 64660 6260 64700
rect 18028 64660 18068 64700
rect 18124 64660 18164 64700
rect 19852 64660 19892 64700
rect 2092 64576 2132 64616
rect 2188 64576 2228 64616
rect 2572 64576 2612 64616
rect 3148 64576 3188 64616
rect 3628 64590 3668 64630
rect 4012 64576 4052 64616
rect 5260 64576 5300 64616
rect 5740 64576 5780 64616
rect 5836 64576 5876 64616
rect 6316 64576 6356 64616
rect 6796 64576 6836 64616
rect 7276 64581 7316 64621
rect 7852 64576 7892 64616
rect 9100 64576 9140 64616
rect 9484 64599 9524 64639
rect 9580 64576 9620 64616
rect 9772 64576 9812 64616
rect 9868 64576 9908 64616
rect 10023 64576 10063 64616
rect 10252 64576 10292 64616
rect 10348 64576 10388 64616
rect 10828 64576 10868 64616
rect 12076 64576 12116 64616
rect 12652 64576 12692 64616
rect 13900 64576 13940 64616
rect 14476 64576 14516 64616
rect 15724 64576 15764 64616
rect 17548 64576 17588 64616
rect 17644 64576 17684 64616
rect 18604 64576 18644 64616
rect 19132 64585 19172 64625
rect 3820 64492 3860 64532
rect 9484 64492 9524 64532
rect 5452 64408 5492 64448
rect 7468 64366 7508 64406
rect 10636 64408 10676 64448
rect 14092 64408 14132 64448
rect 15916 64408 15956 64448
rect 19276 64408 19316 64448
rect 20044 64408 20084 64448
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 8236 64072 8276 64112
rect 15724 63988 15764 64028
rect 1420 63904 1460 63944
rect 2668 63904 2708 63944
rect 3820 63904 3860 63944
rect 5068 63904 5108 63944
rect 6028 63904 6068 63944
rect 7276 63904 7316 63944
rect 8428 63904 8468 63944
rect 8524 63904 8564 63944
rect 8716 63904 8756 63944
rect 9964 63904 10004 63944
rect 10348 63904 10388 63944
rect 11596 63904 11636 63944
rect 12268 63904 12308 63944
rect 13516 63904 13556 63944
rect 13996 63904 14036 63944
rect 14092 63904 14132 63944
rect 14572 63904 14612 63944
rect 15052 63904 15092 63944
rect 15532 63899 15572 63939
rect 16300 63904 16340 63944
rect 17548 63904 17588 63944
rect 18124 63904 18164 63944
rect 19372 63904 19412 63944
rect 14476 63820 14516 63860
rect 19756 63820 19796 63860
rect 2860 63652 2900 63692
rect 5260 63652 5300 63692
rect 7468 63652 7508 63692
rect 10156 63652 10196 63692
rect 11788 63652 11828 63692
rect 13708 63652 13748 63692
rect 17740 63652 17780 63692
rect 17932 63652 17972 63692
rect 19948 63652 19988 63692
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 1516 63232 1556 63272
rect 1900 63232 1940 63272
rect 2284 63232 2324 63272
rect 1708 63148 1748 63188
rect 2092 63148 2132 63188
rect 2476 63148 2516 63188
rect 6508 63148 6548 63188
rect 5548 63106 5588 63146
rect 6604 63148 6644 63188
rect 10252 63148 10292 63188
rect 10348 63148 10388 63188
rect 12268 63148 12308 63188
rect 12364 63148 12404 63188
rect 18412 63148 18452 63188
rect 18508 63148 18548 63188
rect 19852 63148 19892 63188
rect 2860 63064 2900 63104
rect 4108 63064 4148 63104
rect 4300 63064 4340 63104
rect 6028 63064 6068 63104
rect 6124 63064 6164 63104
rect 7084 63064 7124 63104
rect 7564 63078 7604 63118
rect 8044 63064 8084 63104
rect 9292 63064 9332 63104
rect 9772 63064 9812 63104
rect 9868 63064 9908 63104
rect 10828 63064 10868 63104
rect 11308 63069 11348 63109
rect 11788 63083 11828 63123
rect 11884 63064 11924 63104
rect 12844 63064 12884 63104
rect 13324 63078 13364 63118
rect 14860 63064 14900 63104
rect 16108 63064 16148 63104
rect 17932 63064 17972 63104
rect 19516 63106 19556 63146
rect 18028 63064 18068 63104
rect 18988 63064 19028 63104
rect 2668 62980 2708 63020
rect 5740 62980 5780 63020
rect 7756 62896 7796 62936
rect 9484 62896 9524 62936
rect 11500 62896 11540 62936
rect 13516 62896 13556 62936
rect 16300 62896 16340 62936
rect 19660 62896 19700 62936
rect 20044 62896 20084 62936
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 5068 62560 5108 62600
rect 16108 62560 16148 62600
rect 16876 62560 16916 62600
rect 19660 62560 19700 62600
rect 9964 62476 10004 62516
rect 1324 62392 1364 62432
rect 2572 62392 2612 62432
rect 3340 62412 3380 62452
rect 3436 62392 3476 62432
rect 4396 62392 4436 62432
rect 4876 62387 4916 62427
rect 6508 62392 6548 62432
rect 7756 62392 7796 62432
rect 8236 62392 8276 62432
rect 8332 62392 8372 62432
rect 8716 62392 8756 62432
rect 8812 62392 8852 62432
rect 9292 62392 9332 62432
rect 9772 62387 9812 62427
rect 11116 62392 11156 62432
rect 12364 62392 12404 62432
rect 14380 62392 14420 62432
rect 14476 62392 14516 62432
rect 14860 62392 14900 62432
rect 15436 62392 15476 62432
rect 15964 62382 16004 62422
rect 17932 62392 17972 62432
rect 18028 62392 18068 62432
rect 18412 62392 18452 62432
rect 18508 62392 18548 62432
rect 18988 62392 19028 62432
rect 19468 62387 19508 62427
rect 3820 62308 3860 62348
rect 3916 62308 3956 62348
rect 13228 62308 13268 62348
rect 14956 62308 14996 62348
rect 16684 62308 16724 62348
rect 19852 62308 19892 62348
rect 2764 62140 2804 62180
rect 7948 62140 7988 62180
rect 12556 62140 12596 62180
rect 13036 62140 13076 62180
rect 20044 62140 20084 62180
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 14668 61804 14708 61844
rect 16108 61720 16148 61760
rect 4108 61636 4148 61676
rect 4204 61636 4244 61676
rect 14860 61636 14900 61676
rect 15916 61636 15956 61676
rect 19756 61636 19796 61676
rect 1324 61552 1364 61592
rect 2572 61552 2612 61592
rect 3148 61566 3188 61606
rect 3628 61552 3668 61592
rect 4588 61552 4628 61592
rect 4684 61552 4724 61592
rect 6508 61552 6548 61592
rect 7756 61552 7796 61592
rect 8908 61552 8948 61592
rect 10156 61552 10196 61592
rect 11020 61552 11060 61592
rect 12268 61552 12308 61592
rect 13228 61552 13268 61592
rect 14476 61552 14516 61592
rect 16300 61552 16340 61592
rect 17548 61552 17588 61592
rect 18124 61552 18164 61592
rect 19372 61552 19412 61592
rect 2956 61468 2996 61508
rect 2764 61384 2804 61424
rect 7948 61384 7988 61424
rect 10348 61384 10388 61424
rect 12460 61384 12500 61424
rect 15052 61384 15092 61424
rect 17740 61384 17780 61424
rect 19564 61384 19604 61424
rect 19948 61384 19988 61424
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 14956 61048 14996 61088
rect 15532 61048 15572 61088
rect 10252 60964 10292 61004
rect 12268 60964 12308 61004
rect 1900 60880 1940 60920
rect 3148 60880 3188 60920
rect 3532 60880 3572 60920
rect 4780 60880 4820 60920
rect 5164 60880 5204 60920
rect 6412 60880 6452 60920
rect 6892 60880 6932 60920
rect 8140 60880 8180 60920
rect 8812 60880 8852 60920
rect 10060 60880 10100 60920
rect 10540 60880 10580 60920
rect 10636 60880 10676 60920
rect 11116 60880 11156 60920
rect 11596 60880 11636 60920
rect 12076 60875 12116 60915
rect 12844 60880 12884 60920
rect 14092 60880 14132 60920
rect 14476 60880 14516 60920
rect 14572 60880 14612 60920
rect 14764 60880 14804 60920
rect 14860 60880 14900 60920
rect 15017 60865 15057 60905
rect 15244 60880 15284 60920
rect 16300 60922 16340 60962
rect 15340 60880 15380 60920
rect 17548 60880 17588 60920
rect 18124 60880 18164 60920
rect 19372 60880 19412 60920
rect 1708 60796 1748 60836
rect 11020 60796 11060 60836
rect 20044 60796 20084 60836
rect 1516 60628 1556 60668
rect 3340 60628 3380 60668
rect 4972 60628 5012 60668
rect 6604 60628 6644 60668
rect 8332 60628 8372 60668
rect 14284 60628 14324 60668
rect 17740 60628 17780 60668
rect 19564 60628 19604 60668
rect 20236 60628 20276 60668
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 2956 60292 2996 60332
rect 14092 60292 14132 60332
rect 17164 60292 17204 60332
rect 17548 60292 17588 60332
rect 7084 60124 7124 60164
rect 7180 60124 7220 60164
rect 1516 60040 1556 60080
rect 2764 60040 2804 60080
rect 3244 60040 3284 60080
rect 3340 60040 3380 60080
rect 3724 60040 3764 60080
rect 3820 60040 3860 60080
rect 4300 60040 4340 60080
rect 4780 60054 4820 60094
rect 6604 60040 6644 60080
rect 8188 60082 8228 60122
rect 11020 60124 11060 60164
rect 11116 60124 11156 60164
rect 16588 60124 16628 60164
rect 16972 60124 17012 60164
rect 17356 60124 17396 60164
rect 18316 60124 18356 60164
rect 6700 60040 6740 60080
rect 7660 60040 7700 60080
rect 10540 60040 10580 60080
rect 12124 60082 12164 60122
rect 18412 60124 18452 60164
rect 19756 60124 19796 60164
rect 10636 60040 10676 60080
rect 11596 60040 11636 60080
rect 12652 60040 12692 60080
rect 13900 60040 13940 60080
rect 14380 60040 14420 60080
rect 14476 60040 14516 60080
rect 14860 60040 14900 60080
rect 14956 60040 14996 60080
rect 15436 60040 15476 60080
rect 15916 60045 15956 60085
rect 17836 60040 17876 60080
rect 19420 60082 19460 60122
rect 17932 60040 17972 60080
rect 18892 60040 18932 60080
rect 8332 59956 8372 59996
rect 12268 59956 12308 59996
rect 4972 59872 5012 59912
rect 14092 59872 14132 59912
rect 16108 59872 16148 59912
rect 16780 59872 16820 59912
rect 19564 59872 19604 59912
rect 19948 59872 19988 59912
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 12748 59536 12788 59576
rect 13036 59536 13076 59576
rect 14764 59536 14804 59576
rect 16396 59536 16436 59576
rect 2956 59452 2996 59492
rect 8044 59452 8084 59492
rect 9772 59452 9812 59492
rect 11788 59452 11828 59492
rect 19564 59452 19604 59492
rect 1228 59368 1268 59408
rect 2476 59368 2516 59408
rect 3148 59363 3188 59403
rect 3628 59368 3668 59408
rect 4108 59368 4148 59408
rect 4588 59368 4628 59408
rect 4684 59368 4724 59408
rect 6316 59368 6356 59408
rect 6412 59368 6452 59408
rect 6892 59368 6932 59408
rect 7372 59368 7412 59408
rect 7852 59363 7892 59403
rect 8332 59368 8372 59408
rect 9580 59368 9620 59408
rect 10060 59368 10100 59408
rect 10156 59368 10196 59408
rect 10540 59368 10580 59408
rect 10636 59368 10676 59408
rect 11116 59368 11156 59408
rect 11596 59354 11636 59394
rect 12556 59368 12596 59408
rect 12652 59368 12692 59408
rect 12844 59368 12884 59408
rect 13228 59368 13268 59408
rect 14476 59368 14516 59408
rect 14668 59368 14708 59408
rect 14956 59368 14996 59408
rect 16204 59368 16244 59408
rect 17836 59368 17876 59408
rect 17932 59368 17972 59408
rect 18316 59368 18356 59408
rect 18412 59368 18452 59408
rect 18892 59368 18932 59408
rect 19420 59358 19460 59398
rect 4204 59284 4244 59324
rect 5164 59284 5204 59324
rect 6796 59284 6836 59324
rect 16972 59284 17012 59324
rect 17356 59284 17396 59324
rect 19756 59284 19796 59324
rect 4972 59200 5012 59240
rect 17164 59200 17204 59240
rect 2668 59116 2708 59156
rect 17548 59116 17588 59156
rect 19948 59116 19988 59156
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 11500 58780 11540 58820
rect 9868 58612 9908 58652
rect 12940 58612 12980 58652
rect 17260 58612 17300 58652
rect 17644 58612 17684 58652
rect 19660 58612 19700 58652
rect 20044 58612 20084 58652
rect 1420 58528 1460 58568
rect 2668 58528 2708 58568
rect 3052 58528 3092 58568
rect 4300 58528 4340 58568
rect 4684 58528 4724 58568
rect 5932 58528 5972 58568
rect 6316 58528 6356 58568
rect 7564 58528 7604 58568
rect 8044 58528 8084 58568
rect 9292 58528 9332 58568
rect 10060 58528 10100 58568
rect 11308 58528 11348 58568
rect 13708 58528 13748 58568
rect 14956 58528 14996 58568
rect 15340 58528 15380 58568
rect 16588 58528 16628 58568
rect 18028 58528 18068 58568
rect 19276 58528 19316 58568
rect 2860 58360 2900 58400
rect 4492 58360 4532 58400
rect 6124 58360 6164 58400
rect 7756 58360 7796 58400
rect 9484 58360 9524 58400
rect 9676 58360 9716 58400
rect 12748 58360 12788 58400
rect 15148 58360 15188 58400
rect 16780 58360 16820 58400
rect 17452 58360 17492 58400
rect 17836 58360 17876 58400
rect 19468 58360 19508 58400
rect 19852 58360 19892 58400
rect 20236 58360 20276 58400
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 9676 58024 9716 58064
rect 3148 57940 3188 57980
rect 5260 57940 5300 57980
rect 1708 57856 1748 57896
rect 2956 57856 2996 57896
rect 3532 57856 3572 57896
rect 3628 57856 3668 57896
rect 4012 57856 4052 57896
rect 4108 57856 4148 57896
rect 4588 57856 4628 57896
rect 5068 57851 5108 57891
rect 6220 57856 6260 57896
rect 7468 57856 7508 57896
rect 7948 57856 7988 57896
rect 8044 57856 8084 57896
rect 8428 57856 8468 57896
rect 8524 57856 8564 57896
rect 9004 57856 9044 57896
rect 9484 57851 9524 57891
rect 10156 57856 10196 57896
rect 11404 57856 11444 57896
rect 11884 57856 11924 57896
rect 13132 57856 13172 57896
rect 14092 57856 14132 57896
rect 15340 57856 15380 57896
rect 15724 57856 15764 57896
rect 16972 57856 17012 57896
rect 17548 57856 17588 57896
rect 18796 57856 18836 57896
rect 19084 57856 19124 57896
rect 1516 57772 1556 57812
rect 1324 57688 1364 57728
rect 7660 57604 7700 57644
rect 11596 57604 11636 57644
rect 13324 57604 13364 57644
rect 15532 57604 15572 57644
rect 17164 57604 17204 57644
rect 17356 57604 17396 57644
rect 19564 57604 19604 57644
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 1708 57100 1748 57140
rect 2092 57100 2132 57140
rect 3532 57100 3572 57140
rect 3628 57100 3668 57140
rect 11980 57100 12020 57140
rect 2572 57030 2612 57070
rect 3052 57016 3092 57056
rect 4012 57016 4052 57056
rect 4108 57016 4148 57056
rect 4396 57016 4436 57056
rect 5644 57016 5684 57056
rect 6220 57016 6260 57056
rect 6316 57016 6356 57056
rect 6700 57016 6740 57056
rect 6796 57016 6836 57056
rect 7276 57016 7316 57056
rect 7756 57030 7796 57070
rect 8140 57016 8180 57056
rect 9388 57016 9428 57056
rect 9772 57016 9812 57056
rect 11020 57016 11060 57056
rect 11500 57035 11540 57075
rect 11596 57016 11636 57056
rect 13084 57058 13124 57098
rect 14092 57100 14132 57140
rect 16012 57100 16052 57140
rect 19756 57100 19796 57140
rect 12076 57016 12116 57056
rect 12556 57016 12596 57056
rect 13516 57016 13556 57056
rect 13612 57016 13652 57056
rect 13996 57016 14036 57056
rect 14572 57016 14612 57056
rect 15052 57025 15092 57065
rect 15628 57016 15668 57056
rect 15724 57016 15764 57056
rect 15916 57016 15956 57056
rect 16204 57016 16244 57056
rect 16396 57016 16436 57056
rect 16492 57016 16532 57056
rect 16684 57016 16724 57056
rect 16876 57016 16916 57056
rect 16972 57016 17012 57056
rect 17068 57016 17108 57056
rect 17356 57016 17396 57056
rect 17548 57016 17588 57056
rect 17836 57016 17876 57056
rect 17932 57016 17972 57056
rect 18316 57016 18356 57056
rect 18412 57016 18452 57056
rect 18892 57016 18932 57056
rect 19372 57030 19412 57070
rect 7948 56932 7988 56972
rect 13228 56932 13268 56972
rect 1516 56848 1556 56888
rect 1900 56848 1940 56888
rect 2380 56848 2420 56888
rect 5836 56848 5876 56888
rect 9580 56848 9620 56888
rect 11212 56848 11252 56888
rect 15244 56848 15284 56888
rect 16588 56848 16628 56888
rect 17164 56848 17204 56888
rect 17452 56848 17492 56888
rect 19564 56848 19604 56888
rect 19948 56848 19988 56888
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 1228 56512 1268 56552
rect 5356 56512 5396 56552
rect 16972 56512 17012 56552
rect 17452 56512 17492 56552
rect 3052 56428 3092 56468
rect 10156 56428 10196 56468
rect 13804 56428 13844 56468
rect 1612 56344 1652 56384
rect 2860 56344 2900 56384
rect 3628 56344 3668 56384
rect 3724 56344 3764 56384
rect 4684 56344 4724 56384
rect 5164 56339 5204 56379
rect 6028 56344 6068 56384
rect 7276 56344 7316 56384
rect 8524 56344 8564 56384
rect 9772 56344 9812 56384
rect 10348 56339 10388 56379
rect 10828 56344 10868 56384
rect 11308 56344 11348 56384
rect 11404 56344 11444 56384
rect 11788 56344 11828 56384
rect 11884 56344 11924 56384
rect 12364 56344 12404 56384
rect 13612 56344 13652 56384
rect 15244 56344 15284 56384
rect 15340 56344 15380 56384
rect 15724 56344 15764 56384
rect 16300 56344 16340 56384
rect 16780 56339 16820 56379
rect 17164 56344 17204 56384
rect 17644 56344 17684 56384
rect 1420 56260 1460 56300
rect 4108 56260 4148 56300
rect 4204 56260 4244 56300
rect 17260 56302 17300 56342
rect 17356 56302 17396 56342
rect 17836 56344 17876 56384
rect 18124 56344 18164 56384
rect 19372 56344 19412 56384
rect 15820 56260 15860 56300
rect 19756 56260 19796 56300
rect 7468 56092 7508 56132
rect 9964 56092 10004 56132
rect 17644 56092 17684 56132
rect 19564 56092 19604 56132
rect 19948 56092 19988 56132
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 3244 55672 3284 55712
rect 3052 55588 3092 55628
rect 3436 55588 3476 55628
rect 8812 55588 8852 55628
rect 13612 55588 13652 55628
rect 19372 55588 19412 55628
rect 19756 55588 19796 55628
rect 1228 55504 1268 55544
rect 2476 55504 2516 55544
rect 4684 55504 4724 55544
rect 5932 55504 5972 55544
rect 6508 55504 6548 55544
rect 7756 55504 7796 55544
rect 8236 55504 8276 55544
rect 8332 55504 8372 55544
rect 8716 55504 8756 55544
rect 9292 55504 9332 55544
rect 9820 55513 9860 55553
rect 11500 55504 11540 55544
rect 11596 55504 11636 55544
rect 11980 55504 12020 55544
rect 12076 55504 12116 55544
rect 12556 55504 12596 55544
rect 13084 55513 13124 55553
rect 15820 55504 15860 55544
rect 17068 55504 17108 55544
rect 17452 55504 17492 55544
rect 18700 55504 18740 55544
rect 7948 55420 7988 55460
rect 13228 55420 13268 55460
rect 17260 55420 17300 55460
rect 2668 55336 2708 55376
rect 2860 55336 2900 55376
rect 6124 55336 6164 55376
rect 9964 55336 10004 55376
rect 13420 55336 13460 55376
rect 18892 55336 18932 55376
rect 19564 55336 19604 55376
rect 19948 55336 19988 55376
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 11500 55000 11540 55040
rect 13228 55000 13268 55040
rect 13420 55000 13460 55040
rect 2476 54916 2516 54956
rect 7756 54916 7796 54956
rect 16108 54916 16148 54956
rect 19564 54916 19604 54956
rect 2668 54818 2708 54858
rect 3148 54832 3188 54872
rect 3628 54832 3668 54872
rect 4108 54832 4148 54872
rect 4204 54832 4244 54872
rect 6028 54832 6068 54872
rect 6124 54832 6164 54872
rect 6604 54832 6644 54872
rect 7084 54832 7124 54872
rect 7564 54827 7604 54867
rect 8428 54832 8468 54872
rect 9676 54832 9716 54872
rect 10060 54832 10100 54872
rect 11308 54832 11348 54872
rect 11788 54832 11828 54872
rect 13036 54832 13076 54872
rect 14380 54832 14420 54872
rect 14476 54832 14516 54872
rect 14956 54832 14996 54872
rect 15436 54832 15476 54872
rect 15916 54818 15956 54858
rect 16396 54832 16436 54872
rect 16684 54832 16724 54872
rect 16780 54832 16820 54872
rect 17836 54832 17876 54872
rect 17932 54832 17972 54872
rect 18412 54832 18452 54872
rect 18892 54832 18932 54872
rect 19372 54827 19412 54867
rect 1708 54748 1748 54788
rect 2092 54748 2132 54788
rect 3724 54748 3764 54788
rect 6508 54748 6548 54788
rect 13612 54748 13652 54788
rect 14860 54748 14900 54788
rect 18316 54748 18356 54788
rect 19756 54748 19796 54788
rect 17068 54664 17108 54704
rect 1516 54580 1556 54620
rect 1900 54580 1940 54620
rect 9868 54580 9908 54620
rect 19948 54580 19988 54620
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 14668 54244 14708 54284
rect 16300 54244 16340 54284
rect 4012 54160 4052 54200
rect 17836 54160 17876 54200
rect 1708 54076 1748 54116
rect 2092 54076 2132 54116
rect 11404 54076 11444 54116
rect 17644 54076 17684 54116
rect 19660 54076 19700 54116
rect 20044 54076 20084 54116
rect 2572 53992 2612 54032
rect 3820 53992 3860 54032
rect 4396 53992 4436 54032
rect 5644 53992 5684 54032
rect 6316 53992 6356 54032
rect 7564 53992 7604 54032
rect 8044 53992 8084 54032
rect 8140 53992 8180 54032
rect 8524 53992 8564 54032
rect 9628 54034 9668 54074
rect 8620 53992 8660 54032
rect 9100 53992 9140 54032
rect 11596 53992 11636 54032
rect 12844 53992 12884 54032
rect 13228 53992 13268 54032
rect 14476 53992 14516 54032
rect 14860 53992 14900 54032
rect 16108 53992 16148 54032
rect 18028 53992 18068 54032
rect 19276 53992 19316 54032
rect 9772 53908 9812 53948
rect 1516 53824 1556 53864
rect 1900 53824 1940 53864
rect 5836 53824 5876 53864
rect 7756 53824 7796 53864
rect 11212 53824 11252 53864
rect 13036 53824 13076 53864
rect 19468 53824 19508 53864
rect 19852 53824 19892 53864
rect 20236 53824 20276 53864
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 5740 53488 5780 53528
rect 13324 53488 13364 53528
rect 3532 53404 3572 53444
rect 11308 53404 11348 53444
rect 15436 53404 15476 53444
rect 2092 53320 2132 53360
rect 3340 53320 3380 53360
rect 4012 53320 4052 53360
rect 4108 53320 4148 53360
rect 5068 53320 5108 53360
rect 5596 53310 5636 53350
rect 8236 53320 8276 53360
rect 9484 53320 9524 53360
rect 9868 53320 9908 53360
rect 11116 53320 11156 53360
rect 11596 53320 11636 53360
rect 11692 53320 11732 53360
rect 12076 53320 12116 53360
rect 12652 53320 12692 53360
rect 13132 53315 13172 53355
rect 13708 53320 13748 53360
rect 13804 53320 13844 53360
rect 14188 53320 14228 53360
rect 14764 53320 14804 53360
rect 15244 53306 15284 53346
rect 15628 53320 15668 53360
rect 15916 53320 15956 53360
rect 17164 53320 17204 53360
rect 18316 53320 18356 53360
rect 19564 53320 19604 53360
rect 1516 53236 1556 53276
rect 1900 53236 1940 53276
rect 4492 53236 4532 53276
rect 4588 53236 4628 53276
rect 12172 53236 12212 53276
rect 14284 53236 14324 53276
rect 19948 53236 19988 53276
rect 1324 53068 1364 53108
rect 1708 53068 1748 53108
rect 9676 53068 9716 53108
rect 15724 53068 15764 53108
rect 17356 53068 17396 53108
rect 19756 53068 19796 53108
rect 20140 53068 20180 53108
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 14380 52648 14420 52688
rect 15532 52648 15572 52688
rect 17932 52564 17972 52604
rect 18028 52564 18068 52604
rect 19372 52564 19412 52604
rect 19756 52564 19796 52604
rect 1516 52480 1556 52520
rect 2764 52480 2804 52520
rect 3244 52480 3284 52520
rect 3340 52480 3380 52520
rect 3724 52480 3764 52520
rect 3820 52480 3860 52520
rect 4300 52480 4340 52520
rect 4780 52485 4820 52525
rect 6604 52480 6644 52520
rect 7852 52480 7892 52520
rect 8332 52480 8372 52520
rect 8428 52480 8468 52520
rect 8812 52480 8852 52520
rect 8908 52480 8948 52520
rect 9388 52480 9428 52520
rect 9868 52494 9908 52534
rect 12940 52480 12980 52520
rect 14188 52480 14228 52520
rect 14860 52480 14900 52520
rect 15148 52480 15188 52520
rect 15244 52480 15284 52520
rect 15724 52480 15764 52520
rect 16972 52480 17012 52520
rect 17452 52480 17492 52520
rect 17548 52480 17588 52520
rect 18508 52480 18548 52520
rect 18988 52494 19028 52534
rect 2956 52396 2996 52436
rect 4972 52396 5012 52436
rect 8044 52396 8084 52436
rect 10060 52396 10100 52436
rect 17164 52396 17204 52436
rect 19180 52312 19220 52352
rect 19564 52312 19604 52352
rect 19948 52312 19988 52352
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 4588 51976 4628 52016
rect 6220 51976 6260 52016
rect 13708 51976 13748 52016
rect 8236 51892 8276 51932
rect 11692 51892 11732 51932
rect 16012 51892 16052 51932
rect 19084 51892 19124 51932
rect 1516 51808 1556 51848
rect 2764 51808 2804 51848
rect 3148 51808 3188 51848
rect 4396 51808 4436 51848
rect 4780 51808 4820 51848
rect 6028 51808 6068 51848
rect 6508 51808 6548 51848
rect 6604 51808 6644 51848
rect 6988 51808 7028 51848
rect 7084 51808 7124 51848
rect 7564 51808 7604 51848
rect 8044 51794 8084 51834
rect 9292 51808 9332 51848
rect 9580 51808 9620 51848
rect 9964 51808 10004 51848
rect 10060 51808 10100 51848
rect 10540 51808 10580 51848
rect 11020 51808 11060 51848
rect 11500 51794 11540 51834
rect 12268 51808 12308 51848
rect 13516 51808 13556 51848
rect 14092 51808 14132 51848
rect 14380 51808 14420 51848
rect 14572 51808 14612 51848
rect 15820 51808 15860 51848
rect 16204 51808 16244 51848
rect 16396 51808 16436 51848
rect 16589 51819 16629 51859
rect 16780 51808 16820 51848
rect 17356 51808 17396 51848
rect 17452 51808 17492 51848
rect 17836 51808 17876 51848
rect 17932 51808 17972 51848
rect 18412 51808 18452 51848
rect 18892 51803 18932 51843
rect 8620 51724 8660 51764
rect 10444 51724 10484 51764
rect 14188 51724 14228 51764
rect 16300 51724 16340 51764
rect 19372 51724 19412 51764
rect 19756 51724 19796 51764
rect 2956 51640 2996 51680
rect 19564 51640 19604 51680
rect 19948 51640 19988 51680
rect 8428 51556 8468 51596
rect 9292 51556 9332 51596
rect 16588 51556 16628 51596
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 7948 51220 7988 51260
rect 9964 51220 10004 51260
rect 11788 51220 11828 51260
rect 15436 51220 15476 51260
rect 3052 51052 3092 51092
rect 4588 51052 4628 51092
rect 1228 50968 1268 51008
rect 2476 50968 2516 51008
rect 4012 50968 4052 51008
rect 4108 50968 4148 51008
rect 4492 50968 4532 51008
rect 5068 50968 5108 51008
rect 5548 50973 5588 51013
rect 6508 50968 6548 51008
rect 7756 50968 7796 51008
rect 8524 50968 8564 51008
rect 9772 50968 9812 51008
rect 10348 50968 10388 51008
rect 11596 50968 11636 51008
rect 12748 50968 12788 51008
rect 13996 50968 14036 51008
rect 14476 50968 14516 51008
rect 14572 50968 14612 51008
rect 14668 50968 14708 51008
rect 14764 50968 14804 51008
rect 14956 50968 14996 51008
rect 15052 50968 15092 51008
rect 15148 50968 15188 51008
rect 15244 50968 15284 51008
rect 15436 50968 15476 51008
rect 15628 50968 15668 51008
rect 15724 50968 15764 51008
rect 16300 50968 16340 51008
rect 17548 50968 17588 51008
rect 18316 50968 18356 51008
rect 19564 50968 19604 51008
rect 5740 50884 5780 50924
rect 2668 50800 2708 50840
rect 2860 50800 2900 50840
rect 14188 50800 14228 50840
rect 17740 50800 17780 50840
rect 20140 50842 20180 50882
rect 19756 50800 19796 50840
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 5740 50464 5780 50504
rect 9196 50380 9236 50420
rect 14284 50380 14324 50420
rect 2668 50296 2708 50336
rect 3916 50296 3956 50336
rect 4300 50296 4340 50336
rect 5548 50296 5588 50336
rect 5932 50296 5972 50336
rect 7180 50296 7220 50336
rect 7756 50296 7796 50336
rect 9004 50296 9044 50336
rect 9484 50296 9524 50336
rect 9964 50296 10004 50336
rect 10060 50296 10100 50336
rect 10348 50296 10388 50336
rect 10828 50296 10868 50336
rect 12076 50296 12116 50336
rect 12556 50296 12596 50336
rect 12652 50296 12692 50336
rect 13612 50296 13652 50336
rect 1708 50212 1748 50252
rect 2092 50212 2132 50252
rect 2476 50212 2516 50252
rect 13036 50212 13076 50252
rect 13132 50254 13172 50294
rect 14140 50286 14180 50326
rect 14476 50296 14516 50336
rect 15724 50296 15764 50336
rect 16108 50296 16148 50336
rect 17356 50275 17396 50315
rect 17932 50296 17972 50336
rect 19180 50296 19220 50336
rect 19372 50212 19412 50252
rect 12268 50128 12308 50168
rect 19564 50128 19604 50168
rect 19948 50128 19988 50168
rect 1516 50044 1556 50084
rect 1900 50044 1940 50084
rect 2284 50044 2324 50084
rect 4108 50044 4148 50084
rect 7372 50044 7412 50084
rect 9388 50044 9428 50084
rect 9676 50044 9716 50084
rect 15916 50044 15956 50084
rect 17548 50044 17588 50084
rect 17740 50044 17780 50084
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 8140 49708 8180 49748
rect 8908 49540 8948 49580
rect 9004 49540 9044 49580
rect 18604 49540 18644 49580
rect 2764 49456 2804 49496
rect 2860 49456 2900 49496
rect 3244 49456 3284 49496
rect 3340 49456 3380 49496
rect 3820 49456 3860 49496
rect 4300 49470 4340 49510
rect 4684 49456 4724 49496
rect 5932 49456 5972 49496
rect 6700 49456 6740 49496
rect 7948 49456 7988 49496
rect 8428 49456 8468 49496
rect 8524 49456 8564 49496
rect 9484 49456 9524 49496
rect 9964 49470 10004 49510
rect 10348 49456 10388 49496
rect 10444 49456 10484 49496
rect 10540 49464 10580 49504
rect 10828 49456 10868 49496
rect 11020 49456 11060 49496
rect 11212 49456 11252 49496
rect 12460 49456 12500 49496
rect 12940 49456 12980 49496
rect 13036 49456 13076 49496
rect 13420 49456 13460 49496
rect 13516 49456 13556 49496
rect 13996 49456 14036 49496
rect 14524 49465 14564 49505
rect 15052 49456 15092 49496
rect 16300 49456 16340 49496
rect 18028 49456 18068 49496
rect 18124 49456 18164 49496
rect 19612 49498 19652 49538
rect 18508 49456 18548 49496
rect 19084 49456 19124 49496
rect 10156 49372 10196 49412
rect 12652 49372 12692 49412
rect 14860 49372 14900 49412
rect 4492 49288 4532 49328
rect 6124 49288 6164 49328
rect 10636 49288 10676 49328
rect 10924 49288 10964 49328
rect 14668 49288 14708 49328
rect 19756 49246 19796 49286
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 1900 48952 1940 48992
rect 9868 48952 9908 48992
rect 10348 48952 10388 48992
rect 7660 48868 7700 48908
rect 17260 48868 17300 48908
rect 19756 48868 19796 48908
rect 2572 48784 2612 48824
rect 3820 48784 3860 48824
rect 4204 48784 4244 48824
rect 5452 48784 5492 48824
rect 5932 48784 5972 48824
rect 6028 48784 6068 48824
rect 6508 48784 6548 48824
rect 6988 48784 7028 48824
rect 7468 48779 7508 48819
rect 7948 48784 7988 48824
rect 8044 48784 8084 48824
rect 8236 48784 8276 48824
rect 8428 48784 8468 48824
rect 9676 48784 9716 48824
rect 10060 48784 10100 48824
rect 10156 48784 10196 48824
rect 10252 48784 10292 48824
rect 10636 48784 10676 48824
rect 11884 48784 11924 48824
rect 13132 48784 13172 48824
rect 14380 48784 14420 48824
rect 15532 48784 15572 48824
rect 15628 48784 15668 48824
rect 16108 48784 16148 48824
rect 16588 48784 16628 48824
rect 17116 48774 17156 48814
rect 18028 48784 18068 48824
rect 18124 48784 18164 48824
rect 18508 48784 18548 48824
rect 18604 48784 18644 48824
rect 19084 48784 19124 48824
rect 19612 48774 19652 48814
rect 1708 48700 1748 48740
rect 2092 48700 2132 48740
rect 6412 48700 6452 48740
rect 16012 48700 16052 48740
rect 1516 48532 1556 48572
rect 4012 48532 4052 48572
rect 5644 48532 5684 48572
rect 8236 48532 8276 48572
rect 12076 48532 12116 48572
rect 14572 48532 14612 48572
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 1516 48196 1556 48236
rect 1708 48028 1748 48068
rect 2092 48028 2132 48068
rect 2476 48028 2516 48068
rect 3340 48028 3380 48068
rect 8716 48028 8756 48068
rect 2764 47944 2804 47984
rect 2860 47944 2900 47984
rect 3244 47944 3284 47984
rect 3820 47944 3860 47984
rect 4300 47958 4340 47998
rect 4780 47944 4820 47984
rect 6028 47944 6068 47984
rect 6412 47944 6452 47984
rect 7660 47944 7700 47984
rect 8620 47944 8660 47984
rect 10252 47986 10292 48026
rect 8812 47944 8852 47984
rect 9004 47944 9044 47984
rect 11020 47944 11060 47984
rect 12268 47944 12308 47984
rect 12748 47944 12788 47984
rect 12844 47944 12884 47984
rect 13228 47944 13268 47984
rect 13324 47944 13364 47984
rect 13804 47944 13844 47984
rect 14284 47958 14324 47998
rect 14668 47944 14708 47984
rect 15916 47944 15956 47984
rect 16492 47944 16532 47984
rect 17740 47944 17780 47984
rect 18124 47944 18164 47984
rect 19372 47944 19412 47984
rect 4492 47860 4532 47900
rect 12460 47860 12500 47900
rect 1900 47776 1940 47816
rect 2284 47776 2324 47816
rect 6220 47776 6260 47816
rect 7852 47776 7892 47816
rect 10444 47776 10484 47816
rect 14476 47776 14516 47816
rect 16108 47776 16148 47816
rect 16300 47776 16340 47816
rect 17932 47776 17972 47816
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 7948 47440 7988 47480
rect 12076 47440 12116 47480
rect 3340 47356 3380 47396
rect 5548 47356 5588 47396
rect 17164 47356 17204 47396
rect 20044 47356 20084 47396
rect 1900 47272 1940 47312
rect 3148 47272 3188 47312
rect 3820 47272 3860 47312
rect 3916 47272 3956 47312
rect 4300 47272 4340 47312
rect 4396 47272 4436 47312
rect 4876 47272 4916 47312
rect 5404 47262 5444 47302
rect 6220 47272 6260 47312
rect 6316 47272 6356 47312
rect 6700 47272 6740 47312
rect 6796 47272 6836 47312
rect 7276 47272 7316 47312
rect 7804 47262 7844 47302
rect 8524 47272 8564 47312
rect 9772 47272 9812 47312
rect 10348 47272 10388 47312
rect 10444 47272 10484 47312
rect 10924 47272 10964 47312
rect 11404 47272 11444 47312
rect 11932 47262 11972 47302
rect 12940 47272 12980 47312
rect 14188 47272 14228 47312
rect 15436 47272 15476 47312
rect 15532 47272 15572 47312
rect 15916 47272 15956 47312
rect 16012 47272 16052 47312
rect 16492 47272 16532 47312
rect 16972 47267 17012 47307
rect 18316 47272 18356 47312
rect 18412 47272 18452 47312
rect 18796 47272 18836 47312
rect 18892 47272 18932 47312
rect 19372 47272 19412 47312
rect 19852 47258 19892 47298
rect 1708 47188 1748 47228
rect 10828 47188 10868 47228
rect 1516 47020 1556 47060
rect 9964 47020 10004 47060
rect 14380 47020 14420 47060
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 2668 46600 2708 46640
rect 3052 46516 3092 46556
rect 3436 46516 3476 46556
rect 8716 46516 8756 46556
rect 1228 46432 1268 46472
rect 2476 46432 2516 46472
rect 4108 46432 4148 46472
rect 5356 46432 5396 46472
rect 6412 46432 6452 46472
rect 7660 46432 7700 46472
rect 8140 46432 8180 46472
rect 8236 46432 8276 46472
rect 9724 46474 9764 46514
rect 18892 46516 18932 46556
rect 18988 46516 19028 46556
rect 8620 46432 8660 46472
rect 9196 46432 9236 46472
rect 10924 46432 10964 46472
rect 12172 46432 12212 46472
rect 12652 46432 12692 46472
rect 12748 46432 12788 46472
rect 13132 46432 13172 46472
rect 13228 46432 13268 46472
rect 13708 46432 13748 46472
rect 14188 46446 14228 46486
rect 15724 46432 15764 46472
rect 16972 46432 17012 46472
rect 18412 46432 18452 46472
rect 18508 46432 18548 46472
rect 19468 46432 19508 46472
rect 19948 46437 19988 46477
rect 7852 46348 7892 46388
rect 9868 46348 9908 46388
rect 12364 46348 12404 46388
rect 14380 46348 14420 46388
rect 2860 46264 2900 46304
rect 3244 46264 3284 46304
rect 5548 46264 5588 46304
rect 17164 46264 17204 46304
rect 20140 46264 20180 46304
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 2284 45928 2324 45968
rect 18892 45928 18932 45968
rect 4396 45760 4436 45800
rect 5644 45760 5684 45800
rect 8716 45760 8756 45800
rect 9964 45760 10004 45800
rect 10348 45760 10388 45800
rect 11596 45760 11636 45800
rect 14956 45760 14996 45800
rect 15820 45760 15860 45800
rect 17068 45760 17108 45800
rect 17452 45760 17492 45800
rect 18700 45760 18740 45800
rect 13708 45718 13748 45758
rect 1708 45676 1748 45716
rect 2092 45676 2132 45716
rect 2476 45676 2516 45716
rect 2860 45676 2900 45716
rect 19372 45676 19412 45716
rect 19756 45676 19796 45716
rect 1516 45508 1556 45548
rect 1900 45508 1940 45548
rect 2668 45508 2708 45548
rect 5836 45508 5876 45548
rect 10156 45508 10196 45548
rect 11788 45508 11828 45548
rect 15148 45508 15188 45548
rect 17260 45508 17300 45548
rect 19564 45508 19604 45548
rect 19948 45508 19988 45548
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 18316 45172 18356 45212
rect 19948 45172 19988 45212
rect 1420 45004 1460 45044
rect 1804 45004 1844 45044
rect 4204 45004 4244 45044
rect 4300 45004 4340 45044
rect 1996 44920 2036 44960
rect 3244 44920 3284 44960
rect 3724 44920 3764 44960
rect 5308 44962 5348 45002
rect 8428 45004 8468 45044
rect 10732 45004 10772 45044
rect 3820 44920 3860 44960
rect 4780 44920 4820 44960
rect 6124 44920 6164 44960
rect 7372 44920 7412 44960
rect 7852 44920 7892 44960
rect 7948 44920 7988 44960
rect 8332 44920 8372 44960
rect 8908 44920 8948 44960
rect 9436 44929 9476 44969
rect 10156 44920 10196 44960
rect 10252 44920 10292 44960
rect 11740 44962 11780 45002
rect 15916 45004 15956 45044
rect 16012 45004 16052 45044
rect 18124 45004 18164 45044
rect 10636 44920 10676 44960
rect 11212 44920 11252 44960
rect 12172 44920 12212 44960
rect 13420 44920 13460 44960
rect 15436 44920 15476 44960
rect 17020 44962 17060 45002
rect 15532 44920 15572 44960
rect 16492 44920 16532 44960
rect 18508 44920 18548 44960
rect 19756 44920 19796 44960
rect 5452 44836 5492 44876
rect 7564 44836 7604 44876
rect 9580 44836 9620 44876
rect 1228 44752 1268 44792
rect 1612 44752 1652 44792
rect 3436 44752 3476 44792
rect 11884 44752 11924 44792
rect 13612 44752 13652 44792
rect 17164 44752 17204 44792
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 9580 44416 9620 44456
rect 17164 44416 17204 44456
rect 17932 44416 17972 44456
rect 18316 44416 18356 44456
rect 20044 44416 20084 44456
rect 5548 44332 5588 44372
rect 11692 44332 11732 44372
rect 13708 44332 13748 44372
rect 1996 44248 2036 44288
rect 3244 44248 3284 44288
rect 3820 44248 3860 44288
rect 3916 44248 3956 44288
rect 4300 44248 4340 44288
rect 4396 44248 4436 44288
rect 4876 44248 4916 44288
rect 5404 44238 5444 44278
rect 6412 44248 6452 44288
rect 7660 44248 7700 44288
rect 8140 44248 8180 44288
rect 9388 44248 9428 44288
rect 10252 44248 10292 44288
rect 11500 44248 11540 44288
rect 11980 44248 12020 44288
rect 12076 44248 12116 44288
rect 12556 44248 12596 44288
rect 13036 44248 13076 44288
rect 13564 44238 13604 44278
rect 15436 44229 15476 44269
rect 15532 44248 15572 44288
rect 15916 44248 15956 44288
rect 16012 44248 16052 44288
rect 16492 44248 16532 44288
rect 16972 44243 17012 44283
rect 18604 44248 18644 44288
rect 19852 44248 19892 44288
rect 1804 44164 1844 44204
rect 12460 44164 12500 44204
rect 15148 44164 15188 44204
rect 17740 44164 17780 44204
rect 18124 44164 18164 44204
rect 3436 44080 3476 44120
rect 14956 44080 14996 44120
rect 1612 43996 1652 44036
rect 7852 43996 7892 44036
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 15244 43660 15284 43700
rect 17740 43660 17780 43700
rect 18796 43660 18836 43700
rect 19564 43660 19604 43700
rect 19948 43660 19988 43700
rect 13132 43576 13172 43616
rect 11884 43492 11924 43532
rect 13324 43492 13364 43532
rect 17548 43492 17588 43532
rect 17932 43492 17972 43532
rect 18604 43492 18644 43532
rect 18988 43492 19028 43532
rect 19372 43492 19412 43532
rect 19756 43492 19796 43532
rect 2188 43408 2228 43448
rect 3436 43408 3476 43448
rect 3820 43408 3860 43448
rect 3916 43408 3956 43448
rect 4108 43408 4148 43448
rect 6412 43408 6452 43448
rect 6604 43408 6644 43448
rect 6796 43408 6836 43448
rect 6892 43408 6932 43448
rect 7084 43408 7124 43448
rect 7276 43408 7316 43448
rect 7372 43408 7412 43448
rect 7756 43408 7796 43448
rect 7852 43408 7892 43448
rect 8044 43408 8084 43448
rect 8236 43408 8276 43448
rect 8332 43408 8372 43448
rect 9388 43408 9428 43448
rect 13804 43408 13844 43448
rect 15052 43408 15092 43448
rect 6508 43324 6548 43364
rect 3628 43240 3668 43280
rect 4012 43240 4052 43280
rect 6988 43240 7028 43280
rect 7564 43240 7604 43280
rect 8140 43240 8180 43280
rect 9292 43240 9332 43280
rect 11692 43240 11732 43280
rect 18124 43240 18164 43280
rect 19180 43240 19220 43280
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 8524 42904 8564 42944
rect 17356 42904 17396 42944
rect 4780 42820 4820 42860
rect 9484 42820 9524 42860
rect 2764 42736 2804 42776
rect 2956 42736 2996 42776
rect 3052 42736 3092 42776
rect 3244 42736 3284 42776
rect 3436 42736 3476 42776
rect 3532 42736 3572 42776
rect 3724 42736 3764 42776
rect 3820 42736 3860 42776
rect 3916 42736 3956 42776
rect 4012 42736 4052 42776
rect 4204 42757 4244 42797
rect 4300 42757 4340 42797
rect 4396 42736 4436 42776
rect 4492 42736 4532 42776
rect 4684 42736 4724 42776
rect 4876 42736 4916 42776
rect 5260 42736 5300 42776
rect 6508 42736 6548 42776
rect 7372 42736 7412 42776
rect 7756 42736 7796 42776
rect 8140 42736 8180 42776
rect 8332 42736 8372 42776
rect 8428 42736 8468 42776
rect 8620 42736 8660 42776
rect 8716 42736 8756 42776
rect 8873 42721 8913 42761
rect 9100 42736 9140 42776
rect 9292 42736 9332 42776
rect 9676 42736 9716 42776
rect 10924 42736 10964 42776
rect 11500 42736 11540 42776
rect 12748 42736 12788 42776
rect 13132 42736 13172 42776
rect 14380 42736 14420 42776
rect 7852 42652 7892 42692
rect 8044 42652 8084 42692
rect 14956 42652 14996 42692
rect 16108 42652 16148 42692
rect 16588 42652 16628 42692
rect 17164 42652 17204 42692
rect 17740 42652 17780 42692
rect 18124 42652 18164 42692
rect 18796 42652 18836 42692
rect 19372 42652 19412 42692
rect 19756 42652 19796 42692
rect 3340 42568 3380 42608
rect 6988 42568 7028 42608
rect 7372 42568 7412 42608
rect 7948 42568 7988 42608
rect 9196 42568 9236 42608
rect 15148 42568 15188 42608
rect 16300 42568 16340 42608
rect 16780 42568 16820 42608
rect 17932 42568 17972 42608
rect 18316 42568 18356 42608
rect 18988 42568 19028 42608
rect 19564 42568 19604 42608
rect 2764 42484 2804 42524
rect 6700 42484 6740 42524
rect 7564 42484 7604 42524
rect 12940 42484 12980 42524
rect 14572 42484 14612 42524
rect 19948 42484 19988 42524
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 15148 42148 15188 42188
rect 17836 42148 17876 42188
rect 18220 42148 18260 42188
rect 18604 42148 18644 42188
rect 18988 42148 19028 42188
rect 19372 42148 19412 42188
rect 20140 42148 20180 42188
rect 3532 42064 3572 42104
rect 4108 42064 4148 42104
rect 4396 42064 4436 42104
rect 14956 41980 14996 42020
rect 17644 41980 17684 42020
rect 18028 41980 18068 42020
rect 18412 41980 18452 42020
rect 18796 41980 18836 42020
rect 19180 41980 19220 42020
rect 19564 41980 19604 42020
rect 19948 41980 19988 42020
rect 1228 41896 1268 41936
rect 2476 41896 2516 41936
rect 2860 41896 2900 41936
rect 3052 41896 3092 41936
rect 3148 41896 3188 41936
rect 3340 41896 3380 41936
rect 3532 41896 3572 41936
rect 3628 41896 3668 41936
rect 3820 41896 3860 41936
rect 4012 41896 4052 41936
rect 4108 41896 4148 41936
rect 4588 41896 4628 41936
rect 4684 41896 4724 41936
rect 4780 41896 4820 41936
rect 4876 41896 4916 41936
rect 5260 41896 5300 41936
rect 6508 41896 6548 41936
rect 6892 41906 6932 41946
rect 6988 41896 7028 41936
rect 7372 41896 7412 41936
rect 7564 41896 7604 41936
rect 7660 41896 7700 41936
rect 8044 41896 8084 41936
rect 8140 41896 8180 41936
rect 8812 41896 8852 41936
rect 8908 41896 8948 41936
rect 9196 41896 9236 41936
rect 9292 41896 9332 41936
rect 9388 41896 9428 41936
rect 9868 41896 9908 41936
rect 11116 41896 11156 41936
rect 11308 41896 11348 41936
rect 12556 41896 12596 41936
rect 13036 41896 13076 41936
rect 13132 41896 13172 41936
rect 13516 41896 13556 41936
rect 13612 41896 13652 41936
rect 14092 41896 14132 41936
rect 14572 41910 14612 41950
rect 15724 41896 15764 41936
rect 15820 41896 15860 41936
rect 16204 41896 16244 41936
rect 16300 41896 16340 41936
rect 16780 41896 16820 41936
rect 17308 41905 17348 41945
rect 2956 41812 2996 41852
rect 6700 41812 6740 41852
rect 8236 41812 8276 41852
rect 14764 41812 14804 41852
rect 17452 41812 17492 41852
rect 2668 41728 2708 41768
rect 7180 41728 7220 41768
rect 7852 41728 7892 41768
rect 8332 41728 8372 41768
rect 8428 41728 8468 41768
rect 8620 41728 8660 41768
rect 9484 41728 9524 41768
rect 9676 41728 9716 41768
rect 12748 41728 12788 41768
rect 19756 41728 19796 41768
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 2956 41392 2996 41432
rect 4396 41392 4436 41432
rect 6508 41392 6548 41432
rect 8044 41392 8084 41432
rect 8524 41392 8564 41432
rect 9292 41392 9332 41432
rect 10252 41392 10292 41432
rect 15628 41392 15668 41432
rect 17356 41392 17396 41432
rect 19756 41392 19796 41432
rect 20236 41392 20276 41432
rect 7948 41308 7988 41348
rect 10732 41308 10772 41348
rect 1228 41224 1268 41264
rect 2476 41224 2516 41264
rect 2860 41224 2900 41264
rect 3148 41224 3188 41264
rect 3340 41224 3380 41264
rect 3436 41224 3476 41264
rect 3628 41224 3668 41264
rect 4012 41224 4052 41264
rect 4204 41224 4244 41264
rect 4307 41223 4347 41263
rect 4492 41224 4532 41264
rect 4684 41224 4724 41264
rect 4780 41224 4820 41264
rect 4876 41224 4916 41264
rect 5068 41224 5108 41264
rect 6316 41224 6356 41264
rect 6700 41224 6740 41264
rect 6988 41224 7028 41264
rect 7372 41224 7412 41264
rect 7756 41224 7796 41264
rect 3724 41140 3764 41180
rect 3916 41140 3956 41180
rect 6796 41140 6836 41180
rect 7274 41182 7314 41222
rect 7852 41224 7892 41264
rect 8332 41224 8372 41264
rect 8428 41224 8468 41264
rect 8620 41224 8660 41264
rect 8812 41224 8852 41264
rect 8908 41224 8948 41264
rect 9004 41224 9044 41264
rect 9100 41224 9140 41264
rect 9292 41224 9332 41264
rect 9484 41224 9524 41264
rect 9580 41224 9620 41264
rect 9868 41224 9908 41264
rect 9964 41224 10004 41264
rect 10060 41224 10100 41264
rect 10444 41224 10484 41264
rect 10540 41224 10580 41264
rect 10636 41224 10676 41264
rect 10924 41224 10964 41264
rect 11020 41224 11060 41264
rect 11116 41245 11156 41285
rect 11212 41224 11252 41264
rect 13228 41224 13268 41264
rect 13420 41224 13460 41264
rect 13612 41224 13652 41264
rect 13804 41224 13844 41264
rect 13900 41224 13940 41264
rect 14188 41224 14228 41264
rect 15436 41224 15476 41264
rect 15916 41224 15956 41264
rect 17164 41224 17204 41264
rect 17932 41224 17972 41264
rect 19180 41224 19220 41264
rect 19564 41224 19604 41264
rect 19660 41210 19700 41250
rect 19852 41224 19892 41264
rect 7084 41140 7124 41180
rect 17548 41140 17588 41180
rect 20044 41140 20084 41180
rect 2668 41056 2708 41096
rect 3436 41056 3476 41096
rect 3820 41056 3860 41096
rect 2956 40972 2996 41012
rect 7180 41014 7220 41054
rect 8044 40972 8084 41012
rect 13420 40972 13460 41012
rect 13612 40972 13652 41012
rect 17740 40972 17780 41012
rect 19372 40972 19412 41012
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 6220 40636 6260 40676
rect 6988 40636 7028 40676
rect 7180 40636 7220 40676
rect 8140 40636 8180 40676
rect 8332 40636 8372 40676
rect 13324 40636 13364 40676
rect 15436 40636 15476 40676
rect 4972 40552 5012 40592
rect 6028 40552 6068 40592
rect 6796 40552 6836 40592
rect 9100 40552 9140 40592
rect 9772 40552 9812 40592
rect 3052 40468 3092 40508
rect 7276 40468 7316 40508
rect 9676 40468 9716 40508
rect 9868 40468 9908 40508
rect 16204 40468 16244 40508
rect 2188 40384 2228 40424
rect 2284 40384 2324 40424
rect 2572 40384 2612 40424
rect 2668 40384 2708 40424
rect 3148 40384 3188 40424
rect 3628 40384 3668 40424
rect 4108 40398 4148 40438
rect 4492 40384 4532 40424
rect 4588 40384 4628 40424
rect 4684 40384 4724 40424
rect 4780 40384 4820 40424
rect 4972 40384 5012 40424
rect 5260 40384 5300 40424
rect 5836 40384 5876 40424
rect 6220 40384 6260 40424
rect 6412 40384 6452 40424
rect 6508 40384 6548 40424
rect 6796 40384 6836 40424
rect 7173 40401 7213 40441
rect 7468 40384 7508 40424
rect 7852 40384 7892 40424
rect 7948 40384 7988 40424
rect 8140 40384 8180 40424
rect 8332 40384 8372 40424
rect 8524 40384 8564 40424
rect 8620 40384 8660 40424
rect 8908 40384 8948 40424
rect 9100 40384 9140 40424
rect 9580 40384 9620 40424
rect 9964 40384 10004 40424
rect 10156 40384 10196 40424
rect 10252 40384 10292 40424
rect 10348 40384 10388 40424
rect 10444 40384 10484 40424
rect 10636 40384 10676 40424
rect 11500 40426 11540 40466
rect 10828 40384 10868 40424
rect 12748 40384 12788 40424
rect 13324 40384 13364 40424
rect 13516 40384 13556 40424
rect 13612 40384 13652 40424
rect 13996 40384 14036 40424
rect 15244 40384 15284 40424
rect 15724 40384 15764 40424
rect 15820 40384 15860 40424
rect 16300 40384 16340 40424
rect 16780 40384 16820 40424
rect 17260 40389 17300 40429
rect 18220 40384 18260 40424
rect 19468 40384 19508 40424
rect 19852 40384 19892 40424
rect 19948 40384 19988 40424
rect 20044 40384 20084 40424
rect 20140 40384 20180 40424
rect 4300 40300 4340 40340
rect 10732 40300 10772 40340
rect 17452 40300 17492 40340
rect 1996 40216 2036 40256
rect 5740 40216 5780 40256
rect 9292 40216 9332 40256
rect 12940 40216 12980 40256
rect 19660 40216 19700 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 2572 39880 2612 39920
rect 6700 39880 6740 39920
rect 9004 39880 9044 39920
rect 14476 39880 14516 39920
rect 15436 39880 15476 39920
rect 17164 39880 17204 39920
rect 19852 39880 19892 39920
rect 4972 39796 5012 39836
rect 9772 39796 9812 39836
rect 12748 39796 12788 39836
rect 13708 39796 13748 39836
rect 2476 39712 2516 39752
rect 2764 39712 2804 39752
rect 4012 39712 4052 39752
rect 4396 39712 4436 39752
rect 4492 39712 4532 39752
rect 4588 39712 4628 39752
rect 4684 39712 4724 39752
rect 4876 39712 4916 39752
rect 5068 39712 5108 39752
rect 5260 39712 5300 39752
rect 6508 39712 6548 39752
rect 6892 39712 6932 39752
rect 7276 39712 7316 39752
rect 7372 39712 7412 39752
rect 7756 39712 7796 39752
rect 7852 39712 7892 39752
rect 8332 39712 8372 39752
rect 8812 39698 8852 39738
rect 9388 39712 9428 39752
rect 9676 39712 9716 39752
rect 10348 39712 10388 39752
rect 10540 39712 10580 39752
rect 10636 39712 10676 39752
rect 11308 39712 11348 39752
rect 12556 39712 12596 39752
rect 12940 39712 12980 39752
rect 13324 39712 13364 39752
rect 13612 39739 13652 39779
rect 14188 39712 14228 39752
rect 14284 39712 14324 39752
rect 14380 39712 14420 39752
rect 14668 39712 14708 39752
rect 14764 39712 14804 39752
rect 14860 39712 14900 39752
rect 14956 39712 14996 39752
rect 15148 39712 15188 39752
rect 15244 39712 15284 39752
rect 15340 39712 15380 39752
rect 15724 39712 15764 39752
rect 16972 39712 17012 39752
rect 18124 39732 18164 39772
rect 18220 39712 18260 39752
rect 19180 39712 19220 39752
rect 19660 39707 19700 39747
rect 18604 39628 18644 39668
rect 18700 39628 18740 39668
rect 6988 39544 7028 39584
rect 10060 39544 10100 39584
rect 4204 39460 4244 39500
rect 10348 39460 10388 39500
rect 13036 39460 13076 39500
rect 13996 39460 14036 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 12556 39124 12596 39164
rect 14092 39124 14132 39164
rect 17740 39124 17780 39164
rect 9772 39040 9812 39080
rect 12268 39040 12308 39080
rect 3628 38956 3668 38996
rect 5740 38956 5780 38996
rect 7756 38956 7796 38996
rect 3052 38872 3092 38912
rect 3148 38872 3188 38912
rect 3532 38872 3572 38912
rect 4108 38872 4148 38912
rect 4588 38886 4628 38926
rect 5260 38872 5300 38912
rect 5356 38872 5396 38912
rect 5836 38872 5876 38912
rect 6316 38872 6356 38912
rect 6844 38881 6884 38921
rect 7276 38872 7316 38912
rect 7372 38872 7412 38912
rect 7852 38872 7892 38912
rect 8332 38872 8372 38912
rect 8812 38886 8852 38926
rect 9580 38872 9620 38912
rect 9772 38872 9812 38912
rect 9964 38872 10004 38912
rect 11212 38872 11252 38912
rect 11788 38872 11828 38912
rect 11884 38872 11924 38912
rect 11980 38872 12020 38912
rect 12364 38872 12404 38912
rect 12652 38872 12692 38912
rect 12844 38872 12884 38912
rect 12940 38872 12980 38912
rect 13036 38872 13076 38912
rect 13132 38872 13172 38912
rect 13420 38872 13460 38912
rect 13708 38872 13748 38912
rect 14284 38872 14324 38912
rect 14380 38872 14420 38912
rect 14572 38872 14612 38912
rect 16300 38872 16340 38912
rect 17548 38872 17588 38912
rect 18412 38872 18452 38912
rect 18508 38872 18548 38912
rect 18892 38872 18932 38912
rect 18988 38872 19028 38912
rect 19468 38872 19508 38912
rect 19948 38877 19988 38917
rect 6988 38788 7028 38828
rect 9004 38788 9044 38828
rect 13804 38788 13844 38828
rect 14476 38788 14516 38828
rect 20140 38788 20180 38828
rect 2668 38704 2708 38744
rect 4780 38704 4820 38744
rect 11404 38704 11444 38744
rect 11596 38704 11636 38744
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 2668 38368 2708 38408
rect 3052 38368 3092 38408
rect 5356 38368 5396 38408
rect 6988 38368 7028 38408
rect 10732 38368 10772 38408
rect 18892 38368 18932 38408
rect 19564 38368 19604 38408
rect 17260 38284 17300 38324
rect 1228 38200 1268 38240
rect 2476 38200 2516 38240
rect 3916 38200 3956 38240
rect 5164 38200 5204 38240
rect 5548 38200 5588 38240
rect 6796 38200 6836 38240
rect 9292 38200 9332 38240
rect 10540 38200 10580 38240
rect 11116 38200 11156 38240
rect 11212 38200 11252 38240
rect 11308 38200 11348 38240
rect 11404 38200 11444 38240
rect 12652 38200 12692 38240
rect 13900 38200 13940 38240
rect 15532 38200 15572 38240
rect 15628 38200 15668 38240
rect 16108 38200 16148 38240
rect 16588 38200 16628 38240
rect 17452 38200 17492 38240
rect 18700 38200 18740 38240
rect 16012 38116 16052 38156
rect 17116 38158 17156 38198
rect 19372 38116 19412 38156
rect 19756 38116 19796 38156
rect 2956 38032 2996 38072
rect 14092 38032 14132 38072
rect 19948 38032 19988 38072
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 2668 37612 2708 37652
rect 15724 37612 15764 37652
rect 17356 37612 17396 37652
rect 19948 37612 19988 37652
rect 1228 37360 1268 37400
rect 2476 37360 2516 37400
rect 3004 37369 3044 37409
rect 3532 37360 3572 37400
rect 4012 37360 4052 37400
rect 4108 37360 4148 37400
rect 4492 37360 4532 37400
rect 4588 37360 4628 37400
rect 5452 37360 5492 37400
rect 5740 37360 5780 37400
rect 5836 37360 5876 37400
rect 5932 37360 5972 37400
rect 6028 37360 6068 37400
rect 6316 37360 6356 37400
rect 6412 37360 6452 37400
rect 6508 37360 6548 37400
rect 6700 37360 6740 37400
rect 7948 37360 7988 37400
rect 8332 37360 8372 37400
rect 9580 37360 9620 37400
rect 10540 37360 10580 37400
rect 11788 37360 11828 37400
rect 12268 37360 12308 37400
rect 12364 37360 12404 37400
rect 12748 37360 12788 37400
rect 12844 37360 12884 37400
rect 13324 37360 13364 37400
rect 13804 37374 13844 37414
rect 14284 37360 14324 37400
rect 15532 37360 15572 37400
rect 15916 37360 15956 37400
rect 17164 37360 17204 37400
rect 18508 37360 18548 37400
rect 19756 37360 19796 37400
rect 13996 37276 14036 37316
rect 2860 37192 2900 37232
rect 5548 37192 5588 37232
rect 6220 37192 6260 37232
rect 8140 37192 8180 37232
rect 9772 37192 9812 37232
rect 11980 37192 12020 37232
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 2668 36856 2708 36896
rect 4300 36856 4340 36896
rect 5932 36856 5972 36896
rect 6796 36856 6836 36896
rect 7660 36856 7700 36896
rect 10060 36856 10100 36896
rect 12268 36856 12308 36896
rect 14476 36856 14516 36896
rect 6220 36772 6260 36812
rect 17356 36772 17396 36812
rect 20044 36772 20084 36812
rect 1228 36688 1268 36728
rect 2476 36688 2516 36728
rect 2860 36688 2900 36728
rect 4108 36688 4148 36728
rect 4492 36688 4532 36728
rect 5740 36688 5780 36728
rect 6124 36688 6164 36728
rect 6316 36688 6356 36728
rect 6412 36669 6452 36709
rect 6604 36688 6644 36728
rect 6700 36688 6740 36728
rect 6892 36688 6932 36728
rect 7084 36688 7124 36728
rect 7276 36688 7316 36728
rect 7372 36688 7412 36728
rect 7564 36688 7604 36728
rect 7756 36688 7796 36728
rect 8332 36688 8372 36728
rect 8428 36688 8468 36728
rect 9388 36688 9428 36728
rect 9868 36683 9908 36723
rect 10828 36688 10868 36728
rect 12076 36688 12116 36728
rect 12748 36688 12788 36728
rect 12844 36688 12884 36728
rect 13804 36688 13844 36728
rect 8812 36604 8852 36644
rect 8908 36604 8948 36644
rect 13228 36604 13268 36644
rect 13324 36604 13364 36644
rect 14332 36646 14372 36686
rect 15628 36688 15668 36728
rect 15724 36688 15764 36728
rect 16684 36688 16724 36728
rect 17164 36674 17204 36714
rect 18316 36688 18356 36728
rect 18412 36688 18452 36728
rect 18892 36688 18932 36728
rect 19372 36688 19412 36728
rect 19852 36674 19892 36714
rect 16108 36604 16148 36644
rect 16204 36604 16244 36644
rect 18796 36604 18836 36644
rect 7084 36520 7124 36560
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 2668 36100 2708 36140
rect 5452 36100 5492 36140
rect 6988 36100 7028 36140
rect 9196 36100 9236 36140
rect 18316 36100 18356 36140
rect 19948 36100 19988 36140
rect 1228 35848 1268 35888
rect 2476 35848 2516 35888
rect 4012 35848 4052 35888
rect 5260 35848 5300 35888
rect 5740 35848 5780 35888
rect 5836 35848 5876 35888
rect 5932 35848 5972 35888
rect 6028 35848 6068 35888
rect 6316 35848 6356 35888
rect 6604 35848 6644 35888
rect 7180 35848 7220 35888
rect 7276 35848 7316 35888
rect 7468 35848 7508 35888
rect 7564 35848 7604 35888
rect 7756 35848 7796 35888
rect 9004 35848 9044 35888
rect 9484 35848 9524 35888
rect 9580 35848 9620 35888
rect 9964 35848 10004 35888
rect 10060 35848 10100 35888
rect 10540 35848 10580 35888
rect 11068 35857 11108 35897
rect 11404 35848 11444 35888
rect 12652 35848 12692 35888
rect 13420 35848 13460 35888
rect 14668 35848 14708 35888
rect 15052 35848 15092 35888
rect 16300 35848 16340 35888
rect 16876 35848 16916 35888
rect 18124 35848 18164 35888
rect 18508 35848 18548 35888
rect 19756 35848 19796 35888
rect 6700 35764 6740 35804
rect 11212 35764 11252 35804
rect 5452 35680 5492 35720
rect 12844 35680 12884 35720
rect 14860 35680 14900 35720
rect 16492 35680 16532 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 11116 35344 11156 35384
rect 3724 35260 3764 35300
rect 6028 35260 6068 35300
rect 13996 35260 14036 35300
rect 1996 35176 2036 35216
rect 2092 35176 2132 35216
rect 2572 35176 2612 35216
rect 3052 35176 3092 35216
rect 3532 35162 3572 35202
rect 5260 35176 5300 35216
rect 5356 35176 5396 35216
rect 5452 35176 5492 35216
rect 5548 35176 5588 35216
rect 5740 35176 5780 35216
rect 5836 35176 5876 35216
rect 5932 35176 5972 35216
rect 6316 35176 6356 35216
rect 6604 35176 6644 35216
rect 6700 35176 6740 35216
rect 7180 35176 7220 35216
rect 9676 35176 9716 35216
rect 10924 35176 10964 35216
rect 12268 35176 12308 35216
rect 12364 35176 12404 35216
rect 13324 35176 13364 35216
rect 13804 35162 13844 35202
rect 15628 35176 15668 35216
rect 16876 35176 16916 35216
rect 17260 35176 17300 35216
rect 18508 35176 18548 35216
rect 2476 35092 2516 35132
rect 12748 35092 12788 35132
rect 12844 35092 12884 35132
rect 6988 35008 7028 35048
rect 7276 34924 7316 34964
rect 17068 34924 17108 34964
rect 18700 34924 18740 34964
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 3244 34588 3284 34628
rect 13804 34588 13844 34628
rect 5452 34504 5492 34544
rect 1804 34336 1844 34376
rect 3052 34336 3092 34376
rect 4012 34336 4052 34376
rect 5260 34336 5300 34376
rect 5740 34336 5780 34376
rect 5836 34336 5876 34376
rect 6124 34336 6164 34376
rect 6220 34336 6260 34376
rect 6316 34336 6356 34376
rect 6508 34336 6548 34376
rect 6604 34336 6644 34376
rect 6796 34336 6836 34376
rect 6988 34336 7028 34376
rect 7084 34336 7124 34376
rect 7180 34336 7220 34376
rect 7276 34336 7316 34376
rect 7564 34336 7604 34376
rect 8812 34336 8852 34376
rect 9292 34316 9332 34356
rect 9388 34336 9428 34376
rect 9772 34336 9812 34376
rect 9868 34336 9908 34376
rect 10348 34336 10388 34376
rect 10828 34341 10868 34381
rect 12364 34336 12404 34376
rect 13612 34336 13652 34376
rect 14188 34336 14228 34376
rect 15436 34336 15476 34376
rect 15820 34336 15860 34376
rect 17068 34336 17108 34376
rect 17836 34336 17876 34376
rect 17932 34336 17972 34376
rect 18316 34336 18356 34376
rect 18412 34336 18452 34376
rect 18892 34336 18932 34376
rect 19372 34341 19412 34381
rect 6700 34252 6740 34292
rect 11020 34252 11060 34292
rect 19564 34252 19604 34292
rect 6028 34168 6068 34208
rect 9004 34168 9044 34208
rect 13996 34168 14036 34208
rect 15628 34168 15668 34208
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 4012 33832 4052 33872
rect 7372 33832 7412 33872
rect 9004 33832 9044 33872
rect 10636 33832 10676 33872
rect 12652 33832 12692 33872
rect 16396 33832 16436 33872
rect 18028 33832 18068 33872
rect 20236 33832 20276 33872
rect 5740 33748 5780 33788
rect 2284 33664 2324 33704
rect 2380 33664 2420 33704
rect 3340 33664 3380 33704
rect 3820 33650 3860 33690
rect 4300 33664 4340 33704
rect 5548 33664 5588 33704
rect 5932 33664 5972 33704
rect 6028 33664 6068 33704
rect 6316 33664 6356 33704
rect 6604 33664 6644 33704
rect 6700 33664 6740 33704
rect 7180 33664 7220 33704
rect 7276 33664 7316 33704
rect 7468 33664 7508 33704
rect 7660 33664 7700 33704
rect 7852 33664 7892 33704
rect 7948 33664 7988 33704
rect 8236 33664 8276 33704
rect 8428 33664 8468 33704
rect 8524 33664 8564 33704
rect 8716 33664 8756 33704
rect 8812 33664 8852 33704
rect 9196 33664 9236 33704
rect 10444 33664 10484 33704
rect 10924 33664 10964 33704
rect 11020 33664 11060 33704
rect 11404 33664 11444 33704
rect 11980 33664 12020 33704
rect 12460 33650 12500 33690
rect 12940 33664 12980 33704
rect 14188 33664 14228 33704
rect 14668 33664 14708 33704
rect 14764 33664 14804 33704
rect 15724 33664 15764 33704
rect 16204 33659 16244 33699
rect 16588 33664 16628 33704
rect 17836 33664 17876 33704
rect 18508 33664 18548 33704
rect 18604 33664 18644 33704
rect 19564 33664 19604 33704
rect 20044 33650 20084 33690
rect 2764 33580 2804 33620
rect 2860 33580 2900 33620
rect 11500 33580 11540 33620
rect 15148 33580 15188 33620
rect 15244 33580 15284 33620
rect 18988 33580 19028 33620
rect 19084 33580 19124 33620
rect 6988 33496 7028 33536
rect 7660 33496 7700 33536
rect 8524 33496 8564 33536
rect 14380 33412 14420 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 2668 33076 2708 33116
rect 5644 33076 5684 33116
rect 6988 33076 7028 33116
rect 12460 33076 12500 33116
rect 19372 33076 19412 33116
rect 9196 32992 9236 33032
rect 10828 32992 10868 33032
rect 5932 32908 5972 32948
rect 1228 32824 1268 32864
rect 2476 32824 2516 32864
rect 4204 32824 4244 32864
rect 5452 32824 5492 32864
rect 5836 32824 5876 32864
rect 6028 32824 6068 32864
rect 6316 32824 6356 32864
rect 6604 32824 6644 32864
rect 7180 32824 7220 32864
rect 7276 32824 7316 32864
rect 7372 32824 7412 32864
rect 7468 32824 7508 32864
rect 7756 32824 7796 32864
rect 9004 32824 9044 32864
rect 9388 32824 9428 32864
rect 10636 32824 10676 32864
rect 12268 32824 12308 32864
rect 14764 32824 14804 32864
rect 11020 32782 11060 32822
rect 14860 32824 14900 32864
rect 15244 32824 15284 32864
rect 15340 32824 15380 32864
rect 15820 32824 15860 32864
rect 16348 32833 16388 32873
rect 17932 32824 17972 32864
rect 19180 32824 19220 32864
rect 6700 32740 6740 32780
rect 16492 32740 16532 32780
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 5452 32320 5492 32360
rect 9100 32320 9140 32360
rect 9484 32320 9524 32360
rect 16492 32320 16532 32360
rect 3724 32236 3764 32276
rect 12172 32236 12212 32276
rect 14188 32236 14228 32276
rect 19468 32236 19508 32276
rect 1996 32152 2036 32192
rect 2092 32152 2132 32192
rect 2572 32152 2612 32192
rect 3052 32152 3092 32192
rect 3532 32138 3572 32178
rect 5740 32152 5780 32192
rect 6988 32152 7028 32192
rect 7660 32152 7700 32192
rect 8908 32152 8948 32192
rect 9292 32152 9332 32192
rect 9388 32152 9428 32192
rect 9580 32152 9620 32192
rect 9676 32152 9716 32192
rect 9777 32152 9817 32192
rect 10060 32152 10100 32192
rect 10156 32152 10196 32192
rect 10732 32152 10772 32192
rect 11980 32152 12020 32192
rect 12460 32152 12500 32192
rect 12556 32152 12596 32192
rect 13516 32152 13556 32192
rect 13996 32138 14036 32178
rect 15052 32152 15092 32192
rect 16300 32152 16340 32192
rect 17740 32152 17780 32192
rect 17836 32152 17876 32192
rect 18220 32152 18260 32192
rect 18796 32152 18836 32192
rect 19276 32138 19316 32178
rect 2476 32068 2516 32108
rect 12940 32068 12980 32108
rect 13036 32068 13076 32108
rect 18316 32068 18356 32108
rect 7180 31900 7220 31940
rect 9292 31900 9332 31940
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 14092 31564 14132 31604
rect 18124 31564 18164 31604
rect 3052 31480 3092 31520
rect 8044 31396 8084 31436
rect 10060 31396 10100 31436
rect 10156 31396 10196 31436
rect 15340 31396 15380 31436
rect 18988 31396 19028 31436
rect 1612 31312 1652 31352
rect 2860 31312 2900 31352
rect 3340 31312 3380 31352
rect 3436 31312 3476 31352
rect 3820 31312 3860 31352
rect 3916 31312 3956 31352
rect 4396 31312 4436 31352
rect 4876 31317 4916 31357
rect 5548 31312 5588 31352
rect 5644 31312 5684 31352
rect 6028 31312 6068 31352
rect 6124 31312 6164 31352
rect 6604 31312 6644 31352
rect 7084 31326 7124 31366
rect 7564 31312 7604 31352
rect 7660 31312 7700 31352
rect 8140 31312 8180 31352
rect 8620 31312 8660 31352
rect 9100 31317 9140 31357
rect 9580 31312 9620 31352
rect 9676 31312 9716 31352
rect 10636 31312 10676 31352
rect 11164 31321 11204 31361
rect 12652 31312 12692 31352
rect 13900 31312 13940 31352
rect 14380 31312 14420 31352
rect 14764 31312 14804 31352
rect 14860 31312 14900 31352
rect 15244 31312 15284 31352
rect 15820 31312 15860 31352
rect 16300 31317 16340 31357
rect 16684 31312 16724 31352
rect 17932 31312 17972 31352
rect 18412 31312 18452 31352
rect 18508 31312 18548 31352
rect 18892 31312 18932 31352
rect 19468 31312 19508 31352
rect 19948 31317 19988 31357
rect 5068 31228 5108 31268
rect 7276 31228 7316 31268
rect 9292 31144 9332 31184
rect 11308 31144 11348 31184
rect 14284 31144 14324 31184
rect 16492 31144 16532 31184
rect 20140 31144 20180 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 2668 30808 2708 30848
rect 5260 30808 5300 30848
rect 5452 30808 5492 30848
rect 7468 30808 7508 30848
rect 9676 30808 9716 30848
rect 11308 30808 11348 30848
rect 15052 30808 15092 30848
rect 16684 30808 16724 30848
rect 18316 30808 18356 30848
rect 20236 30808 20276 30848
rect 1228 30640 1268 30680
rect 2476 30640 2516 30680
rect 3820 30640 3860 30680
rect 5068 30640 5108 30680
rect 6028 30640 6068 30680
rect 7276 30640 7316 30680
rect 8236 30640 8276 30680
rect 9484 30640 9524 30680
rect 9868 30640 9908 30680
rect 11116 30640 11156 30680
rect 11500 30640 11540 30680
rect 12748 30640 12788 30680
rect 13132 30640 13172 30680
rect 13228 30640 13268 30680
rect 13324 30640 13364 30680
rect 13420 30640 13460 30680
rect 13612 30640 13652 30680
rect 14860 30640 14900 30680
rect 15244 30640 15284 30680
rect 16492 30640 16532 30680
rect 16876 30640 16916 30680
rect 18124 30640 18164 30680
rect 18796 30640 18836 30680
rect 20044 30640 20084 30680
rect 12940 30388 12980 30428
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 5740 30052 5780 30092
rect 9004 30052 9044 30092
rect 17452 30052 17492 30092
rect 14092 29968 14132 30008
rect 2956 29884 2996 29924
rect 2380 29800 2420 29840
rect 2476 29800 2516 29840
rect 2860 29800 2900 29840
rect 3436 29800 3476 29840
rect 3964 29809 4004 29849
rect 4300 29800 4340 29840
rect 5548 29800 5588 29840
rect 6316 29800 6356 29840
rect 6412 29800 6452 29840
rect 12844 29842 12884 29882
rect 6508 29800 6548 29840
rect 6700 29800 6740 29840
rect 7564 29800 7604 29840
rect 8812 29800 8852 29840
rect 11404 29800 11444 29840
rect 11596 29800 11636 29840
rect 13420 29800 13460 29840
rect 13708 29800 13748 29840
rect 13804 29800 13844 29840
rect 14380 29800 14420 29840
rect 15628 29800 15668 29840
rect 16012 29800 16052 29840
rect 17260 29800 17300 29840
rect 17740 29800 17780 29840
rect 17836 29800 17876 29840
rect 18220 29800 18260 29840
rect 18316 29800 18356 29840
rect 18796 29800 18836 29840
rect 19276 29805 19316 29845
rect 13036 29716 13076 29756
rect 19468 29716 19508 29756
rect 4108 29632 4148 29672
rect 6220 29632 6260 29672
rect 6796 29632 6836 29672
rect 11308 29632 11348 29672
rect 15820 29632 15860 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 3148 29296 3188 29336
rect 4300 29296 4340 29336
rect 9004 29296 9044 29336
rect 12748 29296 12788 29336
rect 17452 29296 17492 29336
rect 19660 29296 19700 29336
rect 6604 29212 6644 29252
rect 11020 29212 11060 29252
rect 1708 29128 1748 29168
rect 2956 29128 2996 29168
rect 4492 29128 4532 29168
rect 5740 29128 5780 29168
rect 6028 29128 6068 29168
rect 6124 29128 6164 29168
rect 6700 29128 6740 29168
rect 6988 29111 7028 29151
rect 7276 29128 7316 29168
rect 7564 29128 7604 29168
rect 8812 29128 8852 29168
rect 9292 29128 9332 29168
rect 9388 29128 9428 29168
rect 9868 29128 9908 29168
rect 10348 29128 10388 29168
rect 10828 29114 10868 29154
rect 11308 29128 11348 29168
rect 12556 29128 12596 29168
rect 12940 29139 12980 29179
rect 13132 29128 13172 29168
rect 13420 29128 13460 29168
rect 13708 29128 13748 29168
rect 13804 29128 13844 29168
rect 14284 29149 14324 29189
rect 14380 29128 14420 29168
rect 14476 29149 14516 29189
rect 14572 29128 14612 29168
rect 14764 29128 14804 29168
rect 14860 29128 14900 29168
rect 14956 29128 14996 29168
rect 15052 29128 15092 29168
rect 15244 29128 15284 29168
rect 15436 29128 15476 29168
rect 15532 29128 15572 29168
rect 16012 29128 16052 29168
rect 17260 29128 17300 29168
rect 17932 29128 17972 29168
rect 18028 29128 18068 29168
rect 18508 29128 18548 29168
rect 18988 29128 19028 29168
rect 19516 29118 19556 29158
rect 9772 29044 9812 29084
rect 18412 29044 18452 29084
rect 14092 28960 14132 29000
rect 6316 28876 6356 28916
rect 7372 28876 7412 28916
rect 12940 28876 12980 28916
rect 15244 28876 15284 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 7084 28540 7124 28580
rect 10828 28540 10868 28580
rect 12364 28540 12404 28580
rect 18220 28540 18260 28580
rect 2668 28288 2708 28328
rect 3916 28288 3956 28328
rect 4300 28288 4340 28328
rect 5548 28288 5588 28328
rect 6412 28288 6452 28328
rect 6700 28288 6740 28328
rect 7276 28288 7316 28328
rect 7468 28288 7508 28328
rect 7564 28288 7604 28328
rect 7756 28288 7796 28328
rect 7852 28288 7892 28328
rect 7948 28288 7988 28328
rect 9388 28288 9428 28328
rect 10636 28288 10676 28328
rect 12460 28288 12500 28328
rect 12748 28288 12788 28328
rect 12844 28288 12884 28328
rect 12940 28288 12980 28328
rect 13132 28288 13172 28328
rect 14380 28288 14420 28328
rect 14860 28288 14900 28328
rect 14956 28288 14996 28328
rect 15340 28288 15380 28328
rect 15436 28288 15476 28328
rect 15916 28288 15956 28328
rect 16444 28297 16484 28337
rect 16780 28288 16820 28328
rect 18028 28288 18068 28328
rect 18508 28288 18548 28328
rect 18604 28288 18644 28328
rect 18988 28288 19028 28328
rect 19084 28288 19124 28328
rect 19564 28288 19604 28328
rect 20044 28293 20084 28333
rect 4108 28204 4148 28244
rect 6796 28204 6836 28244
rect 14572 28204 14612 28244
rect 20236 28204 20276 28244
rect 5740 28120 5780 28160
rect 7372 28120 7412 28160
rect 8044 28120 8084 28160
rect 12652 28120 12692 28160
rect 16588 28120 16628 28160
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 11980 27784 12020 27824
rect 12844 27784 12884 27824
rect 14476 27784 14516 27824
rect 16588 27784 16628 27824
rect 18220 27784 18260 27824
rect 4588 27700 4628 27740
rect 8908 27700 8948 27740
rect 10924 27700 10964 27740
rect 20236 27700 20276 27740
rect 2860 27616 2900 27656
rect 2956 27616 2996 27656
rect 3436 27616 3476 27656
rect 3916 27616 3956 27656
rect 4396 27602 4436 27642
rect 4876 27616 4916 27656
rect 6124 27616 6164 27656
rect 6508 27616 6548 27656
rect 6700 27616 6740 27656
rect 6892 27616 6932 27656
rect 6988 27616 7028 27656
rect 7180 27616 7220 27656
rect 7468 27616 7508 27656
rect 8716 27616 8756 27656
rect 9196 27616 9236 27656
rect 9292 27616 9332 27656
rect 9772 27616 9812 27656
rect 10252 27616 10292 27656
rect 10732 27602 10772 27642
rect 11500 27616 11540 27656
rect 11596 27616 11636 27656
rect 11822 27601 11862 27641
rect 11980 27616 12020 27656
rect 12076 27616 12116 27656
rect 12268 27616 12308 27656
rect 12364 27616 12404 27656
rect 12556 27616 12596 27656
rect 12652 27616 12692 27656
rect 13228 27616 13268 27656
rect 13324 27616 13364 27656
rect 13516 27616 13556 27656
rect 13708 27616 13748 27656
rect 13900 27616 13940 27656
rect 13996 27616 14036 27656
rect 14471 27616 14511 27656
rect 14572 27616 14612 27656
rect 18796 27658 18836 27698
rect 14668 27616 14708 27656
rect 14860 27616 14900 27656
rect 14956 27616 14996 27656
rect 15148 27616 15188 27656
rect 16396 27616 16436 27656
rect 16780 27616 16820 27656
rect 18028 27616 18068 27656
rect 20044 27616 20084 27656
rect 3340 27532 3380 27572
rect 9676 27532 9716 27572
rect 13708 27448 13748 27488
rect 6316 27364 6356 27404
rect 6508 27364 6548 27404
rect 7180 27364 7220 27404
rect 12364 27364 12404 27404
rect 13516 27364 13556 27404
rect 14956 27364 14996 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 6220 27028 6260 27068
rect 10444 27028 10484 27068
rect 14764 27028 14804 27068
rect 4300 26944 4340 26984
rect 7468 26944 7508 26984
rect 12460 26944 12500 26984
rect 15052 26944 15092 26984
rect 16972 26944 17012 26984
rect 2956 26860 2996 26900
rect 2380 26776 2420 26816
rect 2476 26776 2516 26816
rect 3964 26818 4004 26858
rect 17740 26860 17780 26900
rect 2860 26776 2900 26816
rect 3436 26776 3476 26816
rect 4492 26776 4532 26816
rect 5740 26776 5780 26816
rect 5932 26776 5972 26816
rect 6028 26776 6068 26816
rect 6220 26776 6260 26816
rect 6508 26776 6548 26816
rect 6604 26776 6644 26816
rect 6700 26776 6740 26816
rect 6796 26776 6836 26816
rect 6988 26776 7028 26816
rect 7084 26776 7124 26816
rect 7276 26776 7316 26816
rect 7468 26776 7508 26816
rect 7756 26776 7796 26816
rect 8524 26776 8564 26816
rect 8716 26776 8756 26816
rect 8812 26776 8852 26816
rect 9004 26776 9044 26816
rect 10252 26776 10292 26816
rect 10636 26776 10676 26816
rect 11884 26776 11924 26816
rect 12268 26776 12308 26816
rect 12364 26776 12404 26816
rect 12556 26776 12596 26816
rect 13324 26776 13364 26816
rect 14572 26776 14612 26816
rect 14956 26776 14996 26816
rect 15052 26776 15092 26816
rect 15244 26776 15284 26816
rect 15532 26776 15572 26816
rect 16780 26776 16820 26816
rect 17260 26776 17300 26816
rect 17356 26776 17396 26816
rect 17836 26776 17876 26816
rect 18316 26776 18356 26816
rect 18796 26781 18836 26821
rect 18988 26692 19028 26732
rect 4108 26608 4148 26648
rect 7180 26608 7220 26648
rect 8620 26608 8660 26648
rect 12076 26608 12116 26648
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 2668 26272 2708 26312
rect 4492 26272 4532 26312
rect 7564 26272 7604 26312
rect 9964 26272 10004 26312
rect 12076 26272 12116 26312
rect 15052 26272 15092 26312
rect 15532 26272 15572 26312
rect 15724 26272 15764 26312
rect 17932 26272 17972 26312
rect 19948 26272 19988 26312
rect 6124 26188 6164 26228
rect 9292 26188 9332 26228
rect 10444 26188 10484 26228
rect 16108 26188 16148 26228
rect 1228 26104 1268 26144
rect 2476 26104 2516 26144
rect 3052 26104 3092 26144
rect 4300 26104 4340 26144
rect 4684 26104 4724 26144
rect 5932 26104 5972 26144
rect 6412 26104 6452 26144
rect 6508 26062 6548 26102
rect 6604 26089 6644 26129
rect 7372 26104 7412 26144
rect 7660 26104 7700 26144
rect 7852 26104 7892 26144
rect 9100 26104 9140 26144
rect 9580 26104 9620 26144
rect 9676 26104 9716 26144
rect 9772 26104 9812 26144
rect 10156 26104 10196 26144
rect 10252 26104 10292 26144
rect 10348 26104 10388 26144
rect 10636 26104 10676 26144
rect 11884 26104 11924 26144
rect 13612 26104 13652 26144
rect 14860 26104 14900 26144
rect 15244 26104 15284 26144
rect 15345 26094 15385 26134
rect 15820 26104 15860 26144
rect 16012 26104 16052 26144
rect 16204 26104 16244 26144
rect 16300 26104 16340 26144
rect 16492 26104 16532 26144
rect 17740 26104 17780 26144
rect 18220 26104 18260 26144
rect 18316 26104 18356 26144
rect 18700 26104 18740 26144
rect 18796 26104 18836 26144
rect 19276 26104 19316 26144
rect 19804 26094 19844 26134
rect 6796 25852 6836 25892
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 2668 25516 2708 25556
rect 2860 25516 2900 25556
rect 5932 25516 5972 25556
rect 8524 25516 8564 25556
rect 18124 25516 18164 25556
rect 19756 25516 19796 25556
rect 13036 25348 13076 25388
rect 1228 25264 1268 25304
rect 2476 25264 2516 25304
rect 3052 25264 3092 25304
rect 4300 25264 4340 25304
rect 4492 25264 4532 25304
rect 5740 25264 5780 25304
rect 6124 25264 6164 25304
rect 6220 25264 6260 25304
rect 6316 25264 6356 25304
rect 6412 25264 6452 25304
rect 6604 25264 6644 25304
rect 6700 25264 6740 25304
rect 6796 25264 6836 25304
rect 7084 25264 7124 25304
rect 8332 25264 8372 25304
rect 8908 25264 8948 25304
rect 10156 25264 10196 25304
rect 10828 25264 10868 25304
rect 12076 25264 12116 25304
rect 12556 25264 12596 25304
rect 12652 25264 12692 25304
rect 13132 25264 13172 25304
rect 13612 25264 13652 25304
rect 14140 25273 14180 25313
rect 15148 25264 15188 25304
rect 15340 25264 15380 25304
rect 15532 25264 15572 25304
rect 15628 25264 15668 25304
rect 15724 25264 15764 25304
rect 15820 25264 15860 25304
rect 16012 25264 16052 25304
rect 16108 25264 16148 25304
rect 16204 25264 16244 25304
rect 16300 25264 16340 25304
rect 16684 25264 16724 25304
rect 17932 25264 17972 25304
rect 18316 25264 18356 25304
rect 19564 25264 19604 25304
rect 8716 25180 8756 25220
rect 12268 25180 12308 25220
rect 15244 25180 15284 25220
rect 6892 25096 6932 25136
rect 14284 25096 14324 25136
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 3916 24760 3956 24800
rect 11884 24760 11924 24800
rect 14188 24760 14228 24800
rect 16396 24760 16436 24800
rect 7564 24676 7604 24716
rect 9580 24676 9620 24716
rect 18220 24676 18260 24716
rect 20236 24676 20276 24716
rect 1612 24592 1652 24632
rect 1900 24592 1940 24632
rect 2188 24592 2228 24632
rect 2284 24592 2324 24632
rect 2764 24592 2804 24632
rect 3244 24592 3284 24632
rect 3724 24578 3764 24618
rect 4300 24592 4340 24632
rect 5548 24592 5588 24632
rect 6124 24592 6164 24632
rect 7372 24592 7412 24632
rect 7852 24592 7892 24632
rect 7948 24592 7988 24632
rect 8332 24592 8372 24632
rect 8428 24592 8468 24632
rect 8908 24592 8948 24632
rect 9388 24587 9428 24627
rect 9964 24592 10004 24632
rect 10252 24592 10292 24632
rect 10444 24592 10484 24632
rect 11692 24592 11732 24632
rect 12268 24604 12308 24644
rect 12364 24592 12404 24632
rect 12460 24592 12500 24632
rect 12748 24592 12788 24632
rect 13996 24592 14036 24632
rect 14668 24592 14708 24632
rect 15916 24592 15956 24632
rect 16300 24592 16340 24632
rect 16492 24592 16532 24632
rect 16588 24592 16628 24632
rect 16780 24592 16820 24632
rect 18028 24592 18068 24632
rect 18508 24592 18548 24632
rect 18604 24592 18644 24632
rect 18988 24592 19028 24632
rect 19564 24592 19604 24632
rect 20044 24578 20084 24618
rect 2668 24508 2708 24548
rect 19084 24508 19124 24548
rect 1900 24340 1940 24380
rect 5740 24340 5780 24380
rect 10252 24340 10292 24380
rect 11884 24340 11924 24380
rect 12076 24340 12116 24380
rect 16108 24340 16148 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 16012 24004 16052 24044
rect 5644 23920 5684 23960
rect 15820 23920 15860 23960
rect 18604 23920 18644 23960
rect 20236 23920 20276 23960
rect 2764 23836 2804 23876
rect 13228 23836 13268 23876
rect 2284 23752 2324 23792
rect 2380 23752 2420 23792
rect 2860 23752 2900 23792
rect 3340 23752 3380 23792
rect 3868 23761 3908 23801
rect 5932 23794 5972 23834
rect 4204 23752 4244 23792
rect 5452 23752 5492 23792
rect 6028 23752 6068 23792
rect 6124 23752 6164 23792
rect 6508 23752 6548 23792
rect 7756 23752 7796 23792
rect 8332 23752 8372 23792
rect 8428 23752 8468 23792
rect 8812 23752 8852 23792
rect 8908 23752 8948 23792
rect 9388 23752 9428 23792
rect 9868 23757 9908 23797
rect 10444 23752 10484 23792
rect 10636 23752 10676 23792
rect 10732 23752 10772 23792
rect 10924 23752 10964 23792
rect 12172 23752 12212 23792
rect 12652 23752 12692 23792
rect 12748 23752 12788 23792
rect 13132 23752 13172 23792
rect 13708 23752 13748 23792
rect 14236 23761 14276 23801
rect 14572 23752 14612 23792
rect 14668 23731 14708 23771
rect 14764 23731 14804 23771
rect 15148 23752 15188 23792
rect 15436 23752 15476 23792
rect 16300 23752 16340 23792
rect 16396 23752 16436 23792
rect 16684 23752 16724 23792
rect 17164 23752 17204 23792
rect 18412 23752 18452 23792
rect 18796 23752 18836 23792
rect 20044 23752 20084 23792
rect 7948 23668 7988 23708
rect 10060 23668 10100 23708
rect 12364 23668 12404 23708
rect 14380 23668 14420 23708
rect 15532 23668 15572 23708
rect 4012 23584 4052 23624
rect 6316 23584 6356 23624
rect 10540 23584 10580 23624
rect 14860 23584 14900 23624
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 2668 23248 2708 23288
rect 5452 23248 5492 23288
rect 6124 23248 6164 23288
rect 9868 23248 9908 23288
rect 11500 23248 11540 23288
rect 12076 23248 12116 23288
rect 14380 23248 14420 23288
rect 14860 23248 14900 23288
rect 15052 23248 15092 23288
rect 16780 23248 16820 23288
rect 17452 23248 17492 23288
rect 17740 23248 17780 23288
rect 20140 23248 20180 23288
rect 18028 23164 18068 23204
rect 1228 23080 1268 23120
rect 2476 23080 2516 23120
rect 3724 23080 3764 23120
rect 4972 23080 5012 23120
rect 5356 23080 5396 23120
rect 5548 23080 5588 23120
rect 5644 23080 5684 23120
rect 5836 23080 5876 23120
rect 5932 23080 5972 23120
rect 6028 23080 6068 23120
rect 6316 23080 6356 23120
rect 7564 23080 7604 23120
rect 8428 23080 8468 23120
rect 9676 23080 9716 23120
rect 10060 23080 10100 23120
rect 11308 23080 11348 23120
rect 11788 23080 11828 23120
rect 11884 23080 11924 23120
rect 11980 23080 12020 23120
rect 12940 23080 12980 23120
rect 14188 23080 14228 23120
rect 14764 23080 14804 23120
rect 15244 23080 15284 23120
rect 16684 23080 16724 23120
rect 16492 23038 16532 23078
rect 16876 23080 16916 23120
rect 16972 23080 17012 23120
rect 17164 23080 17204 23120
rect 17260 23080 17300 23120
rect 17356 23080 17396 23120
rect 17644 23080 17684 23120
rect 17932 23080 17972 23120
rect 18700 23080 18740 23120
rect 19948 23080 19988 23120
rect 5164 22828 5204 22868
rect 7756 22828 7796 22868
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 2668 22492 2708 22532
rect 4300 22492 4340 22532
rect 15148 22492 15188 22532
rect 18220 22408 18260 22448
rect 5260 22324 5300 22364
rect 5356 22324 5396 22364
rect 8332 22324 8372 22364
rect 12844 22324 12884 22364
rect 18988 22324 19028 22364
rect 19084 22324 19124 22364
rect 1228 22240 1268 22280
rect 2476 22240 2516 22280
rect 2860 22240 2900 22280
rect 4108 22240 4148 22280
rect 4780 22259 4820 22299
rect 4876 22240 4916 22280
rect 5836 22240 5876 22280
rect 6316 22245 6356 22285
rect 7756 22240 7796 22280
rect 7852 22240 7892 22280
rect 8236 22240 8276 22280
rect 8812 22240 8852 22280
rect 9292 22245 9332 22285
rect 10540 22240 10580 22280
rect 11788 22240 11828 22280
rect 12268 22240 12308 22280
rect 12364 22240 12404 22280
rect 12748 22240 12788 22280
rect 13324 22240 13364 22280
rect 13804 22245 13844 22285
rect 14375 22253 14415 22293
rect 14668 22240 14708 22280
rect 14860 22240 14900 22280
rect 14956 22240 14996 22280
rect 15340 22240 15380 22280
rect 16588 22240 16628 22280
rect 16780 22240 16820 22280
rect 18028 22240 18068 22280
rect 18508 22240 18548 22280
rect 18604 22240 18644 22280
rect 19564 22240 19604 22280
rect 20044 22245 20084 22285
rect 11980 22156 12020 22196
rect 20236 22156 20276 22196
rect 6508 22072 6548 22112
rect 9484 22072 9524 22112
rect 13996 22072 14036 22112
rect 14476 22072 14516 22112
rect 14764 22072 14804 22112
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 9292 21736 9332 21776
rect 13708 21736 13748 21776
rect 15340 21736 15380 21776
rect 15724 21736 15764 21776
rect 20140 21736 20180 21776
rect 2476 21652 2516 21692
rect 6220 21652 6260 21692
rect 18124 21652 18164 21692
rect 2668 21554 2708 21594
rect 3148 21568 3188 21608
rect 4108 21568 4148 21608
rect 4204 21568 4244 21608
rect 4780 21568 4820 21608
rect 6028 21568 6068 21608
rect 7852 21568 7892 21608
rect 9100 21568 9140 21608
rect 9484 21568 9524 21608
rect 10732 21568 10772 21608
rect 12268 21568 12308 21608
rect 13516 21568 13556 21608
rect 13900 21568 13940 21608
rect 15148 21568 15188 21608
rect 15532 21568 15572 21608
rect 15628 21568 15668 21608
rect 15820 21568 15860 21608
rect 15916 21568 15956 21608
rect 16017 21568 16057 21608
rect 16684 21568 16724 21608
rect 17932 21568 17972 21608
rect 18412 21568 18452 21608
rect 18508 21568 18548 21608
rect 18892 21568 18932 21608
rect 18988 21568 19028 21608
rect 19468 21568 19508 21608
rect 19948 21554 19988 21594
rect 2092 21484 2132 21524
rect 3628 21484 3668 21524
rect 3724 21484 3764 21524
rect 1900 21316 1940 21356
rect 10924 21316 10964 21356
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 15148 20980 15188 21020
rect 6316 20812 6356 20852
rect 9100 20812 9140 20852
rect 11116 20812 11156 20852
rect 1228 20728 1268 20768
rect 2476 20728 2516 20768
rect 4012 20728 4052 20768
rect 5260 20728 5300 20768
rect 5740 20728 5780 20768
rect 5836 20728 5876 20768
rect 6220 20728 6260 20768
rect 6796 20728 6836 20768
rect 7276 20733 7316 20773
rect 8524 20728 8564 20768
rect 8620 20728 8660 20768
rect 9004 20728 9044 20768
rect 9580 20728 9620 20768
rect 10108 20737 10148 20777
rect 10540 20728 10580 20768
rect 10636 20728 10676 20768
rect 11020 20728 11060 20768
rect 11596 20728 11636 20768
rect 12124 20737 12164 20777
rect 13708 20728 13748 20768
rect 14956 20728 14996 20768
rect 15340 20728 15380 20768
rect 15436 20728 15476 20768
rect 16108 20728 16148 20768
rect 16300 20728 16340 20768
rect 16396 20728 16436 20768
rect 16492 20728 16532 20768
rect 16780 20728 16820 20768
rect 16876 20728 16916 20768
rect 17068 20728 17108 20768
rect 18508 20728 18548 20768
rect 19756 20728 19796 20768
rect 2668 20644 2708 20684
rect 5452 20644 5492 20684
rect 10252 20644 10292 20684
rect 7468 20560 7508 20600
rect 12268 20560 12308 20600
rect 15628 20560 15668 20600
rect 16012 20560 16052 20600
rect 16588 20560 16628 20600
rect 16972 20560 17012 20600
rect 19948 20560 19988 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 2668 20224 2708 20264
rect 6796 20224 6836 20264
rect 8428 20224 8468 20264
rect 10156 20224 10196 20264
rect 12268 20224 12308 20264
rect 16972 20140 17012 20180
rect 20236 20140 20276 20180
rect 1228 20056 1268 20096
rect 2476 20056 2516 20096
rect 3724 20056 3764 20096
rect 4972 20056 5012 20096
rect 5356 20056 5396 20096
rect 6604 20056 6644 20096
rect 6988 20056 7028 20096
rect 8236 20056 8276 20096
rect 8716 20056 8756 20096
rect 9964 20056 10004 20096
rect 10828 20056 10868 20096
rect 12076 20056 12116 20096
rect 12844 20056 12884 20096
rect 14092 20056 14132 20096
rect 14860 20056 14900 20096
rect 16108 20056 16148 20096
rect 16588 20056 16628 20096
rect 16876 20056 16916 20096
rect 17452 20056 17492 20096
rect 17644 20056 17684 20096
rect 17740 20056 17780 20096
rect 17932 20056 17972 20096
rect 18508 20056 18548 20096
rect 18604 20056 18644 20096
rect 18988 20056 19028 20096
rect 19564 20056 19604 20096
rect 20044 20042 20084 20082
rect 19084 19972 19124 20012
rect 17260 19888 17300 19928
rect 5164 19804 5204 19844
rect 14284 19804 14324 19844
rect 16300 19804 16340 19844
rect 17452 19804 17492 19844
rect 18028 19804 18068 19844
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 2668 19468 2708 19508
rect 16780 19468 16820 19508
rect 18412 19468 18452 19508
rect 20044 19468 20084 19508
rect 1228 19216 1268 19256
rect 2476 19216 2516 19256
rect 2956 19216 2996 19256
rect 3052 19216 3092 19256
rect 3436 19216 3476 19256
rect 3532 19216 3572 19256
rect 4012 19216 4052 19256
rect 4492 19230 4532 19270
rect 5356 19216 5396 19256
rect 6604 19216 6644 19256
rect 6988 19216 7028 19256
rect 8236 19216 8276 19256
rect 8716 19216 8756 19256
rect 8812 19216 8852 19256
rect 9196 19216 9236 19256
rect 9292 19216 9332 19256
rect 9772 19216 9812 19256
rect 10252 19221 10292 19261
rect 10828 19216 10868 19256
rect 12076 19216 12116 19256
rect 12556 19216 12596 19256
rect 12652 19216 12692 19256
rect 13036 19216 13076 19256
rect 13132 19216 13172 19256
rect 13612 19216 13652 19256
rect 14140 19225 14180 19265
rect 14668 19216 14708 19256
rect 14860 19216 14900 19256
rect 15052 19216 15092 19256
rect 15148 19216 15188 19256
rect 15340 19216 15380 19256
rect 15628 19216 15668 19256
rect 15724 19216 15764 19256
rect 15820 19216 15860 19256
rect 16108 19216 16148 19256
rect 16396 19216 16436 19256
rect 16492 19216 16532 19256
rect 16972 19216 17012 19256
rect 18220 19216 18260 19256
rect 18604 19216 18644 19256
rect 19852 19216 19892 19256
rect 8428 19132 8468 19172
rect 12268 19132 12308 19172
rect 4684 19048 4724 19088
rect 6796 19048 6836 19088
rect 10444 19006 10484 19046
rect 14284 19048 14324 19088
rect 14764 19048 14804 19088
rect 15244 19048 15284 19088
rect 15532 19048 15572 19088
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 10540 18712 10580 18752
rect 16492 18712 16532 18752
rect 17452 18712 17492 18752
rect 17740 18712 17780 18752
rect 20236 18712 20276 18752
rect 2476 18628 2516 18668
rect 7372 18628 7412 18668
rect 12460 18628 12500 18668
rect 14476 18628 14516 18668
rect 2668 18530 2708 18570
rect 3148 18544 3188 18584
rect 3628 18544 3668 18584
rect 4108 18544 4148 18584
rect 4204 18544 4244 18584
rect 5644 18544 5684 18584
rect 5740 18544 5780 18584
rect 6700 18544 6740 18584
rect 7180 18539 7220 18579
rect 9100 18544 9140 18584
rect 10348 18544 10388 18584
rect 11020 18544 11060 18584
rect 12268 18544 12308 18584
rect 12748 18544 12788 18584
rect 12844 18544 12884 18584
rect 13804 18544 13844 18584
rect 14284 18530 14324 18570
rect 15052 18544 15092 18584
rect 16300 18544 16340 18584
rect 16684 18544 16724 18584
rect 16780 18544 16820 18584
rect 16876 18544 16916 18584
rect 16972 18544 17012 18584
rect 17164 18565 17204 18605
rect 17260 18544 17300 18584
rect 17356 18544 17396 18584
rect 17644 18544 17684 18584
rect 18412 18544 18452 18584
rect 18604 18544 18644 18584
rect 18796 18544 18836 18584
rect 20044 18544 20084 18584
rect 3724 18460 3764 18500
rect 6124 18460 6164 18500
rect 6220 18460 6260 18500
rect 13228 18460 13268 18500
rect 13324 18460 13364 18500
rect 18508 18460 18548 18500
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 2668 17956 2708 17996
rect 5836 17956 5876 17996
rect 14860 17956 14900 17996
rect 16876 17956 16916 17996
rect 17644 17956 17684 17996
rect 1228 17704 1268 17744
rect 2476 17704 2516 17744
rect 4396 17704 4436 17744
rect 5644 17704 5684 17744
rect 7084 17704 7124 17744
rect 8332 17704 8372 17744
rect 8812 17704 8852 17744
rect 8908 17704 8948 17744
rect 9292 17704 9332 17744
rect 9388 17704 9428 17744
rect 9868 17704 9908 17744
rect 10396 17713 10436 17753
rect 13420 17704 13460 17744
rect 14668 17704 14708 17744
rect 15436 17704 15476 17744
rect 16684 17704 16724 17744
rect 17740 17704 17780 17744
rect 17932 17704 17972 17744
rect 19180 17704 19220 17744
rect 19564 17704 19604 17744
rect 19660 17704 19700 17744
rect 19756 17704 19796 17744
rect 20044 17704 20084 17744
rect 20140 17704 20180 17744
rect 8524 17620 8564 17660
rect 19372 17620 19412 17660
rect 10540 17536 10580 17576
rect 19852 17536 19892 17576
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 10636 17200 10676 17240
rect 18796 17200 18836 17240
rect 20236 17200 20276 17240
rect 2188 17116 2228 17156
rect 6988 17116 7028 17156
rect 19468 17116 19508 17156
rect 2380 17018 2420 17058
rect 2860 17032 2900 17072
rect 3340 16990 3380 17030
rect 3436 17032 3476 17072
rect 3820 17032 3860 17072
rect 3916 17032 3956 17072
rect 5260 17032 5300 17072
rect 5356 17032 5396 17072
rect 6316 17032 6356 17072
rect 6796 17018 6836 17058
rect 7372 17032 7412 17072
rect 8620 17032 8660 17072
rect 9196 17032 9236 17072
rect 10444 17032 10484 17072
rect 11308 17032 11348 17072
rect 12556 17032 12596 17072
rect 13324 17032 13364 17072
rect 14572 17032 14612 17072
rect 15724 17032 15764 17072
rect 16972 17032 17012 17072
rect 17356 17032 17396 17072
rect 18604 17032 18644 17072
rect 19084 17032 19124 17072
rect 19372 17032 19412 17072
rect 19948 17032 19988 17072
rect 20044 17032 20084 17072
rect 5740 16948 5780 16988
rect 20140 16990 20180 17030
rect 5836 16948 5876 16988
rect 7180 16780 7220 16820
rect 12748 16780 12788 16820
rect 14764 16780 14804 16820
rect 17164 16780 17204 16820
rect 19756 16780 19796 16820
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 19564 16360 19604 16400
rect 1420 16276 1460 16316
rect 3244 16276 3284 16316
rect 6124 16276 6164 16316
rect 6220 16276 6260 16316
rect 10828 16276 10868 16316
rect 17644 16276 17684 16316
rect 2668 16192 2708 16232
rect 2764 16192 2804 16232
rect 3148 16192 3188 16232
rect 3724 16192 3764 16232
rect 4252 16201 4292 16241
rect 5644 16192 5684 16232
rect 5740 16192 5780 16232
rect 6700 16192 6740 16232
rect 7228 16201 7268 16241
rect 8236 16192 8276 16232
rect 8332 16192 8372 16232
rect 8716 16192 8756 16232
rect 8812 16192 8852 16232
rect 9292 16192 9332 16232
rect 9820 16201 9860 16241
rect 10252 16192 10292 16232
rect 10348 16192 10388 16232
rect 10732 16192 10772 16232
rect 11308 16192 11348 16232
rect 11836 16201 11876 16241
rect 12748 16192 12788 16232
rect 12844 16192 12884 16232
rect 13228 16192 13268 16232
rect 13324 16192 13364 16232
rect 13804 16192 13844 16232
rect 14284 16206 14324 16246
rect 15532 16192 15572 16232
rect 15628 16192 15668 16232
rect 16012 16192 16052 16232
rect 16108 16192 16148 16232
rect 16588 16192 16628 16232
rect 17068 16206 17108 16246
rect 17836 16192 17876 16232
rect 17932 16192 17972 16232
rect 18124 16192 18164 16232
rect 18316 16192 18356 16232
rect 18412 16192 18452 16232
rect 18508 16192 18548 16232
rect 18604 16192 18644 16232
rect 18892 16192 18932 16232
rect 19180 16192 19220 16232
rect 19756 16192 19796 16232
rect 19852 16192 19892 16232
rect 19948 16192 19988 16232
rect 9964 16108 10004 16148
rect 17260 16108 17300 16148
rect 19276 16108 19316 16148
rect 1228 16024 1268 16064
rect 4396 16024 4436 16064
rect 7372 16024 7412 16064
rect 11980 16024 12020 16064
rect 14476 16024 14516 16064
rect 17452 16024 17492 16064
rect 18028 16024 18068 16064
rect 20044 16024 20084 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 2668 15688 2708 15728
rect 5164 15688 5204 15728
rect 6796 15688 6836 15728
rect 8428 15688 8468 15728
rect 10252 15688 10292 15728
rect 12460 15604 12500 15644
rect 14476 15604 14516 15644
rect 16108 15604 16148 15644
rect 19564 15604 19604 15644
rect 1228 15520 1268 15560
rect 2476 15520 2516 15560
rect 3724 15520 3764 15560
rect 4972 15520 5012 15560
rect 5356 15520 5396 15560
rect 6604 15520 6644 15560
rect 8236 15520 8276 15560
rect 8812 15520 8852 15560
rect 10060 15520 10100 15560
rect 11020 15520 11060 15560
rect 12268 15520 12308 15560
rect 12748 15520 12788 15560
rect 6988 15478 7028 15518
rect 12844 15520 12884 15560
rect 13228 15520 13268 15560
rect 13804 15520 13844 15560
rect 14332 15510 14372 15550
rect 14668 15520 14708 15560
rect 15916 15520 15956 15560
rect 16492 15520 16532 15560
rect 17740 15520 17780 15560
rect 18124 15520 18164 15560
rect 19372 15520 19412 15560
rect 19756 15520 19796 15560
rect 19852 15520 19892 15560
rect 20044 15520 20084 15560
rect 3052 15436 3092 15476
rect 13324 15436 13364 15476
rect 2860 15352 2900 15392
rect 20044 15352 20084 15392
rect 16300 15268 16340 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 3436 14932 3476 14972
rect 5644 14932 5684 14972
rect 7468 14932 7508 14972
rect 9868 14932 9908 14972
rect 11980 14932 12020 14972
rect 14572 14932 14612 14972
rect 19180 14932 19220 14972
rect 19660 14932 19700 14972
rect 1708 14764 1748 14804
rect 3820 14764 3860 14804
rect 15628 14764 15668 14804
rect 15724 14764 15764 14804
rect 17260 14764 17300 14804
rect 1996 14680 2036 14720
rect 3244 14680 3284 14720
rect 4204 14680 4244 14720
rect 5452 14680 5492 14720
rect 6028 14680 6068 14720
rect 7276 14680 7316 14720
rect 8428 14680 8468 14720
rect 9676 14680 9716 14720
rect 10540 14680 10580 14720
rect 11788 14680 11828 14720
rect 13132 14680 13172 14720
rect 14380 14680 14420 14720
rect 15148 14680 15188 14720
rect 15244 14680 15284 14720
rect 16204 14680 16244 14720
rect 16684 14694 16724 14734
rect 17548 14680 17588 14720
rect 18796 14680 18836 14720
rect 19180 14680 19220 14720
rect 19372 14680 19412 14720
rect 19468 14680 19508 14720
rect 19756 14680 19796 14720
rect 16876 14596 16916 14636
rect 1516 14512 1556 14552
rect 3628 14512 3668 14552
rect 17068 14512 17108 14552
rect 18988 14512 19028 14552
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 2668 14176 2708 14216
rect 7948 14176 7988 14216
rect 15148 14176 15188 14216
rect 20140 14176 20180 14216
rect 4684 14092 4724 14132
rect 10348 14092 10388 14132
rect 12940 14092 12980 14132
rect 14956 14092 14996 14132
rect 1228 14008 1268 14048
rect 2476 14008 2516 14048
rect 2956 14008 2996 14048
rect 3052 14008 3092 14048
rect 3436 14008 3476 14048
rect 3532 14008 3572 14048
rect 4012 14008 4052 14048
rect 4492 13994 4532 14034
rect 6220 14008 6260 14048
rect 6316 14008 6356 14048
rect 6700 14008 6740 14048
rect 6796 14008 6836 14048
rect 7276 14008 7316 14048
rect 7756 13994 7796 14034
rect 8620 14008 8660 14048
rect 8716 14008 8756 14048
rect 9100 14008 9140 14048
rect 9196 14008 9236 14048
rect 9676 14008 9716 14048
rect 10156 13994 10196 14034
rect 11212 14008 11252 14048
rect 11308 14008 11348 14048
rect 11788 14008 11828 14048
rect 12268 14008 12308 14048
rect 12748 13994 12788 14034
rect 13228 14008 13268 14048
rect 13324 14008 13364 14048
rect 14284 14008 14324 14048
rect 14764 13994 14804 14034
rect 15340 14008 15380 14048
rect 16588 14008 16628 14048
rect 18412 14008 18452 14048
rect 18508 14008 18548 14048
rect 18988 14008 19028 14048
rect 19468 14008 19508 14048
rect 19996 13998 20036 14038
rect 11692 13924 11732 13964
rect 13708 13924 13748 13964
rect 13804 13924 13844 13964
rect 18892 13924 18932 13964
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 1804 13420 1844 13460
rect 4396 13420 4436 13460
rect 8908 13420 8948 13460
rect 10924 13420 10964 13460
rect 12556 13420 12596 13460
rect 14572 13420 14612 13460
rect 20236 13420 20276 13460
rect 1612 13252 1652 13292
rect 1996 13252 2036 13292
rect 2764 13252 2804 13292
rect 4204 13252 4244 13292
rect 5932 13252 5972 13292
rect 16492 13252 16532 13292
rect 16588 13252 16628 13292
rect 18124 13252 18164 13292
rect 2284 13168 2324 13208
rect 2380 13168 2420 13208
rect 2860 13168 2900 13208
rect 3340 13168 3380 13208
rect 3820 13173 3860 13213
rect 5452 13168 5492 13208
rect 5548 13168 5588 13208
rect 6028 13168 6068 13208
rect 6508 13168 6548 13208
rect 7036 13177 7076 13217
rect 7468 13168 7508 13208
rect 8716 13168 8756 13208
rect 9484 13168 9524 13208
rect 10732 13168 10772 13208
rect 11116 13168 11156 13208
rect 12364 13168 12404 13208
rect 13132 13168 13172 13208
rect 14380 13168 14420 13208
rect 16012 13168 16052 13208
rect 16108 13168 16148 13208
rect 17068 13168 17108 13208
rect 17596 13177 17636 13217
rect 18796 13168 18836 13208
rect 20044 13168 20084 13208
rect 7180 13084 7220 13124
rect 17740 13084 17780 13124
rect 1420 13000 1460 13040
rect 4012 13000 4052 13040
rect 17932 13000 17972 13040
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 10252 12664 10292 12704
rect 10444 12664 10484 12704
rect 16012 12664 16052 12704
rect 4204 12580 4244 12620
rect 6124 12580 6164 12620
rect 8236 12580 8276 12620
rect 12940 12580 12980 12620
rect 17740 12580 17780 12620
rect 20044 12580 20084 12620
rect 2764 12496 2804 12536
rect 4012 12496 4052 12536
rect 4684 12496 4724 12536
rect 5932 12496 5972 12536
rect 6796 12496 6836 12536
rect 8044 12496 8084 12536
rect 8812 12496 8852 12536
rect 10060 12496 10100 12536
rect 11500 12496 11540 12536
rect 12748 12496 12788 12536
rect 14572 12496 14612 12536
rect 15820 12496 15860 12536
rect 16300 12496 16340 12536
rect 17548 12496 17588 12536
rect 18316 12496 18356 12536
rect 18412 12496 18452 12536
rect 18796 12496 18836 12536
rect 18892 12496 18932 12536
rect 19372 12496 19412 12536
rect 19900 12454 19940 12494
rect 1708 12412 1748 12452
rect 2092 12412 2132 12452
rect 2476 12412 2516 12452
rect 10636 12412 10676 12452
rect 11308 12412 11348 12452
rect 14188 12412 14228 12452
rect 11116 12328 11156 12368
rect 13996 12328 14036 12368
rect 1516 12244 1556 12284
rect 1900 12244 1940 12284
rect 2284 12244 2324 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 2668 11908 2708 11948
rect 5548 11908 5588 11948
rect 12172 11908 12212 11948
rect 18700 11908 18740 11948
rect 3244 11824 3284 11864
rect 3052 11740 3092 11780
rect 3436 11740 3476 11780
rect 3820 11740 3860 11780
rect 6412 11740 6452 11780
rect 9004 11740 9044 11780
rect 9100 11740 9140 11780
rect 12364 11740 12404 11780
rect 15052 11740 15092 11780
rect 1228 11656 1268 11696
rect 2476 11656 2516 11696
rect 4108 11656 4148 11696
rect 5356 11656 5396 11696
rect 5836 11656 5876 11696
rect 5932 11656 5972 11696
rect 6316 11656 6356 11696
rect 6892 11656 6932 11696
rect 7372 11661 7412 11701
rect 8524 11656 8564 11696
rect 8620 11656 8660 11696
rect 9580 11656 9620 11696
rect 10060 11661 10100 11701
rect 10540 11656 10580 11696
rect 11788 11656 11828 11696
rect 12652 11656 12692 11696
rect 13900 11656 13940 11696
rect 14572 11656 14612 11696
rect 14668 11656 14708 11696
rect 15148 11656 15188 11696
rect 15628 11656 15668 11696
rect 16108 11661 16148 11701
rect 17260 11656 17300 11696
rect 18508 11656 18548 11696
rect 7564 11572 7604 11612
rect 10252 11572 10292 11612
rect 16300 11572 16340 11612
rect 2860 11488 2900 11528
rect 3628 11488 3668 11528
rect 11980 11488 12020 11528
rect 14092 11488 14132 11528
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 1900 11152 1940 11192
rect 9964 11152 10004 11192
rect 11980 11152 12020 11192
rect 14284 11152 14324 11192
rect 20140 11152 20180 11192
rect 4300 11068 4340 11108
rect 7180 11068 7220 11108
rect 17452 11068 17492 11108
rect 2572 10984 2612 11024
rect 2668 10984 2708 11024
rect 3628 10984 3668 11024
rect 4108 10970 4148 11010
rect 5452 10984 5492 11024
rect 5548 10984 5588 11024
rect 5932 10984 5972 11024
rect 6028 10984 6068 11024
rect 6508 10984 6548 11024
rect 6988 10970 7028 11010
rect 8524 10984 8564 11024
rect 9772 10984 9812 11024
rect 10252 10984 10292 11024
rect 10348 10984 10388 11024
rect 10732 10984 10772 11024
rect 11308 10984 11348 11024
rect 11836 10974 11876 11014
rect 12556 10984 12596 11024
rect 12652 10984 12692 11024
rect 13132 10984 13172 11024
rect 13612 10984 13652 11024
rect 14092 10979 14132 11019
rect 15724 10984 15764 11024
rect 15820 10984 15860 11024
rect 16300 10984 16340 11024
rect 16780 10984 16820 11024
rect 17260 10970 17300 11010
rect 18700 10984 18740 11024
rect 19948 10984 19988 11024
rect 1708 10900 1748 10940
rect 2092 10900 2132 10940
rect 3052 10900 3092 10940
rect 3148 10900 3188 10940
rect 4684 10900 4724 10940
rect 4876 10900 4916 10940
rect 10828 10900 10868 10940
rect 13036 10900 13076 10940
rect 14668 10900 14708 10940
rect 16204 10900 16244 10940
rect 14476 10816 14516 10856
rect 1516 10732 1556 10772
rect 4492 10732 4532 10772
rect 5068 10732 5108 10772
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 2668 10396 2708 10436
rect 4972 10396 5012 10436
rect 5164 10396 5204 10436
rect 7084 10396 7124 10436
rect 10156 10396 10196 10436
rect 12748 10396 12788 10436
rect 14476 10396 14516 10436
rect 16204 10396 16244 10436
rect 17836 10396 17876 10436
rect 2860 10312 2900 10352
rect 3052 10228 3092 10268
rect 5356 10228 5396 10268
rect 7468 10228 7508 10268
rect 18700 10228 18740 10268
rect 18796 10228 18836 10268
rect 1228 10144 1268 10184
rect 2476 10144 2516 10184
rect 4780 10144 4820 10184
rect 5644 10144 5684 10184
rect 6892 10144 6932 10184
rect 8716 10144 8756 10184
rect 9964 10144 10004 10184
rect 11308 10144 11348 10184
rect 12556 10144 12596 10184
rect 13036 10144 13076 10184
rect 14284 10144 14324 10184
rect 14764 10144 14804 10184
rect 16012 10144 16052 10184
rect 16396 10144 16436 10184
rect 17644 10144 17684 10184
rect 18220 10144 18260 10184
rect 3532 10102 3572 10142
rect 18316 10144 18356 10184
rect 19276 10144 19316 10184
rect 19804 10153 19844 10193
rect 19948 10060 19988 10100
rect 7276 9976 7316 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 1420 9640 1460 9680
rect 2188 9640 2228 9680
rect 4396 9640 4436 9680
rect 7084 9640 7124 9680
rect 8716 9640 8756 9680
rect 13516 9640 13556 9680
rect 15820 9640 15860 9680
rect 17932 9640 17972 9680
rect 19948 9682 19988 9722
rect 11692 9556 11732 9596
rect 11884 9556 11924 9596
rect 2668 9472 2708 9512
rect 2764 9472 2804 9512
rect 3148 9472 3188 9512
rect 3244 9472 3284 9512
rect 3724 9472 3764 9512
rect 4204 9467 4244 9507
rect 5644 9472 5684 9512
rect 6892 9472 6932 9512
rect 7276 9472 7316 9512
rect 8524 9472 8564 9512
rect 9964 9472 10004 9512
rect 10060 9472 10100 9512
rect 10540 9472 10580 9512
rect 11020 9472 11060 9512
rect 11500 9467 11540 9507
rect 12076 9472 12116 9512
rect 13324 9472 13364 9512
rect 14380 9472 14420 9512
rect 15628 9472 15668 9512
rect 16492 9472 16532 9512
rect 17740 9472 17780 9512
rect 18220 9472 18260 9512
rect 18316 9472 18356 9512
rect 18700 9472 18740 9512
rect 18796 9472 18836 9512
rect 19276 9472 19316 9512
rect 1612 9388 1652 9428
rect 1996 9388 2036 9428
rect 2380 9388 2420 9428
rect 4780 9388 4820 9428
rect 5164 9388 5204 9428
rect 19804 9430 19844 9470
rect 10444 9388 10484 9428
rect 13708 9388 13748 9428
rect 1804 9220 1844 9260
rect 4588 9220 4628 9260
rect 4972 9220 5012 9260
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18316 8884 18356 8924
rect 20140 8884 20180 8924
rect 2668 8800 2708 8840
rect 4300 8800 4340 8840
rect 4684 8716 4724 8756
rect 5644 8716 5684 8756
rect 5740 8716 5780 8756
rect 7852 8716 7892 8756
rect 7948 8716 7988 8756
rect 16108 8716 16148 8756
rect 1228 8632 1268 8672
rect 2476 8632 2516 8672
rect 2860 8632 2900 8672
rect 4108 8632 4148 8672
rect 5164 8632 5204 8672
rect 5260 8632 5300 8672
rect 6220 8632 6260 8672
rect 6700 8637 6740 8677
rect 7372 8632 7412 8672
rect 7468 8632 7508 8672
rect 8428 8632 8468 8672
rect 8956 8641 8996 8681
rect 10636 8632 10676 8672
rect 11884 8632 11924 8672
rect 12364 8632 12404 8672
rect 12460 8632 12500 8672
rect 12844 8632 12884 8672
rect 12940 8632 12980 8672
rect 13420 8632 13460 8672
rect 13900 8637 13940 8677
rect 15052 8637 15092 8677
rect 15532 8632 15572 8672
rect 16012 8632 16052 8672
rect 16492 8632 16532 8672
rect 16588 8632 16628 8672
rect 16876 8632 16916 8672
rect 18124 8632 18164 8672
rect 18700 8632 18740 8672
rect 19948 8632 19988 8672
rect 12076 8548 12116 8588
rect 14092 8548 14132 8588
rect 4876 8464 4916 8504
rect 6892 8464 6932 8504
rect 9100 8464 9140 8504
rect 14860 8464 14900 8504
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 2668 8128 2708 8168
rect 2860 8128 2900 8168
rect 3244 8128 3284 8168
rect 5644 8128 5684 8168
rect 7276 8128 7316 8168
rect 9676 8128 9716 8168
rect 9868 8128 9908 8168
rect 13900 8128 13940 8168
rect 15532 8128 15572 8168
rect 15724 8128 15764 8168
rect 19660 8128 19700 8168
rect 1228 7960 1268 8000
rect 2476 7960 2516 8000
rect 4204 7960 4244 8000
rect 5452 7960 5492 8000
rect 5836 7960 5876 8000
rect 7084 7960 7124 8000
rect 8236 7960 8276 8000
rect 9484 7960 9524 8000
rect 10060 7955 10100 7995
rect 10540 7960 10580 8000
rect 11020 7960 11060 8000
rect 11500 7960 11540 8000
rect 11596 7960 11636 8000
rect 12460 7960 12500 8000
rect 13708 7960 13748 8000
rect 14092 7960 14132 8000
rect 15340 7960 15380 8000
rect 15916 7960 15956 8000
rect 17164 7960 17204 8000
rect 17932 7960 17972 8000
rect 18028 7960 18068 8000
rect 18412 7960 18452 8000
rect 18508 7960 18548 8000
rect 18988 7960 19028 8000
rect 19468 7946 19508 7986
rect 3052 7876 3092 7916
rect 3436 7876 3476 7916
rect 3820 7876 3860 7916
rect 7660 7876 7700 7916
rect 8044 7876 8084 7916
rect 11116 7876 11156 7916
rect 4012 7792 4052 7832
rect 7468 7708 7508 7748
rect 7852 7708 7892 7748
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 2956 7372 2996 7412
rect 9580 7372 9620 7412
rect 11692 7372 11732 7412
rect 20044 7372 20084 7412
rect 18028 7288 18068 7328
rect 3724 7204 3764 7244
rect 3820 7204 3860 7244
rect 8812 7204 8852 7244
rect 9388 7204 9428 7244
rect 9772 7204 9812 7244
rect 15052 7204 15092 7244
rect 1516 7120 1556 7160
rect 2764 7120 2804 7160
rect 3244 7120 3284 7160
rect 3340 7120 3380 7160
rect 4300 7120 4340 7160
rect 4780 7125 4820 7165
rect 5164 7120 5204 7160
rect 6412 7120 6452 7160
rect 6988 7125 7028 7165
rect 7468 7120 7508 7160
rect 7948 7120 7988 7160
rect 8044 7120 8084 7160
rect 8428 7120 8468 7160
rect 8524 7120 8564 7160
rect 10252 7120 10292 7160
rect 11500 7120 11540 7160
rect 12844 7120 12884 7160
rect 14092 7120 14132 7160
rect 14572 7120 14612 7160
rect 14668 7120 14708 7160
rect 15148 7120 15188 7160
rect 15628 7120 15668 7160
rect 16156 7129 16196 7169
rect 16588 7120 16628 7160
rect 17836 7120 17876 7160
rect 18604 7120 18644 7160
rect 19852 7120 19892 7160
rect 4972 7036 5012 7076
rect 14284 7036 14324 7076
rect 6604 6952 6644 6992
rect 6796 6952 6836 6992
rect 9004 6952 9044 6992
rect 9196 6952 9236 6992
rect 16300 6952 16340 6992
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 2668 6616 2708 6656
rect 7468 6616 7508 6656
rect 9100 6616 9140 6656
rect 10732 6616 10772 6656
rect 13804 6616 13844 6656
rect 16300 6616 16340 6656
rect 19948 6616 19988 6656
rect 4780 6532 4820 6572
rect 1228 6448 1268 6488
rect 2476 6448 2516 6488
rect 3052 6448 3092 6488
rect 3148 6448 3188 6488
rect 3532 6448 3572 6488
rect 3628 6448 3668 6488
rect 4108 6448 4148 6488
rect 4588 6434 4628 6474
rect 6028 6448 6068 6488
rect 7276 6448 7316 6488
rect 7660 6448 7700 6488
rect 8908 6448 8948 6488
rect 9292 6448 9332 6488
rect 10540 6448 10580 6488
rect 12076 6448 12116 6488
rect 12172 6448 12212 6488
rect 12556 6448 12596 6488
rect 12652 6448 12692 6488
rect 13132 6448 13172 6488
rect 13612 6434 13652 6474
rect 14860 6448 14900 6488
rect 16108 6448 16148 6488
rect 16492 6448 16532 6488
rect 17740 6448 17780 6488
rect 18508 6448 18548 6488
rect 19756 6448 19796 6488
rect 5164 6364 5204 6404
rect 5356 6364 5396 6404
rect 11116 6364 11156 6404
rect 4972 6280 5012 6320
rect 5548 6280 5588 6320
rect 10924 6280 10964 6320
rect 17932 6196 17972 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 1516 5860 1556 5900
rect 1900 5860 1940 5900
rect 3820 5860 3860 5900
rect 4396 5860 4436 5900
rect 6508 5860 6548 5900
rect 11596 5860 11636 5900
rect 13708 5860 13748 5900
rect 4204 5776 4244 5816
rect 9292 5776 9332 5816
rect 1708 5692 1748 5732
rect 2092 5692 2132 5732
rect 4012 5692 4052 5732
rect 4588 5692 4628 5732
rect 4876 5692 4916 5732
rect 7276 5692 7316 5732
rect 7372 5692 7412 5732
rect 8908 5692 8948 5732
rect 10252 5692 10292 5732
rect 11788 5703 11828 5743
rect 14476 5692 14516 5732
rect 14572 5692 14612 5732
rect 17260 5692 17300 5732
rect 17356 5692 17396 5732
rect 2380 5608 2420 5648
rect 3628 5608 3668 5648
rect 5068 5608 5108 5648
rect 6316 5608 6356 5648
rect 6796 5608 6836 5648
rect 6892 5608 6932 5648
rect 7852 5608 7892 5648
rect 8332 5613 8372 5653
rect 9676 5608 9716 5648
rect 9772 5608 9812 5648
rect 10156 5608 10196 5648
rect 10732 5608 10772 5648
rect 11212 5613 11252 5653
rect 12268 5608 12308 5648
rect 13516 5608 13556 5648
rect 13996 5608 14036 5648
rect 14092 5608 14132 5648
rect 15052 5608 15092 5648
rect 15580 5617 15620 5657
rect 16780 5608 16820 5648
rect 16876 5608 16916 5648
rect 17836 5608 17876 5648
rect 18316 5622 18356 5662
rect 18700 5608 18740 5648
rect 19948 5608 19988 5648
rect 8524 5524 8564 5564
rect 11404 5524 11444 5564
rect 18508 5524 18548 5564
rect 9100 5440 9140 5480
rect 11980 5440 12020 5480
rect 15724 5440 15764 5480
rect 20140 5440 20180 5480
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 4780 5104 4820 5144
rect 7180 5104 7220 5144
rect 9004 5104 9044 5144
rect 13996 5104 14036 5144
rect 15724 5104 15764 5144
rect 17356 5104 17396 5144
rect 2668 5020 2708 5060
rect 4300 5020 4340 5060
rect 12268 5020 12308 5060
rect 18316 5020 18356 5060
rect 1228 4936 1268 4976
rect 2476 4936 2516 4976
rect 2860 4936 2900 4976
rect 4108 4936 4148 4976
rect 5452 4936 5492 4976
rect 4924 4894 4964 4934
rect 6412 4917 6452 4957
rect 6508 4936 6548 4976
rect 7564 4936 7604 4976
rect 8812 4936 8852 4976
rect 9196 4936 9236 4976
rect 10444 4936 10484 4976
rect 10828 4936 10868 4976
rect 12076 4936 12116 4976
rect 12556 4936 12596 4976
rect 13804 4936 13844 4976
rect 14284 4936 14324 4976
rect 15532 4936 15572 4976
rect 15916 4936 15956 4976
rect 17164 4936 17204 4976
rect 18508 4922 18548 4962
rect 18988 4936 19028 4976
rect 19468 4936 19508 4976
rect 19564 4936 19604 4976
rect 19948 4936 19988 4976
rect 20044 4936 20084 4976
rect 5932 4852 5972 4892
rect 6028 4852 6068 4892
rect 6988 4852 7028 4892
rect 7372 4852 7412 4892
rect 4588 4768 4628 4808
rect 6796 4768 6836 4808
rect 10636 4684 10676 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 2668 4348 2708 4388
rect 4588 4348 4628 4388
rect 6796 4348 6836 4388
rect 2860 4264 2900 4304
rect 4972 4180 5012 4220
rect 9772 4180 9812 4220
rect 9868 4180 9908 4220
rect 10828 4180 10868 4220
rect 11212 4180 11252 4220
rect 11596 4180 11636 4220
rect 18316 4180 18356 4220
rect 18412 4180 18452 4220
rect 1228 4096 1268 4136
rect 2476 4096 2516 4136
rect 3148 4096 3188 4136
rect 4396 4096 4436 4136
rect 5356 4096 5396 4136
rect 6604 4096 6644 4136
rect 6988 4096 7028 4136
rect 8236 4096 8276 4136
rect 8764 4105 8804 4145
rect 9292 4096 9332 4136
rect 10252 4096 10292 4136
rect 10348 4076 10388 4116
rect 11884 4096 11924 4136
rect 13132 4096 13172 4136
rect 13708 4096 13748 4136
rect 14956 4096 14996 4136
rect 15340 4096 15380 4136
rect 16588 4096 16628 4136
rect 17836 4096 17876 4136
rect 17932 4096 17972 4136
rect 18892 4096 18932 4136
rect 19420 4105 19460 4145
rect 8428 4012 8468 4052
rect 5164 3928 5204 3968
rect 8620 3928 8660 3968
rect 10636 3928 10676 3968
rect 11020 3928 11060 3968
rect 11404 3928 11444 3968
rect 13324 3928 13364 3968
rect 15148 3928 15188 3968
rect 16780 3928 16820 3968
rect 19564 3928 19604 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 1516 3592 1556 3632
rect 2092 3592 2132 3632
rect 3724 3592 3764 3632
rect 5836 3592 5876 3632
rect 10348 3592 10388 3632
rect 13516 3592 13556 3632
rect 16204 3592 16244 3632
rect 19660 3592 19700 3632
rect 1324 3508 1364 3548
rect 2284 3424 2324 3464
rect 3532 3424 3572 3464
rect 4108 3424 4148 3464
rect 4204 3424 4244 3464
rect 5164 3424 5204 3464
rect 5644 3410 5684 3450
rect 6220 3424 6260 3464
rect 7468 3424 7508 3464
rect 8620 3424 8660 3464
rect 8716 3424 8756 3464
rect 9100 3424 9140 3464
rect 9676 3424 9716 3464
rect 1708 3340 1748 3380
rect 1900 3340 1940 3380
rect 4588 3340 4628 3380
rect 4684 3340 4724 3380
rect 7756 3340 7796 3380
rect 8140 3340 8180 3380
rect 9196 3340 9236 3380
rect 10204 3382 10244 3422
rect 11788 3424 11828 3464
rect 11884 3424 11924 3464
rect 12364 3424 12404 3464
rect 12844 3424 12884 3464
rect 13324 3419 13364 3459
rect 14476 3424 14516 3464
rect 14572 3424 14612 3464
rect 14956 3424 14996 3464
rect 15052 3424 15092 3464
rect 15532 3424 15572 3464
rect 10540 3340 10580 3380
rect 10924 3340 10964 3380
rect 11500 3340 11540 3380
rect 16060 3382 16100 3422
rect 17932 3424 17972 3464
rect 18028 3424 18068 3464
rect 18508 3424 18548 3464
rect 18988 3424 19028 3464
rect 12268 3340 12308 3380
rect 13708 3340 13748 3380
rect 16588 3340 16628 3380
rect 16972 3340 17012 3380
rect 17356 3340 17396 3380
rect 18412 3340 18452 3380
rect 19516 3382 19556 3422
rect 6028 3172 6068 3212
rect 7948 3172 7988 3212
rect 8332 3172 8372 3212
rect 10732 3172 10772 3212
rect 11116 3172 11156 3212
rect 11308 3172 11348 3212
rect 13900 3172 13940 3212
rect 16396 3172 16436 3212
rect 16780 3172 16820 3212
rect 17164 3172 17204 3212
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 3436 2836 3476 2876
rect 5068 2836 5108 2876
rect 6700 2836 6740 2876
rect 9484 2836 9524 2876
rect 11500 2836 11540 2876
rect 18508 2836 18548 2876
rect 20236 2836 20276 2876
rect 2860 2752 2900 2792
rect 9100 2752 9140 2792
rect 9868 2752 9908 2792
rect 13708 2752 13748 2792
rect 3244 2668 3284 2708
rect 7564 2668 7604 2708
rect 3628 2626 3668 2666
rect 8908 2668 8948 2708
rect 9292 2668 9332 2708
rect 9676 2668 9716 2708
rect 12268 2668 12308 2708
rect 12364 2668 12404 2708
rect 14188 2668 14228 2708
rect 14572 2668 14612 2708
rect 15628 2668 15668 2708
rect 15724 2668 15764 2708
rect 1420 2584 1460 2624
rect 2668 2584 2708 2624
rect 4876 2584 4916 2624
rect 5260 2584 5300 2624
rect 6508 2584 6548 2624
rect 6988 2584 7028 2624
rect 7084 2584 7124 2624
rect 7468 2584 7508 2624
rect 8044 2584 8084 2624
rect 8524 2598 8564 2638
rect 10060 2584 10100 2624
rect 11308 2584 11348 2624
rect 11788 2584 11828 2624
rect 11884 2584 11924 2624
rect 12844 2584 12884 2624
rect 13324 2589 13364 2629
rect 15148 2584 15188 2624
rect 15244 2584 15284 2624
rect 16204 2584 16244 2624
rect 16684 2598 16724 2638
rect 17068 2584 17108 2624
rect 18316 2584 18356 2624
rect 18796 2584 18836 2624
rect 20044 2584 20084 2624
rect 8716 2500 8756 2540
rect 13516 2500 13556 2540
rect 16876 2500 16916 2540
rect 13996 2416 14036 2456
rect 14380 2416 14420 2456
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 2668 2080 2708 2120
rect 2860 2080 2900 2120
rect 5068 2080 5108 2120
rect 6700 2080 6740 2120
rect 6988 2080 7028 2120
rect 8620 2080 8660 2120
rect 11308 2080 11348 2120
rect 12940 2080 12980 2120
rect 14572 2080 14612 2120
rect 16204 2080 16244 2120
rect 17932 2080 17972 2120
rect 19852 2080 19892 2120
rect 8812 1996 8852 2036
rect 1228 1912 1268 1952
rect 2476 1912 2516 1952
rect 3340 1912 3380 1952
rect 3436 1912 3476 1952
rect 3916 1912 3956 1952
rect 4396 1912 4436 1952
rect 4876 1898 4916 1938
rect 5260 1912 5300 1952
rect 6508 1912 6548 1952
rect 7180 1912 7220 1952
rect 8428 1912 8468 1952
rect 9868 1912 9908 1952
rect 11116 1912 11156 1952
rect 11500 1912 11540 1952
rect 12748 1912 12788 1952
rect 13132 1912 13172 1952
rect 14380 1912 14420 1952
rect 14764 1912 14804 1952
rect 16012 1912 16052 1952
rect 16492 1912 16532 1952
rect 17740 1912 17780 1952
rect 18412 1912 18452 1952
rect 19660 1912 19700 1952
rect 3052 1828 3092 1868
rect 3820 1828 3860 1868
rect 9100 1828 9140 1868
rect 9484 1828 9524 1868
rect 20236 1828 20276 1868
rect 9292 1660 9332 1700
rect 9676 1660 9716 1700
rect 20044 1660 20084 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 2764 1240 2804 1280
rect 4972 1240 5012 1280
rect 6700 1240 6740 1280
rect 6988 1240 7028 1280
rect 8620 1240 8660 1280
rect 10252 1240 10292 1280
rect 12076 1240 12116 1280
rect 13708 1240 13748 1280
rect 15340 1240 15380 1280
rect 19852 1240 19892 1280
rect 3148 1156 3188 1196
rect 17164 1156 17204 1196
rect 17548 1156 17588 1196
rect 18220 1156 18260 1196
rect 1324 1072 1364 1112
rect 2572 1072 2612 1112
rect 3532 1072 3572 1112
rect 4780 1072 4820 1112
rect 5260 1072 5300 1112
rect 6508 1072 6548 1112
rect 7180 1072 7220 1112
rect 8428 1072 8468 1112
rect 8812 1072 8852 1112
rect 10060 1072 10100 1112
rect 10636 1072 10676 1112
rect 11884 1072 11924 1112
rect 12268 1072 12308 1112
rect 13516 1072 13556 1112
rect 13900 1072 13940 1112
rect 15148 1072 15188 1112
rect 15532 1072 15572 1112
rect 16780 1072 16820 1112
rect 18412 1072 18452 1112
rect 19660 1072 19700 1112
rect 2956 904 2996 944
rect 10444 904 10484 944
rect 16972 904 17012 944
rect 17356 904 17396 944
rect 18028 904 18068 944
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
<< metal2 >>
rect 1784 85936 1864 86016
rect 1976 85936 2056 86016
rect 2168 85936 2248 86016
rect 2360 85936 2440 86016
rect 2552 85936 2632 86016
rect 2744 85936 2824 86016
rect 2936 85936 3016 86016
rect 3128 85936 3208 86016
rect 3320 85936 3400 86016
rect 3512 85936 3592 86016
rect 3704 85936 3784 86016
rect 3896 85936 3976 86016
rect 4088 85936 4168 86016
rect 4280 85936 4360 86016
rect 4472 85936 4552 86016
rect 4664 85936 4744 86016
rect 4856 85936 4936 86016
rect 5048 85936 5128 86016
rect 5240 85936 5320 86016
rect 5432 85936 5512 86016
rect 5624 85936 5704 86016
rect 5816 85936 5896 86016
rect 6008 85936 6088 86016
rect 6200 85936 6280 86016
rect 6392 85936 6472 86016
rect 6584 85936 6664 86016
rect 6776 85936 6856 86016
rect 6968 85936 7048 86016
rect 7160 85936 7240 86016
rect 7352 85936 7432 86016
rect 7544 85936 7624 86016
rect 7736 85936 7816 86016
rect 7928 85936 8008 86016
rect 8120 85936 8200 86016
rect 8312 85936 8392 86016
rect 8504 85936 8584 86016
rect 8696 85936 8776 86016
rect 8888 85936 8968 86016
rect 9080 85936 9160 86016
rect 9272 85936 9352 86016
rect 9464 85936 9544 86016
rect 9656 85936 9736 86016
rect 9848 85936 9928 86016
rect 10040 85936 10120 86016
rect 10232 85936 10312 86016
rect 10424 85936 10504 86016
rect 10616 85936 10696 86016
rect 10808 85936 10888 86016
rect 11000 85936 11080 86016
rect 11192 85936 11272 86016
rect 11384 85936 11464 86016
rect 11576 85936 11656 86016
rect 11768 85936 11848 86016
rect 11960 85936 12040 86016
rect 12152 85936 12232 86016
rect 12344 85936 12424 86016
rect 12536 85936 12616 86016
rect 12728 85936 12808 86016
rect 12920 85936 13000 86016
rect 13112 85936 13192 86016
rect 13304 85936 13384 86016
rect 13496 85936 13576 86016
rect 13688 85936 13768 86016
rect 13880 85936 13960 86016
rect 14072 85936 14152 86016
rect 14264 85936 14344 86016
rect 14456 85936 14536 86016
rect 14648 85936 14728 86016
rect 14840 85936 14920 86016
rect 15032 85936 15112 86016
rect 15224 85936 15304 86016
rect 15416 85936 15496 86016
rect 15608 85936 15688 86016
rect 15800 85936 15880 86016
rect 15992 85936 16072 86016
rect 16184 85936 16264 86016
rect 16376 85936 16456 86016
rect 16568 85936 16648 86016
rect 16760 85936 16840 86016
rect 16952 85936 17032 86016
rect 17144 85936 17224 86016
rect 17336 85936 17416 86016
rect 17528 85936 17608 86016
rect 17720 85936 17800 86016
rect 17912 85936 17992 86016
rect 18104 85936 18184 86016
rect 18296 85936 18376 86016
rect 18488 85936 18568 86016
rect 18680 85936 18760 86016
rect 18872 85936 18952 86016
rect 19064 85936 19144 86016
rect 19256 85936 19336 86016
rect 19448 85936 19528 86016
rect 1515 84608 1557 84617
rect 1515 84568 1516 84608
rect 1556 84568 1557 84608
rect 1515 84559 1557 84568
rect 1516 84440 1556 84559
rect 1516 84391 1556 84400
rect 1323 84356 1365 84365
rect 1323 84316 1324 84356
rect 1364 84316 1365 84356
rect 1323 84307 1365 84316
rect 1707 84356 1749 84365
rect 1707 84316 1708 84356
rect 1748 84316 1749 84356
rect 1707 84307 1749 84316
rect 1324 84222 1364 84307
rect 1708 84222 1748 84307
rect 1515 83852 1557 83861
rect 1515 83812 1516 83852
rect 1556 83812 1557 83852
rect 1515 83803 1557 83812
rect 1516 83768 1556 83803
rect 1516 83717 1556 83728
rect 1708 83600 1748 83609
rect 1323 83516 1365 83525
rect 1323 83476 1324 83516
rect 1364 83476 1365 83516
rect 1323 83467 1365 83476
rect 1324 83382 1364 83467
rect 1324 82760 1364 82769
rect 1324 82265 1364 82720
rect 1323 82256 1365 82265
rect 1323 82216 1324 82256
rect 1364 82216 1365 82256
rect 1323 82207 1365 82216
rect 1228 82088 1268 82097
rect 1268 82048 1556 82088
rect 1228 82039 1268 82048
rect 1516 81509 1556 82048
rect 1708 81920 1748 83560
rect 1804 81929 1844 85936
rect 1899 84944 1941 84953
rect 1899 84904 1900 84944
rect 1940 84904 1941 84944
rect 1899 84895 1941 84904
rect 1900 84440 1940 84895
rect 1900 84391 1940 84400
rect 1612 81880 1748 81920
rect 1803 81920 1845 81929
rect 1803 81880 1804 81920
rect 1844 81880 1845 81920
rect 1515 81500 1557 81509
rect 1515 81460 1516 81500
rect 1556 81460 1557 81500
rect 1515 81451 1557 81460
rect 1228 81248 1268 81257
rect 1268 81208 1556 81248
rect 1228 81199 1268 81208
rect 1323 80576 1365 80585
rect 1323 80536 1324 80576
rect 1364 80536 1365 80576
rect 1323 80527 1365 80536
rect 1420 80576 1460 80585
rect 1324 80442 1364 80527
rect 1035 79988 1077 79997
rect 1420 79988 1460 80536
rect 1035 79948 1036 79988
rect 1076 79948 1077 79988
rect 1035 79939 1077 79948
rect 1324 79948 1460 79988
rect 747 79400 789 79409
rect 747 79360 748 79400
rect 788 79360 789 79400
rect 747 79351 789 79360
rect 171 75620 213 75629
rect 171 75580 172 75620
rect 212 75580 213 75620
rect 171 75571 213 75580
rect 75 67808 117 67817
rect 75 67768 76 67808
rect 116 67768 117 67808
rect 75 67759 117 67768
rect 76 67313 116 67759
rect 75 67304 117 67313
rect 75 67264 76 67304
rect 116 67264 117 67304
rect 75 67255 117 67264
rect 75 66296 117 66305
rect 75 66256 76 66296
rect 116 66256 117 66296
rect 75 66247 117 66256
rect 76 55460 116 66247
rect 172 61937 212 75571
rect 459 74948 501 74957
rect 459 74908 460 74948
rect 500 74908 501 74948
rect 459 74899 501 74908
rect 267 71924 309 71933
rect 267 71884 268 71924
rect 308 71884 309 71924
rect 267 71875 309 71884
rect 171 61928 213 61937
rect 171 61888 172 61928
rect 212 61888 213 61928
rect 171 61879 213 61888
rect 268 60593 308 71875
rect 363 69740 405 69749
rect 363 69700 364 69740
rect 404 69700 405 69740
rect 363 69691 405 69700
rect 267 60584 309 60593
rect 267 60544 268 60584
rect 308 60544 309 60584
rect 267 60535 309 60544
rect 364 60257 404 69691
rect 460 64289 500 74899
rect 748 73781 788 79351
rect 747 73772 789 73781
rect 747 73732 748 73772
rect 788 73732 789 73772
rect 747 73723 789 73732
rect 1036 73697 1076 79939
rect 1227 79064 1269 79073
rect 1227 79024 1228 79064
rect 1268 79024 1269 79064
rect 1227 79015 1269 79024
rect 1228 78930 1268 79015
rect 1131 78728 1173 78737
rect 1131 78688 1132 78728
rect 1172 78688 1173 78728
rect 1131 78679 1173 78688
rect 1132 74873 1172 78679
rect 1324 78308 1364 79948
rect 1516 79913 1556 81208
rect 1612 80333 1652 81880
rect 1803 81871 1845 81880
rect 1804 80492 1844 80501
rect 1708 80452 1804 80492
rect 1611 80324 1653 80333
rect 1611 80284 1612 80324
rect 1652 80284 1653 80324
rect 1611 80275 1653 80284
rect 1515 79904 1557 79913
rect 1515 79864 1516 79904
rect 1556 79864 1557 79904
rect 1515 79855 1557 79864
rect 1419 79820 1461 79829
rect 1415 79780 1420 79820
rect 1460 79780 1461 79820
rect 1415 79771 1461 79780
rect 1415 79736 1455 79771
rect 1415 79687 1455 79696
rect 1516 79736 1556 79747
rect 1516 79661 1556 79696
rect 1611 79736 1653 79745
rect 1611 79696 1612 79736
rect 1652 79696 1653 79736
rect 1611 79687 1653 79696
rect 1515 79652 1557 79661
rect 1515 79612 1516 79652
rect 1556 79612 1557 79652
rect 1515 79603 1557 79612
rect 1612 79602 1652 79687
rect 1419 79568 1461 79577
rect 1419 79528 1420 79568
rect 1460 79528 1461 79568
rect 1419 79519 1461 79528
rect 1420 79434 1460 79519
rect 1324 78268 1652 78308
rect 1228 78224 1268 78233
rect 1228 77561 1268 78184
rect 1419 78140 1461 78149
rect 1419 78100 1420 78140
rect 1460 78100 1461 78140
rect 1419 78091 1461 78100
rect 1227 77552 1269 77561
rect 1227 77512 1228 77552
rect 1268 77512 1269 77552
rect 1227 77503 1269 77512
rect 1228 77418 1268 77503
rect 1324 76796 1364 76805
rect 1227 75956 1269 75965
rect 1227 75916 1228 75956
rect 1268 75916 1269 75956
rect 1227 75907 1269 75916
rect 1228 75822 1268 75907
rect 1131 74864 1173 74873
rect 1131 74824 1132 74864
rect 1172 74824 1173 74864
rect 1131 74815 1173 74824
rect 1035 73688 1077 73697
rect 1035 73648 1036 73688
rect 1076 73648 1077 73688
rect 1035 73639 1077 73648
rect 1227 73184 1269 73193
rect 1227 73144 1228 73184
rect 1268 73144 1269 73184
rect 1227 73135 1269 73144
rect 1228 73016 1268 73135
rect 1228 72967 1268 72976
rect 1324 71849 1364 76756
rect 1420 76376 1460 78091
rect 1515 76796 1557 76805
rect 1515 76756 1516 76796
rect 1556 76756 1557 76796
rect 1515 76747 1557 76756
rect 1516 76544 1556 76747
rect 1612 76544 1652 78268
rect 1708 76964 1748 80452
rect 1804 80443 1844 80452
rect 1900 80492 1940 80501
rect 1900 79997 1940 80452
rect 1996 80165 2036 85936
rect 2091 85784 2133 85793
rect 2091 85744 2092 85784
rect 2132 85744 2133 85784
rect 2091 85735 2133 85744
rect 2092 84272 2132 85735
rect 2092 84029 2132 84232
rect 2091 84020 2133 84029
rect 2091 83980 2092 84020
rect 2132 83980 2133 84020
rect 2091 83971 2133 83980
rect 2091 81500 2133 81509
rect 2091 81460 2092 81500
rect 2132 81460 2133 81500
rect 2091 81451 2133 81460
rect 1995 80156 2037 80165
rect 1995 80116 1996 80156
rect 2036 80116 2037 80156
rect 1995 80107 2037 80116
rect 1899 79988 1941 79997
rect 1899 79948 1900 79988
rect 1940 79948 1941 79988
rect 1899 79939 1941 79948
rect 2092 79913 2132 81451
rect 1803 79904 1845 79913
rect 1803 79864 1804 79904
rect 1844 79864 1845 79904
rect 1803 79855 1845 79864
rect 2091 79904 2133 79913
rect 2091 79864 2092 79904
rect 2132 79864 2133 79904
rect 2091 79855 2133 79864
rect 1804 79736 1844 79855
rect 1804 77225 1844 79696
rect 1900 79736 1940 79745
rect 2091 79736 2133 79745
rect 1940 79696 2036 79736
rect 1900 79687 1940 79696
rect 1899 79568 1941 79577
rect 1899 79528 1900 79568
rect 1940 79528 1941 79568
rect 1899 79519 1941 79528
rect 1900 78485 1940 79519
rect 1899 78476 1941 78485
rect 1899 78436 1900 78476
rect 1940 78436 1941 78476
rect 1899 78427 1941 78436
rect 1803 77216 1845 77225
rect 1803 77176 1804 77216
rect 1844 77176 1845 77216
rect 1803 77167 1845 77176
rect 1708 76924 1844 76964
rect 1707 76796 1749 76805
rect 1707 76756 1708 76796
rect 1748 76756 1749 76796
rect 1707 76747 1749 76756
rect 1708 76662 1748 76747
rect 1612 76504 1748 76544
rect 1516 76495 1556 76504
rect 1611 76376 1653 76385
rect 1420 76336 1556 76376
rect 1419 76208 1461 76217
rect 1419 76168 1420 76208
rect 1460 76168 1461 76208
rect 1419 76159 1461 76168
rect 1420 76074 1460 76159
rect 1419 75284 1461 75293
rect 1419 75244 1420 75284
rect 1460 75244 1461 75284
rect 1419 75235 1461 75244
rect 1420 75150 1460 75235
rect 1516 75200 1556 76336
rect 1611 76336 1612 76376
rect 1652 76336 1653 76376
rect 1611 76327 1653 76336
rect 1612 76040 1652 76327
rect 1612 75797 1652 76000
rect 1611 75788 1653 75797
rect 1611 75748 1612 75788
rect 1652 75748 1653 75788
rect 1611 75739 1653 75748
rect 1611 75452 1653 75461
rect 1611 75412 1612 75452
rect 1652 75412 1653 75452
rect 1611 75403 1653 75412
rect 1612 75318 1652 75403
rect 1516 75160 1652 75200
rect 1515 74444 1557 74453
rect 1515 74404 1516 74444
rect 1556 74404 1557 74444
rect 1515 74395 1557 74404
rect 1419 72848 1461 72857
rect 1419 72808 1420 72848
rect 1460 72808 1461 72848
rect 1419 72799 1461 72808
rect 1323 71840 1365 71849
rect 1323 71800 1324 71840
rect 1364 71800 1365 71840
rect 1323 71791 1365 71800
rect 1420 71681 1460 72799
rect 1419 71672 1461 71681
rect 1419 71632 1420 71672
rect 1460 71632 1461 71672
rect 1419 71623 1461 71632
rect 1323 71588 1365 71597
rect 1323 71548 1324 71588
rect 1364 71548 1365 71588
rect 1323 71539 1365 71548
rect 1035 70664 1077 70673
rect 1035 70624 1036 70664
rect 1076 70624 1077 70664
rect 1035 70615 1077 70624
rect 1227 70664 1269 70673
rect 1227 70624 1228 70664
rect 1268 70624 1269 70664
rect 1227 70615 1269 70624
rect 939 70328 981 70337
rect 939 70288 940 70328
rect 980 70288 981 70328
rect 939 70279 981 70288
rect 940 66557 980 70279
rect 939 66548 981 66557
rect 939 66508 940 66548
rect 980 66508 981 66548
rect 939 66499 981 66508
rect 1036 66473 1076 70615
rect 1228 70530 1268 70615
rect 1324 70001 1364 71539
rect 1516 71504 1556 74395
rect 1612 73688 1652 75160
rect 1612 73639 1652 73648
rect 1708 73688 1748 76504
rect 1804 75788 1844 76924
rect 1900 76712 1940 78427
rect 1996 76880 2036 79696
rect 2091 79696 2092 79736
rect 2132 79696 2133 79736
rect 2091 79687 2133 79696
rect 2092 79602 2132 79687
rect 2188 76889 2228 85936
rect 2380 85037 2420 85936
rect 2379 85028 2421 85037
rect 2379 84988 2380 85028
rect 2420 84988 2421 85028
rect 2379 84979 2421 84988
rect 2283 84356 2325 84365
rect 2283 84316 2284 84356
rect 2324 84316 2325 84356
rect 2283 84307 2325 84316
rect 2284 80417 2324 84307
rect 2572 83945 2612 85936
rect 2667 84524 2709 84533
rect 2667 84484 2668 84524
rect 2708 84484 2709 84524
rect 2667 84475 2709 84484
rect 2571 83936 2613 83945
rect 2571 83896 2572 83936
rect 2612 83896 2613 83936
rect 2571 83887 2613 83896
rect 2572 82760 2612 82769
rect 2572 82265 2612 82720
rect 2668 82601 2708 84475
rect 2764 83861 2804 85936
rect 2859 85364 2901 85373
rect 2859 85324 2860 85364
rect 2900 85324 2901 85364
rect 2859 85315 2901 85324
rect 2860 84365 2900 85315
rect 2859 84356 2901 84365
rect 2859 84316 2860 84356
rect 2900 84316 2901 84356
rect 2859 84307 2901 84316
rect 2956 83936 2996 85936
rect 3051 85196 3093 85205
rect 3051 85156 3052 85196
rect 3092 85156 3093 85196
rect 3051 85147 3093 85156
rect 3052 84449 3092 85147
rect 3051 84440 3093 84449
rect 3051 84400 3052 84440
rect 3092 84400 3093 84440
rect 3051 84391 3093 84400
rect 3148 83936 3188 85936
rect 3340 85373 3380 85936
rect 3339 85364 3381 85373
rect 3339 85324 3340 85364
rect 3380 85324 3381 85364
rect 3339 85315 3381 85324
rect 3243 85028 3285 85037
rect 3243 84988 3244 85028
rect 3284 84988 3285 85028
rect 3243 84979 3285 84988
rect 3244 84785 3284 84979
rect 3243 84776 3285 84785
rect 3243 84736 3244 84776
rect 3284 84736 3285 84776
rect 3243 84727 3285 84736
rect 3532 84701 3572 85936
rect 3724 84953 3764 85936
rect 3916 85037 3956 85936
rect 3915 85028 3957 85037
rect 3915 84988 3916 85028
rect 3956 84988 3957 85028
rect 3915 84979 3957 84988
rect 3723 84944 3765 84953
rect 3723 84904 3724 84944
rect 3764 84904 3765 84944
rect 3723 84895 3765 84904
rect 3531 84692 3573 84701
rect 3531 84652 3532 84692
rect 3572 84652 3573 84692
rect 3531 84643 3573 84652
rect 3688 84692 4056 84701
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 3688 84643 4056 84652
rect 3435 84440 3477 84449
rect 3435 84400 3436 84440
rect 3476 84400 3477 84440
rect 3435 84391 3477 84400
rect 2860 83896 2996 83936
rect 3052 83896 3188 83936
rect 3340 84272 3380 84281
rect 2763 83852 2805 83861
rect 2763 83812 2764 83852
rect 2804 83812 2805 83852
rect 2763 83803 2805 83812
rect 2763 83516 2805 83525
rect 2763 83476 2764 83516
rect 2804 83476 2805 83516
rect 2763 83467 2805 83476
rect 2764 82937 2804 83467
rect 2763 82928 2805 82937
rect 2763 82888 2764 82928
rect 2804 82888 2805 82928
rect 2763 82879 2805 82888
rect 2667 82592 2709 82601
rect 2667 82552 2668 82592
rect 2708 82552 2709 82592
rect 2667 82543 2709 82552
rect 2764 82592 2804 82601
rect 2764 82433 2804 82552
rect 2763 82424 2805 82433
rect 2763 82384 2764 82424
rect 2804 82384 2805 82424
rect 2763 82375 2805 82384
rect 2860 82349 2900 83896
rect 2956 83600 2996 83609
rect 2956 83273 2996 83560
rect 2955 83264 2997 83273
rect 2955 83224 2956 83264
rect 2996 83224 2997 83264
rect 2955 83215 2997 83224
rect 3052 83012 3092 83896
rect 3340 83861 3380 84232
rect 3339 83852 3381 83861
rect 3339 83812 3340 83852
rect 3380 83812 3381 83852
rect 3339 83803 3381 83812
rect 3340 83600 3380 83611
rect 3340 83525 3380 83560
rect 3339 83516 3381 83525
rect 3339 83476 3340 83516
rect 3380 83476 3381 83516
rect 3339 83467 3381 83476
rect 3148 83348 3188 83357
rect 3148 83180 3188 83308
rect 3148 83140 3380 83180
rect 2956 82972 3092 83012
rect 3147 83012 3189 83021
rect 3147 82972 3148 83012
rect 3188 82972 3189 83012
rect 2859 82340 2901 82349
rect 2859 82300 2860 82340
rect 2900 82300 2901 82340
rect 2859 82291 2901 82300
rect 2571 82256 2613 82265
rect 2571 82216 2572 82256
rect 2612 82216 2613 82256
rect 2956 82256 2996 82972
rect 3147 82963 3189 82972
rect 3051 82844 3093 82853
rect 3051 82804 3052 82844
rect 3092 82804 3093 82844
rect 3051 82795 3093 82804
rect 3052 82710 3092 82795
rect 3052 82256 3092 82265
rect 2956 82216 3052 82256
rect 2571 82207 2613 82216
rect 3052 82207 3092 82216
rect 2476 82088 2516 82097
rect 2572 82088 2612 82207
rect 2859 82172 2901 82181
rect 2859 82132 2860 82172
rect 2900 82132 2901 82172
rect 2859 82123 2901 82132
rect 2516 82048 2612 82088
rect 2476 82039 2516 82048
rect 2860 82004 2900 82123
rect 2860 81955 2900 81964
rect 2668 81836 2708 81845
rect 2708 81796 2804 81836
rect 2668 81787 2708 81796
rect 2764 81509 2804 81796
rect 2763 81500 2805 81509
rect 2763 81460 2764 81500
rect 2804 81460 2805 81500
rect 2763 81451 2805 81460
rect 3051 81500 3093 81509
rect 3051 81460 3052 81500
rect 3092 81460 3093 81500
rect 3051 81451 3093 81460
rect 3052 81416 3092 81451
rect 3052 81365 3092 81376
rect 3148 81257 3188 82963
rect 3243 82592 3285 82601
rect 3243 82552 3244 82592
rect 3284 82552 3285 82592
rect 3243 82543 3285 82552
rect 3244 82458 3284 82543
rect 3243 82340 3285 82349
rect 3243 82300 3244 82340
rect 3284 82300 3285 82340
rect 3243 82291 3285 82300
rect 2476 81248 2516 81257
rect 2379 80828 2421 80837
rect 2379 80788 2380 80828
rect 2420 80788 2421 80828
rect 2379 80779 2421 80788
rect 2380 80576 2420 80779
rect 2380 80527 2420 80536
rect 2283 80408 2325 80417
rect 2283 80368 2284 80408
rect 2324 80368 2325 80408
rect 2283 80359 2325 80368
rect 2283 80156 2325 80165
rect 2283 80116 2284 80156
rect 2324 80116 2325 80156
rect 2283 80107 2325 80116
rect 2092 76880 2132 76889
rect 1996 76840 2092 76880
rect 2092 76831 2132 76840
rect 2187 76880 2229 76889
rect 2187 76840 2188 76880
rect 2228 76840 2229 76880
rect 2187 76831 2229 76840
rect 2092 76712 2132 76721
rect 1900 76672 2092 76712
rect 2092 76663 2132 76672
rect 2188 76712 2228 76723
rect 2188 76637 2228 76672
rect 2187 76628 2229 76637
rect 2187 76588 2188 76628
rect 2228 76588 2229 76628
rect 2187 76579 2229 76588
rect 1899 76544 1941 76553
rect 1899 76504 1900 76544
rect 1940 76504 1941 76544
rect 1899 76495 1941 76504
rect 1900 76410 1940 76495
rect 1804 75748 2132 75788
rect 1803 75536 1845 75545
rect 1803 75496 1804 75536
rect 1844 75496 1845 75536
rect 1803 75487 1845 75496
rect 1708 73100 1748 73648
rect 1612 73060 1748 73100
rect 1612 71672 1652 73060
rect 1708 72176 1748 72185
rect 1804 72176 1844 75487
rect 1899 74864 1941 74873
rect 1899 74824 1900 74864
rect 1940 74824 1941 74864
rect 1899 74815 1941 74824
rect 1900 74528 1940 74815
rect 1900 74479 1940 74488
rect 2092 73772 2132 75748
rect 2188 75452 2228 75461
rect 2284 75452 2324 80107
rect 2476 79064 2516 81208
rect 2859 81248 2901 81257
rect 2859 81208 2860 81248
rect 2900 81208 2901 81248
rect 2859 81199 2901 81208
rect 3147 81248 3189 81257
rect 3147 81208 3148 81248
rect 3188 81208 3189 81248
rect 3147 81199 3189 81208
rect 2668 81080 2708 81089
rect 2571 79736 2613 79745
rect 2571 79696 2572 79736
rect 2612 79696 2613 79736
rect 2571 79687 2613 79696
rect 2380 79024 2476 79064
rect 2380 77552 2420 79024
rect 2476 79015 2516 79024
rect 2572 78896 2612 79687
rect 2668 79400 2708 81040
rect 2860 80571 2900 81199
rect 3147 81080 3189 81089
rect 3147 81040 3148 81080
rect 3188 81040 3189 81080
rect 3147 81031 3189 81040
rect 3148 80946 3188 81031
rect 3052 80660 3092 80669
rect 3092 80620 3188 80660
rect 3052 80611 3092 80620
rect 2860 80522 2900 80531
rect 3051 80492 3093 80501
rect 3051 80452 3052 80492
rect 3092 80452 3093 80492
rect 3051 80443 3093 80452
rect 2859 80240 2901 80249
rect 2859 80200 2860 80240
rect 2900 80200 2901 80240
rect 2859 80191 2901 80200
rect 2668 79360 2804 79400
rect 2476 78856 2612 78896
rect 2476 78233 2516 78856
rect 2668 78812 2708 78821
rect 2572 78772 2668 78812
rect 2475 78224 2517 78233
rect 2475 78184 2476 78224
rect 2516 78184 2517 78224
rect 2475 78175 2517 78184
rect 2476 78090 2516 78175
rect 2475 77552 2517 77561
rect 2380 77512 2476 77552
rect 2516 77512 2517 77552
rect 2475 77503 2517 77512
rect 2476 77418 2516 77503
rect 2380 76712 2420 76752
rect 2380 76637 2420 76672
rect 2379 76628 2421 76637
rect 2379 76588 2380 76628
rect 2420 76588 2421 76628
rect 2379 76579 2421 76588
rect 2380 75629 2420 76579
rect 2379 75620 2421 75629
rect 2379 75580 2380 75620
rect 2420 75580 2421 75620
rect 2379 75571 2421 75580
rect 2228 75412 2324 75452
rect 2188 75403 2228 75412
rect 2475 75368 2517 75377
rect 2475 75328 2476 75368
rect 2516 75328 2517 75368
rect 2475 75319 2517 75328
rect 2380 75284 2420 75293
rect 2283 74696 2325 74705
rect 2283 74656 2284 74696
rect 2324 74656 2325 74696
rect 2283 74647 2325 74656
rect 2187 74024 2229 74033
rect 2187 73984 2188 74024
rect 2228 73984 2229 74024
rect 2187 73975 2229 73984
rect 2092 73100 2132 73732
rect 2188 73772 2228 73975
rect 2188 73723 2228 73732
rect 1748 72136 1844 72176
rect 1900 73060 2132 73100
rect 1708 72127 1748 72136
rect 1803 71840 1845 71849
rect 1803 71800 1804 71840
rect 1844 71800 1845 71840
rect 1803 71791 1845 71800
rect 1612 71632 1748 71672
rect 1516 71455 1556 71464
rect 1612 71504 1652 71513
rect 1419 71168 1461 71177
rect 1419 71128 1420 71168
rect 1460 71128 1461 71168
rect 1419 71119 1461 71128
rect 1228 69992 1268 70001
rect 1228 69824 1268 69952
rect 1323 69992 1365 70001
rect 1323 69952 1324 69992
rect 1364 69952 1365 69992
rect 1323 69943 1365 69952
rect 1420 69824 1460 71119
rect 1228 69784 1460 69824
rect 1227 69152 1269 69161
rect 1227 69112 1228 69152
rect 1268 69112 1269 69152
rect 1227 69103 1269 69112
rect 1228 69018 1268 69103
rect 1227 68396 1269 68405
rect 1227 68356 1228 68396
rect 1268 68356 1269 68396
rect 1227 68347 1269 68356
rect 1131 66800 1173 66809
rect 1131 66760 1132 66800
rect 1172 66760 1173 66800
rect 1131 66751 1173 66760
rect 1035 66464 1077 66473
rect 1035 66424 1036 66464
rect 1076 66424 1077 66464
rect 1035 66415 1077 66424
rect 747 65204 789 65213
rect 747 65164 748 65204
rect 788 65164 789 65204
rect 747 65155 789 65164
rect 459 64280 501 64289
rect 459 64240 460 64280
rect 500 64240 501 64280
rect 459 64231 501 64240
rect 651 61340 693 61349
rect 651 61300 652 61340
rect 692 61300 693 61340
rect 651 61291 693 61300
rect 363 60248 405 60257
rect 363 60208 364 60248
rect 404 60208 405 60248
rect 363 60199 405 60208
rect 652 57644 692 61291
rect 748 59249 788 65155
rect 939 63020 981 63029
rect 939 62980 940 63020
rect 980 62980 981 63020
rect 939 62971 981 62980
rect 843 61004 885 61013
rect 843 60964 844 61004
rect 884 60964 885 61004
rect 843 60955 885 60964
rect 747 59240 789 59249
rect 747 59200 748 59240
rect 788 59200 789 59240
rect 747 59191 789 59200
rect 844 57728 884 60955
rect 940 58913 980 62971
rect 1035 61760 1077 61769
rect 1035 61720 1036 61760
rect 1076 61720 1077 61760
rect 1035 61711 1077 61720
rect 939 58904 981 58913
rect 939 58864 940 58904
rect 980 58864 981 58904
rect 939 58855 981 58864
rect 844 57688 980 57728
rect 652 57604 884 57644
rect 76 55420 212 55460
rect 172 51773 212 55420
rect 651 55376 693 55385
rect 651 55336 652 55376
rect 692 55336 693 55376
rect 651 55327 693 55336
rect 555 55292 597 55301
rect 555 55252 556 55292
rect 596 55252 597 55292
rect 555 55243 597 55252
rect 171 51764 213 51773
rect 171 51724 172 51764
rect 212 51724 213 51764
rect 171 51715 213 51724
rect 556 50933 596 55243
rect 555 50924 597 50933
rect 555 50884 556 50924
rect 596 50884 597 50924
rect 555 50875 597 50884
rect 652 47153 692 55327
rect 747 51680 789 51689
rect 747 51640 748 51680
rect 788 51640 789 51680
rect 747 51631 789 51640
rect 651 47144 693 47153
rect 651 47104 652 47144
rect 692 47104 693 47144
rect 651 47095 693 47104
rect 748 41600 788 51631
rect 844 51344 884 57604
rect 940 55217 980 57688
rect 939 55208 981 55217
rect 939 55168 940 55208
rect 980 55168 981 55208
rect 939 55159 981 55168
rect 844 51304 980 51344
rect 843 50924 885 50933
rect 843 50884 844 50924
rect 884 50884 885 50924
rect 843 50875 885 50884
rect 652 41560 788 41600
rect 555 39752 597 39761
rect 555 39712 556 39752
rect 596 39712 597 39752
rect 555 39703 597 39712
rect 556 34049 596 39703
rect 555 34040 597 34049
rect 555 34000 556 34040
rect 596 34000 597 34040
rect 555 33991 597 34000
rect 652 33209 692 41560
rect 747 33536 789 33545
rect 747 33496 748 33536
rect 788 33496 789 33536
rect 747 33487 789 33496
rect 651 33200 693 33209
rect 651 33160 652 33200
rect 692 33160 693 33200
rect 651 33151 693 33160
rect 171 33032 213 33041
rect 171 32992 172 33032
rect 212 32992 213 33032
rect 171 32983 213 32992
rect 75 32192 117 32201
rect 75 32152 76 32192
rect 116 32152 117 32192
rect 75 32143 117 32152
rect 76 19265 116 32143
rect 172 23213 212 32983
rect 555 32444 597 32453
rect 555 32404 556 32444
rect 596 32404 597 32444
rect 555 32395 597 32404
rect 363 31016 405 31025
rect 363 30976 364 31016
rect 404 30976 405 31016
rect 363 30967 405 30976
rect 364 23717 404 30967
rect 556 25313 596 32395
rect 748 28925 788 33487
rect 747 28916 789 28925
rect 747 28876 748 28916
rect 788 28876 789 28916
rect 747 28867 789 28876
rect 844 27077 884 50875
rect 940 30941 980 51304
rect 1036 33545 1076 61711
rect 1132 33629 1172 66751
rect 1228 62273 1268 68347
rect 1324 64028 1364 69784
rect 1419 69572 1461 69581
rect 1419 69532 1420 69572
rect 1460 69532 1461 69572
rect 1419 69523 1461 69532
rect 1420 66464 1460 69523
rect 1612 68732 1652 71464
rect 1516 68692 1652 68732
rect 1516 68405 1556 68692
rect 1708 68648 1748 71632
rect 1804 71429 1844 71791
rect 1803 71420 1845 71429
rect 1803 71380 1804 71420
rect 1844 71380 1845 71420
rect 1803 71371 1845 71380
rect 1900 69581 1940 73060
rect 2091 71672 2133 71681
rect 2091 71632 2092 71672
rect 2132 71632 2133 71672
rect 2091 71623 2133 71632
rect 2092 71504 2132 71623
rect 2092 71455 2132 71464
rect 1996 71420 2036 71429
rect 1996 70832 2036 71380
rect 1996 70792 2228 70832
rect 2091 70664 2133 70673
rect 2091 70624 2092 70664
rect 2132 70624 2133 70664
rect 2091 70615 2133 70624
rect 1899 69572 1941 69581
rect 1899 69532 1900 69572
rect 1940 69532 1941 69572
rect 1899 69523 1941 69532
rect 1899 69404 1941 69413
rect 1899 69364 1900 69404
rect 1940 69364 1941 69404
rect 1899 69355 1941 69364
rect 1612 68608 1748 68648
rect 1515 68396 1557 68405
rect 1515 68356 1516 68396
rect 1556 68356 1557 68396
rect 1515 68347 1557 68356
rect 1420 66424 1556 66464
rect 1419 66296 1461 66305
rect 1419 66256 1420 66296
rect 1460 66256 1461 66296
rect 1419 66247 1461 66256
rect 1420 66128 1460 66247
rect 1420 64280 1460 66088
rect 1516 65633 1556 66424
rect 1515 65624 1557 65633
rect 1515 65584 1516 65624
rect 1556 65584 1557 65624
rect 1515 65575 1557 65584
rect 1420 64240 1556 64280
rect 1419 64028 1461 64037
rect 1324 63988 1420 64028
rect 1460 63988 1461 64028
rect 1419 63979 1461 63988
rect 1420 63944 1460 63979
rect 1420 63893 1460 63904
rect 1419 63776 1461 63785
rect 1419 63736 1420 63776
rect 1460 63736 1461 63776
rect 1419 63727 1461 63736
rect 1323 63692 1365 63701
rect 1323 63652 1324 63692
rect 1364 63652 1365 63692
rect 1323 63643 1365 63652
rect 1324 62432 1364 63643
rect 1420 62777 1460 63727
rect 1516 63440 1556 64240
rect 1612 63785 1652 68608
rect 1707 68480 1749 68489
rect 1707 68440 1708 68480
rect 1748 68440 1749 68480
rect 1707 68431 1749 68440
rect 1804 68480 1844 68491
rect 1708 68346 1748 68431
rect 1804 68405 1844 68440
rect 1803 68396 1845 68405
rect 1803 68356 1804 68396
rect 1844 68356 1845 68396
rect 1803 68347 1845 68356
rect 1804 67640 1844 67649
rect 1900 67640 1940 69355
rect 2092 68480 2132 70615
rect 1844 67600 1940 67640
rect 1996 68440 2132 68480
rect 1611 63776 1653 63785
rect 1611 63736 1612 63776
rect 1652 63736 1653 63776
rect 1611 63727 1653 63736
rect 1516 63400 1652 63440
rect 1515 63272 1557 63281
rect 1515 63232 1516 63272
rect 1556 63232 1557 63272
rect 1515 63223 1557 63232
rect 1516 63138 1556 63223
rect 1515 62852 1557 62861
rect 1515 62812 1516 62852
rect 1556 62812 1557 62852
rect 1515 62803 1557 62812
rect 1419 62768 1461 62777
rect 1419 62728 1420 62768
rect 1460 62728 1461 62768
rect 1419 62719 1461 62728
rect 1227 62264 1269 62273
rect 1227 62224 1228 62264
rect 1268 62224 1269 62264
rect 1227 62215 1269 62224
rect 1324 61592 1364 62392
rect 1324 61543 1364 61552
rect 1516 61265 1556 62803
rect 1515 61256 1557 61265
rect 1515 61216 1516 61256
rect 1556 61216 1557 61256
rect 1515 61207 1557 61216
rect 1612 60929 1652 63400
rect 1707 63188 1749 63197
rect 1707 63148 1708 63188
rect 1748 63148 1749 63188
rect 1707 63139 1749 63148
rect 1708 63054 1748 63139
rect 1804 61928 1844 67600
rect 1996 66221 2036 68440
rect 2188 68396 2228 70792
rect 2091 68228 2133 68237
rect 2091 68188 2092 68228
rect 2132 68188 2133 68228
rect 2091 68179 2133 68188
rect 1995 66212 2037 66221
rect 1995 66172 1996 66212
rect 2036 66172 2037 66212
rect 1995 66163 2037 66172
rect 2092 64616 2132 68179
rect 2188 64961 2228 68356
rect 2284 68480 2324 74647
rect 2380 73949 2420 75244
rect 2379 73940 2421 73949
rect 2379 73900 2380 73940
rect 2420 73900 2421 73940
rect 2379 73891 2421 73900
rect 2476 73772 2516 75319
rect 2572 75200 2612 78772
rect 2668 78763 2708 78772
rect 2667 78140 2709 78149
rect 2667 78100 2668 78140
rect 2708 78100 2709 78140
rect 2667 78091 2709 78100
rect 2668 78006 2708 78091
rect 2668 77309 2708 77394
rect 2667 77300 2709 77309
rect 2667 77260 2668 77300
rect 2708 77260 2709 77300
rect 2667 77251 2709 77260
rect 2764 77132 2804 79360
rect 2860 79148 2900 80191
rect 3052 79577 3092 80443
rect 3051 79568 3093 79577
rect 3051 79528 3052 79568
rect 3092 79528 3093 79568
rect 3051 79519 3093 79528
rect 2955 79400 2997 79409
rect 2955 79360 2956 79400
rect 2996 79360 2997 79400
rect 2955 79351 2997 79360
rect 2956 79232 2996 79351
rect 3052 79232 3092 79241
rect 2956 79192 3052 79232
rect 3052 79183 3092 79192
rect 2860 79108 2996 79148
rect 2859 78980 2901 78989
rect 2859 78940 2860 78980
rect 2900 78940 2901 78980
rect 2859 78931 2901 78940
rect 2860 78846 2900 78931
rect 2956 78224 2996 79108
rect 3148 78392 3188 80620
rect 3244 79232 3284 82291
rect 3340 81248 3380 83140
rect 3436 82844 3476 84391
rect 3723 84272 3765 84281
rect 3723 84232 3724 84272
rect 3764 84232 3765 84272
rect 3723 84223 3765 84232
rect 3724 84138 3764 84223
rect 3532 84104 3572 84113
rect 3532 83021 3572 84064
rect 4108 83945 4148 85936
rect 4300 84449 4340 85936
rect 4299 84440 4341 84449
rect 4299 84400 4300 84440
rect 4340 84400 4341 84440
rect 4299 84391 4341 84400
rect 4395 84104 4437 84113
rect 4395 84064 4396 84104
rect 4436 84064 4437 84104
rect 4395 84055 4437 84064
rect 4107 83936 4149 83945
rect 4107 83896 4108 83936
rect 4148 83896 4149 83936
rect 4107 83887 4149 83896
rect 4299 83600 4341 83609
rect 4299 83560 4300 83600
rect 4340 83560 4341 83600
rect 4299 83551 4341 83560
rect 3688 83180 4056 83189
rect 4203 83180 4245 83189
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 3688 83131 4056 83140
rect 4108 83140 4204 83180
rect 4244 83140 4245 83180
rect 3531 83012 3573 83021
rect 3531 82972 3532 83012
rect 3572 82972 3573 83012
rect 3531 82963 3573 82972
rect 4011 83012 4053 83021
rect 4011 82972 4012 83012
rect 4052 82972 4053 83012
rect 4011 82963 4053 82972
rect 3436 82804 3668 82844
rect 3436 82718 3476 82727
rect 3436 82340 3476 82678
rect 3436 82300 3572 82340
rect 3436 82013 3476 82098
rect 3435 82004 3477 82013
rect 3435 81964 3436 82004
rect 3476 81964 3477 82004
rect 3435 81955 3477 81964
rect 3532 81416 3572 82300
rect 3628 82256 3668 82804
rect 3628 82207 3668 82216
rect 4012 82256 4052 82963
rect 4012 82207 4052 82216
rect 3820 82013 3860 82098
rect 3819 82004 3861 82013
rect 3819 81964 3820 82004
rect 3860 81964 3861 82004
rect 3819 81955 3861 81964
rect 3688 81668 4056 81677
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 3688 81619 4056 81628
rect 4011 81500 4053 81509
rect 4011 81460 4012 81500
rect 4052 81460 4053 81500
rect 4011 81451 4053 81460
rect 3532 81376 3668 81416
rect 3436 81248 3476 81257
rect 3340 81208 3436 81248
rect 3436 81199 3476 81208
rect 3531 81248 3573 81257
rect 3531 81208 3532 81248
rect 3572 81208 3573 81248
rect 3531 81199 3573 81208
rect 3532 81114 3572 81199
rect 3339 81080 3381 81089
rect 3339 81040 3340 81080
rect 3380 81040 3381 81080
rect 3339 81031 3381 81040
rect 3340 80744 3380 81031
rect 3628 80996 3668 81376
rect 4012 81332 4052 81451
rect 4012 81283 4052 81292
rect 3915 81248 3957 81257
rect 3915 81208 3916 81248
rect 3956 81208 3957 81248
rect 3915 81199 3957 81208
rect 3916 81114 3956 81199
rect 3532 80956 3668 80996
rect 3435 80912 3477 80921
rect 3435 80872 3436 80912
rect 3476 80872 3477 80912
rect 3435 80863 3477 80872
rect 3340 80081 3380 80704
rect 3339 80072 3381 80081
rect 3339 80032 3340 80072
rect 3380 80032 3381 80072
rect 3339 80023 3381 80032
rect 3340 79736 3380 79745
rect 3436 79736 3476 80863
rect 3532 80501 3572 80956
rect 4108 80921 4148 83140
rect 4203 83131 4245 83140
rect 4204 82013 4244 82098
rect 4203 82004 4245 82013
rect 4203 81964 4204 82004
rect 4244 81964 4245 82004
rect 4203 81955 4245 81964
rect 4300 81668 4340 83551
rect 4396 82256 4436 84055
rect 4396 82207 4436 82216
rect 4492 82013 4532 85936
rect 4587 84440 4629 84449
rect 4587 84400 4588 84440
rect 4628 84400 4629 84440
rect 4587 84391 4629 84400
rect 4588 83600 4628 84391
rect 4684 83768 4724 85936
rect 4876 84113 4916 85936
rect 5068 84617 5108 85936
rect 5163 84692 5205 84701
rect 5163 84652 5164 84692
rect 5204 84652 5205 84692
rect 5163 84643 5205 84652
rect 5067 84608 5109 84617
rect 5067 84568 5068 84608
rect 5108 84568 5109 84608
rect 5067 84559 5109 84568
rect 5164 84524 5204 84643
rect 5260 84533 5300 85936
rect 5164 84475 5204 84484
rect 5259 84524 5301 84533
rect 5259 84484 5260 84524
rect 5300 84484 5301 84524
rect 5259 84475 5301 84484
rect 4971 84440 5013 84449
rect 4971 84400 4972 84440
rect 5012 84400 5013 84440
rect 4971 84391 5013 84400
rect 4972 84272 5012 84391
rect 5012 84232 5108 84272
rect 4972 84223 5012 84232
rect 5068 84113 5108 84232
rect 4875 84104 4917 84113
rect 4875 84064 4876 84104
rect 4916 84064 4917 84104
rect 4875 84055 4917 84064
rect 5067 84104 5109 84113
rect 5067 84064 5068 84104
rect 5108 84064 5109 84104
rect 5067 84055 5109 84064
rect 5356 84104 5396 84113
rect 4928 83936 5296 83945
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 4928 83887 5296 83896
rect 4684 83728 4916 83768
rect 4588 83348 4628 83560
rect 4779 83348 4821 83357
rect 4588 83308 4724 83348
rect 4684 83189 4724 83308
rect 4779 83308 4780 83348
rect 4820 83308 4821 83348
rect 4876 83348 4916 83728
rect 4971 83600 5013 83609
rect 4971 83560 4972 83600
rect 5012 83560 5013 83600
rect 4971 83551 5013 83560
rect 4972 83466 5012 83551
rect 4876 83308 5012 83348
rect 4779 83299 4821 83308
rect 4780 83214 4820 83299
rect 4683 83180 4725 83189
rect 4683 83140 4684 83180
rect 4724 83140 4725 83180
rect 4683 83131 4725 83140
rect 4875 83180 4917 83189
rect 4875 83140 4876 83180
rect 4916 83140 4917 83180
rect 4875 83131 4917 83140
rect 4587 82760 4629 82769
rect 4587 82720 4588 82760
rect 4628 82720 4629 82760
rect 4587 82711 4629 82720
rect 4684 82760 4724 83131
rect 4876 82937 4916 83131
rect 4875 82928 4917 82937
rect 4875 82888 4876 82928
rect 4916 82888 4917 82928
rect 4875 82879 4917 82888
rect 4972 82769 5012 83308
rect 5356 83273 5396 84064
rect 5355 83264 5397 83273
rect 5355 83224 5356 83264
rect 5396 83224 5397 83264
rect 5355 83215 5397 83224
rect 5452 83021 5492 85936
rect 5644 84953 5684 85936
rect 5836 85289 5876 85936
rect 5835 85280 5877 85289
rect 5835 85240 5836 85280
rect 5876 85240 5877 85280
rect 5835 85231 5877 85240
rect 5643 84944 5685 84953
rect 5643 84904 5644 84944
rect 5684 84904 5685 84944
rect 5643 84895 5685 84904
rect 5643 84524 5685 84533
rect 5643 84484 5644 84524
rect 5684 84484 5685 84524
rect 5643 84475 5685 84484
rect 5547 84272 5589 84281
rect 5547 84232 5548 84272
rect 5588 84232 5589 84272
rect 5547 84223 5589 84232
rect 5548 83861 5588 84223
rect 5547 83852 5589 83861
rect 5547 83812 5548 83852
rect 5588 83812 5589 83852
rect 5547 83803 5589 83812
rect 5547 83264 5589 83273
rect 5547 83224 5548 83264
rect 5588 83224 5589 83264
rect 5547 83215 5589 83224
rect 5451 83012 5493 83021
rect 5451 82972 5452 83012
rect 5492 82972 5493 83012
rect 5451 82963 5493 82972
rect 5163 82928 5205 82937
rect 5163 82888 5164 82928
rect 5204 82888 5205 82928
rect 5163 82879 5205 82888
rect 5164 82794 5204 82879
rect 5451 82844 5493 82853
rect 5451 82804 5452 82844
rect 5492 82804 5493 82844
rect 5451 82795 5493 82804
rect 4684 82711 4724 82720
rect 4971 82760 5013 82769
rect 4971 82720 4972 82760
rect 5012 82720 5013 82760
rect 4971 82711 5013 82720
rect 4491 82004 4533 82013
rect 4491 81964 4492 82004
rect 4532 81964 4533 82004
rect 4491 81955 4533 81964
rect 4588 81920 4628 82711
rect 5452 82710 5492 82795
rect 4876 82592 4916 82601
rect 4780 82552 4876 82592
rect 4780 82256 4820 82552
rect 4876 82543 4916 82552
rect 4928 82424 5296 82433
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 4928 82375 5296 82384
rect 4780 82216 5012 82256
rect 4683 82172 4725 82181
rect 4683 82132 4684 82172
rect 4724 82132 4725 82172
rect 4683 82123 4725 82132
rect 4684 82088 4724 82123
rect 4684 82037 4724 82048
rect 4780 82088 4820 82097
rect 4780 81929 4820 82048
rect 4779 81920 4821 81929
rect 4588 81880 4724 81920
rect 4491 81752 4533 81761
rect 4491 81712 4492 81752
rect 4532 81712 4533 81752
rect 4491 81703 4533 81712
rect 4204 81628 4340 81668
rect 4204 81425 4244 81628
rect 4299 81500 4341 81509
rect 4299 81460 4300 81500
rect 4340 81460 4341 81500
rect 4299 81451 4341 81460
rect 4203 81416 4245 81425
rect 4203 81376 4204 81416
rect 4244 81376 4245 81416
rect 4203 81367 4245 81376
rect 4204 81005 4244 81367
rect 4203 80996 4245 81005
rect 4203 80956 4204 80996
rect 4244 80956 4245 80996
rect 4203 80947 4245 80956
rect 4107 80912 4149 80921
rect 4107 80872 4108 80912
rect 4148 80872 4149 80912
rect 4107 80863 4149 80872
rect 3723 80828 3765 80837
rect 3723 80788 3724 80828
rect 3764 80788 3765 80828
rect 3723 80779 3765 80788
rect 3724 80744 3764 80779
rect 3724 80693 3764 80704
rect 3868 80534 3908 80543
rect 3531 80492 3573 80501
rect 3868 80492 3908 80494
rect 3531 80452 3532 80492
rect 3572 80452 3573 80492
rect 3531 80443 3573 80452
rect 3628 80452 3908 80492
rect 3628 80324 3668 80452
rect 3532 80284 3668 80324
rect 3532 79988 3572 80284
rect 3688 80156 4056 80165
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 3688 80107 4056 80116
rect 3532 79939 3572 79948
rect 4012 79745 4052 79830
rect 3380 79696 3476 79736
rect 4011 79736 4053 79745
rect 4011 79696 4012 79736
rect 4052 79696 4053 79736
rect 3340 79687 3380 79696
rect 4011 79687 4053 79696
rect 3531 79568 3573 79577
rect 3531 79528 3532 79568
rect 3572 79528 3573 79568
rect 3531 79519 3573 79528
rect 3820 79568 3860 79577
rect 3244 79192 3380 79232
rect 3244 79064 3284 79073
rect 3244 78569 3284 79024
rect 3243 78560 3285 78569
rect 3243 78520 3244 78560
rect 3284 78520 3285 78560
rect 3243 78511 3285 78520
rect 3148 78352 3284 78392
rect 2956 78175 2996 78184
rect 3052 78224 3092 78233
rect 2955 77720 2997 77729
rect 2955 77680 2956 77720
rect 2996 77680 2997 77720
rect 2955 77671 2997 77680
rect 2859 77552 2901 77561
rect 2859 77512 2860 77552
rect 2900 77512 2901 77552
rect 2859 77503 2901 77512
rect 2956 77552 2996 77671
rect 2956 77503 2996 77512
rect 2668 77092 2804 77132
rect 2668 76712 2708 77092
rect 2668 76663 2708 76672
rect 2764 76712 2804 76723
rect 2764 76637 2804 76672
rect 2763 76628 2805 76637
rect 2763 76588 2764 76628
rect 2804 76588 2805 76628
rect 2763 76579 2805 76588
rect 2860 76040 2900 77503
rect 2955 77300 2997 77309
rect 2955 77260 2956 77300
rect 2996 77260 2997 77300
rect 2955 77251 2997 77260
rect 2668 75200 2708 75209
rect 2572 75160 2668 75200
rect 2668 75151 2708 75160
rect 2763 75200 2805 75209
rect 2763 75160 2764 75200
rect 2804 75160 2805 75200
rect 2763 75151 2805 75160
rect 2764 75066 2804 75151
rect 2571 75032 2613 75041
rect 2571 74992 2572 75032
rect 2612 74992 2613 75032
rect 2571 74983 2613 74992
rect 2380 73732 2516 73772
rect 2380 70673 2420 73732
rect 2476 73016 2516 73025
rect 2572 73016 2612 74983
rect 2860 74789 2900 76000
rect 2859 74780 2901 74789
rect 2859 74740 2860 74780
rect 2900 74740 2901 74780
rect 2859 74731 2901 74740
rect 2956 74453 2996 77251
rect 3052 76637 3092 78184
rect 3147 78224 3189 78233
rect 3147 78184 3148 78224
rect 3188 78184 3189 78224
rect 3147 78175 3189 78184
rect 3148 76805 3188 78175
rect 3244 76889 3284 78352
rect 3340 77225 3380 79192
rect 3532 78737 3572 79519
rect 3820 78821 3860 79528
rect 4300 79232 4340 81451
rect 4492 81248 4532 81703
rect 4492 81199 4532 81208
rect 4491 80828 4533 80837
rect 4491 80788 4492 80828
rect 4532 80788 4533 80828
rect 4491 80779 4533 80788
rect 4396 80576 4436 80585
rect 4396 80417 4436 80536
rect 4395 80408 4437 80417
rect 4395 80368 4396 80408
rect 4436 80368 4437 80408
rect 4395 80359 4437 80368
rect 4492 80249 4532 80779
rect 4587 80744 4629 80753
rect 4587 80704 4588 80744
rect 4628 80704 4629 80744
rect 4587 80695 4629 80704
rect 4491 80240 4533 80249
rect 4491 80200 4492 80240
rect 4532 80200 4533 80240
rect 4491 80191 4533 80200
rect 4588 79913 4628 80695
rect 4587 79904 4629 79913
rect 4587 79864 4588 79904
rect 4628 79864 4629 79904
rect 4587 79855 4629 79864
rect 4108 79192 4340 79232
rect 3819 78812 3861 78821
rect 3819 78772 3820 78812
rect 3860 78772 3861 78812
rect 3819 78763 3861 78772
rect 3531 78728 3573 78737
rect 3531 78688 3532 78728
rect 3572 78688 3573 78728
rect 3531 78679 3573 78688
rect 3688 78644 4056 78653
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 3688 78595 4056 78604
rect 3531 78392 3573 78401
rect 3531 78352 3532 78392
rect 3572 78352 3573 78392
rect 3531 78343 3573 78352
rect 3532 78308 3572 78343
rect 3532 78257 3572 78268
rect 3435 78224 3477 78233
rect 3435 78184 3436 78224
rect 3476 78184 3477 78224
rect 3435 78175 3477 78184
rect 4012 78224 4052 78233
rect 4108 78224 4148 79192
rect 4492 79073 4532 79158
rect 4684 79148 4724 81880
rect 4779 81880 4780 81920
rect 4820 81880 4821 81920
rect 4779 81871 4821 81880
rect 4972 81262 5012 82216
rect 5163 82172 5205 82181
rect 5163 82132 5164 82172
rect 5204 82132 5205 82172
rect 5163 82123 5205 82132
rect 5164 82088 5204 82123
rect 5164 82037 5204 82048
rect 5260 82004 5300 82013
rect 5163 81500 5205 81509
rect 5163 81460 5164 81500
rect 5204 81460 5205 81500
rect 5163 81451 5205 81460
rect 4972 81213 5012 81222
rect 5164 81164 5204 81451
rect 5164 81115 5204 81124
rect 5260 81080 5300 81964
rect 5355 81920 5397 81929
rect 5355 81880 5356 81920
rect 5396 81880 5397 81920
rect 5548 81920 5588 83215
rect 5644 83012 5684 84475
rect 6028 84449 6068 85936
rect 6123 85280 6165 85289
rect 6123 85240 6124 85280
rect 6164 85240 6165 85280
rect 6123 85231 6165 85240
rect 6027 84440 6069 84449
rect 6027 84400 6028 84440
rect 6068 84400 6069 84440
rect 6027 84391 6069 84400
rect 5931 84188 5973 84197
rect 5931 84148 5932 84188
rect 5972 84148 5973 84188
rect 5931 84139 5973 84148
rect 5644 82963 5684 82972
rect 5836 82844 5876 82853
rect 5739 82340 5781 82349
rect 5739 82300 5740 82340
rect 5780 82300 5781 82340
rect 5739 82291 5781 82300
rect 5740 82088 5780 82291
rect 5740 82039 5780 82048
rect 5836 81920 5876 82804
rect 5932 82181 5972 84139
rect 6028 83012 6068 83021
rect 6124 83012 6164 85231
rect 6220 85037 6260 85936
rect 6219 85028 6261 85037
rect 6219 84988 6220 85028
rect 6260 84988 6261 85028
rect 6219 84979 6261 84988
rect 6412 84449 6452 85936
rect 6604 84449 6644 85936
rect 6796 85625 6836 85936
rect 6988 85709 7028 85936
rect 6987 85700 7029 85709
rect 6987 85660 6988 85700
rect 7028 85660 7029 85700
rect 6987 85651 7029 85660
rect 6795 85616 6837 85625
rect 6795 85576 6796 85616
rect 6836 85576 6837 85616
rect 6795 85567 6837 85576
rect 6795 85448 6837 85457
rect 6795 85408 6796 85448
rect 6836 85408 6837 85448
rect 6795 85399 6837 85408
rect 6796 84617 6836 85399
rect 6795 84608 6837 84617
rect 6795 84568 6796 84608
rect 6836 84568 6837 84608
rect 6795 84559 6837 84568
rect 6411 84440 6453 84449
rect 6411 84400 6412 84440
rect 6452 84400 6453 84440
rect 6411 84391 6453 84400
rect 6603 84440 6645 84449
rect 6603 84400 6604 84440
rect 6644 84400 6645 84440
rect 6603 84391 6645 84400
rect 6796 84272 6836 84559
rect 6987 84356 7029 84365
rect 6987 84316 6988 84356
rect 7028 84316 7029 84356
rect 6987 84307 7029 84316
rect 7084 84356 7124 84365
rect 6796 84223 6836 84232
rect 6219 84104 6261 84113
rect 6219 84064 6220 84104
rect 6260 84064 6261 84104
rect 6219 84055 6261 84064
rect 6220 83609 6260 84055
rect 6699 83936 6741 83945
rect 6699 83896 6700 83936
rect 6740 83896 6741 83936
rect 6699 83887 6741 83896
rect 6700 83768 6740 83887
rect 6700 83719 6740 83728
rect 6219 83600 6261 83609
rect 6219 83560 6220 83600
rect 6260 83560 6261 83600
rect 6219 83551 6261 83560
rect 6220 83466 6260 83551
rect 6604 83432 6644 83441
rect 6412 83348 6452 83357
rect 6068 82972 6164 83012
rect 6316 83308 6412 83348
rect 6028 82963 6068 82972
rect 6220 82853 6260 82938
rect 6219 82844 6261 82853
rect 6219 82804 6220 82844
rect 6260 82804 6261 82844
rect 6219 82795 6261 82804
rect 6316 82676 6356 83308
rect 6412 83299 6452 83308
rect 6411 83180 6453 83189
rect 6411 83140 6412 83180
rect 6452 83140 6453 83180
rect 6411 83131 6453 83140
rect 6412 83012 6452 83131
rect 6412 82963 6452 82972
rect 6220 82636 6356 82676
rect 5931 82172 5973 82181
rect 5931 82132 5932 82172
rect 5972 82132 5973 82172
rect 5931 82123 5973 82132
rect 6220 82083 6260 82636
rect 6604 82256 6644 83392
rect 6699 83348 6741 83357
rect 6699 83308 6700 83348
rect 6740 83308 6741 83348
rect 6699 83299 6741 83308
rect 6700 82760 6740 83299
rect 6891 83012 6933 83021
rect 6891 82972 6892 83012
rect 6932 82972 6933 83012
rect 6891 82963 6933 82972
rect 6700 82711 6740 82720
rect 6795 82760 6837 82769
rect 6795 82720 6796 82760
rect 6836 82720 6837 82760
rect 6795 82711 6837 82720
rect 6796 82626 6836 82711
rect 6795 82424 6837 82433
rect 6795 82384 6796 82424
rect 6836 82384 6837 82424
rect 6795 82375 6837 82384
rect 6604 82181 6644 82216
rect 6220 82034 6260 82043
rect 6412 82172 6452 82181
rect 6412 81920 6452 82132
rect 6603 82172 6645 82181
rect 6603 82132 6604 82172
rect 6644 82132 6645 82172
rect 6603 82123 6645 82132
rect 6604 82092 6644 82123
rect 6699 82004 6741 82013
rect 6699 81964 6700 82004
rect 6740 81964 6741 82004
rect 6699 81955 6741 81964
rect 5548 81880 5684 81920
rect 5836 81880 5972 81920
rect 5355 81871 5397 81880
rect 5356 81500 5396 81871
rect 5356 81451 5396 81460
rect 5547 81332 5589 81341
rect 5547 81292 5548 81332
rect 5588 81292 5589 81332
rect 5547 81283 5589 81292
rect 5548 81198 5588 81283
rect 5451 81080 5493 81089
rect 5260 81040 5396 81080
rect 4779 80912 4821 80921
rect 4779 80872 4780 80912
rect 4820 80872 4821 80912
rect 4779 80863 4821 80872
rect 4928 80912 5296 80921
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 4928 80863 5296 80872
rect 4780 80753 4820 80863
rect 4779 80744 4821 80753
rect 5356 80744 5396 81040
rect 5451 81040 5452 81080
rect 5492 81040 5493 81080
rect 5451 81031 5493 81040
rect 4779 80704 4780 80744
rect 4820 80704 4821 80744
rect 4779 80695 4821 80704
rect 5260 80704 5396 80744
rect 4971 80576 5013 80585
rect 4971 80536 4972 80576
rect 5012 80536 5013 80576
rect 4971 80527 5013 80536
rect 4875 80492 4917 80501
rect 4875 80452 4876 80492
rect 4916 80452 4917 80492
rect 4875 80443 4917 80452
rect 4876 80358 4916 80443
rect 4779 80324 4821 80333
rect 4779 80284 4780 80324
rect 4820 80284 4821 80324
rect 4779 80275 4821 80284
rect 4780 79325 4820 80275
rect 4972 79577 5012 80527
rect 5163 80240 5205 80249
rect 5163 80200 5164 80240
rect 5204 80200 5205 80240
rect 5163 80191 5205 80200
rect 5164 79736 5204 80191
rect 5260 79904 5300 80704
rect 5356 80576 5396 80585
rect 5356 80081 5396 80536
rect 5452 80576 5492 81031
rect 5644 80669 5684 81880
rect 5739 81248 5781 81257
rect 5739 81208 5740 81248
rect 5780 81208 5876 81248
rect 5739 81199 5781 81208
rect 5740 81114 5780 81199
rect 5643 80660 5685 80669
rect 5643 80620 5644 80660
rect 5684 80620 5685 80660
rect 5643 80611 5685 80620
rect 5452 80527 5492 80536
rect 5739 80492 5781 80501
rect 5739 80452 5740 80492
rect 5780 80452 5781 80492
rect 5739 80443 5781 80452
rect 5740 80358 5780 80443
rect 5643 80240 5685 80249
rect 5643 80200 5644 80240
rect 5684 80200 5685 80240
rect 5643 80191 5685 80200
rect 5355 80072 5397 80081
rect 5355 80032 5356 80072
rect 5396 80032 5397 80072
rect 5355 80023 5397 80032
rect 5260 79864 5492 79904
rect 5260 79736 5300 79745
rect 5164 79696 5260 79736
rect 5260 79687 5300 79696
rect 5355 79652 5397 79661
rect 5355 79612 5356 79652
rect 5396 79612 5397 79652
rect 5355 79603 5397 79612
rect 4971 79568 5013 79577
rect 4971 79528 4972 79568
rect 5012 79528 5013 79568
rect 4971 79519 5013 79528
rect 4928 79400 5296 79409
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 4928 79351 5296 79360
rect 4779 79316 4821 79325
rect 4779 79276 4780 79316
rect 4820 79276 4821 79316
rect 4779 79267 4821 79276
rect 4971 79232 5013 79241
rect 5356 79232 5396 79603
rect 5452 79577 5492 79864
rect 5547 79820 5589 79829
rect 5547 79780 5548 79820
rect 5588 79780 5589 79820
rect 5547 79771 5589 79780
rect 5451 79568 5493 79577
rect 5451 79528 5452 79568
rect 5492 79528 5493 79568
rect 5451 79519 5493 79528
rect 5452 79434 5492 79519
rect 4971 79192 4972 79232
rect 5012 79192 5013 79232
rect 4971 79183 5013 79192
rect 5164 79192 5396 79232
rect 4684 79108 4820 79148
rect 4491 79064 4533 79073
rect 4052 78184 4148 78224
rect 4012 78175 4052 78184
rect 3436 78090 3476 78175
rect 3435 77972 3477 77981
rect 3435 77932 3436 77972
rect 3476 77932 3477 77972
rect 3435 77923 3477 77932
rect 3339 77216 3381 77225
rect 3339 77176 3340 77216
rect 3380 77176 3381 77216
rect 3339 77167 3381 77176
rect 3243 76880 3285 76889
rect 3243 76840 3244 76880
rect 3284 76840 3285 76880
rect 3243 76831 3285 76840
rect 3147 76796 3189 76805
rect 3147 76756 3148 76796
rect 3188 76756 3189 76796
rect 3147 76747 3189 76756
rect 3148 76662 3188 76747
rect 3243 76712 3285 76721
rect 3243 76672 3244 76712
rect 3284 76672 3285 76712
rect 3243 76663 3285 76672
rect 3051 76628 3093 76637
rect 3051 76588 3052 76628
rect 3092 76588 3093 76628
rect 3051 76579 3093 76588
rect 3244 76578 3284 76663
rect 3436 76040 3476 77923
rect 3723 77720 3765 77729
rect 3723 77680 3724 77720
rect 3764 77680 3765 77720
rect 3723 77671 3765 77680
rect 3724 77309 3764 77671
rect 3723 77300 3765 77309
rect 3723 77260 3724 77300
rect 3764 77260 3765 77300
rect 3723 77251 3765 77260
rect 3688 77132 4056 77141
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 3688 77083 4056 77092
rect 4108 76721 4148 78184
rect 4396 79024 4492 79064
rect 4532 79024 4533 79064
rect 4204 77561 4244 77646
rect 4203 77552 4245 77561
rect 4396 77552 4436 79024
rect 4491 79015 4533 79024
rect 4491 78812 4533 78821
rect 4684 78812 4724 78821
rect 4491 78772 4492 78812
rect 4532 78772 4533 78812
rect 4491 78763 4533 78772
rect 4588 78772 4684 78812
rect 4492 78238 4532 78763
rect 4492 78189 4532 78198
rect 4203 77512 4204 77552
rect 4244 77512 4436 77552
rect 4203 77503 4245 77512
rect 4588 77468 4628 78772
rect 4684 78763 4724 78772
rect 4683 78140 4725 78149
rect 4683 78100 4684 78140
rect 4724 78100 4725 78140
rect 4683 78091 4725 78100
rect 4684 78006 4724 78091
rect 4780 77720 4820 79108
rect 4972 79064 5012 79183
rect 4972 79015 5012 79024
rect 5067 78980 5109 78989
rect 5067 78940 5068 78980
rect 5108 78940 5109 78980
rect 5067 78931 5109 78940
rect 4875 78476 4917 78485
rect 4875 78436 4876 78476
rect 4916 78436 4917 78476
rect 4875 78427 4917 78436
rect 4876 78224 4916 78427
rect 4876 78175 4916 78184
rect 4971 78224 5013 78233
rect 4971 78184 4972 78224
rect 5012 78184 5013 78224
rect 4971 78175 5013 78184
rect 4972 78090 5012 78175
rect 5068 78149 5108 78931
rect 5067 78140 5109 78149
rect 5067 78100 5068 78140
rect 5108 78100 5109 78140
rect 5067 78091 5109 78100
rect 5164 78056 5204 79192
rect 5259 78560 5301 78569
rect 5259 78520 5260 78560
rect 5300 78520 5301 78560
rect 5259 78511 5301 78520
rect 5260 78056 5300 78511
rect 5356 78476 5396 78485
rect 5548 78476 5588 79771
rect 5644 79157 5684 80191
rect 5836 80081 5876 81208
rect 5932 80408 5972 81880
rect 6316 81880 6452 81920
rect 6028 80576 6068 80585
rect 6219 80576 6261 80585
rect 6068 80536 6164 80576
rect 6028 80527 6068 80536
rect 6028 80408 6068 80417
rect 5932 80368 6028 80408
rect 6028 80359 6068 80368
rect 5835 80072 5877 80081
rect 5835 80032 5836 80072
rect 5876 80032 5877 80072
rect 5835 80023 5877 80032
rect 5739 79904 5781 79913
rect 5739 79864 5740 79904
rect 5780 79864 5781 79904
rect 5739 79855 5781 79864
rect 5740 79736 5780 79855
rect 5740 79661 5780 79696
rect 5739 79652 5781 79661
rect 5739 79612 5740 79652
rect 5780 79612 5781 79652
rect 5739 79603 5781 79612
rect 5643 79148 5685 79157
rect 5643 79108 5644 79148
rect 5684 79108 5685 79148
rect 5643 79099 5685 79108
rect 5643 78728 5685 78737
rect 5643 78688 5644 78728
rect 5684 78688 5685 78728
rect 5643 78679 5685 78688
rect 5396 78436 5588 78476
rect 5356 78427 5396 78436
rect 5644 78392 5684 78679
rect 5452 78352 5684 78392
rect 5452 78224 5492 78352
rect 5260 78016 5396 78056
rect 5164 78007 5204 78016
rect 4928 77888 5296 77897
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 4928 77839 5296 77848
rect 4972 77720 5012 77729
rect 4780 77680 4972 77720
rect 4972 77671 5012 77680
rect 4875 77552 4917 77561
rect 4875 77512 4876 77552
rect 4916 77512 4917 77552
rect 4875 77503 4917 77512
rect 4300 77428 4628 77468
rect 4780 77468 4820 77477
rect 4300 77384 4340 77428
rect 4204 77344 4340 77384
rect 4204 76726 4244 77344
rect 4396 77300 4436 77309
rect 3723 76712 3765 76721
rect 3723 76672 3724 76712
rect 3764 76672 3765 76712
rect 3723 76663 3765 76672
rect 4107 76712 4149 76721
rect 4107 76672 4108 76712
rect 4148 76672 4149 76712
rect 4204 76677 4244 76686
rect 4300 77260 4396 77300
rect 4107 76663 4149 76672
rect 3724 76578 3764 76663
rect 4108 76049 4148 76663
rect 3052 75788 3092 75797
rect 2955 74444 2997 74453
rect 2955 74404 2956 74444
rect 2996 74404 2997 74444
rect 2955 74395 2997 74404
rect 2859 74192 2901 74201
rect 2859 74152 2860 74192
rect 2900 74152 2901 74192
rect 2859 74143 2901 74152
rect 2668 73688 2708 73699
rect 2668 73613 2708 73648
rect 2667 73604 2709 73613
rect 2667 73564 2668 73604
rect 2708 73564 2709 73604
rect 2667 73555 2709 73564
rect 2516 72976 2612 73016
rect 2476 72437 2516 72976
rect 2668 72932 2708 73555
rect 2572 72892 2708 72932
rect 2475 72428 2517 72437
rect 2475 72388 2476 72428
rect 2516 72388 2517 72428
rect 2475 72379 2517 72388
rect 2476 71000 2516 72379
rect 2572 71765 2612 72892
rect 2668 72764 2708 72773
rect 2708 72724 2804 72764
rect 2668 72715 2708 72724
rect 2571 71756 2613 71765
rect 2571 71716 2572 71756
rect 2612 71716 2613 71756
rect 2571 71707 2613 71716
rect 2571 71588 2613 71597
rect 2571 71548 2572 71588
rect 2612 71548 2613 71588
rect 2571 71539 2613 71548
rect 2572 71504 2612 71539
rect 2572 71453 2612 71464
rect 2476 70960 2612 71000
rect 2475 70832 2517 70841
rect 2475 70792 2476 70832
rect 2516 70792 2517 70832
rect 2475 70783 2517 70792
rect 2379 70664 2421 70673
rect 2379 70624 2380 70664
rect 2420 70624 2421 70664
rect 2379 70615 2421 70624
rect 2476 70664 2516 70783
rect 2476 70615 2516 70624
rect 2379 70496 2421 70505
rect 2572 70496 2612 70960
rect 2379 70456 2380 70496
rect 2420 70456 2421 70496
rect 2379 70447 2421 70456
rect 2476 70456 2612 70496
rect 2667 70496 2709 70505
rect 2667 70456 2668 70496
rect 2708 70456 2709 70496
rect 2284 67733 2324 68440
rect 2283 67724 2325 67733
rect 2283 67684 2284 67724
rect 2324 67684 2325 67724
rect 2283 67675 2325 67684
rect 2380 66968 2420 70447
rect 2476 69992 2516 70456
rect 2667 70447 2709 70456
rect 2668 70362 2708 70447
rect 2476 69943 2516 69952
rect 2764 69908 2804 72724
rect 2860 72353 2900 74143
rect 2955 72428 2997 72437
rect 2955 72388 2956 72428
rect 2996 72388 2997 72428
rect 2955 72379 2997 72388
rect 2859 72344 2901 72353
rect 2859 72304 2860 72344
rect 2900 72304 2901 72344
rect 2859 72295 2901 72304
rect 2956 72176 2996 72379
rect 2956 72127 2996 72136
rect 2955 71756 2997 71765
rect 2955 71716 2956 71756
rect 2996 71716 2997 71756
rect 2955 71707 2997 71716
rect 2572 69868 2804 69908
rect 2475 69236 2517 69245
rect 2475 69196 2476 69236
rect 2516 69196 2517 69236
rect 2475 69187 2517 69196
rect 2476 69152 2516 69187
rect 2476 69101 2516 69112
rect 2572 68489 2612 69868
rect 2668 69740 2708 69749
rect 2668 69161 2708 69700
rect 2667 69152 2709 69161
rect 2667 69112 2668 69152
rect 2708 69112 2709 69152
rect 2667 69103 2709 69112
rect 2860 69152 2900 69161
rect 2668 68984 2708 68993
rect 2571 68480 2613 68489
rect 2571 68440 2572 68480
rect 2612 68440 2613 68480
rect 2571 68431 2613 68440
rect 2668 68237 2708 68944
rect 2860 68732 2900 69112
rect 2956 68909 2996 71707
rect 3052 71499 3092 75748
rect 3244 75788 3284 75797
rect 3284 75748 3380 75788
rect 3244 75739 3284 75748
rect 3148 75200 3188 75209
rect 3148 74957 3188 75160
rect 3243 75200 3285 75209
rect 3243 75160 3244 75200
rect 3284 75160 3285 75200
rect 3243 75151 3285 75160
rect 3244 75066 3284 75151
rect 3147 74948 3189 74957
rect 3147 74908 3148 74948
rect 3188 74908 3189 74948
rect 3147 74899 3189 74908
rect 3147 74780 3189 74789
rect 3147 74740 3148 74780
rect 3188 74740 3189 74780
rect 3147 74731 3189 74740
rect 3148 74528 3188 74731
rect 3148 74453 3188 74488
rect 3340 74518 3380 75748
rect 3436 75041 3476 76000
rect 4107 76040 4149 76049
rect 4107 76000 4108 76040
rect 4148 76000 4149 76040
rect 4107 75991 4149 76000
rect 3688 75620 4056 75629
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 3688 75571 4056 75580
rect 4107 75284 4149 75293
rect 4300 75284 4340 77260
rect 4396 77251 4436 77260
rect 4588 77300 4628 77311
rect 4588 77225 4628 77260
rect 4587 77216 4629 77225
rect 4587 77176 4588 77216
rect 4628 77176 4629 77216
rect 4587 77167 4629 77176
rect 4780 77057 4820 77428
rect 4779 77048 4821 77057
rect 4779 77008 4780 77048
rect 4820 77008 4821 77048
rect 4779 76999 4821 77008
rect 4395 76964 4437 76973
rect 4395 76924 4396 76964
rect 4436 76924 4437 76964
rect 4395 76915 4437 76924
rect 4396 76628 4436 76915
rect 4587 76880 4629 76889
rect 4587 76840 4588 76880
rect 4628 76840 4629 76880
rect 4587 76831 4629 76840
rect 4588 76746 4628 76831
rect 4779 76796 4821 76805
rect 4779 76756 4780 76796
rect 4820 76756 4821 76796
rect 4779 76747 4821 76756
rect 4780 76662 4820 76747
rect 4396 76579 4436 76588
rect 4587 76544 4629 76553
rect 4876 76544 4916 77503
rect 5163 77468 5205 77477
rect 5163 77428 5164 77468
rect 5204 77428 5205 77468
rect 5163 77419 5205 77428
rect 5164 77334 5204 77419
rect 5068 76712 5108 76721
rect 5356 76712 5396 78016
rect 5108 76672 5396 76712
rect 5068 76663 5108 76672
rect 4587 76504 4588 76544
rect 4628 76504 4629 76544
rect 4587 76495 4629 76504
rect 4780 76504 4916 76544
rect 4395 76292 4437 76301
rect 4395 76252 4396 76292
rect 4436 76252 4437 76292
rect 4395 76243 4437 76252
rect 4107 75244 4108 75284
rect 4148 75244 4149 75284
rect 4107 75235 4149 75244
rect 4252 75244 4340 75284
rect 4252 75242 4292 75244
rect 3627 75200 3669 75209
rect 3627 75160 3628 75200
rect 3668 75160 3669 75200
rect 3627 75151 3669 75160
rect 3724 75200 3764 75211
rect 3435 75032 3477 75041
rect 3435 74992 3436 75032
rect 3476 74992 3477 75032
rect 3435 74983 3477 74992
rect 3340 74478 3572 74518
rect 3147 74444 3189 74453
rect 3147 74404 3148 74444
rect 3188 74404 3189 74444
rect 3147 74395 3189 74404
rect 3340 74285 3380 74370
rect 3339 74276 3381 74285
rect 3339 74236 3340 74276
rect 3380 74236 3381 74276
rect 3339 74227 3381 74236
rect 3532 73865 3572 74478
rect 3628 74285 3668 75151
rect 3724 75125 3764 75160
rect 3723 75116 3765 75125
rect 3723 75076 3724 75116
rect 3764 75076 3765 75116
rect 3723 75067 3765 75076
rect 4108 74360 4148 75235
rect 4252 75193 4292 75202
rect 4396 75116 4436 76243
rect 4588 76040 4628 76495
rect 4684 76040 4724 76049
rect 4588 76000 4684 76040
rect 4588 75797 4628 76000
rect 4684 75991 4724 76000
rect 4587 75788 4629 75797
rect 4587 75748 4588 75788
rect 4628 75748 4629 75788
rect 4587 75739 4629 75748
rect 4587 75284 4629 75293
rect 4587 75244 4588 75284
rect 4628 75244 4629 75284
rect 4587 75235 4629 75244
rect 4491 75200 4533 75209
rect 4491 75160 4492 75200
rect 4532 75160 4533 75200
rect 4491 75151 4533 75160
rect 4588 75200 4628 75235
rect 4396 75067 4436 75076
rect 4492 74873 4532 75151
rect 4588 75149 4628 75160
rect 4780 75032 4820 76504
rect 4928 76376 5296 76385
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 4928 76327 5296 76336
rect 4971 76124 5013 76133
rect 4971 76084 4972 76124
rect 5012 76084 5013 76124
rect 4971 76075 5013 76084
rect 4875 76040 4917 76049
rect 4875 76000 4876 76040
rect 4916 76000 4917 76040
rect 4875 75991 4917 76000
rect 4972 76040 5012 76075
rect 4876 75293 4916 75991
rect 4972 75881 5012 76000
rect 4971 75872 5013 75881
rect 4971 75832 4972 75872
rect 5012 75832 5013 75872
rect 4971 75823 5013 75832
rect 4875 75284 4917 75293
rect 4875 75244 4876 75284
rect 4916 75244 4917 75284
rect 4875 75235 4917 75244
rect 4876 75041 4916 75235
rect 5452 75125 5492 78184
rect 5643 78224 5685 78233
rect 5643 78184 5644 78224
rect 5684 78184 5685 78224
rect 5643 78175 5685 78184
rect 5547 78140 5589 78149
rect 5547 78100 5548 78140
rect 5588 78100 5589 78140
rect 5547 78091 5589 78100
rect 5451 75116 5493 75125
rect 5451 75076 5452 75116
rect 5492 75076 5493 75116
rect 5451 75067 5493 75076
rect 4588 74992 4820 75032
rect 4875 75032 4917 75041
rect 4875 74992 4876 75032
rect 4916 74992 4917 75032
rect 4491 74864 4533 74873
rect 4491 74824 4492 74864
rect 4532 74824 4533 74864
rect 4491 74815 4533 74824
rect 4204 74528 4244 74537
rect 4204 74444 4244 74488
rect 4299 74444 4341 74453
rect 4204 74404 4300 74444
rect 4340 74404 4341 74444
rect 4299 74395 4341 74404
rect 4492 74360 4532 74815
rect 4108 74320 4244 74360
rect 3627 74276 3669 74285
rect 3627 74236 3628 74276
rect 3668 74236 3669 74276
rect 3627 74227 3669 74236
rect 4012 74276 4052 74285
rect 4052 74236 4148 74276
rect 4012 74227 4052 74236
rect 3688 74108 4056 74117
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 3688 74059 4056 74068
rect 3147 73856 3189 73865
rect 3147 73816 3148 73856
rect 3188 73816 3189 73856
rect 3147 73807 3189 73816
rect 3531 73856 3573 73865
rect 3531 73816 3532 73856
rect 3572 73816 3573 73856
rect 3531 73807 3573 73816
rect 3148 73702 3188 73807
rect 3148 73653 3188 73662
rect 3531 73688 3573 73697
rect 4108 73688 4148 74236
rect 3531 73648 3532 73688
rect 3572 73648 3573 73688
rect 3531 73639 3573 73648
rect 3820 73648 4148 73688
rect 3532 73554 3572 73639
rect 3340 73478 3380 73487
rect 3339 73438 3340 73445
rect 3380 73438 3381 73445
rect 3339 73436 3381 73438
rect 3339 73396 3340 73436
rect 3380 73396 3381 73436
rect 3339 73387 3381 73396
rect 3340 73343 3380 73387
rect 3339 73268 3381 73277
rect 3339 73228 3340 73268
rect 3380 73228 3381 73268
rect 3339 73219 3381 73228
rect 3052 71450 3092 71459
rect 3148 72008 3188 72017
rect 3148 70832 3188 71968
rect 3243 71840 3285 71849
rect 3243 71800 3244 71840
rect 3284 71800 3285 71840
rect 3243 71791 3285 71800
rect 3244 71672 3284 71791
rect 3340 71765 3380 73219
rect 3628 73100 3668 73140
rect 3628 73025 3668 73060
rect 3627 73016 3669 73025
rect 3627 72976 3628 73016
rect 3668 72976 3669 73016
rect 3627 72967 3669 72976
rect 3820 73011 3860 73648
rect 3628 72965 3668 72967
rect 3820 72962 3860 72971
rect 3688 72596 4056 72605
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 3688 72547 4056 72556
rect 3435 72344 3477 72353
rect 3435 72304 3436 72344
rect 3476 72304 3477 72344
rect 3435 72295 3477 72304
rect 4011 72344 4053 72353
rect 4011 72304 4012 72344
rect 4052 72304 4053 72344
rect 4011 72295 4053 72304
rect 3339 71756 3381 71765
rect 3339 71716 3340 71756
rect 3380 71716 3381 71756
rect 3339 71707 3381 71716
rect 3244 71623 3284 71632
rect 3339 71588 3381 71597
rect 3339 71548 3340 71588
rect 3380 71548 3381 71588
rect 3339 71539 3381 71548
rect 3148 70792 3284 70832
rect 3051 70664 3093 70673
rect 3051 70624 3052 70664
rect 3092 70624 3093 70664
rect 3051 70615 3093 70624
rect 3148 70664 3188 70675
rect 3052 70412 3092 70615
rect 3148 70589 3188 70624
rect 3147 70580 3189 70589
rect 3147 70540 3148 70580
rect 3188 70540 3189 70580
rect 3147 70531 3189 70540
rect 3148 70500 3188 70531
rect 3052 70372 3188 70412
rect 3051 69236 3093 69245
rect 3051 69196 3052 69236
rect 3092 69196 3093 69236
rect 3051 69187 3093 69196
rect 2955 68900 2997 68909
rect 2955 68860 2956 68900
rect 2996 68860 2997 68900
rect 2955 68851 2997 68860
rect 2860 68692 2996 68732
rect 2763 68480 2805 68489
rect 2763 68440 2764 68480
rect 2804 68440 2805 68480
rect 2763 68431 2805 68440
rect 2764 68346 2804 68431
rect 2667 68228 2709 68237
rect 2667 68188 2668 68228
rect 2708 68188 2709 68228
rect 2667 68179 2709 68188
rect 2956 67229 2996 68692
rect 3052 67640 3092 69187
rect 3052 67591 3092 67600
rect 2955 67220 2997 67229
rect 2955 67180 2956 67220
rect 2996 67180 2997 67220
rect 2955 67171 2997 67180
rect 2476 66968 2516 66977
rect 2380 66928 2476 66968
rect 2476 66919 2516 66928
rect 2572 66968 2612 66977
rect 2379 66548 2421 66557
rect 2379 66508 2380 66548
rect 2420 66508 2421 66548
rect 2379 66499 2421 66508
rect 2187 64952 2229 64961
rect 2187 64912 2188 64952
rect 2228 64912 2229 64952
rect 2187 64903 2229 64912
rect 2092 64567 2132 64576
rect 2188 64616 2228 64625
rect 1995 64028 2037 64037
rect 1995 63988 1996 64028
rect 2036 63988 2037 64028
rect 1995 63979 2037 63988
rect 1899 63272 1941 63281
rect 1899 63232 1900 63272
rect 1940 63232 1941 63272
rect 1899 63223 1941 63232
rect 1900 63138 1940 63223
rect 1708 61888 1844 61928
rect 1708 61844 1748 61888
rect 1697 61804 1748 61844
rect 1697 61760 1737 61804
rect 1697 61720 1748 61760
rect 1708 61508 1748 61720
rect 1697 61468 1748 61508
rect 1697 61340 1737 61468
rect 1697 61300 1748 61340
rect 1708 61004 1748 61300
rect 1708 60964 1844 61004
rect 1611 60920 1653 60929
rect 1611 60880 1612 60920
rect 1652 60880 1653 60920
rect 1611 60871 1653 60880
rect 1323 60836 1365 60845
rect 1323 60796 1324 60836
rect 1364 60796 1365 60836
rect 1323 60787 1365 60796
rect 1228 59408 1268 59417
rect 1324 59408 1364 60787
rect 1516 60668 1556 60677
rect 1268 59368 1364 59408
rect 1420 60628 1516 60668
rect 1228 59359 1268 59368
rect 1420 58988 1460 60628
rect 1516 60619 1556 60628
rect 1516 60080 1556 60089
rect 1612 60080 1652 60871
rect 1708 60836 1748 60845
rect 1708 60593 1748 60796
rect 1707 60584 1749 60593
rect 1707 60544 1708 60584
rect 1748 60544 1749 60584
rect 1707 60535 1749 60544
rect 1556 60040 1652 60080
rect 1516 60031 1556 60040
rect 1420 58948 1556 58988
rect 1419 58820 1461 58829
rect 1419 58780 1420 58820
rect 1460 58780 1461 58820
rect 1419 58771 1461 58780
rect 1323 58568 1365 58577
rect 1323 58528 1324 58568
rect 1364 58528 1365 58568
rect 1323 58519 1365 58528
rect 1420 58568 1460 58771
rect 1420 58519 1460 58528
rect 1324 57728 1364 58519
rect 1516 57980 1556 58948
rect 1324 57679 1364 57688
rect 1420 57940 1556 57980
rect 1420 57569 1460 57940
rect 1708 57896 1748 57905
rect 1515 57812 1557 57821
rect 1515 57772 1516 57812
rect 1556 57772 1557 57812
rect 1515 57763 1557 57772
rect 1516 57678 1556 57763
rect 1419 57560 1461 57569
rect 1419 57520 1420 57560
rect 1460 57520 1461 57560
rect 1419 57511 1461 57520
rect 1708 57317 1748 57856
rect 1707 57308 1749 57317
rect 1707 57268 1708 57308
rect 1748 57268 1749 57308
rect 1707 57259 1749 57268
rect 1227 57224 1269 57233
rect 1227 57184 1228 57224
rect 1268 57184 1269 57224
rect 1227 57175 1269 57184
rect 1228 56552 1268 57175
rect 1707 57140 1749 57149
rect 1707 57100 1708 57140
rect 1748 57100 1749 57140
rect 1707 57091 1749 57100
rect 1708 57006 1748 57091
rect 1228 56503 1268 56512
rect 1516 56888 1556 56897
rect 1420 56300 1460 56309
rect 1323 56048 1365 56057
rect 1323 56008 1324 56048
rect 1364 56008 1365 56048
rect 1323 55999 1365 56008
rect 1228 55544 1268 55553
rect 1324 55544 1364 55999
rect 1268 55504 1364 55544
rect 1228 55495 1268 55504
rect 1323 55040 1365 55049
rect 1323 55000 1324 55040
rect 1364 55000 1365 55040
rect 1323 54991 1365 55000
rect 1324 53276 1364 54991
rect 1420 54041 1460 56260
rect 1516 55469 1556 56848
rect 1707 56804 1749 56813
rect 1707 56764 1708 56804
rect 1748 56764 1749 56804
rect 1707 56755 1749 56764
rect 1612 56384 1652 56393
rect 1515 55460 1557 55469
rect 1515 55420 1516 55460
rect 1556 55420 1557 55460
rect 1515 55411 1557 55420
rect 1612 55217 1652 56344
rect 1611 55208 1653 55217
rect 1611 55168 1612 55208
rect 1652 55168 1653 55208
rect 1611 55159 1653 55168
rect 1708 54788 1748 56755
rect 1708 54739 1748 54748
rect 1804 54713 1844 60964
rect 1899 60920 1941 60929
rect 1899 60880 1900 60920
rect 1940 60880 1941 60920
rect 1899 60871 1941 60880
rect 1900 60786 1940 60871
rect 1899 56888 1941 56897
rect 1899 56848 1900 56888
rect 1940 56848 1941 56888
rect 1899 56839 1941 56848
rect 1900 56754 1940 56839
rect 1996 56057 2036 63979
rect 2092 63188 2132 63197
rect 2092 60425 2132 63148
rect 2188 62861 2228 64576
rect 2284 63272 2324 63281
rect 2284 63029 2324 63232
rect 2283 63020 2325 63029
rect 2283 62980 2284 63020
rect 2324 62980 2325 63020
rect 2283 62971 2325 62980
rect 2187 62852 2229 62861
rect 2187 62812 2188 62852
rect 2228 62812 2229 62852
rect 2187 62803 2229 62812
rect 2091 60416 2133 60425
rect 2091 60376 2092 60416
rect 2132 60376 2133 60416
rect 2091 60367 2133 60376
rect 2380 59156 2420 66499
rect 2572 65465 2612 66928
rect 3052 66968 3092 66977
rect 3148 66968 3188 70372
rect 3244 68475 3284 70792
rect 3340 68489 3380 71539
rect 3436 69992 3476 72295
rect 3531 71756 3573 71765
rect 3531 71716 3532 71756
rect 3572 71716 3573 71756
rect 3531 71707 3573 71716
rect 3532 71177 3572 71707
rect 4012 71261 4052 72295
rect 4011 71252 4053 71261
rect 4011 71212 4012 71252
rect 4052 71212 4053 71252
rect 4011 71203 4053 71212
rect 3531 71168 3573 71177
rect 3531 71128 3532 71168
rect 3572 71128 3573 71168
rect 3531 71119 3573 71128
rect 3532 70673 3572 71119
rect 3688 71084 4056 71093
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 3688 71035 4056 71044
rect 3531 70664 3573 70673
rect 3531 70624 3532 70664
rect 3572 70624 3573 70664
rect 3531 70615 3573 70624
rect 4204 70505 4244 74320
rect 4396 74320 4532 74360
rect 4300 73016 4340 73025
rect 4300 72353 4340 72976
rect 4299 72344 4341 72353
rect 4299 72304 4300 72344
rect 4340 72304 4341 72344
rect 4299 72295 4341 72304
rect 4299 72176 4341 72185
rect 4299 72136 4300 72176
rect 4340 72136 4341 72176
rect 4299 72127 4341 72136
rect 4300 72042 4340 72127
rect 4396 71765 4436 74320
rect 4588 73100 4628 74992
rect 4875 74983 4917 74992
rect 4928 74864 5296 74873
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 4928 74815 5296 74824
rect 5452 74528 5492 74537
rect 5548 74528 5588 78091
rect 5492 74488 5588 74528
rect 5452 74479 5492 74488
rect 5355 74444 5397 74453
rect 5355 74404 5356 74444
rect 5396 74404 5397 74444
rect 5355 74395 5397 74404
rect 4779 73856 4821 73865
rect 4779 73816 4780 73856
rect 4820 73816 4821 73856
rect 4779 73807 4821 73816
rect 4780 73688 4820 73807
rect 5356 73781 5396 74395
rect 5355 73772 5397 73781
rect 5355 73732 5356 73772
rect 5396 73732 5397 73772
rect 5355 73723 5397 73732
rect 4780 73639 4820 73648
rect 5356 73688 5396 73723
rect 5356 73639 5396 73648
rect 4972 73520 5012 73529
rect 4492 73060 4628 73100
rect 4684 73480 4972 73520
rect 4395 71756 4437 71765
rect 4395 71716 4396 71756
rect 4436 71716 4437 71756
rect 4395 71707 4437 71716
rect 4299 71504 4341 71513
rect 4299 71464 4300 71504
rect 4340 71464 4341 71504
rect 4299 71455 4341 71464
rect 4396 71504 4436 71513
rect 4300 71370 4340 71455
rect 4299 71252 4341 71261
rect 4299 71212 4300 71252
rect 4340 71212 4341 71252
rect 4299 71203 4341 71212
rect 4300 70589 4340 71203
rect 4396 70925 4436 71464
rect 4395 70916 4437 70925
rect 4395 70876 4396 70916
rect 4436 70876 4437 70916
rect 4395 70867 4437 70876
rect 4492 70841 4532 73060
rect 4587 71756 4629 71765
rect 4587 71716 4588 71756
rect 4628 71716 4629 71756
rect 4587 71707 4629 71716
rect 4491 70832 4533 70841
rect 4491 70792 4492 70832
rect 4532 70792 4533 70832
rect 4491 70783 4533 70792
rect 4395 70748 4437 70757
rect 4395 70708 4396 70748
rect 4436 70708 4437 70748
rect 4395 70699 4437 70708
rect 4396 70664 4436 70699
rect 4588 70664 4628 71707
rect 4684 71513 4724 73480
rect 4972 73471 5012 73480
rect 5164 73520 5204 73529
rect 5204 73480 5396 73520
rect 5164 73471 5204 73480
rect 4928 73352 5296 73361
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 4928 73303 5296 73312
rect 4876 73025 4916 73056
rect 4875 73016 4917 73025
rect 4875 72976 4876 73016
rect 4916 72976 4917 73016
rect 4875 72967 4917 72976
rect 5260 73016 5300 73025
rect 4780 72932 4820 72943
rect 4780 72857 4820 72892
rect 4876 72932 4916 72967
rect 4779 72848 4821 72857
rect 4779 72808 4780 72848
rect 4820 72808 4821 72848
rect 4779 72799 4821 72808
rect 4876 72101 4916 72892
rect 5260 72773 5300 72976
rect 5356 73016 5396 73480
rect 5548 73352 5588 74488
rect 5644 74117 5684 78175
rect 5740 77561 5780 79603
rect 5739 77552 5781 77561
rect 5739 77512 5740 77552
rect 5780 77512 5781 77552
rect 5739 77503 5781 77512
rect 5836 77384 5876 80023
rect 5931 79820 5973 79829
rect 5931 79780 5932 79820
rect 5972 79780 5973 79820
rect 5931 79771 5973 79780
rect 5740 77344 5876 77384
rect 5643 74108 5685 74117
rect 5643 74068 5644 74108
rect 5684 74068 5685 74108
rect 5643 74059 5685 74068
rect 5643 73856 5685 73865
rect 5643 73816 5644 73856
rect 5684 73816 5685 73856
rect 5643 73807 5685 73816
rect 5356 72967 5396 72976
rect 5452 73312 5588 73352
rect 5259 72764 5301 72773
rect 5259 72724 5260 72764
rect 5300 72724 5301 72764
rect 5259 72715 5301 72724
rect 4875 72092 4917 72101
rect 4875 72052 4876 72092
rect 4916 72052 4917 72092
rect 4875 72043 4917 72052
rect 5260 72017 5300 72715
rect 5452 72185 5492 73312
rect 5644 73277 5684 73807
rect 5643 73268 5685 73277
rect 5548 73228 5644 73268
rect 5684 73228 5685 73268
rect 5451 72176 5493 72185
rect 5451 72136 5452 72176
rect 5492 72136 5493 72176
rect 5451 72127 5493 72136
rect 5548 72176 5588 73228
rect 5643 73219 5685 73228
rect 5643 73100 5685 73109
rect 5643 73060 5644 73100
rect 5684 73060 5685 73100
rect 5643 73051 5685 73060
rect 5259 72008 5301 72017
rect 5259 71968 5260 72008
rect 5300 71968 5301 72008
rect 5259 71959 5301 71968
rect 4928 71840 5296 71849
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 4928 71791 5296 71800
rect 5355 71756 5397 71765
rect 5355 71716 5356 71756
rect 5396 71716 5397 71756
rect 5355 71707 5397 71716
rect 4683 71504 4725 71513
rect 4683 71464 4684 71504
rect 4724 71464 4725 71504
rect 4683 71455 4725 71464
rect 5356 71504 5396 71707
rect 5356 71455 5396 71464
rect 4780 71420 4820 71429
rect 4780 70841 4820 71380
rect 4876 71420 4916 71431
rect 4876 71345 4916 71380
rect 4875 71336 4917 71345
rect 4875 71296 4876 71336
rect 4916 71296 4917 71336
rect 4875 71287 4917 71296
rect 5355 71336 5397 71345
rect 5355 71296 5356 71336
rect 5396 71296 5397 71336
rect 5355 71287 5397 71296
rect 4779 70832 4821 70841
rect 4779 70792 4780 70832
rect 4820 70792 4821 70832
rect 4779 70783 4821 70792
rect 4299 70580 4341 70589
rect 4299 70540 4300 70580
rect 4340 70540 4341 70580
rect 4299 70531 4341 70540
rect 4203 70496 4245 70505
rect 4203 70456 4204 70496
rect 4244 70456 4245 70496
rect 4203 70447 4245 70456
rect 3916 70036 4148 70076
rect 3436 69943 3476 69952
rect 3532 69992 3572 70001
rect 3435 68564 3477 68573
rect 3435 68524 3436 68564
rect 3476 68524 3477 68564
rect 3435 68515 3477 68524
rect 3244 68426 3284 68435
rect 3339 68480 3381 68489
rect 3339 68440 3340 68480
rect 3380 68440 3381 68480
rect 3339 68431 3381 68440
rect 3436 68430 3476 68515
rect 3092 66928 3188 66968
rect 3244 67472 3284 67481
rect 3052 66919 3092 66928
rect 2956 66884 2996 66893
rect 2956 66212 2996 66844
rect 2956 66172 3188 66212
rect 2668 66128 2708 66137
rect 2571 65456 2613 65465
rect 2571 65416 2572 65456
rect 2612 65416 2613 65456
rect 2571 65407 2613 65416
rect 2668 65204 2708 66088
rect 2860 65960 2900 65969
rect 2900 65920 3092 65960
rect 2860 65911 2900 65920
rect 2859 65624 2901 65633
rect 2859 65584 2860 65624
rect 2900 65584 2901 65624
rect 2859 65575 2901 65584
rect 2860 65456 2900 65575
rect 2860 65407 2900 65416
rect 2955 65456 2997 65465
rect 2955 65416 2956 65456
rect 2996 65416 2997 65456
rect 2955 65407 2997 65416
rect 2668 65164 2804 65204
rect 2667 64700 2709 64709
rect 2667 64660 2668 64700
rect 2708 64660 2709 64700
rect 2667 64651 2709 64660
rect 2572 64616 2612 64625
rect 2572 63953 2612 64576
rect 2668 64566 2708 64651
rect 2764 64280 2804 65164
rect 2668 64240 2804 64280
rect 2668 64037 2708 64240
rect 2667 64028 2709 64037
rect 2667 63988 2668 64028
rect 2708 63988 2709 64028
rect 2667 63979 2709 63988
rect 2571 63944 2613 63953
rect 2571 63904 2572 63944
rect 2612 63904 2613 63944
rect 2571 63895 2613 63904
rect 2668 63944 2708 63979
rect 2476 63188 2516 63197
rect 2476 62609 2516 63148
rect 2571 63188 2613 63197
rect 2571 63148 2572 63188
rect 2612 63148 2613 63188
rect 2668 63188 2708 63904
rect 2860 63692 2900 63701
rect 2860 63281 2900 63652
rect 2859 63272 2901 63281
rect 2859 63232 2860 63272
rect 2900 63232 2901 63272
rect 2859 63223 2901 63232
rect 2668 63148 2804 63188
rect 2571 63139 2613 63148
rect 2572 62684 2612 63139
rect 2764 63104 2804 63148
rect 2860 63104 2900 63113
rect 2764 63064 2860 63104
rect 2860 63055 2900 63064
rect 2667 63020 2709 63029
rect 2667 62980 2668 63020
rect 2708 62980 2709 63020
rect 2667 62971 2709 62980
rect 2668 62886 2708 62971
rect 2956 62693 2996 65407
rect 2955 62684 2997 62693
rect 2572 62644 2900 62684
rect 2475 62600 2517 62609
rect 2475 62560 2476 62600
rect 2516 62560 2517 62600
rect 2475 62551 2517 62560
rect 2572 62432 2612 62443
rect 2572 62357 2612 62392
rect 2571 62348 2613 62357
rect 2571 62308 2572 62348
rect 2612 62308 2613 62348
rect 2571 62299 2613 62308
rect 2763 62180 2805 62189
rect 2763 62140 2764 62180
rect 2804 62140 2805 62180
rect 2763 62131 2805 62140
rect 2764 62046 2804 62131
rect 2572 61592 2612 61601
rect 2612 61552 2708 61592
rect 2572 61543 2612 61552
rect 2668 60080 2708 61552
rect 2860 61508 2900 62644
rect 2955 62644 2956 62684
rect 2996 62644 2997 62684
rect 2955 62635 2997 62644
rect 3052 62525 3092 65920
rect 3148 65297 3188 66172
rect 3147 65288 3189 65297
rect 3147 65248 3148 65288
rect 3188 65248 3189 65288
rect 3147 65239 3189 65248
rect 3244 65204 3284 67432
rect 3532 67136 3572 69952
rect 3916 69992 3956 70036
rect 3916 69943 3956 69952
rect 4011 69908 4053 69917
rect 4011 69868 4012 69908
rect 4052 69868 4053 69908
rect 4011 69859 4053 69868
rect 4012 69774 4052 69859
rect 3688 69572 4056 69581
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 3688 69523 4056 69532
rect 4108 69413 4148 70036
rect 4107 69404 4149 69413
rect 4107 69364 4108 69404
rect 4148 69364 4149 69404
rect 4107 69355 4149 69364
rect 4107 69236 4149 69245
rect 4107 69196 4108 69236
rect 4148 69196 4149 69236
rect 4107 69187 4149 69196
rect 4108 69152 4148 69187
rect 4108 69101 4148 69112
rect 4107 68984 4149 68993
rect 4107 68944 4108 68984
rect 4148 68944 4149 68984
rect 4107 68935 4149 68944
rect 3688 68060 4056 68069
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 3688 68011 4056 68020
rect 3436 67096 3572 67136
rect 3339 66128 3381 66137
rect 3339 66088 3340 66128
rect 3380 66088 3381 66128
rect 3339 66079 3381 66088
rect 3340 65994 3380 66079
rect 3436 65624 3476 67096
rect 3532 66968 3572 66977
rect 4108 66968 4148 68935
rect 4204 68909 4244 70447
rect 4396 69572 4436 70624
rect 4492 70624 4628 70664
rect 4780 70706 4820 70715
rect 4780 70664 4820 70666
rect 4875 70664 4917 70673
rect 4780 70624 4876 70664
rect 4916 70624 4917 70664
rect 4492 70328 4532 70624
rect 4875 70615 4917 70624
rect 4588 70496 4628 70505
rect 4628 70456 4724 70496
rect 4588 70447 4628 70456
rect 4492 70288 4628 70328
rect 4491 70076 4533 70085
rect 4491 70036 4492 70076
rect 4532 70036 4533 70076
rect 4588 70076 4628 70288
rect 4684 70160 4724 70456
rect 4928 70328 5296 70337
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 4928 70279 5296 70288
rect 5163 70160 5205 70169
rect 4684 70120 5012 70160
rect 4588 70036 4820 70076
rect 4491 70027 4533 70036
rect 4492 69992 4532 70027
rect 4492 69941 4532 69952
rect 4396 69532 4532 69572
rect 4395 69404 4437 69413
rect 4395 69364 4396 69404
rect 4436 69364 4437 69404
rect 4395 69355 4437 69364
rect 4300 68993 4340 69078
rect 4299 68984 4341 68993
rect 4299 68944 4300 68984
rect 4340 68944 4341 68984
rect 4299 68935 4341 68944
rect 4203 68900 4245 68909
rect 4203 68860 4204 68900
rect 4244 68860 4245 68900
rect 4203 68851 4245 68860
rect 4203 67136 4245 67145
rect 4203 67096 4204 67136
rect 4244 67096 4245 67136
rect 4203 67087 4245 67096
rect 4204 67002 4244 67087
rect 3532 66809 3572 66928
rect 4060 66958 4148 66968
rect 4100 66928 4148 66958
rect 4060 66909 4100 66918
rect 3531 66800 3573 66809
rect 3531 66760 3532 66800
rect 3572 66760 3573 66800
rect 3531 66751 3573 66760
rect 4107 66800 4149 66809
rect 4107 66760 4108 66800
rect 4148 66760 4149 66800
rect 4107 66751 4149 66760
rect 3688 66548 4056 66557
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 3688 66499 4056 66508
rect 3436 65584 3572 65624
rect 3340 65381 3380 65466
rect 3435 65456 3477 65465
rect 3435 65416 3436 65456
rect 3476 65416 3477 65456
rect 3435 65407 3477 65416
rect 3339 65372 3381 65381
rect 3339 65332 3340 65372
rect 3380 65332 3381 65372
rect 3339 65323 3381 65332
rect 3436 65322 3476 65407
rect 3532 65381 3572 65584
rect 3916 65456 3956 65465
rect 4108 65456 4148 66751
rect 4203 66128 4245 66137
rect 4203 66088 4204 66128
rect 4244 66088 4245 66128
rect 4203 66079 4245 66088
rect 3956 65416 4148 65456
rect 3916 65407 3956 65416
rect 3531 65372 3573 65381
rect 3531 65332 3532 65372
rect 3572 65332 3573 65372
rect 3531 65323 3573 65332
rect 3532 65204 3572 65323
rect 3244 65164 3380 65204
rect 3243 64952 3285 64961
rect 3243 64912 3244 64952
rect 3284 64912 3285 64952
rect 3243 64903 3285 64912
rect 3147 64784 3189 64793
rect 3147 64744 3148 64784
rect 3188 64744 3189 64784
rect 3147 64735 3189 64744
rect 3148 64616 3188 64735
rect 3148 64567 3188 64576
rect 3147 63020 3189 63029
rect 3147 62980 3148 63020
rect 3188 62980 3189 63020
rect 3147 62971 3189 62980
rect 3051 62516 3093 62525
rect 3051 62476 3052 62516
rect 3092 62476 3093 62516
rect 3051 62467 3093 62476
rect 3051 62348 3093 62357
rect 3051 62308 3052 62348
rect 3092 62308 3093 62348
rect 3051 62299 3093 62308
rect 2956 61508 2996 61517
rect 2860 61468 2956 61508
rect 2956 61459 2996 61468
rect 2764 61424 2804 61433
rect 2764 60257 2804 61384
rect 3052 61172 3092 62299
rect 3148 61606 3188 62971
rect 3148 61557 3188 61566
rect 3147 61172 3189 61181
rect 3052 61132 3148 61172
rect 3188 61132 3189 61172
rect 3147 61123 3189 61132
rect 3148 60920 3188 61123
rect 3244 61097 3284 64903
rect 3340 64709 3380 65164
rect 3531 65164 3572 65204
rect 3531 65120 3571 65164
rect 3531 65080 3572 65120
rect 3532 64961 3572 65080
rect 3688 65036 4056 65045
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 3688 64987 4056 64996
rect 3531 64952 3573 64961
rect 3531 64912 3532 64952
rect 3572 64912 3573 64952
rect 3531 64903 3573 64912
rect 3339 64700 3381 64709
rect 3339 64660 3340 64700
rect 3380 64660 3381 64700
rect 3339 64651 3381 64660
rect 3627 64700 3669 64709
rect 3627 64660 3628 64700
rect 3668 64660 3669 64700
rect 3627 64651 3669 64660
rect 3628 64630 3668 64651
rect 3628 64565 3668 64590
rect 4012 64616 4052 64625
rect 3819 64532 3861 64541
rect 3819 64492 3820 64532
rect 3860 64492 3861 64532
rect 3819 64483 3861 64492
rect 3820 64398 3860 64483
rect 4012 64280 4052 64576
rect 4012 64240 4148 64280
rect 3819 64196 3861 64205
rect 3819 64156 3820 64196
rect 3860 64156 3861 64196
rect 3819 64147 3861 64156
rect 3820 63944 3860 64147
rect 3820 63701 3860 63904
rect 3819 63692 3861 63701
rect 3819 63652 3820 63692
rect 3860 63652 3861 63692
rect 3819 63643 3861 63652
rect 3688 63524 4056 63533
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 3688 63475 4056 63484
rect 4108 63272 4148 64240
rect 4012 63232 4148 63272
rect 3340 62525 3380 62547
rect 4012 62525 4052 63232
rect 4204 63113 4244 66079
rect 4396 65540 4436 69355
rect 4492 69245 4532 69532
rect 4491 69236 4533 69245
rect 4491 69196 4492 69236
rect 4532 69196 4533 69236
rect 4491 69187 4533 69196
rect 4684 69161 4724 69246
rect 4683 69152 4725 69161
rect 4683 69112 4684 69152
rect 4724 69112 4725 69152
rect 4683 69103 4725 69112
rect 4492 68984 4532 68993
rect 4492 68396 4532 68944
rect 4780 68480 4820 70036
rect 4972 69987 5012 70120
rect 5163 70120 5164 70160
rect 5204 70120 5205 70160
rect 5163 70111 5205 70120
rect 5164 70026 5204 70111
rect 4972 69938 5012 69947
rect 4928 68816 5296 68825
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 4928 68767 5296 68776
rect 4820 68440 4916 68480
rect 4780 68431 4820 68440
rect 4491 68356 4532 68396
rect 4491 68312 4531 68356
rect 4491 68272 4532 68312
rect 4492 67817 4532 68272
rect 4491 67808 4533 67817
rect 4491 67768 4492 67808
rect 4532 67768 4533 67808
rect 4491 67759 4533 67768
rect 4683 67808 4725 67817
rect 4683 67768 4684 67808
rect 4724 67768 4725 67808
rect 4683 67759 4725 67768
rect 4684 67640 4724 67759
rect 4780 67649 4820 67734
rect 4684 67591 4724 67600
rect 4779 67640 4821 67649
rect 4779 67600 4780 67640
rect 4820 67600 4821 67640
rect 4779 67591 4821 67600
rect 4876 67472 4916 68440
rect 5163 67808 5205 67817
rect 5163 67768 5164 67808
rect 5204 67768 5205 67808
rect 5163 67759 5205 67768
rect 5164 67724 5204 67759
rect 5164 67673 5204 67684
rect 5259 67640 5301 67649
rect 5259 67600 5260 67640
rect 5300 67600 5301 67640
rect 5259 67591 5301 67600
rect 5260 67506 5300 67591
rect 4684 67432 4916 67472
rect 4587 66380 4629 66389
rect 4587 66340 4588 66380
rect 4628 66340 4629 66380
rect 4587 66331 4629 66340
rect 4588 66128 4628 66331
rect 4588 66079 4628 66088
rect 4491 65960 4533 65969
rect 4491 65920 4492 65960
rect 4532 65920 4533 65960
rect 4491 65911 4533 65920
rect 4300 65500 4436 65540
rect 4300 65288 4340 65500
rect 4492 65456 4532 65911
rect 4444 65446 4532 65456
rect 4484 65416 4532 65446
rect 4588 65540 4628 65549
rect 4444 65397 4484 65406
rect 4300 65248 4532 65288
rect 4492 64625 4532 65248
rect 4491 64616 4533 64625
rect 4491 64576 4492 64616
rect 4532 64576 4533 64616
rect 4491 64567 4533 64576
rect 4492 63617 4532 64567
rect 4588 64373 4628 65500
rect 4684 65129 4724 67432
rect 4928 67304 5296 67313
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 4928 67255 5296 67264
rect 5163 67136 5205 67145
rect 5163 67096 5164 67136
rect 5204 67096 5205 67136
rect 5163 67087 5205 67096
rect 5164 66968 5204 67087
rect 5164 66919 5204 66928
rect 5067 66212 5109 66221
rect 5067 66172 5068 66212
rect 5108 66172 5109 66212
rect 5067 66163 5109 66172
rect 5068 66128 5108 66163
rect 5068 66077 5108 66088
rect 4780 65969 4820 66054
rect 4779 65960 4821 65969
rect 4779 65920 4780 65960
rect 4820 65920 4821 65960
rect 4779 65911 4821 65920
rect 4928 65792 5296 65801
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 4928 65743 5296 65752
rect 4683 65120 4725 65129
rect 4683 65080 4684 65120
rect 4724 65080 4725 65120
rect 4683 65071 4725 65080
rect 5260 64616 5300 64627
rect 5260 64541 5300 64576
rect 5259 64532 5301 64541
rect 5259 64492 5260 64532
rect 5300 64492 5301 64532
rect 5259 64483 5301 64492
rect 4587 64364 4629 64373
rect 4587 64324 4588 64364
rect 4628 64324 4629 64364
rect 4587 64315 4629 64324
rect 4928 64280 5296 64289
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 4928 64231 5296 64240
rect 5067 64028 5109 64037
rect 5067 63988 5068 64028
rect 5108 63988 5109 64028
rect 5067 63979 5109 63988
rect 5068 63944 5108 63979
rect 4587 63776 4629 63785
rect 4587 63736 4588 63776
rect 4628 63736 4629 63776
rect 4587 63727 4629 63736
rect 4491 63608 4533 63617
rect 4491 63568 4492 63608
rect 4532 63568 4533 63608
rect 4491 63559 4533 63568
rect 4108 63104 4148 63113
rect 4203 63104 4245 63113
rect 4148 63064 4204 63104
rect 4244 63064 4245 63104
rect 4108 63055 4148 63064
rect 4203 63055 4245 63064
rect 4300 63104 4340 63115
rect 4204 62970 4244 63055
rect 4300 63029 4340 63064
rect 4299 63020 4341 63029
rect 4299 62980 4300 63020
rect 4340 62980 4341 63020
rect 4299 62971 4341 62980
rect 4395 62684 4437 62693
rect 4395 62644 4396 62684
rect 4436 62644 4437 62684
rect 4395 62635 4437 62644
rect 3339 62516 3381 62525
rect 3339 62476 3340 62516
rect 3380 62476 3381 62516
rect 3339 62467 3381 62476
rect 4011 62516 4053 62525
rect 4011 62476 4012 62516
rect 4052 62476 4053 62516
rect 4011 62467 4053 62476
rect 3340 62452 3380 62467
rect 3340 62403 3380 62412
rect 3436 62432 3476 62441
rect 3436 62348 3476 62392
rect 4396 62432 4436 62635
rect 4396 62383 4436 62392
rect 3340 62308 3476 62348
rect 3819 62348 3861 62357
rect 3819 62308 3820 62348
rect 3860 62308 3861 62348
rect 3340 61433 3380 62308
rect 3819 62299 3861 62308
rect 3916 62348 3956 62359
rect 3820 62214 3860 62299
rect 3916 62273 3956 62308
rect 3915 62264 3957 62273
rect 3915 62224 3916 62264
rect 3956 62224 3957 62264
rect 3915 62215 3957 62224
rect 4107 62264 4149 62273
rect 4107 62224 4108 62264
rect 4148 62224 4149 62264
rect 4107 62215 4149 62224
rect 3435 62096 3477 62105
rect 3435 62056 3436 62096
rect 3476 62056 3477 62096
rect 3435 62047 3477 62056
rect 3339 61424 3381 61433
rect 3339 61384 3340 61424
rect 3380 61384 3381 61424
rect 3339 61375 3381 61384
rect 3243 61088 3285 61097
rect 3243 61048 3244 61088
rect 3284 61048 3285 61088
rect 3243 61039 3285 61048
rect 3148 60871 3188 60880
rect 3051 60668 3093 60677
rect 3340 60668 3380 60677
rect 3051 60628 3052 60668
rect 3092 60628 3093 60668
rect 3051 60619 3093 60628
rect 3148 60628 3340 60668
rect 2955 60332 2997 60341
rect 2955 60292 2956 60332
rect 2996 60292 2997 60332
rect 2955 60283 2997 60292
rect 2763 60248 2805 60257
rect 2763 60208 2764 60248
rect 2804 60208 2805 60248
rect 2763 60199 2805 60208
rect 2956 60198 2996 60283
rect 2764 60080 2804 60089
rect 2476 60040 2764 60080
rect 2476 59408 2516 60040
rect 2764 60031 2804 60040
rect 2476 59240 2516 59368
rect 2956 59492 2996 59501
rect 2476 59200 2612 59240
rect 2380 59116 2516 59156
rect 2091 57560 2133 57569
rect 2091 57520 2092 57560
rect 2132 57520 2133 57560
rect 2091 57511 2133 57520
rect 2092 57140 2132 57511
rect 2092 57091 2132 57100
rect 2380 56888 2420 56897
rect 1995 56048 2037 56057
rect 1995 56008 1996 56048
rect 2036 56008 2037 56048
rect 1995 55999 2037 56008
rect 2380 55460 2420 56848
rect 2476 56645 2516 59116
rect 2572 58568 2612 59200
rect 2667 59156 2709 59165
rect 2667 59116 2668 59156
rect 2708 59116 2709 59156
rect 2667 59107 2709 59116
rect 2668 59022 2708 59107
rect 2668 58568 2708 58577
rect 2572 58528 2668 58568
rect 2668 57989 2708 58528
rect 2860 58400 2900 58409
rect 2764 58360 2860 58400
rect 2667 57980 2709 57989
rect 2667 57940 2668 57980
rect 2708 57940 2709 57980
rect 2667 57931 2709 57940
rect 2764 57728 2804 58360
rect 2860 58351 2900 58360
rect 2956 58148 2996 59452
rect 3052 58736 3092 60619
rect 3148 59403 3188 60628
rect 3340 60619 3380 60628
rect 3339 60500 3381 60509
rect 3339 60460 3340 60500
rect 3380 60460 3381 60500
rect 3339 60451 3381 60460
rect 3243 60248 3285 60257
rect 3243 60208 3244 60248
rect 3284 60208 3285 60248
rect 3243 60199 3285 60208
rect 3244 60080 3284 60199
rect 3244 60031 3284 60040
rect 3340 60080 3380 60451
rect 3148 59354 3188 59363
rect 3340 58829 3380 60040
rect 3339 58820 3381 58829
rect 3339 58780 3340 58820
rect 3380 58780 3381 58820
rect 3339 58771 3381 58780
rect 3052 58696 3188 58736
rect 3051 58568 3093 58577
rect 3051 58528 3052 58568
rect 3092 58528 3093 58568
rect 3051 58519 3093 58528
rect 3052 58434 3092 58519
rect 3148 58148 3188 58696
rect 3436 58577 3476 62047
rect 3531 62012 3573 62021
rect 3531 61972 3532 62012
rect 3572 61972 3573 62012
rect 3531 61963 3573 61972
rect 3688 62012 4056 62021
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 3688 61963 4056 61972
rect 3532 61760 3572 61963
rect 3532 61720 3668 61760
rect 3628 61601 3668 61720
rect 4108 61676 4148 62215
rect 4491 62180 4533 62189
rect 4491 62140 4492 62180
rect 4532 62140 4533 62180
rect 4491 62131 4533 62140
rect 4203 61928 4245 61937
rect 4203 61888 4204 61928
rect 4244 61888 4245 61928
rect 4203 61879 4245 61888
rect 4395 61928 4437 61937
rect 4395 61888 4396 61928
rect 4436 61888 4439 61928
rect 4395 61879 4439 61888
rect 4108 61627 4148 61636
rect 4204 61676 4244 61879
rect 4299 61760 4341 61769
rect 4399 61760 4439 61879
rect 4299 61720 4300 61760
rect 4340 61720 4341 61760
rect 4299 61711 4341 61720
rect 4396 61720 4439 61760
rect 4204 61625 4244 61636
rect 3627 61592 3669 61601
rect 3627 61552 3628 61592
rect 3668 61552 3669 61592
rect 3627 61543 3669 61552
rect 3627 61424 3669 61433
rect 3627 61384 3628 61424
rect 3668 61384 3669 61424
rect 3627 61375 3669 61384
rect 3532 60929 3572 61014
rect 3531 60920 3573 60929
rect 3531 60880 3532 60920
rect 3572 60880 3573 60920
rect 3531 60871 3573 60880
rect 3628 60752 3668 61375
rect 3532 60712 3668 60752
rect 3532 60509 3572 60712
rect 4300 60677 4340 61711
rect 4299 60668 4341 60677
rect 4299 60628 4300 60668
rect 4340 60628 4341 60668
rect 4299 60619 4341 60628
rect 3531 60500 3573 60509
rect 3531 60460 3532 60500
rect 3572 60460 3573 60500
rect 3531 60451 3573 60460
rect 3688 60500 4056 60509
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 3688 60451 4056 60460
rect 4107 60164 4149 60173
rect 4107 60124 4108 60164
rect 4148 60124 4149 60164
rect 4107 60115 4149 60124
rect 3724 60080 3764 60089
rect 3627 59996 3669 60005
rect 3627 59956 3628 59996
rect 3668 59956 3669 59996
rect 3627 59947 3669 59956
rect 3628 59408 3668 59947
rect 3628 59359 3668 59368
rect 3724 59333 3764 60040
rect 3819 60080 3861 60089
rect 3819 60040 3820 60080
rect 3860 60040 3861 60080
rect 3819 60031 3861 60040
rect 3820 59946 3860 60031
rect 4108 59408 4148 60115
rect 4300 60080 4340 60091
rect 4300 60005 4340 60040
rect 4299 59996 4341 60005
rect 4299 59956 4300 59996
rect 4340 59956 4341 59996
rect 4299 59947 4341 59956
rect 4108 59359 4148 59368
rect 4204 59333 4244 59418
rect 3723 59324 3765 59333
rect 3723 59284 3724 59324
rect 3764 59284 3765 59324
rect 3723 59275 3765 59284
rect 4203 59324 4245 59333
rect 4203 59284 4204 59324
rect 4244 59284 4245 59324
rect 4203 59275 4245 59284
rect 4203 59156 4245 59165
rect 4203 59116 4204 59156
rect 4244 59116 4245 59156
rect 4203 59107 4245 59116
rect 3688 58988 4056 58997
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 3688 58939 4056 58948
rect 3627 58820 3669 58829
rect 3627 58780 3628 58820
rect 3668 58780 3669 58820
rect 3627 58771 3669 58780
rect 3435 58568 3477 58577
rect 3435 58528 3436 58568
rect 3476 58528 3477 58568
rect 3435 58519 3477 58528
rect 2572 57688 2804 57728
rect 2860 58108 2996 58148
rect 3052 58108 3188 58148
rect 2572 57070 2612 57688
rect 2572 57021 2612 57030
rect 2763 56972 2805 56981
rect 2763 56932 2764 56972
rect 2804 56932 2805 56972
rect 2763 56923 2805 56932
rect 2475 56636 2517 56645
rect 2475 56596 2476 56636
rect 2516 56596 2517 56636
rect 2475 56587 2517 56596
rect 2284 55420 2420 55460
rect 2476 55544 2516 55553
rect 2091 55124 2133 55133
rect 2091 55084 2092 55124
rect 2132 55084 2133 55124
rect 2091 55075 2133 55084
rect 2092 54788 2132 55075
rect 2187 54956 2229 54965
rect 2187 54916 2188 54956
rect 2228 54916 2229 54956
rect 2187 54907 2229 54916
rect 2092 54739 2132 54748
rect 1803 54704 1845 54713
rect 1803 54664 1804 54704
rect 1844 54664 1845 54704
rect 1803 54655 1845 54664
rect 1516 54620 1556 54629
rect 1899 54620 1941 54629
rect 1556 54580 1652 54620
rect 1516 54571 1556 54580
rect 1419 54032 1461 54041
rect 1419 53992 1420 54032
rect 1460 53992 1461 54032
rect 1419 53983 1461 53992
rect 1516 53864 1556 53873
rect 1516 53453 1556 53824
rect 1515 53444 1557 53453
rect 1515 53404 1516 53444
rect 1556 53404 1557 53444
rect 1515 53395 1557 53404
rect 1516 53276 1556 53285
rect 1324 53236 1516 53276
rect 1516 53227 1556 53236
rect 1324 53108 1364 53117
rect 1324 51185 1364 53068
rect 1515 52688 1557 52697
rect 1515 52648 1516 52688
rect 1556 52648 1557 52688
rect 1515 52639 1557 52648
rect 1516 52520 1556 52639
rect 1612 52529 1652 54580
rect 1899 54580 1900 54620
rect 1940 54580 1941 54620
rect 1899 54571 1941 54580
rect 1900 54486 1940 54571
rect 1708 54116 1748 54125
rect 2092 54116 2132 54125
rect 1748 54076 2036 54116
rect 1708 54067 1748 54076
rect 1900 53864 1940 53873
rect 1804 53824 1900 53864
rect 1708 53108 1748 53117
rect 1420 52480 1516 52520
rect 1323 51176 1365 51185
rect 1323 51136 1324 51176
rect 1364 51136 1365 51176
rect 1323 51127 1365 51136
rect 1228 51008 1268 51017
rect 1420 51008 1460 52480
rect 1516 52471 1556 52480
rect 1611 52520 1653 52529
rect 1611 52480 1612 52520
rect 1652 52480 1653 52520
rect 1611 52471 1653 52480
rect 1611 52352 1653 52361
rect 1611 52312 1612 52352
rect 1652 52312 1653 52352
rect 1611 52303 1653 52312
rect 1516 51848 1556 51859
rect 1516 51773 1556 51808
rect 1515 51764 1557 51773
rect 1515 51724 1516 51764
rect 1556 51724 1557 51764
rect 1515 51715 1557 51724
rect 1515 51596 1557 51605
rect 1515 51556 1516 51596
rect 1556 51556 1557 51596
rect 1515 51547 1557 51556
rect 1268 50968 1460 51008
rect 1228 50959 1268 50968
rect 1516 50924 1556 51547
rect 1420 50884 1556 50924
rect 1420 49589 1460 50884
rect 1516 50084 1556 50093
rect 1516 49841 1556 50044
rect 1612 49925 1652 52303
rect 1708 51857 1748 53068
rect 1804 52865 1844 53824
rect 1900 53815 1940 53824
rect 1899 53276 1941 53285
rect 1899 53236 1900 53276
rect 1940 53236 1941 53276
rect 1899 53227 1941 53236
rect 1900 53142 1940 53227
rect 1996 52865 2036 54076
rect 2092 53957 2132 54076
rect 2091 53948 2133 53957
rect 2091 53908 2092 53948
rect 2132 53908 2133 53948
rect 2091 53899 2133 53908
rect 2092 53360 2132 53369
rect 1803 52856 1845 52865
rect 1803 52816 1804 52856
rect 1844 52816 1845 52856
rect 1803 52807 1845 52816
rect 1995 52856 2037 52865
rect 1995 52816 1996 52856
rect 2036 52816 2037 52856
rect 1995 52807 2037 52816
rect 1707 51848 1749 51857
rect 1707 51808 1708 51848
rect 1748 51808 1749 51848
rect 1707 51799 1749 51808
rect 2092 51773 2132 53320
rect 2091 51764 2133 51773
rect 2091 51724 2092 51764
rect 2132 51724 2133 51764
rect 2091 51715 2133 51724
rect 1995 51512 2037 51521
rect 1995 51472 1996 51512
rect 2036 51472 2037 51512
rect 1995 51463 2037 51472
rect 1803 50504 1845 50513
rect 1803 50464 1804 50504
rect 1844 50464 1845 50504
rect 1803 50455 1845 50464
rect 1707 50252 1749 50261
rect 1707 50212 1708 50252
rect 1748 50212 1749 50252
rect 1707 50203 1749 50212
rect 1708 50118 1748 50203
rect 1611 49916 1653 49925
rect 1611 49876 1612 49916
rect 1652 49876 1653 49916
rect 1611 49867 1653 49876
rect 1515 49832 1557 49841
rect 1515 49792 1516 49832
rect 1556 49792 1557 49832
rect 1515 49783 1557 49792
rect 1419 49580 1461 49589
rect 1419 49540 1420 49580
rect 1460 49540 1461 49580
rect 1419 49531 1461 49540
rect 1707 49328 1749 49337
rect 1707 49288 1708 49328
rect 1748 49288 1749 49328
rect 1707 49279 1749 49288
rect 1323 49160 1365 49169
rect 1323 49120 1324 49160
rect 1364 49120 1365 49160
rect 1323 49111 1365 49120
rect 1324 47648 1364 49111
rect 1611 48824 1653 48833
rect 1611 48784 1612 48824
rect 1652 48784 1653 48824
rect 1611 48775 1653 48784
rect 1516 48572 1556 48581
rect 1420 48532 1516 48572
rect 1420 47825 1460 48532
rect 1516 48523 1556 48532
rect 1516 48236 1556 48245
rect 1612 48236 1652 48775
rect 1708 48740 1748 49279
rect 1804 48992 1844 50455
rect 1900 50084 1940 50093
rect 1996 50084 2036 51463
rect 2092 50252 2132 50261
rect 2188 50252 2228 54907
rect 2132 50212 2228 50252
rect 2284 50252 2324 55420
rect 2476 55124 2516 55504
rect 2667 55376 2709 55385
rect 2667 55336 2668 55376
rect 2708 55336 2709 55376
rect 2667 55327 2709 55336
rect 2668 55242 2708 55327
rect 2476 55084 2612 55124
rect 2475 54956 2517 54965
rect 2475 54916 2476 54956
rect 2516 54916 2517 54956
rect 2475 54907 2517 54916
rect 2476 54822 2516 54907
rect 2379 54620 2421 54629
rect 2379 54580 2380 54620
rect 2420 54580 2421 54620
rect 2379 54571 2421 54580
rect 2380 52193 2420 54571
rect 2572 54377 2612 55084
rect 2668 54858 2708 54867
rect 2571 54368 2613 54377
rect 2571 54328 2572 54368
rect 2612 54328 2613 54368
rect 2571 54319 2613 54328
rect 2668 54209 2708 54818
rect 2667 54200 2709 54209
rect 2667 54160 2668 54200
rect 2708 54160 2709 54200
rect 2667 54151 2709 54160
rect 2572 54032 2612 54041
rect 2572 53369 2612 53992
rect 2571 53360 2613 53369
rect 2571 53320 2572 53360
rect 2612 53320 2613 53360
rect 2571 53311 2613 53320
rect 2764 52856 2804 56923
rect 2860 56552 2900 58108
rect 2955 57980 2997 57989
rect 2955 57940 2956 57980
rect 2996 57940 2997 57980
rect 2955 57931 2997 57940
rect 2956 57896 2996 57931
rect 2956 57845 2996 57856
rect 3052 57056 3092 58108
rect 3628 58073 3668 58771
rect 4107 58316 4149 58325
rect 4107 58276 4108 58316
rect 4148 58276 4149 58316
rect 4107 58267 4149 58276
rect 3627 58064 3669 58073
rect 3627 58024 3628 58064
rect 3668 58024 3669 58064
rect 3627 58015 3669 58024
rect 3148 57980 3188 57989
rect 3188 57940 3572 57980
rect 3148 57931 3188 57940
rect 3532 57896 3572 57940
rect 3532 57847 3572 57856
rect 3628 57896 3668 58015
rect 3628 57847 3668 57856
rect 4011 57896 4053 57905
rect 4011 57856 4012 57896
rect 4052 57856 4053 57896
rect 4011 57847 4053 57856
rect 4108 57896 4148 58267
rect 4108 57847 4148 57856
rect 4012 57762 4052 57847
rect 3531 57728 3573 57737
rect 3531 57688 3532 57728
rect 3572 57688 3573 57728
rect 3531 57679 3573 57688
rect 3532 57140 3572 57679
rect 3688 57476 4056 57485
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 3688 57427 4056 57436
rect 3627 57224 3669 57233
rect 3627 57184 3628 57224
rect 3668 57184 3669 57224
rect 3627 57175 3669 57184
rect 3819 57224 3861 57233
rect 3819 57184 3820 57224
rect 3860 57184 3861 57224
rect 3819 57175 3861 57184
rect 3092 57016 3188 57056
rect 3052 57007 3092 57016
rect 2860 56512 2996 56552
rect 2956 56393 2996 56512
rect 3052 56477 3092 56562
rect 3051 56468 3093 56477
rect 3051 56428 3052 56468
rect 3092 56428 3093 56468
rect 3051 56419 3093 56428
rect 2860 56384 2900 56393
rect 2860 56216 2900 56344
rect 2955 56384 2997 56393
rect 2955 56344 2956 56384
rect 2996 56344 2997 56384
rect 2955 56335 2997 56344
rect 3148 56379 3188 57016
rect 3435 56384 3477 56393
rect 3148 56339 3189 56379
rect 3149 56216 3189 56339
rect 3435 56344 3436 56384
rect 3476 56344 3477 56384
rect 3435 56335 3477 56344
rect 2860 56176 2996 56216
rect 2860 55376 2900 55385
rect 2860 54293 2900 55336
rect 2956 54713 2996 56176
rect 3148 56176 3189 56216
rect 3051 55796 3093 55805
rect 3051 55756 3052 55796
rect 3092 55756 3093 55796
rect 3051 55747 3093 55756
rect 3052 55628 3092 55747
rect 3052 55579 3092 55588
rect 3148 55553 3188 56176
rect 3339 56132 3381 56141
rect 3339 56092 3340 56132
rect 3380 56092 3381 56132
rect 3339 56083 3381 56092
rect 3243 55712 3285 55721
rect 3243 55672 3244 55712
rect 3284 55672 3285 55712
rect 3243 55663 3285 55672
rect 3244 55578 3284 55663
rect 3147 55544 3189 55553
rect 3147 55504 3148 55544
rect 3188 55504 3189 55544
rect 3147 55495 3189 55504
rect 3148 54872 3188 55495
rect 3340 55460 3380 56083
rect 3436 55628 3476 56335
rect 3532 55796 3572 57100
rect 3628 57140 3668 57175
rect 3628 57089 3668 57100
rect 3627 56468 3669 56477
rect 3627 56428 3628 56468
rect 3668 56428 3669 56468
rect 3627 56419 3669 56428
rect 3628 56384 3668 56419
rect 3628 56333 3668 56344
rect 3724 56384 3764 56393
rect 3820 56384 3860 57175
rect 4012 57056 4052 57065
rect 4012 56888 4052 57016
rect 4108 57056 4148 57065
rect 4204 57056 4244 59107
rect 4300 59072 4340 59947
rect 4396 59333 4436 61720
rect 4492 60752 4532 62131
rect 4588 62105 4628 63727
rect 4779 63692 4821 63701
rect 4779 63652 4780 63692
rect 4820 63652 4821 63692
rect 4779 63643 4821 63652
rect 4683 63272 4725 63281
rect 4683 63232 4684 63272
rect 4724 63232 4725 63272
rect 4683 63223 4725 63232
rect 4587 62096 4629 62105
rect 4587 62056 4588 62096
rect 4628 62056 4629 62096
rect 4587 62047 4629 62056
rect 4588 61592 4628 61601
rect 4588 61433 4628 61552
rect 4684 61592 4724 63223
rect 4780 62600 4820 63643
rect 5068 63113 5108 63904
rect 5259 63692 5301 63701
rect 5259 63652 5260 63692
rect 5300 63652 5301 63692
rect 5259 63643 5301 63652
rect 5260 63558 5300 63643
rect 5067 63104 5109 63113
rect 5067 63064 5068 63104
rect 5108 63064 5109 63104
rect 5067 63055 5109 63064
rect 4928 62768 5296 62777
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 4928 62719 5296 62728
rect 5067 62600 5109 62609
rect 4780 62560 4916 62600
rect 4876 62427 4916 62560
rect 5067 62560 5068 62600
rect 5108 62560 5109 62600
rect 5067 62551 5109 62560
rect 5068 62466 5108 62551
rect 4876 62378 4916 62387
rect 4684 61543 4724 61552
rect 4587 61424 4629 61433
rect 4587 61384 4588 61424
rect 4628 61384 4629 61424
rect 4587 61375 4629 61384
rect 4928 61256 5296 61265
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 4928 61207 5296 61216
rect 4779 61172 4821 61181
rect 4779 61132 4780 61172
rect 4820 61132 4821 61172
rect 4779 61123 4821 61132
rect 4780 60920 4820 61123
rect 4780 60871 4820 60880
rect 5163 60920 5205 60929
rect 5163 60880 5164 60920
rect 5204 60880 5205 60920
rect 5163 60871 5205 60880
rect 5164 60786 5204 60871
rect 4492 60712 4724 60752
rect 4587 59408 4629 59417
rect 4587 59368 4588 59408
rect 4628 59368 4629 59408
rect 4587 59359 4629 59368
rect 4684 59408 4724 60712
rect 4971 60668 5013 60677
rect 4971 60628 4972 60668
rect 5012 60628 5013 60668
rect 4971 60619 5013 60628
rect 4972 60534 5012 60619
rect 4779 60332 4821 60341
rect 4779 60292 4780 60332
rect 4820 60292 4821 60332
rect 4779 60283 4821 60292
rect 4780 60094 4820 60283
rect 4780 60045 4820 60054
rect 4972 59912 5012 59921
rect 4684 59359 4724 59368
rect 4780 59872 4972 59912
rect 4395 59324 4437 59333
rect 4395 59284 4396 59324
rect 4436 59284 4437 59324
rect 4395 59275 4437 59284
rect 4588 59274 4628 59359
rect 4780 59333 4820 59872
rect 4972 59863 5012 59872
rect 4928 59744 5296 59753
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 4928 59695 5296 59704
rect 5356 59333 5396 71287
rect 5452 64709 5492 72127
rect 5548 69161 5588 72136
rect 5547 69152 5589 69161
rect 5547 69112 5548 69152
rect 5588 69112 5589 69152
rect 5547 69103 5589 69112
rect 5547 68816 5589 68825
rect 5547 68776 5548 68816
rect 5588 68776 5589 68816
rect 5547 68767 5589 68776
rect 5548 65204 5588 68767
rect 5644 67817 5684 73051
rect 5740 72521 5780 77344
rect 5932 75461 5972 79771
rect 6124 79493 6164 80536
rect 6219 80536 6220 80576
rect 6260 80536 6261 80576
rect 6219 80527 6261 80536
rect 6220 80442 6260 80527
rect 6123 79484 6165 79493
rect 6123 79444 6124 79484
rect 6164 79444 6165 79484
rect 6123 79435 6165 79444
rect 6219 79064 6261 79073
rect 6219 79024 6220 79064
rect 6260 79024 6261 79064
rect 6219 79015 6261 79024
rect 6220 78930 6260 79015
rect 6027 78644 6069 78653
rect 6027 78604 6028 78644
rect 6068 78604 6069 78644
rect 6316 78644 6356 81880
rect 6604 80576 6644 80585
rect 6508 80536 6604 80576
rect 6508 79073 6548 80536
rect 6604 80527 6644 80536
rect 6700 79241 6740 81955
rect 6796 81920 6836 82375
rect 6892 82256 6932 82963
rect 6988 82256 7028 84307
rect 7084 83768 7124 84316
rect 7180 83861 7220 85936
rect 7276 84440 7316 84449
rect 7372 84440 7412 85936
rect 7564 84533 7604 85936
rect 7659 85196 7701 85205
rect 7659 85156 7660 85196
rect 7700 85156 7701 85196
rect 7659 85147 7701 85156
rect 7563 84524 7605 84533
rect 7563 84484 7564 84524
rect 7604 84484 7605 84524
rect 7660 84524 7700 85147
rect 7756 84701 7796 85936
rect 7948 85289 7988 85936
rect 7947 85280 7989 85289
rect 7947 85240 7948 85280
rect 7988 85240 7989 85280
rect 7947 85231 7989 85240
rect 8140 84944 8180 85936
rect 7948 84904 8180 84944
rect 7755 84692 7797 84701
rect 7755 84652 7756 84692
rect 7796 84652 7797 84692
rect 7755 84643 7797 84652
rect 7660 84484 7796 84524
rect 7563 84475 7605 84484
rect 7316 84400 7412 84440
rect 7276 84391 7316 84400
rect 7659 84356 7701 84365
rect 7659 84316 7660 84356
rect 7700 84316 7701 84356
rect 7659 84307 7701 84316
rect 7660 84222 7700 84307
rect 7275 83936 7317 83945
rect 7275 83896 7276 83936
rect 7316 83896 7317 83936
rect 7275 83887 7317 83896
rect 7179 83852 7221 83861
rect 7179 83812 7180 83852
rect 7220 83812 7221 83852
rect 7179 83803 7221 83812
rect 7084 83719 7124 83728
rect 7083 83600 7125 83609
rect 7083 83560 7084 83600
rect 7124 83560 7125 83600
rect 7083 83551 7125 83560
rect 7084 82433 7124 83551
rect 7179 83432 7221 83441
rect 7179 83392 7180 83432
rect 7220 83392 7221 83432
rect 7179 83383 7221 83392
rect 7180 83298 7220 83383
rect 7276 83180 7316 83887
rect 7180 83140 7316 83180
rect 7372 83600 7412 83609
rect 7180 82844 7220 83140
rect 7180 82795 7220 82804
rect 7275 82760 7317 82769
rect 7275 82720 7276 82760
rect 7316 82720 7317 82760
rect 7275 82711 7317 82720
rect 7276 82626 7316 82711
rect 7372 82517 7412 83560
rect 7563 83348 7605 83357
rect 7563 83308 7564 83348
rect 7604 83308 7605 83348
rect 7563 83299 7605 83308
rect 7371 82508 7413 82517
rect 7371 82468 7372 82508
rect 7412 82468 7413 82508
rect 7371 82459 7413 82468
rect 7083 82424 7125 82433
rect 7083 82384 7084 82424
rect 7124 82384 7125 82424
rect 7083 82375 7125 82384
rect 7180 82256 7220 82265
rect 6988 82216 7180 82256
rect 6892 82207 6932 82216
rect 7180 82207 7220 82216
rect 7372 82181 7412 82459
rect 7371 82172 7413 82181
rect 7371 82132 7372 82172
rect 7412 82132 7413 82172
rect 7371 82123 7413 82132
rect 7083 82088 7125 82097
rect 7083 82048 7084 82088
rect 7124 82048 7125 82088
rect 7083 82039 7125 82048
rect 7564 82088 7604 83299
rect 7756 83096 7796 84484
rect 7851 84440 7893 84449
rect 7851 84400 7852 84440
rect 7892 84400 7893 84440
rect 7851 84391 7893 84400
rect 7852 84306 7892 84391
rect 7948 83189 7988 84904
rect 8043 84776 8085 84785
rect 8043 84736 8044 84776
rect 8084 84736 8085 84776
rect 8043 84727 8085 84736
rect 8044 84440 8084 84727
rect 8044 84391 8084 84400
rect 8236 84356 8276 84365
rect 8140 84316 8236 84356
rect 7947 83180 7989 83189
rect 7947 83140 7948 83180
rect 7988 83140 7989 83180
rect 7947 83131 7989 83140
rect 7660 83056 7796 83096
rect 7660 82517 7700 83056
rect 7755 82760 7797 82769
rect 7755 82720 7756 82760
rect 7796 82720 7797 82760
rect 7755 82711 7797 82720
rect 7756 82626 7796 82711
rect 7659 82508 7701 82517
rect 7659 82468 7660 82508
rect 7700 82468 7701 82508
rect 7659 82459 7701 82468
rect 6796 81880 7028 81920
rect 6988 81248 7028 81880
rect 6988 81199 7028 81208
rect 6891 80744 6933 80753
rect 6891 80704 6892 80744
rect 6932 80704 6933 80744
rect 6891 80695 6933 80704
rect 6892 80576 6932 80695
rect 7084 80660 7124 82039
rect 7372 82004 7412 82013
rect 7412 81964 7508 82004
rect 7372 81955 7412 81964
rect 7371 81248 7413 81257
rect 7371 81208 7372 81248
rect 7412 81208 7413 81248
rect 7371 81199 7413 81208
rect 7372 81114 7412 81199
rect 7180 81080 7220 81089
rect 7220 81040 7316 81080
rect 7180 81031 7220 81040
rect 7084 80620 7220 80660
rect 6796 80492 6836 80501
rect 6699 79232 6741 79241
rect 6699 79192 6700 79232
rect 6740 79192 6741 79232
rect 6699 79183 6741 79192
rect 6507 79064 6549 79073
rect 6507 79024 6508 79064
rect 6548 79024 6549 79064
rect 6507 79015 6549 79024
rect 6412 78812 6452 78821
rect 6508 78812 6548 79015
rect 6452 78772 6548 78812
rect 6412 78763 6452 78772
rect 6316 78604 6452 78644
rect 6027 78595 6069 78604
rect 6028 78233 6068 78595
rect 6027 78224 6069 78233
rect 6027 78184 6028 78224
rect 6068 78184 6069 78224
rect 6027 78175 6069 78184
rect 6123 77552 6165 77561
rect 6123 77512 6124 77552
rect 6164 77512 6165 77552
rect 6123 77503 6165 77512
rect 6220 77552 6260 77561
rect 6124 77418 6164 77503
rect 6220 76637 6260 77512
rect 6316 76805 6356 76836
rect 6315 76796 6357 76805
rect 6315 76756 6316 76796
rect 6356 76756 6357 76796
rect 6315 76747 6357 76756
rect 6316 76712 6356 76747
rect 6219 76628 6261 76637
rect 6124 76588 6220 76628
rect 6260 76588 6261 76628
rect 5931 75452 5973 75461
rect 5931 75412 5932 75452
rect 5972 75412 5973 75452
rect 5931 75403 5973 75412
rect 5836 75200 5876 75209
rect 5836 74285 5876 75160
rect 5932 74360 5972 75403
rect 6028 75032 6068 75041
rect 6028 74528 6068 74992
rect 6028 74479 6068 74488
rect 6124 74528 6164 76588
rect 6219 76579 6261 76588
rect 6220 76040 6260 76049
rect 6316 76040 6356 76672
rect 6412 76376 6452 78604
rect 6508 78149 6548 78772
rect 6700 78233 6740 79183
rect 6699 78224 6741 78233
rect 6699 78184 6700 78224
rect 6740 78184 6741 78224
rect 6699 78175 6741 78184
rect 6507 78140 6549 78149
rect 6507 78100 6508 78140
rect 6548 78100 6549 78140
rect 6507 78091 6549 78100
rect 6508 77561 6548 78091
rect 6507 77552 6549 77561
rect 6507 77512 6508 77552
rect 6548 77512 6549 77552
rect 6507 77503 6549 77512
rect 6604 77468 6644 77477
rect 6604 76628 6644 77428
rect 6700 77468 6740 77477
rect 6700 76964 6740 77428
rect 6796 77393 6836 80452
rect 6892 79409 6932 80536
rect 7180 80501 7220 80620
rect 6987 80492 7029 80501
rect 7084 80492 7124 80501
rect 6987 80452 6988 80492
rect 7028 80452 7084 80492
rect 6987 80443 7029 80452
rect 7084 80443 7124 80452
rect 7179 80492 7221 80501
rect 7179 80452 7180 80492
rect 7220 80452 7221 80492
rect 7179 80443 7221 80452
rect 7276 80333 7316 81040
rect 7468 80744 7508 81964
rect 7564 80753 7604 82048
rect 7660 81920 7700 82459
rect 7660 81880 7796 81920
rect 7660 81248 7700 81257
rect 7660 81005 7700 81208
rect 7659 80996 7701 81005
rect 7659 80956 7660 80996
rect 7700 80956 7701 80996
rect 7659 80947 7701 80956
rect 7372 80704 7508 80744
rect 7563 80744 7605 80753
rect 7563 80704 7564 80744
rect 7604 80704 7605 80744
rect 7275 80324 7317 80333
rect 7275 80284 7276 80324
rect 7316 80284 7317 80324
rect 7275 80275 7317 80284
rect 6988 79736 7028 79745
rect 6891 79400 6933 79409
rect 6891 79360 6892 79400
rect 6932 79360 6933 79400
rect 6891 79351 6933 79360
rect 6988 79241 7028 79696
rect 7180 79568 7220 79577
rect 7180 79241 7220 79528
rect 6987 79232 7029 79241
rect 6987 79192 6988 79232
rect 7028 79192 7029 79232
rect 6987 79183 7029 79192
rect 7179 79232 7221 79241
rect 7179 79192 7180 79232
rect 7220 79192 7221 79232
rect 7179 79183 7221 79192
rect 6891 79064 6933 79073
rect 6891 79024 6892 79064
rect 6932 79024 6933 79064
rect 6891 79015 6933 79024
rect 6988 79064 7028 79073
rect 6892 78930 6932 79015
rect 6988 78317 7028 79024
rect 7084 79064 7124 79073
rect 7084 78476 7124 79024
rect 7180 79064 7220 79073
rect 7372 79064 7412 80704
rect 7563 80695 7605 80704
rect 7468 80576 7508 80585
rect 7468 80333 7508 80536
rect 7564 80576 7604 80587
rect 7564 80501 7604 80536
rect 7659 80576 7701 80585
rect 7659 80536 7660 80576
rect 7700 80536 7701 80576
rect 7659 80527 7701 80536
rect 7563 80492 7605 80501
rect 7563 80452 7564 80492
rect 7604 80452 7605 80492
rect 7563 80443 7605 80452
rect 7467 80324 7509 80333
rect 7467 80284 7468 80324
rect 7508 80284 7509 80324
rect 7467 80275 7509 80284
rect 7467 79820 7509 79829
rect 7467 79780 7468 79820
rect 7508 79780 7509 79820
rect 7467 79771 7509 79780
rect 7468 79686 7508 79771
rect 7563 79568 7605 79577
rect 7468 79528 7564 79568
rect 7604 79528 7605 79568
rect 7468 79232 7508 79528
rect 7563 79519 7605 79528
rect 7563 79400 7605 79409
rect 7563 79360 7564 79400
rect 7604 79360 7605 79400
rect 7563 79351 7605 79360
rect 7468 79183 7508 79192
rect 7220 79024 7316 79064
rect 7372 79024 7508 79064
rect 7180 79015 7220 79024
rect 7084 78427 7124 78436
rect 6987 78308 7029 78317
rect 6987 78268 6988 78308
rect 7028 78268 7029 78308
rect 6987 78259 7029 78268
rect 6891 78224 6933 78233
rect 6891 78184 6892 78224
rect 6932 78184 6933 78224
rect 6891 78175 6933 78184
rect 6892 78090 6932 78175
rect 7084 78056 7124 78065
rect 7084 77645 7124 78016
rect 7083 77636 7125 77645
rect 7083 77596 7084 77636
rect 7124 77596 7125 77636
rect 7083 77587 7125 77596
rect 7179 77552 7221 77561
rect 7179 77512 7180 77552
rect 7220 77512 7221 77552
rect 7179 77503 7221 77512
rect 7180 77418 7220 77503
rect 7276 77477 7316 79024
rect 7371 78896 7413 78905
rect 7371 78856 7372 78896
rect 7412 78856 7413 78896
rect 7371 78847 7413 78856
rect 7372 78762 7412 78847
rect 7372 78224 7412 78235
rect 7372 78149 7412 78184
rect 7371 78140 7413 78149
rect 7371 78100 7372 78140
rect 7412 78100 7413 78140
rect 7371 78091 7413 78100
rect 7275 77468 7317 77477
rect 7275 77428 7276 77468
rect 7316 77428 7317 77468
rect 7275 77419 7317 77428
rect 6795 77384 6837 77393
rect 6795 77344 6796 77384
rect 6836 77344 6837 77384
rect 6795 77335 6837 77344
rect 6700 76924 7316 76964
rect 6700 76754 6740 76763
rect 6700 76712 6740 76714
rect 7083 76712 7125 76721
rect 6700 76672 7084 76712
rect 7124 76672 7125 76712
rect 7083 76663 7125 76672
rect 6604 76588 7028 76628
rect 6508 76544 6548 76553
rect 6548 76504 6836 76544
rect 6508 76495 6548 76504
rect 6412 76336 6548 76376
rect 6260 76000 6356 76040
rect 6412 76124 6452 76133
rect 6220 75991 6260 76000
rect 6412 75965 6452 76084
rect 6411 75956 6453 75965
rect 6411 75916 6412 75956
rect 6452 75916 6453 75956
rect 6411 75907 6453 75916
rect 6508 75704 6548 76336
rect 6700 76217 6740 76302
rect 6699 76208 6741 76217
rect 6699 76168 6700 76208
rect 6740 76168 6741 76208
rect 6699 76159 6741 76168
rect 6796 76133 6836 76504
rect 6891 76208 6933 76217
rect 6891 76168 6892 76208
rect 6932 76168 6933 76208
rect 6891 76159 6933 76168
rect 6795 76124 6837 76133
rect 6795 76084 6796 76124
rect 6836 76084 6837 76124
rect 6795 76075 6837 76084
rect 6796 76040 6836 76075
rect 6412 75664 6548 75704
rect 6638 76025 6678 76034
rect 6796 75990 6836 76000
rect 6892 76040 6932 76159
rect 6892 75991 6932 76000
rect 6315 75620 6357 75629
rect 6315 75580 6316 75620
rect 6356 75580 6357 75620
rect 6315 75571 6357 75580
rect 6316 75452 6356 75571
rect 6316 75403 6356 75412
rect 6219 75284 6261 75293
rect 6219 75244 6220 75284
rect 6260 75244 6261 75284
rect 6219 75235 6261 75244
rect 6220 75200 6260 75235
rect 6220 75149 6260 75160
rect 6124 74479 6164 74488
rect 5932 74320 6260 74360
rect 5835 74276 5877 74285
rect 5835 74236 5836 74276
rect 5876 74236 5877 74276
rect 5835 74227 5877 74236
rect 5739 72512 5781 72521
rect 5739 72472 5740 72512
rect 5780 72472 5781 72512
rect 5739 72463 5781 72472
rect 5836 72437 5876 74227
rect 5931 74108 5973 74117
rect 5931 74068 5932 74108
rect 5972 74068 5973 74108
rect 5931 74059 5973 74068
rect 5932 73193 5972 74059
rect 5931 73184 5973 73193
rect 5931 73144 5932 73184
rect 5972 73144 5973 73184
rect 5931 73135 5973 73144
rect 6028 73016 6068 73025
rect 5835 72428 5877 72437
rect 5835 72388 5836 72428
rect 5876 72388 5877 72428
rect 5835 72379 5877 72388
rect 5931 72176 5973 72185
rect 5931 72136 5932 72176
rect 5972 72136 5973 72176
rect 5931 72127 5973 72136
rect 5932 72042 5972 72127
rect 5740 72008 5780 72017
rect 5780 71968 5876 72008
rect 5740 71959 5780 71968
rect 5836 71499 5876 71968
rect 5931 71924 5973 71933
rect 5931 71884 5932 71924
rect 5972 71884 5973 71924
rect 5931 71875 5973 71884
rect 5836 71450 5876 71459
rect 5932 70664 5972 71875
rect 6028 71849 6068 72976
rect 6123 72512 6165 72521
rect 6123 72472 6124 72512
rect 6164 72472 6165 72512
rect 6123 72463 6165 72472
rect 6027 71840 6069 71849
rect 6027 71800 6028 71840
rect 6068 71800 6069 71840
rect 6027 71791 6069 71800
rect 6028 71588 6068 71599
rect 6028 71513 6068 71548
rect 6027 71504 6069 71513
rect 6027 71464 6028 71504
rect 6068 71464 6069 71504
rect 6027 71455 6069 71464
rect 6028 70664 6068 70673
rect 5932 70624 6028 70664
rect 6028 69329 6068 70624
rect 6027 69320 6069 69329
rect 6027 69280 6028 69320
rect 6068 69280 6069 69320
rect 6027 69271 6069 69280
rect 5932 69152 5972 69161
rect 5932 68825 5972 69112
rect 6027 69152 6069 69161
rect 6027 69112 6028 69152
rect 6068 69112 6069 69152
rect 6027 69103 6069 69112
rect 6124 69152 6164 72463
rect 6220 71504 6260 74320
rect 6412 73100 6452 75664
rect 6638 75629 6678 75985
rect 6603 75620 6678 75629
rect 6603 75580 6604 75620
rect 6644 75580 6678 75620
rect 6795 75620 6837 75629
rect 6795 75580 6796 75620
rect 6836 75580 6837 75620
rect 6603 75571 6645 75580
rect 6795 75571 6837 75580
rect 6507 75200 6549 75209
rect 6507 75160 6508 75200
rect 6548 75160 6549 75200
rect 6507 75151 6549 75160
rect 6508 75066 6548 75151
rect 6507 74948 6549 74957
rect 6507 74908 6508 74948
rect 6548 74908 6549 74948
rect 6507 74899 6549 74908
rect 6508 74528 6548 74899
rect 6508 74479 6548 74488
rect 6603 74528 6645 74537
rect 6603 74488 6604 74528
rect 6644 74488 6645 74528
rect 6603 74479 6645 74488
rect 6604 74394 6644 74479
rect 6796 73856 6836 75571
rect 6988 75284 7028 76588
rect 7180 76049 7220 76134
rect 7084 76040 7124 76049
rect 7084 75881 7124 76000
rect 7179 76040 7221 76049
rect 7179 76000 7180 76040
rect 7220 76000 7221 76040
rect 7179 75991 7221 76000
rect 7083 75872 7125 75881
rect 7083 75832 7084 75872
rect 7124 75832 7125 75872
rect 7083 75823 7125 75832
rect 6700 73816 6836 73856
rect 6892 75244 7028 75284
rect 6604 73697 6644 73716
rect 6603 73688 6645 73697
rect 6700 73688 6740 73816
rect 6603 73648 6604 73688
rect 6644 73648 6740 73688
rect 6603 73639 6645 73648
rect 6604 73554 6644 73639
rect 6700 73361 6740 73648
rect 6796 73688 6836 73697
rect 6699 73352 6741 73361
rect 6699 73312 6700 73352
rect 6740 73312 6741 73352
rect 6699 73303 6741 73312
rect 6796 73100 6836 73648
rect 6412 73060 6548 73100
rect 6220 71345 6260 71464
rect 6219 71336 6261 71345
rect 6219 71296 6220 71336
rect 6260 71296 6261 71336
rect 6219 71287 6261 71296
rect 6220 70496 6260 70505
rect 6220 69992 6260 70456
rect 6315 70328 6357 70337
rect 6315 70288 6316 70328
rect 6356 70288 6357 70328
rect 6315 70279 6357 70288
rect 6220 69943 6260 69952
rect 6316 69992 6356 70279
rect 6316 69749 6356 69952
rect 6315 69740 6357 69749
rect 6315 69700 6316 69740
rect 6356 69700 6357 69740
rect 6315 69691 6357 69700
rect 6220 69152 6260 69161
rect 6124 69112 6220 69152
rect 5931 68816 5973 68825
rect 5931 68776 5932 68816
rect 5972 68776 5973 68816
rect 5931 68767 5973 68776
rect 6028 68480 6068 69103
rect 6028 68431 6068 68440
rect 6124 68312 6164 69112
rect 6220 69103 6260 69112
rect 6508 68648 6548 73060
rect 6700 73060 6836 73100
rect 6700 72773 6740 73060
rect 6795 72932 6837 72941
rect 6795 72892 6796 72932
rect 6836 72892 6837 72932
rect 6795 72883 6837 72892
rect 6699 72764 6741 72773
rect 6699 72724 6700 72764
rect 6740 72724 6741 72764
rect 6699 72715 6741 72724
rect 6603 72176 6645 72185
rect 6603 72136 6604 72176
rect 6644 72136 6645 72176
rect 6603 72127 6645 72136
rect 6604 70664 6644 72127
rect 6604 70169 6644 70624
rect 6603 70160 6645 70169
rect 6603 70120 6604 70160
rect 6644 70120 6645 70160
rect 6603 70111 6645 70120
rect 6700 69992 6740 72715
rect 6700 69943 6740 69952
rect 6796 69992 6836 72883
rect 6892 71345 6932 75244
rect 7083 75116 7125 75125
rect 7083 75076 7084 75116
rect 7124 75076 7125 75116
rect 7083 75067 7125 75076
rect 7084 74528 7124 75067
rect 7276 74873 7316 76924
rect 7468 76301 7508 79024
rect 7564 77216 7604 79351
rect 7660 78896 7700 80527
rect 7756 79409 7796 81880
rect 7947 81248 7989 81257
rect 7947 81208 7948 81248
rect 7988 81208 7989 81248
rect 7947 81199 7989 81208
rect 7851 80744 7893 80753
rect 7851 80704 7852 80744
rect 7892 80704 7893 80744
rect 7851 80695 7893 80704
rect 7852 80324 7892 80695
rect 7948 80501 7988 81199
rect 7947 80492 7989 80501
rect 7947 80452 7948 80492
rect 7988 80452 7989 80492
rect 7947 80443 7989 80452
rect 8044 80492 8084 80501
rect 7852 80284 7988 80324
rect 7852 79736 7892 79747
rect 7852 79661 7892 79696
rect 7851 79652 7893 79661
rect 7851 79612 7852 79652
rect 7892 79612 7893 79652
rect 7851 79603 7893 79612
rect 7948 79409 7988 80284
rect 8044 79577 8084 80452
rect 8140 79661 8180 84316
rect 8236 84307 8276 84316
rect 8332 83777 8372 85936
rect 8524 84449 8564 85936
rect 8523 84440 8565 84449
rect 8523 84400 8524 84440
rect 8564 84400 8565 84440
rect 8523 84391 8565 84400
rect 8428 84272 8468 84281
rect 8331 83768 8373 83777
rect 8331 83728 8332 83768
rect 8372 83728 8373 83768
rect 8331 83719 8373 83728
rect 8235 83684 8277 83693
rect 8235 83644 8236 83684
rect 8276 83644 8277 83684
rect 8235 83635 8277 83644
rect 8236 83189 8276 83635
rect 8331 83348 8373 83357
rect 8331 83308 8332 83348
rect 8372 83308 8373 83348
rect 8331 83299 8373 83308
rect 8235 83180 8277 83189
rect 8235 83140 8236 83180
rect 8276 83140 8277 83180
rect 8235 83131 8277 83140
rect 8332 82844 8372 83299
rect 8428 83105 8468 84232
rect 8523 84104 8565 84113
rect 8523 84064 8524 84104
rect 8564 84064 8565 84104
rect 8523 84055 8565 84064
rect 8427 83096 8469 83105
rect 8427 83056 8428 83096
rect 8468 83056 8469 83096
rect 8427 83047 8469 83056
rect 8428 82853 8468 83047
rect 8284 82804 8372 82844
rect 8427 82844 8469 82853
rect 8427 82804 8428 82844
rect 8468 82804 8469 82844
rect 8284 82802 8324 82804
rect 8427 82795 8469 82804
rect 8284 82753 8324 82762
rect 8331 82592 8373 82601
rect 8331 82552 8332 82592
rect 8372 82552 8373 82592
rect 8331 82543 8373 82552
rect 8428 82592 8468 82601
rect 8332 82097 8372 82543
rect 8331 82088 8373 82097
rect 8331 82048 8332 82088
rect 8372 82048 8373 82088
rect 8331 82039 8373 82048
rect 8235 80996 8277 81005
rect 8235 80956 8236 80996
rect 8276 80956 8277 80996
rect 8235 80947 8277 80956
rect 8236 79745 8276 80947
rect 8332 80669 8372 82039
rect 8331 80660 8373 80669
rect 8331 80620 8332 80660
rect 8372 80620 8373 80660
rect 8331 80611 8373 80620
rect 8235 79736 8277 79745
rect 8235 79696 8236 79736
rect 8276 79696 8277 79736
rect 8235 79687 8277 79696
rect 8139 79652 8181 79661
rect 8139 79612 8140 79652
rect 8180 79612 8181 79652
rect 8139 79603 8181 79612
rect 8043 79568 8085 79577
rect 8043 79528 8044 79568
rect 8084 79528 8085 79568
rect 8043 79519 8085 79528
rect 7755 79400 7797 79409
rect 7755 79360 7756 79400
rect 7796 79360 7797 79400
rect 7755 79351 7797 79360
rect 7947 79400 7989 79409
rect 7947 79360 7948 79400
rect 7988 79360 7989 79400
rect 7947 79351 7989 79360
rect 8428 79241 8468 82552
rect 8524 80576 8564 84055
rect 8619 83684 8661 83693
rect 8619 83644 8620 83684
rect 8660 83644 8661 83684
rect 8619 83635 8661 83644
rect 8620 83600 8660 83635
rect 8620 83549 8660 83560
rect 8619 83180 8661 83189
rect 8619 83140 8620 83180
rect 8660 83140 8661 83180
rect 8619 83131 8661 83140
rect 8620 82760 8660 83131
rect 8716 83105 8756 85936
rect 8908 84533 8948 85936
rect 8907 84524 8949 84533
rect 8907 84484 8908 84524
rect 8948 84484 8949 84524
rect 8907 84475 8949 84484
rect 9100 84440 9140 85936
rect 9292 85373 9332 85936
rect 9484 85868 9524 85936
rect 9484 85828 9620 85868
rect 9291 85364 9333 85373
rect 9291 85324 9292 85364
rect 9332 85324 9333 85364
rect 9291 85315 9333 85324
rect 9100 84400 9428 84440
rect 9291 84272 9333 84281
rect 9291 84232 9292 84272
rect 9332 84232 9333 84272
rect 9291 84223 9333 84232
rect 9003 83768 9045 83777
rect 9003 83728 9004 83768
rect 9044 83728 9045 83768
rect 9003 83719 9045 83728
rect 9004 83634 9044 83719
rect 9196 83516 9236 83525
rect 9100 83476 9196 83516
rect 8811 83348 8853 83357
rect 8811 83308 8812 83348
rect 8852 83308 8853 83348
rect 8811 83299 8853 83308
rect 8812 83214 8852 83299
rect 8715 83096 8757 83105
rect 8715 83056 8716 83096
rect 8756 83056 8757 83096
rect 8715 83047 8757 83056
rect 8716 82760 8756 82769
rect 8620 82720 8716 82760
rect 8620 81920 8660 82720
rect 8716 82711 8756 82720
rect 8907 82256 8949 82265
rect 8907 82216 8908 82256
rect 8948 82216 8949 82256
rect 8907 82207 8949 82216
rect 8812 82088 8852 82099
rect 8812 82013 8852 82048
rect 8811 82004 8853 82013
rect 8811 81964 8812 82004
rect 8852 81964 8853 82004
rect 8811 81955 8853 81964
rect 8620 81880 8756 81920
rect 8619 80660 8661 80669
rect 8619 80620 8620 80660
rect 8660 80620 8661 80660
rect 8619 80611 8661 80620
rect 8524 80527 8564 80536
rect 8620 80408 8660 80611
rect 8524 80368 8660 80408
rect 8427 79232 8469 79241
rect 7756 79192 8372 79232
rect 7756 79064 7796 79192
rect 7756 79015 7796 79024
rect 7947 79064 7989 79073
rect 7947 79024 7948 79064
rect 7988 79024 7989 79064
rect 7947 79015 7989 79024
rect 8044 79064 8084 79073
rect 8236 79064 8276 79073
rect 7948 78930 7988 79015
rect 7756 78896 7796 78905
rect 7660 78856 7756 78896
rect 7756 78847 7796 78856
rect 7851 78812 7893 78821
rect 7851 78772 7852 78812
rect 7892 78772 7893 78812
rect 7851 78763 7893 78772
rect 7659 78224 7701 78233
rect 7659 78184 7660 78224
rect 7700 78184 7701 78224
rect 7659 78175 7701 78184
rect 7756 78224 7796 78233
rect 7852 78224 7892 78763
rect 8044 78476 8084 79024
rect 8044 78427 8084 78436
rect 8140 79024 8236 79064
rect 7796 78184 7892 78224
rect 7756 78175 7796 78184
rect 7660 78090 7700 78175
rect 7852 77720 7892 77729
rect 8140 77720 8180 79024
rect 8236 79015 8276 79024
rect 8235 78896 8277 78905
rect 8235 78856 8236 78896
rect 8276 78856 8277 78896
rect 8235 78847 8277 78856
rect 8236 78762 8276 78847
rect 8235 78392 8277 78401
rect 8235 78352 8236 78392
rect 8276 78352 8277 78392
rect 8235 78343 8277 78352
rect 7892 77680 8180 77720
rect 7852 77671 7892 77680
rect 7659 77636 7701 77645
rect 7659 77596 7660 77636
rect 7700 77596 7701 77636
rect 7659 77587 7701 77596
rect 7660 77547 7700 77587
rect 7660 77498 7700 77507
rect 8044 77552 8084 77561
rect 8044 77393 8084 77512
rect 8140 77552 8180 77563
rect 8140 77477 8180 77512
rect 8236 77552 8276 78343
rect 8332 77720 8372 79192
rect 8427 79192 8428 79232
rect 8468 79192 8469 79232
rect 8427 79183 8469 79192
rect 8428 79064 8468 79075
rect 8428 78989 8468 79024
rect 8427 78980 8469 78989
rect 8427 78940 8428 78980
rect 8468 78940 8469 78980
rect 8427 78931 8469 78940
rect 8428 78401 8468 78931
rect 8427 78392 8469 78401
rect 8427 78352 8428 78392
rect 8468 78352 8469 78392
rect 8427 78343 8469 78352
rect 8332 77671 8372 77680
rect 8428 78224 8468 78233
rect 8524 78224 8564 80368
rect 8716 79745 8756 81880
rect 8908 81416 8948 82207
rect 9003 81836 9045 81845
rect 9003 81796 9004 81836
rect 9044 81796 9045 81836
rect 9003 81787 9045 81796
rect 9004 81702 9044 81787
rect 9003 81584 9045 81593
rect 9003 81544 9004 81584
rect 9044 81544 9045 81584
rect 9003 81535 9045 81544
rect 8812 81376 8948 81416
rect 8715 79736 8757 79745
rect 8715 79696 8716 79736
rect 8756 79696 8757 79736
rect 8715 79687 8757 79696
rect 8812 79661 8852 81376
rect 9004 81332 9044 81535
rect 8908 81292 9044 81332
rect 8908 81290 8948 81292
rect 8908 81241 8948 81250
rect 9100 81248 9140 83476
rect 9196 83467 9236 83476
rect 9195 82844 9237 82853
rect 9195 82804 9196 82844
rect 9236 82804 9237 82844
rect 9195 82795 9237 82804
rect 9004 81208 9140 81248
rect 9196 82088 9236 82795
rect 9004 81164 9044 81208
rect 8908 81124 9044 81164
rect 8811 79652 8853 79661
rect 8811 79612 8812 79652
rect 8852 79612 8853 79652
rect 8811 79603 8853 79612
rect 8811 79400 8853 79409
rect 8811 79360 8812 79400
rect 8852 79360 8853 79400
rect 8811 79351 8853 79360
rect 8619 79064 8661 79073
rect 8619 79024 8620 79064
rect 8660 79024 8661 79064
rect 8619 79015 8661 79024
rect 8812 79064 8852 79351
rect 8468 78184 8564 78224
rect 8236 77503 8276 77512
rect 8139 77468 8181 77477
rect 8139 77428 8140 77468
rect 8180 77428 8181 77468
rect 8139 77419 8181 77428
rect 8043 77384 8085 77393
rect 8043 77344 8044 77384
rect 8084 77344 8085 77384
rect 8043 77335 8085 77344
rect 7564 77176 8084 77216
rect 7948 76712 7988 76721
rect 7467 76292 7509 76301
rect 7467 76252 7468 76292
rect 7508 76252 7509 76292
rect 7467 76243 7509 76252
rect 7948 76217 7988 76672
rect 8044 76460 8084 77176
rect 8428 76880 8468 78184
rect 8620 77720 8660 79015
rect 8812 78233 8852 79024
rect 8811 78224 8853 78233
rect 8811 78184 8812 78224
rect 8852 78184 8853 78224
rect 8811 78175 8853 78184
rect 8620 77671 8660 77680
rect 8523 77636 8565 77645
rect 8523 77596 8524 77636
rect 8564 77596 8565 77636
rect 8523 77587 8565 77596
rect 8524 77552 8564 77587
rect 8524 77501 8564 77512
rect 8908 77468 8948 81124
rect 9100 81080 9140 81089
rect 9004 81040 9100 81080
rect 9004 80571 9044 81040
rect 9100 81031 9140 81040
rect 9196 80828 9236 82048
rect 9292 81425 9332 84223
rect 9291 81416 9333 81425
rect 9291 81376 9292 81416
rect 9332 81376 9333 81416
rect 9291 81367 9333 81376
rect 9291 81080 9333 81089
rect 9291 81040 9292 81080
rect 9332 81040 9333 81080
rect 9291 81031 9333 81040
rect 9292 80946 9332 81031
rect 9196 80788 9332 80828
rect 9004 80522 9044 80531
rect 9196 80660 9236 80669
rect 9196 79904 9236 80620
rect 9004 79864 9236 79904
rect 9004 78737 9044 79864
rect 9100 79736 9140 79747
rect 9292 79736 9332 80788
rect 9100 79661 9140 79696
rect 9196 79696 9332 79736
rect 9099 79652 9141 79661
rect 9099 79612 9100 79652
rect 9140 79612 9141 79652
rect 9099 79603 9141 79612
rect 9003 78728 9045 78737
rect 9003 78688 9004 78728
rect 9044 78688 9045 78728
rect 9003 78679 9045 78688
rect 9099 78308 9141 78317
rect 9099 78268 9100 78308
rect 9140 78268 9141 78308
rect 9099 78259 9141 78268
rect 9003 77804 9045 77813
rect 9003 77764 9004 77804
rect 9044 77764 9045 77804
rect 9003 77755 9045 77764
rect 9004 77552 9044 77755
rect 9004 77503 9044 77512
rect 8812 77428 8948 77468
rect 8428 76840 8660 76880
rect 8428 76712 8468 76721
rect 8140 76628 8180 76637
rect 8428 76628 8468 76672
rect 8524 76712 8564 76723
rect 8524 76637 8564 76672
rect 8180 76588 8468 76628
rect 8523 76628 8565 76637
rect 8523 76588 8524 76628
rect 8564 76588 8565 76628
rect 8140 76579 8180 76588
rect 8523 76579 8565 76588
rect 8044 76420 8276 76460
rect 7371 76208 7413 76217
rect 7371 76168 7372 76208
rect 7412 76168 7413 76208
rect 7371 76159 7413 76168
rect 7947 76208 7989 76217
rect 7947 76168 7948 76208
rect 7988 76168 7989 76208
rect 7947 76159 7989 76168
rect 7372 76074 7412 76159
rect 7851 76124 7893 76133
rect 7851 76084 7852 76124
rect 7892 76084 7893 76124
rect 7851 76075 7893 76084
rect 7564 76040 7604 76049
rect 7564 74957 7604 76000
rect 7660 76040 7700 76049
rect 7852 76040 7892 76075
rect 7700 76000 7852 76025
rect 7660 75985 7892 76000
rect 7948 76040 7988 76049
rect 7948 75881 7988 76000
rect 8043 76040 8085 76049
rect 8043 76000 8044 76040
rect 8084 76000 8085 76040
rect 8043 75991 8085 76000
rect 8140 76040 8180 76049
rect 8044 75906 8084 75991
rect 7947 75872 7989 75881
rect 7947 75832 7948 75872
rect 7988 75832 7989 75872
rect 7947 75823 7989 75832
rect 8140 75536 8180 76000
rect 8044 75496 8180 75536
rect 7948 75452 7988 75461
rect 7660 75412 7948 75452
rect 7563 74948 7605 74957
rect 7563 74908 7564 74948
rect 7604 74908 7605 74948
rect 7563 74899 7605 74908
rect 7275 74864 7317 74873
rect 7275 74824 7276 74864
rect 7316 74824 7317 74864
rect 7275 74815 7317 74824
rect 7084 74479 7124 74488
rect 7276 74033 7316 74815
rect 7660 74528 7700 75412
rect 7948 75403 7988 75412
rect 7756 75200 7796 75209
rect 7796 75160 7892 75200
rect 7756 75151 7796 75160
rect 7755 74612 7797 74621
rect 7755 74572 7756 74612
rect 7796 74572 7797 74612
rect 7755 74563 7797 74572
rect 7612 74518 7700 74528
rect 7652 74488 7700 74518
rect 7756 74478 7796 74563
rect 7612 74469 7652 74478
rect 7852 74285 7892 75160
rect 8044 74537 8084 75496
rect 8139 75368 8181 75377
rect 8139 75328 8140 75368
rect 8180 75328 8181 75368
rect 8139 75319 8181 75328
rect 8140 75200 8180 75319
rect 8140 75151 8180 75160
rect 8043 74528 8085 74537
rect 8043 74488 8044 74528
rect 8084 74488 8085 74528
rect 8043 74479 8085 74488
rect 7851 74276 7893 74285
rect 7851 74236 7852 74276
rect 7892 74236 7893 74276
rect 7851 74227 7893 74236
rect 7275 74024 7317 74033
rect 7275 73984 7276 74024
rect 7316 73984 7317 74024
rect 7275 73975 7317 73984
rect 7084 73856 7124 73865
rect 7124 73816 7316 73856
rect 7084 73807 7124 73816
rect 6988 73688 7028 73697
rect 6988 73529 7028 73648
rect 7083 73688 7125 73697
rect 7083 73648 7084 73688
rect 7124 73648 7125 73688
rect 7083 73639 7125 73648
rect 7276 73688 7316 73816
rect 7660 73697 7700 73782
rect 7276 73639 7316 73648
rect 7372 73688 7412 73697
rect 7084 73554 7124 73639
rect 7372 73529 7412 73648
rect 7467 73688 7509 73697
rect 7467 73648 7468 73688
rect 7508 73648 7509 73688
rect 7467 73639 7509 73648
rect 7564 73688 7604 73697
rect 6987 73520 7029 73529
rect 6987 73480 6988 73520
rect 7028 73480 7029 73520
rect 6987 73471 7029 73480
rect 7371 73520 7413 73529
rect 7371 73480 7372 73520
rect 7412 73480 7413 73520
rect 7371 73471 7413 73480
rect 7083 73352 7125 73361
rect 7083 73312 7084 73352
rect 7124 73312 7125 73352
rect 7083 73303 7125 73312
rect 6891 71336 6933 71345
rect 6891 71296 6892 71336
rect 6932 71296 6933 71336
rect 6891 71287 6933 71296
rect 6892 70757 6932 71287
rect 6891 70748 6933 70757
rect 6891 70708 6892 70748
rect 6932 70708 6933 70748
rect 6891 70699 6933 70708
rect 6891 70160 6933 70169
rect 6891 70120 6892 70160
rect 6932 70120 6933 70160
rect 6891 70111 6933 70120
rect 6796 69943 6836 69952
rect 6699 69320 6741 69329
rect 6699 69280 6700 69320
rect 6740 69280 6741 69320
rect 6699 69271 6741 69280
rect 6028 68272 6164 68312
rect 6316 68608 6548 68648
rect 5739 67976 5781 67985
rect 5739 67936 5740 67976
rect 5780 67936 5781 67976
rect 5739 67927 5781 67936
rect 5643 67808 5685 67817
rect 5643 67768 5644 67808
rect 5684 67768 5685 67808
rect 5643 67759 5685 67768
rect 5740 67640 5780 67927
rect 5740 67591 5780 67600
rect 5739 66464 5781 66473
rect 5739 66424 5740 66464
rect 5780 66424 5781 66464
rect 5739 66415 5781 66424
rect 5740 65624 5780 66415
rect 5931 66128 5973 66137
rect 5931 66088 5932 66128
rect 5972 66088 5973 66128
rect 5931 66079 5973 66088
rect 5835 65960 5877 65969
rect 5835 65920 5836 65960
rect 5876 65920 5877 65960
rect 5835 65911 5877 65920
rect 5740 65575 5780 65584
rect 5644 65456 5684 65467
rect 5644 65381 5684 65416
rect 5836 65456 5876 65911
rect 5836 65407 5876 65416
rect 5932 65456 5972 66079
rect 5932 65407 5972 65416
rect 5643 65372 5685 65381
rect 5643 65332 5644 65372
rect 5684 65332 5691 65372
rect 5643 65323 5691 65332
rect 5651 65288 5691 65323
rect 5835 65288 5877 65297
rect 5651 65248 5780 65288
rect 5548 65164 5684 65204
rect 5451 64700 5493 64709
rect 5451 64660 5452 64700
rect 5492 64660 5493 64700
rect 5451 64651 5493 64660
rect 5451 64448 5493 64457
rect 5451 64408 5452 64448
rect 5492 64408 5493 64448
rect 5451 64399 5493 64408
rect 5452 64314 5492 64399
rect 5451 63692 5493 63701
rect 5451 63652 5452 63692
rect 5492 63652 5493 63692
rect 5451 63643 5493 63652
rect 5452 63188 5492 63643
rect 5644 63272 5684 65164
rect 5740 65045 5780 65248
rect 5835 65248 5836 65288
rect 5876 65248 5877 65288
rect 5835 65239 5877 65248
rect 5739 65036 5781 65045
rect 5739 64996 5740 65036
rect 5780 64996 5781 65036
rect 5739 64987 5781 64996
rect 5740 64616 5780 64625
rect 5740 64457 5780 64576
rect 5836 64616 5876 65239
rect 5931 64700 5973 64709
rect 5931 64660 5932 64700
rect 5972 64660 5973 64700
rect 5931 64651 5973 64660
rect 5739 64448 5781 64457
rect 5739 64408 5740 64448
rect 5780 64408 5781 64448
rect 5739 64399 5781 64408
rect 5836 63953 5876 64576
rect 5835 63944 5877 63953
rect 5835 63904 5836 63944
rect 5876 63904 5877 63944
rect 5835 63895 5877 63904
rect 5932 63944 5972 64651
rect 6028 64280 6068 68272
rect 6220 68228 6260 68237
rect 6123 67808 6165 67817
rect 6123 67768 6124 67808
rect 6164 67768 6165 67808
rect 6123 67759 6165 67768
rect 6124 65456 6164 67759
rect 6220 67654 6260 68188
rect 6220 67605 6260 67614
rect 6316 67052 6356 68608
rect 6507 68480 6549 68489
rect 6507 68440 6508 68480
rect 6548 68440 6549 68480
rect 6507 68431 6549 68440
rect 6508 68346 6548 68431
rect 6412 67472 6452 67481
rect 6452 67432 6548 67472
rect 6412 67423 6452 67432
rect 6220 67012 6356 67052
rect 6220 65456 6260 67012
rect 6508 66977 6548 67432
rect 6412 66968 6452 66977
rect 6316 66928 6412 66968
rect 6316 66128 6356 66928
rect 6412 66919 6452 66928
rect 6507 66968 6549 66977
rect 6507 66928 6508 66968
rect 6548 66928 6549 66968
rect 6507 66919 6549 66928
rect 6508 66809 6548 66919
rect 6507 66800 6549 66809
rect 6507 66760 6508 66800
rect 6548 66760 6549 66800
rect 6507 66751 6549 66760
rect 6604 66716 6644 66725
rect 6604 66557 6644 66676
rect 6603 66548 6645 66557
rect 6603 66508 6604 66548
rect 6644 66508 6645 66548
rect 6603 66499 6645 66508
rect 6507 66464 6549 66473
rect 6507 66424 6508 66464
rect 6548 66424 6549 66464
rect 6507 66415 6549 66424
rect 6411 66212 6453 66221
rect 6411 66172 6412 66212
rect 6452 66172 6453 66212
rect 6411 66163 6453 66172
rect 6316 65633 6356 66088
rect 6315 65624 6357 65633
rect 6315 65584 6316 65624
rect 6356 65584 6357 65624
rect 6315 65575 6357 65584
rect 6412 65540 6452 66163
rect 6508 66128 6548 66415
rect 6700 66389 6740 69271
rect 6892 69077 6932 70111
rect 6891 69068 6933 69077
rect 6891 69028 6892 69068
rect 6932 69028 6933 69068
rect 6891 69019 6933 69028
rect 7084 67481 7124 73303
rect 7276 73016 7316 73025
rect 7180 72976 7276 73016
rect 7180 72353 7220 72976
rect 7276 72967 7316 72976
rect 7372 72428 7412 73471
rect 7468 73184 7508 73639
rect 7564 73193 7604 73648
rect 7659 73688 7701 73697
rect 7659 73648 7660 73688
rect 7700 73648 7701 73688
rect 7659 73639 7701 73648
rect 7815 73688 7855 73697
rect 8044 73688 8084 73697
rect 7855 73648 8044 73688
rect 7815 73639 7855 73648
rect 8044 73639 8084 73648
rect 8139 73688 8181 73697
rect 8139 73648 8140 73688
rect 8180 73648 8181 73688
rect 8139 73639 8181 73648
rect 8140 73554 8180 73639
rect 8236 73529 8276 76420
rect 8427 76376 8469 76385
rect 8427 76336 8428 76376
rect 8468 76336 8469 76376
rect 8427 76327 8469 76336
rect 8331 76292 8373 76301
rect 8331 76252 8332 76292
rect 8372 76252 8373 76292
rect 8331 76243 8373 76252
rect 8332 75377 8372 76243
rect 8331 75368 8373 75377
rect 8331 75328 8332 75368
rect 8372 75328 8373 75368
rect 8331 75319 8373 75328
rect 8428 75200 8468 76327
rect 8332 75160 8468 75200
rect 7659 73520 7701 73529
rect 7659 73480 7660 73520
rect 7700 73480 7701 73520
rect 7659 73471 7701 73480
rect 7851 73520 7893 73529
rect 7851 73480 7852 73520
rect 7892 73480 7893 73520
rect 7851 73471 7893 73480
rect 8235 73520 8277 73529
rect 8235 73480 8236 73520
rect 8276 73480 8277 73520
rect 8235 73471 8277 73480
rect 7660 73386 7700 73471
rect 7468 73016 7508 73144
rect 7563 73184 7605 73193
rect 7563 73144 7564 73184
rect 7604 73144 7605 73184
rect 7563 73135 7605 73144
rect 7660 73016 7700 73025
rect 7468 72976 7660 73016
rect 7660 72967 7700 72976
rect 7755 73016 7797 73025
rect 7755 72976 7756 73016
rect 7796 72976 7797 73016
rect 7755 72967 7797 72976
rect 7756 72882 7796 72967
rect 7852 72941 7892 73471
rect 8139 73436 8181 73445
rect 8139 73396 8140 73436
rect 8180 73396 8181 73436
rect 8139 73387 8181 73396
rect 7948 73193 7988 73278
rect 7947 73184 7989 73193
rect 7947 73144 7948 73184
rect 7988 73144 7989 73184
rect 7947 73135 7989 73144
rect 7851 72932 7893 72941
rect 7851 72892 7852 72932
rect 7892 72892 7893 72932
rect 7851 72883 7893 72892
rect 7372 72379 7412 72388
rect 7179 72344 7221 72353
rect 7179 72304 7180 72344
rect 7220 72304 7221 72344
rect 7179 72295 7221 72304
rect 7180 72176 7220 72295
rect 7180 72127 7220 72136
rect 7756 72176 7796 72185
rect 7852 72176 7892 72883
rect 7796 72136 7892 72176
rect 7756 72127 7796 72136
rect 7755 72008 7797 72017
rect 7755 71968 7756 72008
rect 7796 71968 7797 72008
rect 7755 71959 7797 71968
rect 7659 71924 7701 71933
rect 7659 71884 7660 71924
rect 7700 71884 7701 71924
rect 7659 71875 7701 71884
rect 7563 71840 7605 71849
rect 7563 71800 7564 71840
rect 7604 71800 7605 71840
rect 7563 71791 7605 71800
rect 7467 71588 7509 71597
rect 7467 71548 7468 71588
rect 7508 71548 7509 71588
rect 7467 71539 7509 71548
rect 7371 71504 7413 71513
rect 7371 71464 7372 71504
rect 7412 71464 7413 71504
rect 7371 71455 7413 71464
rect 7468 71504 7508 71539
rect 7275 69992 7317 70001
rect 7275 69952 7276 69992
rect 7316 69952 7317 69992
rect 7275 69943 7317 69952
rect 7276 69413 7316 69943
rect 7275 69404 7317 69413
rect 7275 69364 7276 69404
rect 7316 69364 7317 69404
rect 7275 69355 7317 69364
rect 7275 68480 7317 68489
rect 7275 68440 7276 68480
rect 7316 68440 7317 68480
rect 7275 68431 7317 68440
rect 7083 67472 7125 67481
rect 7083 67432 7084 67472
rect 7124 67432 7125 67472
rect 7083 67423 7125 67432
rect 6879 66977 6919 67028
rect 6843 66971 6919 66977
rect 6843 66968 6879 66971
rect 6843 66928 6844 66968
rect 6884 66928 6919 66931
rect 6843 66922 6919 66928
rect 7180 66968 7220 66977
rect 7276 66968 7316 68431
rect 7372 67649 7412 71455
rect 7468 71453 7508 71464
rect 7564 70001 7604 71791
rect 7660 71672 7700 71875
rect 7660 71623 7700 71632
rect 7659 71084 7701 71093
rect 7659 71044 7660 71084
rect 7700 71044 7701 71084
rect 7659 71035 7701 71044
rect 7563 69992 7605 70001
rect 7563 69952 7564 69992
rect 7604 69952 7605 69992
rect 7563 69943 7605 69952
rect 7660 69572 7700 71035
rect 7756 70169 7796 71959
rect 7947 71924 7989 71933
rect 7947 71884 7948 71924
rect 7988 71884 7989 71924
rect 7947 71875 7989 71884
rect 7948 71504 7988 71875
rect 7948 71455 7988 71464
rect 8044 71504 8084 71513
rect 8044 71000 8084 71464
rect 7948 70960 8084 71000
rect 7852 70664 7892 70673
rect 7755 70160 7797 70169
rect 7755 70120 7756 70160
rect 7796 70120 7797 70160
rect 7755 70111 7797 70120
rect 7564 69532 7700 69572
rect 7756 69978 7796 69987
rect 7467 69320 7509 69329
rect 7467 69280 7468 69320
rect 7508 69280 7509 69320
rect 7467 69271 7509 69280
rect 7468 69152 7508 69271
rect 7468 69103 7508 69112
rect 7364 67640 7412 67649
rect 7364 67600 7365 67640
rect 7364 67591 7412 67600
rect 7467 67640 7509 67649
rect 7467 67600 7468 67640
rect 7508 67600 7509 67640
rect 7467 67591 7509 67600
rect 7468 67506 7508 67591
rect 7371 67472 7413 67481
rect 7371 67432 7372 67472
rect 7412 67432 7413 67472
rect 7371 67423 7413 67432
rect 7372 67229 7412 67423
rect 7371 67220 7413 67229
rect 7371 67180 7372 67220
rect 7412 67180 7413 67220
rect 7371 67171 7413 67180
rect 7220 66928 7316 66968
rect 6843 66919 6885 66922
rect 7180 66919 7220 66928
rect 6988 66716 7028 66725
rect 7028 66676 7220 66716
rect 6988 66667 7028 66676
rect 7083 66548 7125 66557
rect 7083 66508 7084 66548
rect 7124 66508 7125 66548
rect 7083 66499 7125 66508
rect 6699 66380 6741 66389
rect 6699 66340 6700 66380
rect 6740 66340 6741 66380
rect 6699 66331 6741 66340
rect 7084 66221 7124 66499
rect 7083 66212 7125 66221
rect 7083 66172 7084 66212
rect 7124 66172 7125 66212
rect 7083 66163 7125 66172
rect 7084 66157 7124 66163
rect 6690 66137 6730 66146
rect 6508 66097 6690 66128
rect 6508 66088 6730 66097
rect 6796 66128 6836 66137
rect 6796 66044 6836 66088
rect 6604 66004 6836 66044
rect 6988 66128 7028 66137
rect 6507 65960 6549 65969
rect 6604 65960 6644 66004
rect 6988 65969 7028 66088
rect 7084 66077 7124 66117
rect 7180 66137 7220 66676
rect 7180 66128 7225 66137
rect 7180 66088 7185 66128
rect 7185 66079 7225 66088
rect 6507 65920 6508 65960
rect 6548 65920 6644 65960
rect 6987 65960 7029 65969
rect 6987 65920 6988 65960
rect 7028 65920 7029 65960
rect 6507 65911 6549 65920
rect 6987 65911 7029 65920
rect 7084 65960 7124 65969
rect 7276 65960 7316 66928
rect 6508 65826 6548 65911
rect 6795 65876 6837 65885
rect 6795 65836 6796 65876
rect 6836 65836 6837 65876
rect 6795 65827 6837 65836
rect 6412 65500 6644 65540
rect 6220 65416 6452 65456
rect 6124 64961 6164 65416
rect 6412 65045 6452 65416
rect 6507 65372 6549 65381
rect 6507 65332 6508 65372
rect 6548 65332 6549 65372
rect 6507 65323 6549 65332
rect 6219 65036 6261 65045
rect 6219 64996 6220 65036
rect 6260 64996 6261 65036
rect 6219 64987 6261 64996
rect 6411 65036 6453 65045
rect 6411 64996 6412 65036
rect 6452 64996 6453 65036
rect 6411 64987 6453 64996
rect 6123 64952 6165 64961
rect 6123 64912 6124 64952
rect 6164 64912 6165 64952
rect 6123 64903 6165 64912
rect 6220 64700 6260 64987
rect 6412 64793 6452 64987
rect 6411 64784 6453 64793
rect 6411 64744 6412 64784
rect 6452 64744 6453 64784
rect 6411 64735 6453 64744
rect 6220 64651 6260 64660
rect 6315 64616 6357 64625
rect 6315 64576 6316 64616
rect 6356 64576 6357 64616
rect 6315 64567 6357 64576
rect 6316 64482 6356 64567
rect 6219 64364 6261 64373
rect 6219 64324 6220 64364
rect 6260 64324 6261 64364
rect 6219 64315 6261 64324
rect 6411 64364 6453 64373
rect 6411 64324 6412 64364
rect 6452 64324 6453 64364
rect 6411 64315 6453 64324
rect 6028 64240 6164 64280
rect 6027 63944 6069 63953
rect 5932 63904 6028 63944
rect 6068 63904 6069 63944
rect 5932 63785 5972 63904
rect 6027 63895 6069 63904
rect 6028 63810 6068 63895
rect 5931 63776 5973 63785
rect 5931 63736 5932 63776
rect 5972 63736 5973 63776
rect 5931 63727 5973 63736
rect 6124 63272 6164 64240
rect 6220 63356 6260 64315
rect 6220 63316 6356 63356
rect 5644 63232 5691 63272
rect 6124 63232 6260 63272
rect 5452 63148 5588 63188
rect 5548 63146 5588 63148
rect 5548 63097 5588 63106
rect 5651 63104 5691 63232
rect 5644 63064 5691 63104
rect 6028 63104 6068 63113
rect 5451 62768 5493 62777
rect 5451 62728 5452 62768
rect 5492 62728 5493 62768
rect 5451 62719 5493 62728
rect 5452 59828 5492 62719
rect 5452 59788 5588 59828
rect 4779 59324 4821 59333
rect 4779 59284 4780 59324
rect 4820 59284 4821 59324
rect 4779 59275 4821 59284
rect 5163 59324 5205 59333
rect 5163 59284 5164 59324
rect 5204 59284 5205 59324
rect 5163 59275 5205 59284
rect 5355 59324 5397 59333
rect 5355 59284 5356 59324
rect 5396 59284 5397 59324
rect 5355 59275 5397 59284
rect 4971 59240 5013 59249
rect 4971 59200 4972 59240
rect 5012 59200 5013 59240
rect 4971 59191 5013 59200
rect 4972 59106 5012 59191
rect 5164 59190 5204 59275
rect 4300 59032 4628 59072
rect 4300 58568 4340 58579
rect 4300 58493 4340 58528
rect 4299 58484 4341 58493
rect 4299 58444 4300 58484
rect 4340 58444 4341 58484
rect 4299 58435 4341 58444
rect 4300 57989 4340 58435
rect 4492 58400 4532 58409
rect 4492 57989 4532 58360
rect 4299 57980 4341 57989
rect 4299 57940 4300 57980
rect 4340 57940 4341 57980
rect 4299 57931 4341 57940
rect 4491 57980 4533 57989
rect 4491 57940 4492 57980
rect 4532 57940 4533 57980
rect 4491 57931 4533 57940
rect 4588 57896 4628 59032
rect 4683 58568 4725 58577
rect 4683 58528 4684 58568
rect 4724 58528 4725 58568
rect 4683 58519 4725 58528
rect 4684 58434 4724 58519
rect 4928 58232 5296 58241
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 4928 58183 5296 58192
rect 5067 57980 5109 57989
rect 5067 57940 5068 57980
rect 5108 57940 5109 57980
rect 5067 57931 5109 57940
rect 5260 57980 5300 57989
rect 4588 57847 4628 57856
rect 5068 57891 5108 57931
rect 5068 57842 5108 57851
rect 4299 57728 4341 57737
rect 4299 57688 4300 57728
rect 4340 57688 4341 57728
rect 4299 57679 4341 57688
rect 4148 57016 4244 57056
rect 4108 57007 4148 57016
rect 4300 56888 4340 57679
rect 4396 57056 4436 57065
rect 4436 57016 4628 57056
rect 4396 57007 4436 57016
rect 4012 56848 4340 56888
rect 3764 56344 3860 56384
rect 3724 56141 3764 56344
rect 4108 56300 4148 56309
rect 4108 56141 4148 56260
rect 4203 56300 4245 56309
rect 4203 56260 4204 56300
rect 4244 56260 4245 56300
rect 4203 56251 4245 56260
rect 4204 56166 4244 56251
rect 3723 56132 3765 56141
rect 3723 56092 3724 56132
rect 3764 56092 3765 56132
rect 3723 56083 3765 56092
rect 4107 56132 4149 56141
rect 4107 56092 4108 56132
rect 4148 56092 4149 56132
rect 4107 56083 4149 56092
rect 3688 55964 4056 55973
rect 4300 55964 4340 56848
rect 4491 56132 4533 56141
rect 4491 56092 4492 56132
rect 4532 56092 4533 56132
rect 4491 56083 4533 56092
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 3688 55915 4056 55924
rect 4108 55924 4340 55964
rect 3532 55756 3668 55796
rect 3436 55579 3476 55588
rect 3148 54823 3188 54832
rect 3244 55420 3380 55460
rect 2955 54704 2997 54713
rect 2955 54664 2956 54704
rect 2996 54664 2997 54704
rect 2955 54655 2997 54664
rect 2859 54284 2901 54293
rect 2859 54244 2860 54284
rect 2900 54244 2901 54284
rect 2859 54235 2901 54244
rect 2668 52816 2804 52856
rect 2571 52772 2613 52781
rect 2571 52732 2572 52772
rect 2612 52732 2613 52772
rect 2571 52723 2613 52732
rect 2379 52184 2421 52193
rect 2379 52144 2380 52184
rect 2420 52144 2421 52184
rect 2379 52135 2421 52144
rect 2379 51932 2421 51941
rect 2379 51892 2380 51932
rect 2420 51892 2421 51932
rect 2379 51883 2421 51892
rect 2380 50336 2420 51883
rect 2476 51008 2516 51017
rect 2476 50513 2516 50968
rect 2475 50504 2517 50513
rect 2475 50464 2476 50504
rect 2516 50464 2517 50504
rect 2475 50455 2517 50464
rect 2380 50296 2516 50336
rect 2476 50252 2516 50296
rect 2284 50212 2420 50252
rect 2092 50203 2132 50212
rect 2284 50084 2324 50093
rect 1996 50044 2284 50084
rect 1900 49505 1940 50044
rect 2284 50035 2324 50044
rect 1995 49916 2037 49925
rect 1995 49876 1996 49916
rect 2036 49876 2037 49916
rect 1995 49867 2037 49876
rect 1899 49496 1941 49505
rect 1899 49456 1900 49496
rect 1940 49456 1941 49496
rect 1899 49447 1941 49456
rect 1900 48992 1940 49001
rect 1804 48952 1900 48992
rect 1900 48943 1940 48952
rect 1708 48691 1748 48700
rect 1556 48196 1652 48236
rect 1516 48187 1556 48196
rect 1707 48068 1749 48077
rect 1707 48028 1708 48068
rect 1748 48028 1749 48068
rect 1707 48019 1749 48028
rect 1708 47934 1748 48019
rect 1803 47900 1845 47909
rect 1803 47860 1804 47900
rect 1844 47860 1845 47900
rect 1803 47851 1845 47860
rect 1419 47816 1461 47825
rect 1419 47776 1420 47816
rect 1460 47776 1461 47816
rect 1419 47767 1461 47776
rect 1324 47608 1652 47648
rect 1516 47060 1556 47069
rect 1228 46472 1268 46481
rect 1268 46432 1364 46472
rect 1228 46423 1268 46432
rect 1324 46313 1364 46432
rect 1419 46388 1461 46397
rect 1419 46348 1420 46388
rect 1460 46348 1461 46388
rect 1419 46339 1461 46348
rect 1323 46304 1365 46313
rect 1323 46264 1324 46304
rect 1364 46264 1365 46304
rect 1323 46255 1365 46264
rect 1420 45044 1460 46339
rect 1516 46145 1556 47020
rect 1515 46136 1557 46145
rect 1515 46096 1516 46136
rect 1556 46096 1557 46136
rect 1515 46087 1557 46096
rect 1516 45548 1556 45557
rect 1612 45548 1652 47608
rect 1707 47228 1749 47237
rect 1707 47188 1708 47228
rect 1748 47188 1749 47228
rect 1707 47179 1749 47188
rect 1708 47094 1748 47179
rect 1708 45716 1748 45725
rect 1804 45716 1844 47851
rect 1900 47816 1940 47825
rect 1900 47489 1940 47776
rect 1899 47480 1941 47489
rect 1899 47440 1900 47480
rect 1940 47440 1941 47480
rect 1899 47431 1941 47440
rect 1899 47312 1941 47321
rect 1899 47272 1900 47312
rect 1940 47272 1941 47312
rect 1899 47263 1941 47272
rect 1900 47178 1940 47263
rect 1996 46556 2036 49867
rect 2092 48740 2132 48749
rect 2132 48700 2228 48740
rect 2092 48691 2132 48700
rect 2092 48068 2132 48077
rect 2092 47741 2132 48028
rect 2091 47732 2133 47741
rect 2091 47692 2092 47732
rect 2132 47692 2133 47732
rect 2091 47683 2133 47692
rect 2188 47489 2228 48700
rect 2380 48068 2420 50212
rect 2476 50203 2516 50212
rect 2475 50000 2517 50009
rect 2475 49960 2476 50000
rect 2516 49960 2517 50000
rect 2475 49951 2517 49960
rect 2476 48665 2516 49951
rect 2572 49496 2612 52723
rect 2668 51092 2708 52816
rect 3244 52781 3284 55420
rect 3531 55208 3573 55217
rect 3531 55168 3532 55208
rect 3572 55168 3573 55208
rect 3531 55159 3573 55168
rect 3532 54713 3572 55159
rect 3628 54965 3668 55756
rect 3627 54956 3669 54965
rect 3627 54916 3628 54956
rect 3668 54916 3669 54956
rect 3627 54907 3669 54916
rect 3628 54872 3668 54907
rect 3628 54822 3668 54832
rect 4108 54872 4148 55924
rect 4203 55376 4245 55385
rect 4203 55336 4204 55376
rect 4244 55336 4245 55376
rect 4203 55327 4245 55336
rect 4108 54823 4148 54832
rect 4204 54872 4244 55327
rect 4204 54823 4244 54832
rect 3724 54788 3764 54797
rect 3339 54704 3381 54713
rect 3531 54704 3573 54713
rect 3339 54664 3340 54704
rect 3380 54664 3381 54704
rect 3339 54655 3381 54664
rect 3436 54664 3532 54704
rect 3572 54664 3573 54704
rect 3340 54041 3380 54655
rect 3339 54032 3381 54041
rect 3339 53992 3340 54032
rect 3380 53992 3381 54032
rect 3339 53983 3381 53992
rect 3340 53360 3380 53983
rect 3340 53311 3380 53320
rect 3243 52772 3285 52781
rect 3243 52732 3244 52772
rect 3284 52732 3285 52772
rect 3243 52723 3285 52732
rect 2764 52520 2804 52529
rect 2764 51848 2804 52480
rect 3244 52520 3284 52529
rect 2956 52436 2996 52445
rect 3244 52436 3284 52480
rect 3339 52520 3381 52529
rect 3339 52480 3340 52520
rect 3380 52480 3381 52520
rect 3339 52471 3381 52480
rect 2996 52396 3284 52436
rect 2956 52387 2996 52396
rect 3340 52386 3380 52471
rect 3436 52268 3476 54664
rect 3531 54655 3573 54664
rect 3724 54629 3764 54748
rect 3723 54620 3765 54629
rect 3723 54580 3724 54620
rect 3764 54580 3765 54620
rect 3723 54571 3765 54580
rect 3688 54452 4056 54461
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 3688 54403 4056 54412
rect 3819 54284 3861 54293
rect 3819 54244 3820 54284
rect 3860 54244 3861 54284
rect 3819 54235 3861 54244
rect 3820 54032 3860 54235
rect 4011 54200 4053 54209
rect 4011 54160 4012 54200
rect 4052 54160 4053 54200
rect 4011 54151 4053 54160
rect 4012 54066 4052 54151
rect 3531 53444 3573 53453
rect 3531 53404 3532 53444
rect 3572 53404 3573 53444
rect 3531 53395 3573 53404
rect 3532 53310 3572 53395
rect 3820 53108 3860 53992
rect 4396 54032 4436 54041
rect 4011 53444 4053 53453
rect 4011 53404 4012 53444
rect 4052 53404 4053 53444
rect 4011 53395 4053 53404
rect 4012 53360 4052 53395
rect 4012 53309 4052 53320
rect 4108 53360 4148 53369
rect 2764 51773 2804 51808
rect 3148 52228 3476 52268
rect 3532 53068 3860 53108
rect 3148 51848 3188 52228
rect 2763 51764 2805 51773
rect 2763 51724 2764 51764
rect 2804 51724 2805 51764
rect 2763 51715 2805 51724
rect 2955 51680 2997 51689
rect 2955 51640 2956 51680
rect 2996 51640 2997 51680
rect 2955 51631 2997 51640
rect 2956 51546 2996 51631
rect 3051 51092 3093 51101
rect 2668 51052 2996 51092
rect 2668 50840 2708 50849
rect 2860 50840 2900 50849
rect 2708 50800 2804 50840
rect 2668 50791 2708 50800
rect 2667 50336 2709 50345
rect 2667 50296 2668 50336
rect 2708 50296 2709 50336
rect 2667 50287 2709 50296
rect 2668 50202 2708 50287
rect 2764 49496 2804 50800
rect 2860 50177 2900 50800
rect 2859 50168 2901 50177
rect 2859 50128 2860 50168
rect 2900 50128 2901 50168
rect 2859 50119 2901 50128
rect 2572 49456 2708 49496
rect 2668 49328 2708 49456
rect 2764 49447 2804 49456
rect 2860 49496 2900 49505
rect 2860 49328 2900 49456
rect 2668 49288 2900 49328
rect 2571 48824 2613 48833
rect 2571 48784 2572 48824
rect 2612 48784 2613 48824
rect 2571 48775 2613 48784
rect 2572 48690 2612 48775
rect 2475 48656 2517 48665
rect 2475 48616 2476 48656
rect 2516 48616 2517 48656
rect 2475 48607 2517 48616
rect 2476 48068 2516 48077
rect 2380 48028 2476 48068
rect 2476 48019 2516 48028
rect 2764 47984 2804 47993
rect 2284 47816 2324 47825
rect 2187 47480 2229 47489
rect 2187 47440 2188 47480
rect 2228 47440 2229 47480
rect 2187 47431 2229 47440
rect 2284 46817 2324 47776
rect 2283 46808 2325 46817
rect 2283 46768 2284 46808
rect 2324 46768 2325 46808
rect 2283 46759 2325 46768
rect 2475 46640 2517 46649
rect 2475 46600 2476 46640
rect 2516 46600 2517 46640
rect 2475 46591 2517 46600
rect 2668 46640 2708 46649
rect 2764 46640 2804 47944
rect 2860 47984 2900 49288
rect 2860 46985 2900 47944
rect 2859 46976 2901 46985
rect 2859 46936 2860 46976
rect 2900 46936 2901 46976
rect 2859 46927 2901 46936
rect 2708 46600 2804 46640
rect 2668 46591 2708 46600
rect 1996 46516 2324 46556
rect 2284 45968 2324 46516
rect 2476 46472 2516 46591
rect 2860 46472 2900 46927
rect 2284 45919 2324 45928
rect 2380 46432 2476 46472
rect 1748 45676 1844 45716
rect 2092 45716 2132 45725
rect 1708 45667 1748 45676
rect 1995 45632 2037 45641
rect 1995 45592 1996 45632
rect 2036 45592 2037 45632
rect 1995 45583 2037 45592
rect 1900 45548 1940 45557
rect 1612 45508 1900 45548
rect 1516 45137 1556 45508
rect 1900 45499 1940 45508
rect 1611 45380 1653 45389
rect 1611 45340 1612 45380
rect 1652 45340 1653 45380
rect 1611 45331 1653 45340
rect 1515 45128 1557 45137
rect 1515 45088 1516 45128
rect 1556 45088 1557 45128
rect 1515 45079 1557 45088
rect 1420 44995 1460 45004
rect 1612 44960 1652 45331
rect 1803 45044 1845 45053
rect 1803 45004 1804 45044
rect 1844 45004 1845 45044
rect 1803 44995 1845 45004
rect 1516 44920 1652 44960
rect 1228 44792 1268 44801
rect 1228 44465 1268 44752
rect 1227 44456 1269 44465
rect 1227 44416 1228 44456
rect 1268 44416 1269 44456
rect 1227 44407 1269 44416
rect 1228 41936 1268 41945
rect 1268 41896 1364 41936
rect 1228 41887 1268 41896
rect 1227 41264 1269 41273
rect 1227 41224 1228 41264
rect 1268 41224 1269 41264
rect 1227 41215 1269 41224
rect 1228 41130 1268 41215
rect 1324 38501 1364 41896
rect 1323 38492 1365 38501
rect 1323 38452 1324 38492
rect 1364 38452 1365 38492
rect 1323 38443 1365 38452
rect 1323 38324 1365 38333
rect 1228 38284 1324 38324
rect 1364 38284 1460 38324
rect 1228 38240 1268 38284
rect 1323 38275 1365 38284
rect 1228 38191 1268 38200
rect 1227 37400 1269 37409
rect 1227 37360 1228 37400
rect 1268 37360 1364 37400
rect 1227 37351 1269 37360
rect 1228 37266 1268 37351
rect 1324 37157 1364 37360
rect 1323 37148 1365 37157
rect 1323 37108 1324 37148
rect 1364 37108 1365 37148
rect 1323 37099 1365 37108
rect 1420 36905 1460 38284
rect 1419 36896 1461 36905
rect 1419 36856 1420 36896
rect 1460 36856 1461 36896
rect 1419 36847 1461 36856
rect 1228 36728 1268 36737
rect 1419 36728 1461 36737
rect 1268 36688 1364 36728
rect 1228 36679 1268 36688
rect 1324 36401 1364 36688
rect 1419 36688 1420 36728
rect 1460 36688 1461 36728
rect 1419 36679 1461 36688
rect 1323 36392 1365 36401
rect 1323 36352 1324 36392
rect 1364 36352 1365 36392
rect 1323 36343 1365 36352
rect 1228 35888 1268 35897
rect 1420 35888 1460 36679
rect 1268 35848 1460 35888
rect 1228 35839 1268 35848
rect 1324 34637 1364 35848
rect 1323 34628 1365 34637
rect 1323 34588 1324 34628
rect 1364 34588 1365 34628
rect 1323 34579 1365 34588
rect 1419 33956 1461 33965
rect 1419 33916 1420 33956
rect 1460 33916 1461 33956
rect 1419 33907 1461 33916
rect 1131 33620 1173 33629
rect 1131 33580 1132 33620
rect 1172 33580 1173 33620
rect 1131 33571 1173 33580
rect 1035 33536 1077 33545
rect 1035 33496 1036 33536
rect 1076 33496 1077 33536
rect 1035 33487 1077 33496
rect 1131 33200 1173 33209
rect 1131 33160 1132 33200
rect 1172 33160 1173 33200
rect 1131 33151 1173 33160
rect 939 30932 981 30941
rect 939 30892 940 30932
rect 980 30892 981 30932
rect 939 30883 981 30892
rect 843 27068 885 27077
rect 843 27028 844 27068
rect 884 27028 885 27068
rect 843 27019 885 27028
rect 939 25724 981 25733
rect 939 25684 940 25724
rect 980 25684 981 25724
rect 939 25675 981 25684
rect 555 25304 597 25313
rect 555 25264 556 25304
rect 596 25264 597 25304
rect 555 25255 597 25264
rect 363 23708 405 23717
rect 363 23668 364 23708
rect 404 23668 405 23708
rect 363 23659 405 23668
rect 171 23204 213 23213
rect 171 23164 172 23204
rect 212 23164 213 23204
rect 171 23155 213 23164
rect 75 19256 117 19265
rect 75 19216 76 19256
rect 116 19216 117 19256
rect 75 19207 117 19216
rect 940 18929 980 25675
rect 1132 23960 1172 33151
rect 1323 32948 1365 32957
rect 1228 32908 1324 32948
rect 1364 32908 1365 32948
rect 1228 32864 1268 32908
rect 1323 32899 1365 32908
rect 1228 32815 1268 32824
rect 1228 30680 1268 30689
rect 1268 30640 1364 30680
rect 1228 30631 1268 30640
rect 1324 29765 1364 30640
rect 1420 30017 1460 33907
rect 1419 30008 1461 30017
rect 1419 29968 1420 30008
rect 1460 29968 1461 30008
rect 1419 29959 1461 29968
rect 1323 29756 1365 29765
rect 1323 29716 1324 29756
rect 1364 29716 1365 29756
rect 1323 29707 1365 29716
rect 1227 29672 1269 29681
rect 1227 29632 1228 29672
rect 1268 29632 1269 29672
rect 1227 29623 1269 29632
rect 1228 27749 1268 29623
rect 1227 27740 1269 27749
rect 1227 27700 1228 27740
rect 1268 27700 1269 27740
rect 1227 27691 1269 27700
rect 1323 26564 1365 26573
rect 1323 26524 1324 26564
rect 1364 26524 1365 26564
rect 1323 26515 1365 26524
rect 1227 26144 1269 26153
rect 1227 26104 1228 26144
rect 1268 26104 1269 26144
rect 1227 26095 1269 26104
rect 1228 26010 1268 26095
rect 1227 25304 1269 25313
rect 1227 25264 1228 25304
rect 1268 25264 1269 25304
rect 1227 25255 1269 25264
rect 1228 25170 1268 25255
rect 1036 23920 1172 23960
rect 939 18920 981 18929
rect 939 18880 940 18920
rect 980 18880 981 18920
rect 939 18871 981 18880
rect 75 16064 117 16073
rect 75 16024 76 16064
rect 116 16024 117 16064
rect 75 16015 117 16024
rect 76 4481 116 16015
rect 1036 13721 1076 23920
rect 1228 23120 1268 23129
rect 1228 22877 1268 23080
rect 1227 22868 1269 22877
rect 1227 22828 1228 22868
rect 1268 22828 1269 22868
rect 1227 22819 1269 22828
rect 1228 22280 1268 22289
rect 1324 22280 1364 26515
rect 1419 25052 1461 25061
rect 1419 25012 1420 25052
rect 1460 25012 1461 25052
rect 1419 25003 1461 25012
rect 1268 22240 1364 22280
rect 1228 22231 1268 22240
rect 1131 22028 1173 22037
rect 1131 21988 1132 22028
rect 1172 21988 1173 22028
rect 1131 21979 1173 21988
rect 1035 13712 1077 13721
rect 1035 13672 1036 13712
rect 1076 13672 1077 13712
rect 1035 13663 1077 13672
rect 843 13208 885 13217
rect 843 13168 844 13208
rect 884 13168 885 13208
rect 843 13159 885 13168
rect 171 10688 213 10697
rect 171 10648 172 10688
rect 212 10648 213 10688
rect 171 10639 213 10648
rect 75 4472 117 4481
rect 75 4432 76 4472
rect 116 4432 117 4472
rect 75 4423 117 4432
rect 172 1793 212 10639
rect 844 6833 884 13159
rect 1132 8765 1172 21979
rect 1420 21617 1460 25003
rect 1419 21608 1461 21617
rect 1419 21568 1420 21608
rect 1460 21568 1461 21608
rect 1419 21559 1461 21568
rect 1323 21440 1365 21449
rect 1323 21400 1324 21440
rect 1364 21400 1365 21440
rect 1323 21391 1365 21400
rect 1228 20768 1268 20777
rect 1324 20768 1364 21391
rect 1268 20728 1364 20768
rect 1228 20719 1268 20728
rect 1228 20096 1268 20105
rect 1268 20056 1364 20096
rect 1228 20047 1268 20056
rect 1324 19433 1364 20056
rect 1323 19424 1365 19433
rect 1323 19384 1324 19424
rect 1364 19384 1365 19424
rect 1323 19375 1365 19384
rect 1228 19256 1268 19265
rect 1228 19172 1268 19216
rect 1323 19172 1365 19181
rect 1228 19132 1324 19172
rect 1364 19132 1365 19172
rect 1323 19123 1365 19132
rect 1227 19004 1269 19013
rect 1227 18964 1228 19004
rect 1268 18964 1269 19004
rect 1227 18955 1269 18964
rect 1228 17744 1268 18955
rect 1419 18668 1461 18677
rect 1419 18628 1420 18668
rect 1460 18628 1461 18668
rect 1419 18619 1461 18628
rect 1228 17660 1268 17704
rect 1228 17620 1364 17660
rect 1227 16064 1269 16073
rect 1227 16024 1228 16064
rect 1268 16024 1269 16064
rect 1227 16015 1269 16024
rect 1228 15930 1268 16015
rect 1227 15728 1269 15737
rect 1227 15688 1228 15728
rect 1268 15688 1269 15728
rect 1227 15679 1269 15688
rect 1228 15560 1268 15679
rect 1228 15511 1268 15520
rect 1228 14048 1268 14057
rect 1324 14048 1364 17620
rect 1420 16316 1460 18619
rect 1420 16267 1460 16276
rect 1516 15401 1556 44920
rect 1804 44910 1844 44995
rect 1996 44960 2036 45583
rect 1611 44792 1653 44801
rect 1611 44752 1612 44792
rect 1652 44752 1653 44792
rect 1611 44743 1653 44752
rect 1612 44658 1652 44743
rect 1996 44288 2036 44920
rect 2092 44885 2132 45676
rect 2380 45389 2420 46432
rect 2476 46423 2516 46432
rect 2764 46432 2900 46472
rect 2476 45716 2516 45725
rect 2379 45380 2421 45389
rect 2379 45340 2380 45380
rect 2420 45340 2421 45380
rect 2379 45331 2421 45340
rect 2091 44876 2133 44885
rect 2091 44836 2092 44876
rect 2132 44836 2133 44876
rect 2091 44827 2133 44836
rect 2476 44381 2516 45676
rect 2667 45548 2709 45557
rect 2667 45508 2668 45548
rect 2708 45508 2709 45548
rect 2667 45499 2709 45508
rect 2668 45414 2708 45499
rect 2764 45221 2804 46432
rect 2860 46304 2900 46313
rect 2860 45893 2900 46264
rect 2859 45884 2901 45893
rect 2859 45844 2860 45884
rect 2900 45844 2901 45884
rect 2859 45835 2901 45844
rect 2860 45716 2900 45725
rect 2956 45716 2996 51052
rect 3051 51052 3052 51092
rect 3092 51052 3093 51092
rect 3051 51043 3093 51052
rect 3052 50958 3092 51043
rect 3148 50345 3188 51808
rect 3532 51773 3572 53068
rect 3688 52940 4056 52949
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 4108 52940 4148 53320
rect 4108 52900 4244 52940
rect 3688 52891 4056 52900
rect 3819 52772 3861 52781
rect 3819 52732 3820 52772
rect 3860 52732 3861 52772
rect 3819 52723 3861 52732
rect 3724 52520 3764 52529
rect 3531 51764 3573 51773
rect 3531 51724 3532 51764
rect 3572 51724 3573 51764
rect 3531 51715 3573 51724
rect 3724 51596 3764 52480
rect 3820 52520 3860 52723
rect 4204 52529 4244 52900
rect 3820 51857 3860 52480
rect 4203 52520 4245 52529
rect 4203 52480 4204 52520
rect 4244 52480 4245 52520
rect 4203 52471 4245 52480
rect 4300 52520 4340 52531
rect 3819 51848 3861 51857
rect 3819 51808 3820 51848
rect 3860 51808 3861 51848
rect 3819 51799 3861 51808
rect 4107 51680 4149 51689
rect 4107 51640 4108 51680
rect 4148 51640 4149 51680
rect 4107 51631 4149 51640
rect 3532 51556 3764 51596
rect 3532 51017 3572 51556
rect 3688 51428 4056 51437
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 3688 51379 4056 51388
rect 4108 51260 4148 51631
rect 4012 51220 4148 51260
rect 3243 51008 3285 51017
rect 3243 50968 3244 51008
rect 3284 50968 3285 51008
rect 3243 50959 3285 50968
rect 3531 51008 3573 51017
rect 3531 50968 3532 51008
rect 3572 50968 3573 51008
rect 3531 50959 3573 50968
rect 4012 51008 4052 51220
rect 4204 51050 4244 52471
rect 4300 52445 4340 52480
rect 4299 52436 4341 52445
rect 4299 52396 4300 52436
rect 4340 52396 4341 52436
rect 4299 52387 4341 52396
rect 4396 52016 4436 53992
rect 4492 53276 4532 56083
rect 4588 53444 4628 57016
rect 5260 56981 5300 57940
rect 5355 57812 5397 57821
rect 5355 57772 5356 57812
rect 5396 57772 5397 57812
rect 5355 57763 5397 57772
rect 5259 56972 5301 56981
rect 5259 56932 5260 56972
rect 5300 56932 5301 56972
rect 5259 56923 5301 56932
rect 4928 56720 5296 56729
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 4928 56671 5296 56680
rect 5356 56552 5396 57763
rect 5356 56503 5396 56512
rect 5163 56468 5205 56477
rect 5163 56428 5164 56468
rect 5204 56428 5205 56468
rect 5163 56419 5205 56428
rect 4683 56384 4725 56393
rect 4683 56344 4684 56384
rect 4724 56344 4725 56384
rect 4683 56335 4725 56344
rect 5164 56379 5204 56419
rect 4684 56250 4724 56335
rect 5164 56330 5204 56339
rect 4684 55544 4724 55553
rect 4684 54881 4724 55504
rect 5451 55460 5493 55469
rect 5451 55420 5452 55460
rect 5492 55420 5493 55460
rect 5451 55411 5493 55420
rect 5452 55301 5492 55411
rect 5451 55292 5493 55301
rect 5451 55252 5452 55292
rect 5492 55252 5493 55292
rect 5451 55243 5493 55252
rect 4928 55208 5296 55217
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 4928 55159 5296 55168
rect 4683 54872 4725 54881
rect 4683 54832 4684 54872
rect 4724 54832 4725 54872
rect 4683 54823 4725 54832
rect 4928 53696 5296 53705
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 4928 53647 5296 53656
rect 5548 53444 5588 59788
rect 5644 57653 5684 63064
rect 5740 63020 5780 63029
rect 6028 63020 6068 63064
rect 5780 62980 6068 63020
rect 6124 63104 6164 63113
rect 5740 62971 5780 62980
rect 5739 62768 5781 62777
rect 5739 62728 5740 62768
rect 5780 62728 5781 62768
rect 5739 62719 5781 62728
rect 5643 57644 5685 57653
rect 5643 57604 5644 57644
rect 5684 57604 5685 57644
rect 5643 57595 5685 57604
rect 5644 57056 5684 57065
rect 5644 54041 5684 57016
rect 5740 55469 5780 62719
rect 5835 62684 5877 62693
rect 5835 62644 5836 62684
rect 5876 62644 5877 62684
rect 5835 62635 5877 62644
rect 5836 59753 5876 62635
rect 6124 61433 6164 63064
rect 6123 61424 6165 61433
rect 6123 61384 6124 61424
rect 6164 61384 6165 61424
rect 6123 61375 6165 61384
rect 6027 61256 6069 61265
rect 6027 61216 6028 61256
rect 6068 61216 6069 61256
rect 6027 61207 6069 61216
rect 5835 59744 5877 59753
rect 5835 59704 5836 59744
rect 5876 59704 5877 59744
rect 5835 59695 5877 59704
rect 5932 58568 5972 58577
rect 5932 58493 5972 58528
rect 5931 58484 5973 58493
rect 5931 58444 5932 58484
rect 5972 58444 5973 58484
rect 5931 58435 5973 58444
rect 5932 58241 5972 58435
rect 5931 58232 5973 58241
rect 5931 58192 5932 58232
rect 5972 58192 5973 58232
rect 5931 58183 5973 58192
rect 5836 56888 5876 56897
rect 5836 56477 5876 56848
rect 5835 56468 5877 56477
rect 5835 56428 5836 56468
rect 5876 56428 5877 56468
rect 5835 56419 5877 56428
rect 5835 56300 5877 56309
rect 5835 56260 5836 56300
rect 5876 56260 5877 56300
rect 5835 56251 5877 56260
rect 5739 55460 5781 55469
rect 5739 55420 5740 55460
rect 5780 55420 5781 55460
rect 5739 55411 5781 55420
rect 5643 54032 5685 54041
rect 5643 53992 5644 54032
rect 5684 53992 5685 54032
rect 5836 54032 5876 56251
rect 5932 55544 5972 58183
rect 6028 56384 6068 61207
rect 6220 60248 6260 63232
rect 6316 62777 6356 63316
rect 6412 63281 6452 64315
rect 6508 63692 6548 65323
rect 6604 64280 6644 65500
rect 6796 64616 6836 65827
rect 7084 65624 7124 65920
rect 6604 64240 6740 64280
rect 6508 63652 6644 63692
rect 6411 63272 6453 63281
rect 6411 63232 6412 63272
rect 6452 63232 6453 63272
rect 6411 63223 6453 63232
rect 6507 63188 6549 63197
rect 6507 63148 6508 63188
rect 6548 63148 6549 63188
rect 6507 63139 6549 63148
rect 6604 63188 6644 63652
rect 6604 63139 6644 63148
rect 6508 63054 6548 63139
rect 6603 63020 6645 63029
rect 6603 62980 6604 63020
rect 6644 62980 6645 63020
rect 6603 62971 6645 62980
rect 6315 62768 6357 62777
rect 6315 62728 6316 62768
rect 6356 62728 6357 62768
rect 6315 62719 6357 62728
rect 6508 62432 6548 62441
rect 6604 62432 6644 62971
rect 6548 62392 6644 62432
rect 6508 62189 6548 62392
rect 6507 62180 6549 62189
rect 6507 62140 6508 62180
rect 6548 62140 6549 62180
rect 6507 62131 6549 62140
rect 6507 61592 6549 61601
rect 6507 61552 6508 61592
rect 6548 61552 6549 61592
rect 6507 61543 6549 61552
rect 6508 61458 6548 61543
rect 6411 61088 6453 61097
rect 6411 61048 6412 61088
rect 6452 61048 6453 61088
rect 6411 61039 6453 61048
rect 6412 60920 6452 61039
rect 6412 60871 6452 60880
rect 6315 60668 6357 60677
rect 6315 60628 6316 60668
rect 6356 60628 6357 60668
rect 6315 60619 6357 60628
rect 6604 60668 6644 60677
rect 6124 60208 6260 60248
rect 6124 58997 6164 60208
rect 6219 60080 6261 60089
rect 6219 60040 6220 60080
rect 6260 60040 6261 60080
rect 6219 60031 6261 60040
rect 6220 59417 6260 60031
rect 6219 59408 6261 59417
rect 6219 59368 6220 59408
rect 6260 59368 6261 59408
rect 6219 59359 6261 59368
rect 6316 59408 6356 60619
rect 6604 60080 6644 60628
rect 6700 60257 6740 64240
rect 6699 60248 6741 60257
rect 6699 60208 6700 60248
rect 6740 60208 6741 60248
rect 6699 60199 6741 60208
rect 6604 60031 6644 60040
rect 6699 60080 6741 60089
rect 6699 60040 6700 60080
rect 6740 60040 6741 60080
rect 6699 60031 6741 60040
rect 6700 59946 6740 60031
rect 6412 59417 6452 59502
rect 6796 59492 6836 64576
rect 6988 65584 7124 65624
rect 7180 65920 7316 65960
rect 6988 63449 7028 65584
rect 7083 65456 7125 65465
rect 7083 65416 7084 65456
rect 7124 65416 7125 65456
rect 7083 65407 7125 65416
rect 7084 64625 7124 65407
rect 7083 64616 7125 64625
rect 7083 64576 7084 64616
rect 7124 64576 7125 64616
rect 7083 64567 7125 64576
rect 6987 63440 7029 63449
rect 6987 63400 6988 63440
rect 7028 63400 7029 63440
rect 6987 63391 7029 63400
rect 6891 63272 6933 63281
rect 6891 63232 6892 63272
rect 6932 63232 6933 63272
rect 6891 63223 6933 63232
rect 6892 61601 6932 63223
rect 7084 63104 7124 63113
rect 6988 63064 7084 63104
rect 6891 61592 6933 61601
rect 6891 61552 6892 61592
rect 6932 61552 6933 61592
rect 6891 61543 6933 61552
rect 6892 60920 6932 61543
rect 6892 60845 6932 60880
rect 6891 60836 6933 60845
rect 6891 60796 6892 60836
rect 6932 60796 6933 60836
rect 6891 60787 6933 60796
rect 6988 60005 7028 63064
rect 7084 63055 7124 63064
rect 7083 62348 7125 62357
rect 7083 62308 7084 62348
rect 7124 62308 7125 62348
rect 7083 62299 7125 62308
rect 7180 62348 7220 65920
rect 7275 65792 7317 65801
rect 7275 65752 7276 65792
rect 7316 65752 7317 65792
rect 7275 65743 7317 65752
rect 7276 65456 7316 65743
rect 7372 65624 7412 67171
rect 7564 66893 7604 69532
rect 7660 69404 7700 69413
rect 7756 69404 7796 69938
rect 7700 69364 7796 69404
rect 7660 69355 7700 69364
rect 7852 69245 7892 70624
rect 7948 70421 7988 70960
rect 8044 70589 8084 70674
rect 8043 70580 8085 70589
rect 8043 70540 8044 70580
rect 8084 70540 8085 70580
rect 8140 70580 8180 73387
rect 8235 73352 8277 73361
rect 8235 73312 8236 73352
rect 8276 73312 8277 73352
rect 8235 73303 8277 73312
rect 8236 71093 8276 73303
rect 8332 73016 8372 75160
rect 8427 73688 8469 73697
rect 8427 73648 8428 73688
rect 8468 73648 8469 73688
rect 8427 73639 8469 73648
rect 8428 73554 8468 73639
rect 8620 73445 8660 76840
rect 8619 73436 8661 73445
rect 8619 73396 8620 73436
rect 8660 73396 8661 73436
rect 8619 73387 8661 73396
rect 8235 71084 8277 71093
rect 8235 71044 8236 71084
rect 8276 71044 8277 71084
rect 8235 71035 8277 71044
rect 8332 70916 8372 72976
rect 8812 71840 8852 77428
rect 9100 77384 9140 78259
rect 8908 77344 9140 77384
rect 8908 76796 8948 77344
rect 8908 76553 8948 76756
rect 9196 76721 9236 79696
rect 9292 79568 9332 79577
rect 9292 78233 9332 79528
rect 9291 78224 9333 78233
rect 9291 78184 9292 78224
rect 9332 78184 9333 78224
rect 9291 78175 9333 78184
rect 9388 77552 9428 84400
rect 9483 83432 9525 83441
rect 9483 83392 9484 83432
rect 9524 83392 9525 83432
rect 9483 83383 9525 83392
rect 9484 83298 9524 83383
rect 9483 82592 9525 82601
rect 9483 82552 9484 82592
rect 9524 82552 9525 82592
rect 9483 82543 9525 82552
rect 9484 81593 9524 82543
rect 9483 81584 9525 81593
rect 9483 81544 9484 81584
rect 9524 81544 9525 81584
rect 9483 81535 9525 81544
rect 9484 81248 9524 81535
rect 9484 80576 9524 81208
rect 9580 80753 9620 85828
rect 9676 84449 9716 85936
rect 9868 84449 9908 85936
rect 9675 84440 9717 84449
rect 9675 84400 9676 84440
rect 9716 84400 9717 84440
rect 9675 84391 9717 84400
rect 9867 84440 9909 84449
rect 9867 84400 9868 84440
rect 9908 84400 9909 84440
rect 9867 84391 9909 84400
rect 10060 84281 10100 85936
rect 10252 85280 10292 85936
rect 10444 85364 10484 85936
rect 10444 85324 10580 85364
rect 10252 85240 10484 85280
rect 9676 84272 9716 84281
rect 9676 83693 9716 84232
rect 10059 84272 10101 84281
rect 10059 84232 10060 84272
rect 10100 84232 10101 84272
rect 10059 84223 10101 84232
rect 10252 84272 10292 84281
rect 10292 84232 10388 84272
rect 10252 84223 10292 84232
rect 9771 84188 9813 84197
rect 9771 84148 9772 84188
rect 9812 84148 9813 84188
rect 9771 84139 9813 84148
rect 9675 83684 9717 83693
rect 9675 83644 9676 83684
rect 9716 83644 9717 83684
rect 9675 83635 9717 83644
rect 9675 83432 9717 83441
rect 9675 83392 9676 83432
rect 9716 83392 9717 83432
rect 9675 83383 9717 83392
rect 9676 83298 9716 83383
rect 9772 83096 9812 84139
rect 9868 84104 9908 84113
rect 10060 84104 10100 84113
rect 9908 84064 10004 84104
rect 9868 84055 9908 84064
rect 9867 83684 9909 83693
rect 9867 83644 9868 83684
rect 9908 83644 9909 83684
rect 9867 83635 9909 83644
rect 9676 83056 9812 83096
rect 9579 80744 9621 80753
rect 9579 80704 9580 80744
rect 9620 80704 9621 80744
rect 9579 80695 9621 80704
rect 9484 80536 9620 80576
rect 9483 80072 9525 80081
rect 9483 80032 9484 80072
rect 9524 80032 9525 80072
rect 9483 80023 9525 80032
rect 9484 79736 9524 80023
rect 9484 79687 9524 79696
rect 9580 79568 9620 80536
rect 9292 77512 9428 77552
rect 9484 79528 9620 79568
rect 9004 76712 9044 76721
rect 9195 76712 9237 76721
rect 9044 76672 9140 76712
rect 9004 76663 9044 76672
rect 8907 76544 8949 76553
rect 8907 76504 8908 76544
rect 8948 76504 8949 76544
rect 8907 76495 8949 76504
rect 9003 76124 9045 76133
rect 9003 76084 9004 76124
rect 9044 76084 9045 76124
rect 9003 76075 9045 76084
rect 9004 72176 9044 76075
rect 9100 72689 9140 76672
rect 9195 76672 9196 76712
rect 9236 76672 9237 76712
rect 9195 76663 9237 76672
rect 9099 72680 9141 72689
rect 9099 72640 9100 72680
rect 9140 72640 9141 72680
rect 9099 72631 9141 72640
rect 9196 72269 9236 76663
rect 9292 74117 9332 77512
rect 9387 77048 9429 77057
rect 9484 77048 9524 79528
rect 9676 79064 9716 83056
rect 9771 82844 9813 82853
rect 9771 82804 9772 82844
rect 9812 82804 9813 82844
rect 9771 82795 9813 82804
rect 9772 82517 9812 82795
rect 9868 82601 9908 83635
rect 9964 83600 10004 84064
rect 10100 84064 10292 84104
rect 10060 84055 10100 84064
rect 10060 83600 10100 83609
rect 9964 83560 10060 83600
rect 10060 83551 10100 83560
rect 10155 83600 10197 83609
rect 10155 83560 10156 83600
rect 10196 83560 10197 83600
rect 10155 83551 10197 83560
rect 10156 83466 10196 83551
rect 10252 83012 10292 84064
rect 10348 83609 10388 84232
rect 10347 83600 10389 83609
rect 10347 83560 10348 83600
rect 10388 83560 10389 83600
rect 10347 83551 10389 83560
rect 10060 82972 10292 83012
rect 9964 82760 10004 82769
rect 9867 82592 9909 82601
rect 9867 82552 9868 82592
rect 9908 82552 9909 82592
rect 9867 82543 9909 82552
rect 9771 82508 9813 82517
rect 9771 82468 9772 82508
rect 9812 82468 9813 82508
rect 9771 82459 9813 82468
rect 9964 82013 10004 82720
rect 9963 82004 10005 82013
rect 9963 81964 9964 82004
rect 10004 81964 10005 82004
rect 9963 81955 10005 81964
rect 9771 81836 9813 81845
rect 9771 81796 9772 81836
rect 9812 81796 9813 81836
rect 9771 81787 9813 81796
rect 9772 81257 9812 81787
rect 9963 81416 10005 81425
rect 9963 81376 9964 81416
rect 10004 81376 10005 81416
rect 9963 81367 10005 81376
rect 9771 81248 9813 81257
rect 9771 81208 9772 81248
rect 9812 81208 9813 81248
rect 9771 81199 9813 81208
rect 9772 80576 9812 81199
rect 9772 80527 9812 80536
rect 9868 80576 9908 80585
rect 9868 80333 9908 80536
rect 9867 80324 9909 80333
rect 9867 80284 9868 80324
rect 9908 80284 9909 80324
rect 9867 80275 9909 80284
rect 9964 79997 10004 81367
rect 10060 80837 10100 82972
rect 10348 82760 10388 82769
rect 10252 82720 10348 82760
rect 10155 82676 10197 82685
rect 10155 82636 10156 82676
rect 10196 82636 10197 82676
rect 10155 82627 10197 82636
rect 10156 82542 10196 82627
rect 10155 82424 10197 82433
rect 10155 82384 10156 82424
rect 10196 82384 10197 82424
rect 10155 82375 10197 82384
rect 10059 80828 10101 80837
rect 10059 80788 10060 80828
rect 10100 80788 10101 80828
rect 10059 80779 10101 80788
rect 9771 79988 9813 79997
rect 9771 79948 9772 79988
rect 9812 79948 9813 79988
rect 9771 79939 9813 79948
rect 9963 79988 10005 79997
rect 9963 79948 9964 79988
rect 10004 79948 10005 79988
rect 9963 79939 10005 79948
rect 9580 79024 9716 79064
rect 9580 77813 9620 79024
rect 9676 78224 9716 78233
rect 9772 78224 9812 79939
rect 10059 79652 10101 79661
rect 10059 79612 10060 79652
rect 10100 79612 10101 79652
rect 10059 79603 10101 79612
rect 10060 79064 10100 79603
rect 9964 79024 10060 79064
rect 9964 78737 10004 79024
rect 10060 79015 10100 79024
rect 9963 78728 10005 78737
rect 9963 78688 9964 78728
rect 10004 78688 10005 78728
rect 9963 78679 10005 78688
rect 9716 78184 9812 78224
rect 9579 77804 9621 77813
rect 9579 77764 9580 77804
rect 9620 77764 9621 77804
rect 9579 77755 9621 77764
rect 9387 77008 9388 77048
rect 9428 77008 9524 77048
rect 9387 76999 9429 77008
rect 9388 75209 9428 76999
rect 9484 76712 9524 76721
rect 9387 75200 9429 75209
rect 9387 75160 9388 75200
rect 9428 75160 9429 75200
rect 9387 75151 9429 75160
rect 9291 74108 9333 74117
rect 9291 74068 9292 74108
rect 9332 74068 9333 74108
rect 9291 74059 9333 74068
rect 9388 73277 9428 75151
rect 9484 74621 9524 76672
rect 9676 76133 9716 78184
rect 9868 78056 9908 78065
rect 9908 78016 10004 78056
rect 9868 78007 9908 78016
rect 9964 76726 10004 78016
rect 10156 76721 10196 82375
rect 10252 82097 10292 82720
rect 10348 82711 10388 82720
rect 10444 82592 10484 85240
rect 10540 83693 10580 85324
rect 10636 83945 10676 85936
rect 10731 84272 10773 84281
rect 10731 84232 10732 84272
rect 10772 84232 10773 84272
rect 10731 84223 10773 84232
rect 10635 83936 10677 83945
rect 10635 83896 10636 83936
rect 10676 83896 10677 83936
rect 10635 83887 10677 83896
rect 10539 83684 10581 83693
rect 10539 83644 10540 83684
rect 10580 83644 10581 83684
rect 10539 83635 10581 83644
rect 10539 83516 10581 83525
rect 10539 83476 10540 83516
rect 10580 83476 10581 83516
rect 10539 83467 10581 83476
rect 10636 83516 10676 83527
rect 10540 83382 10580 83467
rect 10636 83441 10676 83476
rect 10635 83432 10677 83441
rect 10635 83392 10636 83432
rect 10676 83392 10677 83432
rect 10635 83383 10677 83392
rect 10539 83180 10581 83189
rect 10539 83140 10540 83180
rect 10580 83140 10581 83180
rect 10539 83131 10581 83140
rect 10348 82552 10484 82592
rect 10251 82088 10293 82097
rect 10251 82048 10252 82088
rect 10292 82048 10293 82088
rect 10251 82039 10293 82048
rect 10348 81341 10388 82552
rect 10444 82088 10484 82099
rect 10444 82013 10484 82048
rect 10443 82004 10485 82013
rect 10443 81964 10444 82004
rect 10484 81964 10485 82004
rect 10443 81955 10485 81964
rect 10347 81332 10389 81341
rect 10347 81292 10348 81332
rect 10388 81292 10389 81332
rect 10347 81283 10389 81292
rect 10252 80492 10292 80501
rect 10252 79400 10292 80452
rect 10348 80492 10388 80501
rect 10388 80452 10484 80492
rect 10348 80443 10388 80452
rect 10444 79409 10484 80452
rect 10540 80417 10580 83131
rect 10635 82256 10677 82265
rect 10635 82216 10636 82256
rect 10676 82216 10677 82256
rect 10635 82207 10677 82216
rect 10636 82122 10676 82207
rect 10732 81677 10772 84223
rect 10828 83525 10868 85936
rect 10923 83936 10965 83945
rect 10923 83896 10924 83936
rect 10964 83896 10965 83936
rect 10923 83887 10965 83896
rect 10827 83516 10869 83525
rect 10827 83476 10828 83516
rect 10868 83476 10869 83516
rect 10827 83467 10869 83476
rect 10924 83273 10964 83887
rect 10923 83264 10965 83273
rect 10923 83224 10924 83264
rect 10964 83224 10965 83264
rect 10923 83215 10965 83224
rect 11020 83189 11060 85936
rect 11212 84449 11252 85936
rect 11404 84524 11444 85936
rect 11499 85532 11541 85541
rect 11499 85492 11500 85532
rect 11540 85492 11541 85532
rect 11499 85483 11541 85492
rect 11308 84484 11444 84524
rect 11211 84440 11253 84449
rect 11211 84400 11212 84440
rect 11252 84400 11253 84440
rect 11211 84391 11253 84400
rect 11115 83600 11157 83609
rect 11115 83560 11116 83600
rect 11156 83560 11157 83600
rect 11115 83551 11157 83560
rect 11116 83466 11156 83551
rect 11019 83180 11061 83189
rect 11019 83140 11020 83180
rect 11060 83140 11061 83180
rect 11019 83131 11061 83140
rect 10923 83096 10965 83105
rect 10923 83056 10924 83096
rect 10964 83056 10965 83096
rect 10923 83047 10965 83056
rect 10827 82256 10869 82265
rect 10827 82216 10828 82256
rect 10868 82216 10869 82256
rect 10827 82207 10869 82216
rect 10828 82088 10868 82207
rect 10828 82013 10868 82048
rect 10827 82004 10869 82013
rect 10827 81964 10828 82004
rect 10868 81964 10869 82004
rect 10827 81955 10869 81964
rect 10924 81920 10964 83047
rect 11308 82433 11348 84484
rect 11500 84440 11540 85483
rect 11404 84400 11540 84440
rect 11404 82769 11444 84400
rect 11499 84272 11541 84281
rect 11499 84232 11500 84272
rect 11540 84232 11541 84272
rect 11499 84223 11541 84232
rect 11500 84138 11540 84223
rect 11596 83936 11636 85936
rect 11788 85028 11828 85936
rect 11788 84988 11924 85028
rect 11884 84449 11924 84988
rect 11980 84533 12020 85936
rect 12172 85541 12212 85936
rect 12171 85532 12213 85541
rect 12171 85492 12172 85532
rect 12212 85492 12213 85532
rect 12171 85483 12213 85492
rect 12364 85364 12404 85936
rect 12172 85324 12404 85364
rect 11979 84524 12021 84533
rect 11979 84484 11980 84524
rect 12020 84484 12021 84524
rect 11979 84475 12021 84484
rect 11883 84440 11925 84449
rect 11883 84400 11884 84440
rect 11924 84400 11925 84440
rect 11883 84391 11925 84400
rect 11787 84356 11829 84365
rect 11787 84316 11788 84356
rect 11828 84316 11829 84356
rect 11787 84307 11829 84316
rect 11500 83896 11636 83936
rect 11692 84272 11732 84281
rect 11403 82760 11445 82769
rect 11403 82720 11404 82760
rect 11444 82720 11445 82760
rect 11403 82711 11445 82720
rect 11500 82433 11540 83896
rect 11596 83586 11636 83595
rect 11596 83021 11636 83546
rect 11595 83012 11637 83021
rect 11595 82972 11596 83012
rect 11636 82972 11637 83012
rect 11595 82963 11637 82972
rect 11596 82760 11636 82769
rect 11596 82601 11636 82720
rect 11595 82592 11637 82601
rect 11595 82552 11596 82592
rect 11636 82552 11637 82592
rect 11595 82543 11637 82552
rect 11307 82424 11349 82433
rect 11307 82384 11308 82424
rect 11348 82384 11349 82424
rect 11307 82375 11349 82384
rect 11499 82424 11541 82433
rect 11692 82424 11732 84232
rect 11788 84222 11828 84307
rect 11884 84272 11924 84281
rect 11924 84232 12116 84272
rect 11884 84223 11924 84232
rect 11788 83684 11828 83693
rect 11788 83600 11828 83644
rect 11788 83560 12020 83600
rect 11787 83012 11829 83021
rect 11787 82972 11788 83012
rect 11828 82972 11829 83012
rect 11787 82963 11829 82972
rect 11788 82878 11828 82963
rect 11883 82508 11925 82517
rect 11883 82468 11884 82508
rect 11924 82468 11925 82508
rect 11883 82459 11925 82468
rect 11499 82384 11500 82424
rect 11540 82384 11541 82424
rect 11499 82375 11541 82384
rect 11596 82384 11732 82424
rect 11019 82256 11061 82265
rect 11596 82256 11636 82384
rect 11884 82340 11924 82459
rect 11884 82300 11931 82340
rect 11891 82256 11931 82300
rect 11019 82216 11020 82256
rect 11060 82216 11061 82256
rect 11019 82207 11061 82216
rect 11500 82216 11636 82256
rect 11692 82216 11931 82256
rect 11020 82122 11060 82207
rect 11116 82088 11156 82097
rect 11404 82088 11444 82097
rect 10924 81880 11060 81920
rect 10731 81668 10773 81677
rect 10731 81628 10732 81668
rect 10772 81628 10773 81668
rect 10731 81619 10773 81628
rect 10732 81248 10772 81257
rect 10635 80912 10677 80921
rect 10635 80872 10636 80912
rect 10676 80872 10677 80912
rect 10635 80863 10677 80872
rect 10539 80408 10581 80417
rect 10539 80368 10540 80408
rect 10580 80368 10581 80408
rect 10539 80359 10581 80368
rect 10636 79409 10676 80863
rect 10732 80249 10772 81208
rect 10828 80576 10868 80585
rect 10828 80417 10868 80536
rect 10827 80408 10869 80417
rect 10827 80368 10828 80408
rect 10868 80368 10869 80408
rect 10827 80359 10869 80368
rect 10731 80240 10773 80249
rect 10731 80200 10732 80240
rect 10772 80200 10773 80240
rect 10731 80191 10773 80200
rect 10732 79904 10772 80191
rect 10732 79864 10868 79904
rect 10732 79736 10772 79747
rect 10732 79661 10772 79696
rect 10731 79652 10773 79661
rect 10731 79612 10732 79652
rect 10772 79612 10773 79652
rect 10731 79603 10773 79612
rect 10443 79400 10485 79409
rect 10252 79360 10388 79400
rect 10251 79148 10293 79157
rect 10251 79108 10252 79148
rect 10292 79108 10293 79148
rect 10251 79099 10293 79108
rect 10252 79014 10292 79099
rect 10348 78905 10388 79360
rect 10443 79360 10444 79400
rect 10484 79360 10485 79400
rect 10443 79351 10485 79360
rect 10635 79400 10677 79409
rect 10635 79360 10636 79400
rect 10676 79360 10677 79400
rect 10635 79351 10677 79360
rect 10635 79232 10677 79241
rect 10635 79192 10636 79232
rect 10676 79192 10677 79232
rect 10635 79183 10677 79192
rect 10636 79064 10676 79183
rect 10636 79015 10676 79024
rect 10732 79064 10772 79073
rect 10347 78896 10389 78905
rect 10347 78856 10348 78896
rect 10388 78856 10389 78896
rect 10347 78847 10389 78856
rect 10251 78728 10293 78737
rect 10251 78688 10252 78728
rect 10292 78688 10293 78728
rect 10251 78679 10293 78688
rect 10252 77552 10292 78679
rect 10348 78485 10388 78847
rect 10347 78476 10389 78485
rect 10347 78436 10348 78476
rect 10388 78436 10389 78476
rect 10347 78427 10389 78436
rect 10539 78224 10581 78233
rect 10539 78184 10540 78224
rect 10580 78184 10581 78224
rect 10539 78175 10581 78184
rect 10636 78224 10676 78233
rect 10732 78224 10772 79024
rect 10828 78401 10868 79864
rect 10924 79568 10964 79577
rect 10827 78392 10869 78401
rect 10827 78352 10828 78392
rect 10868 78352 10869 78392
rect 10827 78343 10869 78352
rect 10924 78233 10964 79528
rect 11020 79148 11060 81880
rect 11116 81509 11156 82048
rect 11308 82048 11404 82088
rect 11211 82004 11253 82013
rect 11308 82004 11348 82048
rect 11404 82039 11444 82048
rect 11211 81964 11212 82004
rect 11252 81964 11348 82004
rect 11211 81955 11253 81964
rect 11115 81500 11157 81509
rect 11115 81460 11116 81500
rect 11156 81460 11157 81500
rect 11115 81451 11157 81460
rect 11212 81248 11252 81955
rect 11500 81509 11540 82216
rect 11692 82088 11732 82216
rect 11980 82097 12020 83560
rect 12076 82769 12116 84232
rect 12172 83693 12212 85324
rect 12267 85196 12309 85205
rect 12267 85156 12268 85196
rect 12308 85156 12309 85196
rect 12267 85147 12309 85156
rect 12268 84356 12308 85147
rect 12363 84776 12405 84785
rect 12363 84736 12364 84776
rect 12404 84736 12405 84776
rect 12363 84727 12405 84736
rect 12268 84307 12308 84316
rect 12364 83936 12404 84727
rect 12459 84104 12501 84113
rect 12459 84064 12460 84104
rect 12500 84064 12501 84104
rect 12459 84055 12501 84064
rect 12460 83970 12500 84055
rect 12268 83896 12404 83936
rect 12268 83768 12308 83896
rect 12268 83728 12404 83768
rect 12171 83684 12213 83693
rect 12171 83644 12172 83684
rect 12212 83644 12213 83684
rect 12171 83635 12213 83644
rect 12267 83600 12309 83609
rect 12267 83560 12268 83600
rect 12308 83560 12309 83600
rect 12267 83551 12309 83560
rect 12172 83516 12212 83525
rect 12075 82760 12117 82769
rect 12075 82720 12076 82760
rect 12116 82720 12117 82760
rect 12075 82711 12117 82720
rect 12172 82601 12212 83476
rect 12171 82592 12213 82601
rect 12171 82552 12172 82592
rect 12212 82552 12213 82592
rect 12171 82543 12213 82552
rect 12172 82458 12212 82543
rect 12268 82340 12308 83551
rect 12364 83516 12404 83728
rect 12556 83693 12596 85936
rect 12651 84692 12693 84701
rect 12651 84652 12652 84692
rect 12692 84652 12693 84692
rect 12651 84643 12693 84652
rect 12555 83684 12597 83693
rect 12555 83644 12556 83684
rect 12596 83644 12597 83684
rect 12555 83635 12597 83644
rect 12364 83476 12596 83516
rect 12556 83432 12596 83476
rect 12556 83383 12596 83392
rect 12363 83348 12405 83357
rect 12363 83308 12364 83348
rect 12404 83308 12405 83348
rect 12363 83299 12405 83308
rect 12364 83214 12404 83299
rect 12652 82937 12692 84643
rect 12748 84449 12788 85936
rect 12940 84524 12980 85936
rect 13132 85457 13172 85936
rect 13131 85448 13173 85457
rect 13131 85408 13132 85448
rect 13172 85408 13173 85448
rect 13131 85399 13173 85408
rect 13131 85112 13173 85121
rect 13131 85072 13132 85112
rect 13172 85072 13173 85112
rect 13131 85063 13173 85072
rect 13035 85028 13077 85037
rect 13035 84988 13036 85028
rect 13076 84988 13077 85028
rect 13035 84979 13077 84988
rect 12844 84484 12980 84524
rect 12747 84440 12789 84449
rect 12747 84400 12748 84440
rect 12788 84400 12789 84440
rect 12747 84391 12789 84400
rect 12747 84104 12789 84113
rect 12747 84064 12748 84104
rect 12788 84064 12789 84104
rect 12747 84055 12789 84064
rect 12748 83970 12788 84055
rect 12748 83516 12788 83525
rect 12748 83189 12788 83476
rect 12747 83180 12789 83189
rect 12747 83140 12748 83180
rect 12788 83140 12789 83180
rect 12747 83131 12789 83140
rect 12651 82928 12693 82937
rect 12651 82888 12652 82928
rect 12692 82888 12693 82928
rect 12651 82879 12693 82888
rect 12363 82760 12405 82769
rect 12363 82720 12364 82760
rect 12404 82720 12405 82760
rect 12363 82711 12405 82720
rect 12460 82760 12500 82769
rect 12172 82300 12308 82340
rect 11692 82039 11732 82048
rect 11788 82088 11828 82097
rect 11788 81845 11828 82048
rect 11979 82088 12021 82097
rect 11979 82048 11980 82088
rect 12020 82048 12021 82088
rect 11979 82039 12021 82048
rect 11787 81836 11829 81845
rect 11787 81796 11788 81836
rect 11828 81796 11829 81836
rect 11787 81787 11829 81796
rect 12076 81836 12116 81845
rect 11499 81500 11541 81509
rect 11499 81460 11500 81500
rect 11540 81460 11541 81500
rect 11499 81451 11541 81460
rect 11691 81500 11733 81509
rect 11691 81460 11692 81500
rect 11732 81460 11733 81500
rect 11691 81451 11733 81460
rect 11692 81366 11732 81451
rect 11499 81332 11541 81341
rect 11499 81292 11500 81332
rect 11540 81292 11541 81332
rect 11499 81283 11541 81292
rect 11212 80660 11252 81208
rect 11308 81248 11348 81257
rect 11308 80837 11348 81208
rect 11403 81248 11445 81257
rect 11403 81208 11404 81248
rect 11444 81208 11445 81248
rect 11403 81199 11445 81208
rect 11500 81248 11540 81283
rect 11404 81114 11444 81199
rect 11500 81197 11540 81208
rect 11692 81248 11732 81257
rect 11692 81089 11732 81208
rect 11787 81248 11829 81257
rect 11787 81208 11788 81248
rect 11828 81208 11829 81248
rect 11787 81199 11829 81208
rect 11884 81248 11924 81257
rect 11499 81080 11541 81089
rect 11691 81080 11733 81089
rect 11499 81040 11500 81080
rect 11540 81040 11636 81080
rect 11499 81031 11541 81040
rect 11307 80828 11349 80837
rect 11307 80788 11308 80828
rect 11348 80788 11349 80828
rect 11307 80779 11349 80788
rect 11499 80660 11541 80669
rect 11212 80620 11348 80660
rect 11308 80576 11348 80620
rect 11499 80620 11500 80660
rect 11540 80620 11541 80660
rect 11499 80611 11541 80620
rect 11308 80566 11396 80576
rect 11308 80536 11356 80566
rect 11500 80526 11540 80611
rect 11211 80492 11253 80501
rect 11211 80452 11212 80492
rect 11252 80452 11253 80492
rect 11356 80460 11396 80526
rect 11211 80443 11253 80452
rect 11212 80249 11252 80443
rect 11307 80408 11349 80417
rect 11307 80368 11308 80408
rect 11348 80368 11349 80408
rect 11307 80359 11349 80368
rect 11499 80408 11541 80417
rect 11499 80368 11500 80408
rect 11540 80368 11541 80408
rect 11596 80408 11636 81040
rect 11691 81040 11692 81080
rect 11732 81040 11733 81080
rect 11691 81031 11733 81040
rect 11788 80576 11828 81199
rect 11884 80744 11924 81208
rect 11980 81248 12020 81257
rect 12076 81248 12116 81796
rect 12172 81425 12212 82300
rect 12364 82256 12404 82711
rect 12460 82265 12500 82720
rect 12556 82760 12596 82769
rect 12364 82207 12404 82216
rect 12459 82256 12501 82265
rect 12459 82216 12460 82256
rect 12500 82216 12501 82256
rect 12459 82207 12501 82216
rect 12268 82088 12308 82097
rect 12171 81416 12213 81425
rect 12171 81376 12172 81416
rect 12212 81376 12213 81416
rect 12171 81367 12213 81376
rect 12020 81208 12116 81248
rect 12171 81248 12213 81257
rect 12171 81208 12172 81248
rect 12212 81208 12213 81248
rect 11980 81199 12020 81208
rect 12171 81199 12213 81208
rect 12172 81114 12212 81199
rect 11884 80695 11924 80704
rect 12268 80669 12308 82048
rect 12363 82088 12405 82097
rect 12363 82048 12364 82088
rect 12404 82048 12405 82088
rect 12363 82039 12405 82048
rect 12460 82088 12506 82097
rect 12505 82048 12506 82088
rect 12460 82039 12506 82048
rect 12364 81584 12404 82039
rect 12465 81958 12505 82039
rect 12364 81544 12500 81584
rect 12363 81416 12405 81425
rect 12363 81376 12364 81416
rect 12404 81376 12405 81416
rect 12363 81367 12405 81376
rect 12267 80660 12309 80669
rect 12267 80620 12268 80660
rect 12308 80620 12309 80660
rect 12267 80611 12309 80620
rect 11788 80527 11828 80536
rect 12076 80576 12116 80585
rect 11596 80368 11924 80408
rect 11499 80359 11541 80368
rect 11211 80240 11253 80249
rect 11211 80200 11212 80240
rect 11252 80200 11253 80240
rect 11211 80191 11253 80200
rect 11308 80240 11348 80359
rect 11500 80240 11540 80359
rect 11308 80200 11540 80240
rect 11115 79736 11157 79745
rect 11115 79696 11116 79736
rect 11156 79696 11157 79736
rect 11115 79687 11157 79696
rect 11116 79602 11156 79687
rect 11020 79108 11252 79148
rect 11212 79064 11252 79108
rect 11116 78980 11156 78989
rect 11020 78940 11116 78980
rect 10923 78224 10965 78233
rect 10676 78184 10868 78224
rect 10636 78175 10676 78184
rect 10540 78090 10580 78175
rect 10444 77636 10484 77645
rect 10484 77596 10772 77636
rect 10444 77587 10484 77596
rect 10252 77468 10292 77512
rect 10732 77552 10772 77596
rect 10732 77503 10772 77512
rect 10828 77552 10868 78184
rect 10923 78184 10924 78224
rect 10964 78184 10965 78224
rect 10923 78175 10965 78184
rect 11020 78224 11060 78940
rect 11116 78931 11156 78940
rect 10923 78056 10965 78065
rect 10923 78016 10924 78056
rect 10964 78016 10965 78056
rect 10923 78007 10965 78016
rect 10635 77468 10677 77477
rect 10252 77428 10580 77468
rect 10347 77216 10389 77225
rect 10347 77176 10348 77216
rect 10388 77176 10389 77216
rect 10347 77167 10389 77176
rect 9964 76677 10004 76686
rect 10155 76712 10197 76721
rect 10155 76672 10156 76712
rect 10196 76672 10197 76712
rect 10155 76663 10197 76672
rect 10156 76544 10196 76553
rect 10060 76504 10156 76544
rect 9675 76124 9717 76133
rect 9675 76084 9676 76124
rect 9716 76084 9717 76124
rect 9675 76075 9717 76084
rect 10060 75965 10100 76504
rect 10156 76495 10196 76504
rect 10155 76376 10197 76385
rect 10155 76336 10156 76376
rect 10196 76336 10197 76376
rect 10155 76327 10197 76336
rect 10156 76040 10196 76327
rect 10156 75991 10196 76000
rect 10059 75956 10101 75965
rect 10059 75916 10060 75956
rect 10100 75916 10101 75956
rect 10059 75907 10101 75916
rect 9867 75704 9909 75713
rect 9867 75664 9868 75704
rect 9908 75664 9909 75704
rect 9867 75655 9909 75664
rect 9771 75536 9813 75545
rect 9771 75496 9772 75536
rect 9812 75496 9813 75536
rect 9771 75487 9813 75496
rect 9772 75200 9812 75487
rect 9772 75151 9812 75160
rect 9580 75032 9620 75041
rect 9483 74612 9525 74621
rect 9483 74572 9484 74612
rect 9524 74572 9525 74612
rect 9483 74563 9525 74572
rect 9580 74537 9620 74992
rect 9771 74696 9813 74705
rect 9771 74656 9772 74696
rect 9812 74656 9813 74696
rect 9771 74647 9813 74656
rect 9579 74528 9621 74537
rect 9579 74488 9580 74528
rect 9620 74488 9621 74528
rect 9579 74479 9621 74488
rect 9676 74528 9716 74537
rect 9483 74192 9525 74201
rect 9483 74152 9484 74192
rect 9524 74152 9525 74192
rect 9483 74143 9525 74152
rect 9387 73268 9429 73277
rect 9387 73228 9388 73268
rect 9428 73228 9429 73268
rect 9387 73219 9429 73228
rect 9387 72428 9429 72437
rect 9387 72388 9388 72428
rect 9428 72388 9429 72428
rect 9484 72428 9524 74143
rect 9676 73856 9716 74488
rect 9772 74528 9812 74647
rect 9772 74479 9812 74488
rect 9868 74201 9908 75655
rect 9964 74696 10004 74705
rect 9867 74192 9909 74201
rect 9867 74152 9868 74192
rect 9908 74152 9909 74192
rect 9867 74143 9909 74152
rect 9964 73865 10004 74656
rect 10059 74612 10101 74621
rect 10059 74572 10060 74612
rect 10100 74572 10101 74612
rect 10059 74563 10101 74572
rect 10060 73940 10100 74563
rect 10251 74528 10293 74537
rect 10251 74488 10252 74528
rect 10292 74488 10293 74528
rect 10251 74479 10293 74488
rect 10348 74528 10388 77167
rect 10540 76805 10580 77428
rect 10635 77428 10636 77468
rect 10676 77428 10677 77468
rect 10635 77419 10677 77428
rect 10539 76796 10581 76805
rect 10539 76756 10540 76796
rect 10580 76756 10581 76796
rect 10539 76747 10581 76756
rect 10252 74394 10292 74479
rect 10348 74276 10388 74488
rect 10060 73891 10100 73900
rect 10252 74236 10388 74276
rect 9963 73856 10005 73865
rect 9676 73816 9812 73856
rect 9676 73688 9716 73697
rect 9676 73277 9716 73648
rect 9772 73361 9812 73816
rect 9963 73816 9964 73856
rect 10004 73816 10005 73856
rect 9963 73807 10005 73816
rect 10155 73856 10197 73865
rect 10155 73816 10156 73856
rect 10196 73816 10197 73856
rect 10155 73807 10197 73816
rect 10156 73703 10196 73807
rect 10060 73688 10100 73697
rect 10156 73654 10196 73663
rect 9867 73604 9909 73613
rect 9867 73564 9868 73604
rect 9908 73564 9909 73604
rect 9867 73555 9909 73564
rect 9868 73470 9908 73555
rect 9771 73352 9813 73361
rect 9771 73312 9772 73352
rect 9812 73312 9813 73352
rect 9771 73303 9813 73312
rect 9675 73268 9717 73277
rect 9675 73228 9676 73268
rect 9716 73228 9717 73268
rect 9675 73219 9717 73228
rect 9580 73016 9620 73044
rect 9676 73016 9716 73219
rect 9772 73100 9812 73303
rect 10060 73184 10100 73648
rect 10155 73520 10197 73529
rect 10155 73480 10156 73520
rect 10196 73480 10197 73520
rect 10155 73471 10197 73480
rect 10060 73135 10100 73144
rect 9812 73060 10004 73100
rect 9772 73051 9812 73060
rect 9620 72976 9716 73016
rect 9580 72967 9620 72976
rect 9484 72388 9620 72428
rect 9387 72379 9429 72388
rect 9195 72260 9237 72269
rect 9195 72220 9196 72260
rect 9236 72220 9237 72260
rect 9195 72211 9237 72220
rect 9388 72176 9428 72379
rect 9044 72136 9140 72176
rect 9004 72127 9044 72136
rect 8716 71800 8852 71840
rect 8523 71504 8565 71513
rect 8523 71464 8524 71504
rect 8564 71464 8565 71504
rect 8523 71455 8565 71464
rect 8428 71420 8468 71429
rect 8428 71093 8468 71380
rect 8524 71370 8564 71455
rect 8716 71168 8756 71800
rect 8811 71672 8853 71681
rect 8811 71632 8812 71672
rect 8852 71632 8853 71672
rect 8811 71623 8853 71632
rect 8812 71177 8852 71623
rect 9100 71597 9140 72136
rect 9388 72127 9428 72136
rect 9196 72008 9236 72017
rect 9236 71968 9524 72008
rect 9196 71959 9236 71968
rect 9291 71840 9333 71849
rect 9291 71800 9292 71840
rect 9332 71800 9333 71840
rect 9291 71791 9333 71800
rect 9099 71588 9141 71597
rect 9099 71548 9100 71588
rect 9140 71548 9141 71588
rect 9099 71539 9141 71548
rect 8907 71504 8949 71513
rect 8907 71464 8908 71504
rect 8948 71464 8949 71504
rect 8907 71455 8949 71464
rect 9004 71504 9044 71513
rect 8620 71128 8756 71168
rect 8811 71168 8853 71177
rect 8811 71128 8812 71168
rect 8852 71128 8853 71168
rect 8427 71084 8469 71093
rect 8427 71044 8428 71084
rect 8468 71044 8469 71084
rect 8427 71035 8469 71044
rect 8332 70876 8564 70916
rect 8332 70673 8372 70758
rect 8331 70664 8373 70673
rect 8331 70624 8332 70664
rect 8372 70624 8373 70664
rect 8331 70615 8373 70624
rect 8428 70664 8468 70673
rect 8140 70540 8276 70580
rect 8043 70531 8085 70540
rect 8236 70496 8276 70540
rect 8140 70456 8276 70496
rect 7947 70412 7989 70421
rect 7947 70372 7948 70412
rect 7988 70372 7989 70412
rect 7947 70363 7989 70372
rect 7948 70244 7988 70363
rect 7948 70204 8084 70244
rect 7947 70076 7989 70085
rect 7947 70036 7948 70076
rect 7988 70036 7989 70076
rect 7947 70027 7989 70036
rect 7948 69942 7988 70027
rect 7851 69236 7893 69245
rect 7851 69196 7852 69236
rect 7892 69196 7893 69236
rect 7851 69187 7893 69196
rect 7756 68480 7796 68489
rect 7852 68480 7892 69187
rect 7796 68440 7892 68480
rect 7756 68237 7796 68440
rect 7755 68228 7797 68237
rect 7755 68188 7756 68228
rect 7796 68188 7797 68228
rect 7755 68179 7797 68188
rect 7948 68228 7988 68237
rect 7948 68069 7988 68188
rect 7947 68060 7989 68069
rect 7947 68020 7948 68060
rect 7988 68020 7989 68060
rect 7947 68011 7989 68020
rect 7659 67808 7701 67817
rect 7659 67768 7660 67808
rect 7700 67768 7701 67808
rect 7659 67759 7701 67768
rect 7660 67640 7700 67759
rect 7660 67591 7700 67600
rect 7948 67640 7988 68011
rect 7948 67591 7988 67600
rect 8044 67640 8084 70204
rect 7563 66884 7605 66893
rect 7563 66844 7564 66884
rect 7604 66844 7605 66884
rect 7563 66835 7605 66844
rect 7467 66128 7509 66137
rect 7467 66088 7468 66128
rect 7508 66088 7509 66128
rect 7467 66079 7509 66088
rect 7564 66128 7604 66137
rect 7468 65994 7508 66079
rect 7372 65584 7508 65624
rect 7372 65456 7412 65465
rect 7276 65416 7372 65456
rect 7276 64793 7316 65416
rect 7372 65407 7412 65416
rect 7275 64784 7317 64793
rect 7275 64744 7276 64784
rect 7316 64744 7317 64784
rect 7275 64735 7317 64744
rect 7276 64621 7316 64630
rect 7276 64289 7316 64581
rect 7468 64532 7508 65584
rect 7564 65465 7604 66088
rect 7755 65960 7797 65969
rect 7755 65920 7756 65960
rect 7796 65920 7797 65960
rect 7755 65911 7797 65920
rect 7756 65826 7796 65911
rect 7755 65708 7797 65717
rect 7755 65668 7756 65708
rect 7796 65668 7797 65708
rect 7755 65659 7797 65668
rect 7563 65456 7605 65465
rect 7563 65416 7564 65456
rect 7604 65416 7605 65456
rect 7563 65407 7605 65416
rect 7756 65456 7796 65659
rect 7372 64492 7508 64532
rect 7564 65204 7604 65213
rect 7275 64280 7317 64289
rect 7275 64240 7276 64280
rect 7316 64240 7317 64280
rect 7275 64231 7317 64240
rect 7276 63944 7316 63953
rect 7276 63701 7316 63904
rect 7275 63692 7317 63701
rect 7275 63652 7276 63692
rect 7316 63652 7317 63692
rect 7275 63643 7317 63652
rect 7275 62348 7317 62357
rect 7180 62308 7276 62348
rect 7316 62308 7317 62348
rect 7084 62105 7124 62299
rect 7083 62096 7125 62105
rect 7083 62056 7084 62096
rect 7124 62056 7125 62096
rect 7083 62047 7125 62056
rect 7084 60173 7124 62047
rect 7180 60929 7220 62308
rect 7275 62299 7317 62308
rect 7275 62180 7317 62189
rect 7372 62180 7412 64492
rect 7468 64406 7508 64415
rect 7467 64366 7468 64373
rect 7508 64366 7509 64373
rect 7467 64364 7509 64366
rect 7467 64324 7468 64364
rect 7508 64324 7509 64364
rect 7467 64315 7509 64324
rect 7468 64271 7508 64315
rect 7564 64289 7604 65164
rect 7659 64532 7701 64541
rect 7659 64492 7660 64532
rect 7700 64492 7701 64532
rect 7659 64483 7701 64492
rect 7563 64280 7605 64289
rect 7563 64240 7564 64280
rect 7604 64240 7605 64280
rect 7563 64231 7605 64240
rect 7468 63692 7508 63701
rect 7508 63652 7604 63692
rect 7468 63643 7508 63652
rect 7467 63524 7509 63533
rect 7467 63484 7468 63524
rect 7508 63484 7509 63524
rect 7467 63475 7509 63484
rect 7275 62140 7276 62180
rect 7316 62140 7412 62180
rect 7275 62131 7317 62140
rect 7179 60920 7221 60929
rect 7179 60880 7180 60920
rect 7220 60880 7221 60920
rect 7179 60871 7221 60880
rect 7179 60752 7221 60761
rect 7179 60712 7180 60752
rect 7220 60712 7221 60752
rect 7179 60703 7221 60712
rect 7083 60164 7125 60173
rect 7083 60124 7084 60164
rect 7124 60124 7125 60164
rect 7083 60115 7125 60124
rect 7180 60164 7220 60703
rect 7084 60030 7124 60115
rect 6987 59996 7029 60005
rect 6987 59956 6988 59996
rect 7028 59956 7029 59996
rect 6987 59947 7029 59956
rect 7180 59828 7220 60124
rect 6700 59452 6836 59492
rect 6892 59788 7220 59828
rect 6316 59359 6356 59368
rect 6411 59408 6453 59417
rect 6411 59368 6412 59408
rect 6452 59368 6453 59408
rect 6411 59359 6453 59368
rect 6411 59156 6453 59165
rect 6411 59116 6412 59156
rect 6452 59116 6453 59156
rect 6411 59107 6453 59116
rect 6123 58988 6165 58997
rect 6123 58948 6124 58988
rect 6164 58948 6165 58988
rect 6123 58939 6165 58948
rect 6219 58736 6261 58745
rect 6219 58696 6220 58736
rect 6260 58696 6261 58736
rect 6219 58687 6261 58696
rect 6124 58400 6164 58409
rect 6124 57056 6164 58360
rect 6220 57896 6260 58687
rect 6315 58652 6357 58661
rect 6315 58612 6316 58652
rect 6356 58612 6357 58652
rect 6315 58603 6357 58612
rect 6316 58568 6356 58603
rect 6316 58517 6356 58528
rect 6220 57847 6260 57856
rect 6220 57056 6260 57065
rect 6124 57016 6220 57056
rect 6220 57007 6260 57016
rect 6316 57056 6356 57065
rect 6412 57056 6452 59107
rect 6700 59072 6740 59452
rect 6892 59408 6932 59788
rect 7372 59669 7412 62140
rect 7468 61601 7508 63475
rect 7564 63118 7604 63652
rect 7660 63113 7700 64483
rect 7756 63785 7796 65416
rect 8044 65297 8084 67600
rect 8140 68480 8180 70456
rect 8428 70421 8468 70624
rect 8427 70412 8469 70421
rect 8427 70372 8428 70412
rect 8468 70372 8469 70412
rect 8427 70363 8469 70372
rect 8524 70244 8564 70876
rect 8140 66809 8180 68440
rect 8236 70204 8564 70244
rect 8139 66800 8181 66809
rect 8139 66760 8140 66800
rect 8180 66760 8181 66800
rect 8139 66751 8181 66760
rect 8043 65288 8085 65297
rect 8043 65248 8044 65288
rect 8084 65248 8085 65288
rect 8043 65239 8085 65248
rect 7947 65120 7989 65129
rect 7947 65080 7948 65120
rect 7988 65080 7989 65120
rect 7947 65071 7989 65080
rect 7852 64625 7892 64710
rect 7851 64616 7893 64625
rect 7851 64576 7852 64616
rect 7892 64576 7893 64616
rect 7851 64567 7893 64576
rect 7851 64448 7893 64457
rect 7851 64408 7852 64448
rect 7892 64408 7893 64448
rect 7851 64399 7893 64408
rect 7755 63776 7797 63785
rect 7755 63736 7756 63776
rect 7796 63736 7797 63776
rect 7755 63727 7797 63736
rect 7564 63069 7604 63078
rect 7659 63104 7701 63113
rect 7659 63064 7660 63104
rect 7700 63064 7701 63104
rect 7659 63055 7701 63064
rect 7563 62600 7605 62609
rect 7563 62560 7564 62600
rect 7604 62560 7605 62600
rect 7563 62551 7605 62560
rect 7467 61592 7509 61601
rect 7467 61552 7468 61592
rect 7508 61552 7509 61592
rect 7467 61543 7509 61552
rect 7467 60836 7509 60845
rect 7467 60796 7468 60836
rect 7508 60796 7509 60836
rect 7467 60787 7509 60796
rect 7371 59660 7413 59669
rect 7371 59620 7372 59660
rect 7412 59620 7413 59660
rect 7371 59611 7413 59620
rect 6892 59359 6932 59368
rect 7372 59408 7412 59417
rect 6796 59324 6836 59335
rect 6796 59249 6836 59284
rect 6795 59240 6837 59249
rect 6795 59200 6796 59240
rect 6836 59200 6837 59240
rect 6795 59191 6837 59200
rect 7179 59240 7221 59249
rect 7179 59200 7180 59240
rect 7220 59200 7221 59240
rect 7179 59191 7221 59200
rect 6700 59032 7124 59072
rect 6507 58988 6549 58997
rect 6507 58948 6508 58988
rect 6548 58948 6549 58988
rect 6507 58939 6549 58948
rect 6356 57016 6452 57056
rect 6028 56335 6068 56344
rect 5932 54116 5972 55504
rect 6124 55376 6164 55385
rect 6028 55336 6124 55376
rect 6028 54872 6068 55336
rect 6124 55327 6164 55336
rect 6316 55124 6356 57016
rect 6411 56636 6453 56645
rect 6411 56596 6412 56636
rect 6452 56596 6453 56636
rect 6411 56587 6453 56596
rect 6412 56309 6452 56587
rect 6411 56300 6453 56309
rect 6411 56260 6412 56300
rect 6452 56260 6453 56300
rect 6411 56251 6453 56260
rect 6028 54823 6068 54832
rect 6124 55084 6356 55124
rect 6508 55544 6548 58939
rect 6987 58904 7029 58913
rect 6987 58864 6988 58904
rect 7028 58864 7029 58904
rect 6987 58855 7029 58864
rect 6795 58484 6837 58493
rect 6795 58444 6796 58484
rect 6836 58444 6837 58484
rect 6795 58435 6837 58444
rect 6796 57401 6836 58435
rect 6795 57392 6837 57401
rect 6795 57352 6796 57392
rect 6836 57352 6837 57392
rect 6795 57343 6837 57352
rect 6700 57056 6740 57065
rect 6700 56225 6740 57016
rect 6796 57056 6836 57343
rect 6699 56216 6741 56225
rect 6699 56176 6700 56216
rect 6740 56176 6741 56216
rect 6699 56167 6741 56176
rect 6124 54872 6164 55084
rect 6508 54956 6548 55504
rect 6124 54545 6164 54832
rect 6412 54916 6548 54956
rect 6603 54956 6645 54965
rect 6603 54916 6604 54956
rect 6644 54916 6645 54956
rect 6123 54536 6165 54545
rect 6123 54496 6124 54536
rect 6164 54496 6165 54536
rect 6123 54487 6165 54496
rect 6315 54452 6357 54461
rect 6315 54412 6316 54452
rect 6356 54412 6357 54452
rect 6315 54403 6357 54412
rect 5932 54076 6068 54116
rect 5836 53992 5972 54032
rect 5643 53983 5685 53992
rect 5836 53864 5876 53873
rect 4588 53404 4724 53444
rect 4492 52781 4532 53236
rect 4588 53276 4628 53285
rect 4588 53033 4628 53236
rect 4587 53024 4629 53033
rect 4587 52984 4588 53024
rect 4628 52984 4629 53024
rect 4587 52975 4629 52984
rect 4491 52772 4533 52781
rect 4491 52732 4492 52772
rect 4532 52732 4533 52772
rect 4491 52723 4533 52732
rect 4684 52697 4724 53404
rect 5452 53404 5588 53444
rect 5644 53824 5836 53864
rect 5068 53360 5108 53369
rect 5068 52949 5108 53320
rect 5067 52940 5109 52949
rect 5067 52900 5068 52940
rect 5108 52900 5109 52940
rect 5067 52891 5109 52900
rect 5355 52940 5397 52949
rect 5355 52900 5356 52940
rect 5396 52900 5397 52940
rect 5355 52891 5397 52900
rect 4971 52856 5013 52865
rect 4971 52816 4972 52856
rect 5012 52816 5013 52856
rect 4971 52807 5013 52816
rect 4683 52688 4725 52697
rect 4683 52648 4684 52688
rect 4724 52648 4725 52688
rect 4683 52639 4725 52648
rect 4780 52525 4820 52534
rect 4491 52436 4533 52445
rect 4491 52396 4492 52436
rect 4532 52396 4533 52436
rect 4491 52387 4533 52396
rect 4012 50959 4052 50968
rect 4108 51010 4244 51050
rect 4108 51008 4148 51010
rect 4108 50959 4148 50968
rect 3147 50336 3189 50345
rect 3147 50296 3148 50336
rect 3188 50296 3189 50336
rect 3147 50287 3189 50296
rect 3244 49496 3284 50959
rect 4204 50933 4244 51010
rect 4300 51976 4436 52016
rect 4203 50924 4245 50933
rect 4203 50884 4204 50924
rect 4244 50884 4245 50924
rect 4203 50875 4245 50884
rect 3915 50336 3957 50345
rect 3915 50296 3916 50336
rect 3956 50296 3957 50336
rect 3915 50287 3957 50296
rect 4300 50336 4340 51976
rect 4396 51848 4436 51857
rect 4492 51848 4532 52387
rect 4780 52100 4820 52485
rect 4972 52436 5012 52807
rect 4972 52387 5012 52396
rect 4928 52184 5296 52193
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 4928 52135 5296 52144
rect 4588 52060 4820 52100
rect 4588 52016 4628 52060
rect 4588 51967 4628 51976
rect 5067 52016 5109 52025
rect 5067 51976 5068 52016
rect 5108 51976 5109 52016
rect 5067 51967 5109 51976
rect 4780 51848 4820 51857
rect 4492 51808 4724 51848
rect 4396 51773 4436 51808
rect 4395 51764 4437 51773
rect 4395 51724 4396 51764
rect 4436 51724 4437 51764
rect 4395 51715 4437 51724
rect 4396 51185 4436 51715
rect 4395 51176 4437 51185
rect 4395 51136 4396 51176
rect 4436 51136 4437 51176
rect 4395 51127 4437 51136
rect 4587 51176 4629 51185
rect 4587 51136 4588 51176
rect 4628 51136 4629 51176
rect 4587 51127 4629 51136
rect 4588 51092 4628 51127
rect 4588 51041 4628 51052
rect 4491 51008 4533 51017
rect 4491 50968 4492 51008
rect 4532 50968 4533 51008
rect 4491 50959 4533 50968
rect 4395 50924 4437 50933
rect 4395 50884 4396 50924
rect 4436 50884 4437 50924
rect 4395 50875 4437 50884
rect 3916 50202 3956 50287
rect 4300 50261 4340 50296
rect 4299 50252 4341 50261
rect 4299 50212 4300 50252
rect 4340 50212 4341 50252
rect 4299 50203 4341 50212
rect 4108 50084 4148 50093
rect 3688 49916 4056 49925
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 4108 49916 4148 50044
rect 4108 49876 4340 49916
rect 3688 49867 4056 49876
rect 4107 49748 4149 49757
rect 4107 49708 4108 49748
rect 4148 49708 4149 49748
rect 4107 49699 4149 49708
rect 3244 47993 3284 49456
rect 3340 49496 3380 49505
rect 3340 48833 3380 49456
rect 3820 49496 3860 49505
rect 4108 49496 4148 49699
rect 3860 49456 4148 49496
rect 4300 49510 4340 49876
rect 4300 49461 4340 49470
rect 3820 49447 3860 49456
rect 3819 49244 3861 49253
rect 3819 49204 3820 49244
rect 3860 49204 3861 49244
rect 3819 49195 3861 49204
rect 3339 48824 3381 48833
rect 3339 48784 3340 48824
rect 3380 48784 3381 48824
rect 3339 48775 3381 48784
rect 3820 48824 3860 49195
rect 3340 48068 3380 48775
rect 3820 48572 3860 48784
rect 4012 48581 4052 48666
rect 3340 48019 3380 48028
rect 3532 48532 3860 48572
rect 4011 48572 4053 48581
rect 4011 48532 4012 48572
rect 4052 48532 4053 48572
rect 3243 47984 3285 47993
rect 3243 47944 3244 47984
rect 3284 47944 3285 47984
rect 3243 47935 3285 47944
rect 3244 47850 3284 47935
rect 3532 47732 3572 48532
rect 4011 48523 4053 48532
rect 3688 48404 4056 48413
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 3688 48355 4056 48364
rect 3820 47984 3860 47993
rect 3820 47825 3860 47944
rect 4108 47825 4148 49456
rect 4204 48824 4244 48835
rect 4204 48749 4244 48784
rect 4203 48740 4245 48749
rect 4203 48700 4204 48740
rect 4244 48700 4245 48740
rect 4203 48691 4245 48700
rect 4299 48572 4341 48581
rect 4299 48532 4300 48572
rect 4340 48532 4341 48572
rect 4299 48523 4341 48532
rect 4300 47998 4340 48523
rect 4300 47949 4340 47958
rect 3819 47816 3861 47825
rect 3819 47776 3820 47816
rect 3860 47776 3861 47816
rect 3819 47767 3861 47776
rect 4107 47816 4149 47825
rect 4107 47776 4108 47816
rect 4148 47776 4149 47816
rect 4107 47767 4149 47776
rect 3148 47692 3572 47732
rect 3148 47312 3188 47692
rect 3339 47396 3381 47405
rect 3339 47356 3340 47396
rect 3380 47356 3381 47396
rect 3339 47347 3381 47356
rect 3819 47396 3861 47405
rect 3819 47356 3820 47396
rect 3860 47356 3861 47396
rect 3819 47347 3861 47356
rect 3148 46733 3188 47272
rect 3340 47262 3380 47347
rect 3820 47312 3860 47347
rect 3820 47261 3860 47272
rect 3915 47312 3957 47321
rect 3915 47272 3916 47312
rect 3956 47272 3957 47312
rect 3915 47263 3957 47272
rect 4299 47312 4341 47321
rect 4299 47272 4300 47312
rect 4340 47272 4341 47312
rect 4299 47263 4341 47272
rect 4396 47312 4436 50875
rect 4492 50874 4532 50959
rect 4684 49757 4724 51808
rect 4780 51185 4820 51808
rect 4779 51176 4821 51185
rect 4779 51136 4780 51176
rect 4820 51136 4821 51176
rect 4779 51127 4821 51136
rect 4683 49748 4725 49757
rect 4683 49708 4684 49748
rect 4724 49708 4725 49748
rect 4683 49699 4725 49708
rect 4587 49496 4629 49505
rect 4587 49456 4588 49496
rect 4628 49456 4629 49496
rect 4587 49447 4629 49456
rect 4684 49496 4724 49505
rect 4780 49496 4820 51127
rect 5068 51008 5108 51967
rect 5068 50933 5108 50968
rect 5067 50924 5109 50933
rect 5067 50884 5068 50924
rect 5108 50884 5109 50924
rect 5067 50875 5109 50884
rect 5068 50844 5108 50875
rect 4928 50672 5296 50681
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 4928 50623 5296 50632
rect 4875 50252 4917 50261
rect 4875 50212 4876 50252
rect 4916 50212 4917 50252
rect 4875 50203 4917 50212
rect 4724 49456 4820 49496
rect 4684 49447 4724 49456
rect 4491 49328 4533 49337
rect 4491 49288 4492 49328
rect 4532 49288 4533 49328
rect 4491 49279 4533 49288
rect 4492 49194 4532 49279
rect 4491 47900 4533 47909
rect 4491 47860 4492 47900
rect 4532 47860 4533 47900
rect 4491 47851 4533 47860
rect 4492 47766 4532 47851
rect 3916 47178 3956 47263
rect 3688 46892 4056 46901
rect 4300 46892 4340 47263
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 3688 46843 4056 46852
rect 4204 46852 4340 46892
rect 3147 46724 3189 46733
rect 3147 46684 3148 46724
rect 3188 46684 3189 46724
rect 3147 46675 3189 46684
rect 3051 46556 3093 46565
rect 3051 46516 3052 46556
rect 3092 46516 3093 46556
rect 3051 46507 3093 46516
rect 3435 46556 3477 46565
rect 3435 46516 3436 46556
rect 3476 46516 3477 46556
rect 3435 46507 3477 46516
rect 3052 46422 3092 46507
rect 3243 46472 3285 46481
rect 3243 46432 3244 46472
rect 3284 46432 3285 46472
rect 3243 46423 3285 46432
rect 3244 46304 3284 46423
rect 3436 46422 3476 46507
rect 4108 46472 4148 46481
rect 3244 46255 3284 46264
rect 3339 46220 3381 46229
rect 3339 46180 3340 46220
rect 3380 46180 3381 46220
rect 3339 46171 3381 46180
rect 2900 45676 2996 45716
rect 2860 45667 2900 45676
rect 2763 45212 2805 45221
rect 2763 45172 2764 45212
rect 2804 45172 2805 45212
rect 2763 45163 2805 45172
rect 3243 44960 3285 44969
rect 3243 44920 3244 44960
rect 3284 44920 3285 44960
rect 3243 44911 3285 44920
rect 3244 44826 3284 44911
rect 2475 44372 2517 44381
rect 2475 44332 2476 44372
rect 2516 44332 2517 44372
rect 2475 44323 2517 44332
rect 1996 44239 2036 44248
rect 3244 44288 3284 44297
rect 3340 44288 3380 46171
rect 4108 45809 4148 46432
rect 4107 45800 4149 45809
rect 4107 45760 4108 45800
rect 4148 45760 4149 45800
rect 4107 45751 4149 45760
rect 3688 45380 4056 45389
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 3688 45331 4056 45340
rect 3915 45212 3957 45221
rect 3915 45172 3916 45212
rect 3956 45172 3957 45212
rect 3915 45163 3957 45172
rect 3724 44960 3764 44969
rect 3436 44792 3476 44801
rect 3436 44297 3476 44752
rect 3284 44248 3380 44288
rect 3435 44288 3477 44297
rect 3435 44248 3436 44288
rect 3476 44248 3477 44288
rect 3244 44239 3284 44248
rect 3435 44239 3477 44248
rect 1803 44204 1845 44213
rect 1803 44164 1804 44204
rect 1844 44164 1845 44204
rect 1803 44155 1845 44164
rect 1804 44070 1844 44155
rect 3436 44120 3476 44129
rect 3724 44120 3764 44920
rect 3820 44960 3860 44969
rect 3820 44801 3860 44920
rect 3819 44792 3861 44801
rect 3819 44752 3820 44792
rect 3860 44752 3861 44792
rect 3819 44743 3861 44752
rect 3819 44288 3861 44297
rect 3819 44248 3820 44288
rect 3860 44248 3861 44288
rect 3819 44239 3861 44248
rect 3916 44288 3956 45163
rect 4204 45044 4244 46852
rect 4396 46817 4436 47272
rect 4395 46808 4437 46817
rect 4204 44288 4244 45004
rect 4300 46768 4396 46808
rect 4436 46768 4437 46808
rect 4300 45044 4340 46768
rect 4395 46759 4437 46768
rect 4588 46640 4628 49447
rect 4876 49412 4916 50203
rect 4780 49372 4916 49412
rect 4780 48749 4820 49372
rect 4928 49160 5296 49169
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 4928 49111 5296 49120
rect 5356 48833 5396 52891
rect 5452 52781 5492 53404
rect 5644 53360 5684 53824
rect 5836 53815 5876 53824
rect 5739 53696 5781 53705
rect 5739 53656 5740 53696
rect 5780 53656 5781 53696
rect 5739 53647 5781 53656
rect 5740 53528 5780 53647
rect 5740 53479 5780 53488
rect 5835 53444 5877 53453
rect 5835 53404 5836 53444
rect 5876 53404 5877 53444
rect 5835 53395 5877 53404
rect 5596 53350 5684 53360
rect 5636 53320 5684 53350
rect 5596 53301 5636 53310
rect 5739 53276 5781 53285
rect 5739 53236 5740 53276
rect 5780 53236 5781 53276
rect 5739 53227 5781 53236
rect 5451 52772 5493 52781
rect 5451 52732 5452 52772
rect 5492 52732 5493 52772
rect 5451 52723 5493 52732
rect 5548 51013 5588 51022
rect 5452 50973 5548 51008
rect 5452 50968 5588 50973
rect 5452 50513 5492 50968
rect 5548 50964 5588 50968
rect 5740 50924 5780 53227
rect 5836 51521 5876 53395
rect 5835 51512 5877 51521
rect 5835 51472 5836 51512
rect 5876 51472 5877 51512
rect 5835 51463 5877 51472
rect 5835 51344 5877 51353
rect 5835 51304 5836 51344
rect 5876 51304 5877 51344
rect 5835 51295 5877 51304
rect 5740 50875 5780 50884
rect 5547 50756 5589 50765
rect 5547 50716 5548 50756
rect 5588 50716 5589 50756
rect 5547 50707 5589 50716
rect 5451 50504 5493 50513
rect 5451 50464 5452 50504
rect 5492 50464 5493 50504
rect 5451 50455 5493 50464
rect 5548 50336 5588 50707
rect 5740 50513 5780 50598
rect 5739 50504 5781 50513
rect 5739 50464 5740 50504
rect 5780 50464 5781 50504
rect 5739 50455 5781 50464
rect 5548 50168 5588 50296
rect 5548 50128 5780 50168
rect 5643 49748 5685 49757
rect 5643 49708 5644 49748
rect 5684 49708 5685 49748
rect 5643 49699 5685 49708
rect 5644 49253 5684 49699
rect 5643 49244 5685 49253
rect 5643 49204 5644 49244
rect 5684 49204 5685 49244
rect 5643 49195 5685 49204
rect 5355 48824 5397 48833
rect 5355 48784 5356 48824
rect 5396 48784 5397 48824
rect 5355 48775 5397 48784
rect 5452 48824 5492 48833
rect 5644 48824 5684 49195
rect 5492 48784 5684 48824
rect 5452 48775 5492 48784
rect 4779 48740 4821 48749
rect 4779 48700 4780 48740
rect 4820 48700 4821 48740
rect 4779 48691 4821 48700
rect 5644 48572 5684 48581
rect 5452 48532 5644 48572
rect 4779 48404 4821 48413
rect 4779 48364 4780 48404
rect 4820 48364 4821 48404
rect 4779 48355 4821 48364
rect 4780 47984 4820 48355
rect 4780 47935 4820 47944
rect 4928 47648 5296 47657
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 4928 47599 5296 47608
rect 4876 47312 4916 47321
rect 5452 47312 5492 48532
rect 5644 48523 5684 48532
rect 5740 47984 5780 50128
rect 5836 49337 5876 51295
rect 5932 51176 5972 53992
rect 6028 53453 6068 54076
rect 6123 54032 6165 54041
rect 6123 53992 6124 54032
rect 6164 53992 6165 54032
rect 6123 53983 6165 53992
rect 6316 54032 6356 54403
rect 6027 53444 6069 53453
rect 6027 53404 6028 53444
rect 6068 53404 6069 53444
rect 6027 53395 6069 53404
rect 6028 51848 6068 51859
rect 6124 51848 6164 53983
rect 6219 52184 6261 52193
rect 6219 52144 6220 52184
rect 6260 52144 6261 52184
rect 6219 52135 6261 52144
rect 6220 52016 6260 52135
rect 6220 51967 6260 51976
rect 6124 51808 6260 51848
rect 6028 51773 6068 51808
rect 6027 51764 6069 51773
rect 6027 51724 6028 51764
rect 6068 51724 6069 51764
rect 6027 51715 6069 51724
rect 6123 51512 6165 51521
rect 6123 51472 6124 51512
rect 6164 51472 6165 51512
rect 6123 51463 6165 51472
rect 5932 51136 6068 51176
rect 5931 51008 5973 51017
rect 5931 50968 5932 51008
rect 5972 50968 5973 51008
rect 5931 50959 5973 50968
rect 5932 50336 5972 50959
rect 5932 50287 5972 50296
rect 5931 50168 5973 50177
rect 5931 50128 5932 50168
rect 5972 50128 5973 50168
rect 5931 50119 5973 50128
rect 5932 49757 5972 50119
rect 5931 49748 5973 49757
rect 5931 49708 5932 49748
rect 5972 49708 5973 49748
rect 5931 49699 5973 49708
rect 5932 49496 5972 49699
rect 6028 49505 6068 51136
rect 6124 50345 6164 51463
rect 6123 50336 6165 50345
rect 6123 50296 6124 50336
rect 6164 50296 6165 50336
rect 6123 50287 6165 50296
rect 5932 49447 5972 49456
rect 6027 49496 6069 49505
rect 6027 49456 6028 49496
rect 6068 49456 6069 49496
rect 6027 49447 6069 49456
rect 5835 49328 5877 49337
rect 6124 49328 6164 49337
rect 5835 49288 5836 49328
rect 5876 49288 5877 49328
rect 5835 49279 5877 49288
rect 5932 49288 6124 49328
rect 5932 48824 5972 49288
rect 6124 49279 6164 49288
rect 6220 49160 6260 51808
rect 6124 49120 6260 49160
rect 5932 48775 5972 48784
rect 6028 48824 6068 48833
rect 6028 48245 6068 48784
rect 6027 48236 6069 48245
rect 6027 48196 6028 48236
rect 6068 48196 6069 48236
rect 6027 48187 6069 48196
rect 6028 47984 6068 47993
rect 5740 47944 6028 47984
rect 6028 47657 6068 47944
rect 6027 47648 6069 47657
rect 6027 47608 6028 47648
rect 6068 47608 6069 47648
rect 6027 47599 6069 47608
rect 4876 46640 4916 47272
rect 5404 47302 5492 47312
rect 5444 47272 5492 47302
rect 5548 47396 5588 47405
rect 5404 47253 5444 47262
rect 4492 46600 4628 46640
rect 4780 46600 4916 46640
rect 4395 45800 4437 45809
rect 4395 45760 4396 45800
rect 4436 45760 4437 45800
rect 4395 45751 4437 45760
rect 4396 45666 4436 45751
rect 4300 44465 4340 45004
rect 4299 44456 4341 44465
rect 4299 44416 4300 44456
rect 4340 44416 4341 44456
rect 4299 44407 4341 44416
rect 4300 44288 4340 44297
rect 4204 44248 4300 44288
rect 3916 44239 3956 44248
rect 4300 44239 4340 44248
rect 4396 44288 4436 44297
rect 4492 44288 4532 46600
rect 4780 45389 4820 46600
rect 5548 46565 5588 47356
rect 5547 46556 5589 46565
rect 5547 46516 5548 46556
rect 5588 46516 5589 46556
rect 5547 46507 5589 46516
rect 5356 46472 5396 46481
rect 5356 46229 5396 46432
rect 5548 46304 5588 46313
rect 5355 46220 5397 46229
rect 5355 46180 5356 46220
rect 5396 46180 5397 46220
rect 5355 46171 5397 46180
rect 4928 46136 5296 46145
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 4928 46087 5296 46096
rect 4779 45380 4821 45389
rect 4779 45340 4780 45380
rect 4820 45340 4821 45380
rect 4779 45331 4821 45340
rect 4780 44960 4820 45331
rect 5308 45002 5348 45011
rect 5548 45002 5588 46264
rect 6028 46229 6068 47599
rect 6027 46220 6069 46229
rect 6027 46180 6028 46220
rect 6068 46180 6069 46220
rect 6027 46171 6069 46180
rect 6124 46052 6164 49120
rect 6316 48413 6356 53992
rect 6412 51017 6452 54916
rect 6603 54907 6645 54916
rect 6604 54872 6644 54907
rect 6604 54821 6644 54832
rect 6508 54788 6548 54797
rect 6508 54704 6548 54748
rect 6700 54704 6740 56167
rect 6796 54965 6836 57016
rect 6988 56981 7028 58855
rect 6987 56972 7029 56981
rect 6987 56932 6988 56972
rect 7028 56932 7029 56972
rect 6987 56923 7029 56932
rect 6987 56804 7029 56813
rect 6987 56764 6988 56804
rect 7028 56764 7029 56804
rect 6987 56755 7029 56764
rect 6988 55544 7028 56755
rect 7084 56393 7124 59032
rect 7083 56384 7125 56393
rect 7083 56344 7084 56384
rect 7124 56344 7125 56384
rect 7083 56335 7125 56344
rect 7084 56132 7124 56335
rect 7180 56216 7220 59191
rect 7372 58493 7412 59368
rect 7468 58997 7508 60787
rect 7467 58988 7509 58997
rect 7467 58948 7468 58988
rect 7508 58948 7509 58988
rect 7564 58988 7604 62551
rect 7660 62432 7700 63055
rect 7756 62936 7796 62945
rect 7756 62609 7796 62896
rect 7755 62600 7797 62609
rect 7755 62560 7756 62600
rect 7796 62560 7797 62600
rect 7755 62551 7797 62560
rect 7756 62432 7796 62441
rect 7660 62392 7756 62432
rect 7756 62383 7796 62392
rect 7659 61592 7701 61601
rect 7756 61592 7796 61601
rect 7659 61552 7660 61592
rect 7700 61552 7756 61592
rect 7659 61543 7701 61552
rect 7756 61543 7796 61552
rect 7660 61181 7700 61543
rect 7659 61172 7701 61181
rect 7659 61132 7660 61172
rect 7700 61132 7701 61172
rect 7659 61123 7701 61132
rect 7660 60257 7700 61123
rect 7755 61088 7797 61097
rect 7755 61048 7756 61088
rect 7796 61048 7797 61088
rect 7755 61039 7797 61048
rect 7659 60248 7701 60257
rect 7659 60208 7660 60248
rect 7700 60208 7701 60248
rect 7659 60199 7701 60208
rect 7660 60080 7700 60089
rect 7660 59921 7700 60040
rect 7659 59912 7701 59921
rect 7659 59872 7660 59912
rect 7700 59872 7701 59912
rect 7659 59863 7701 59872
rect 7756 59240 7796 61039
rect 7852 60593 7892 64399
rect 7948 62684 7988 65071
rect 8236 64280 8276 70204
rect 8620 70160 8660 71128
rect 8811 71119 8853 71128
rect 8715 70916 8757 70925
rect 8715 70876 8716 70916
rect 8756 70876 8757 70916
rect 8715 70867 8757 70876
rect 8524 70120 8660 70160
rect 8524 69236 8564 70120
rect 8716 70076 8756 70867
rect 8811 70664 8853 70673
rect 8811 70624 8812 70664
rect 8852 70624 8853 70664
rect 8811 70615 8853 70624
rect 8908 70664 8948 71455
rect 9004 70925 9044 71464
rect 9003 70916 9045 70925
rect 9003 70876 9004 70916
rect 9044 70876 9045 70916
rect 9003 70867 9045 70876
rect 9100 70841 9140 71539
rect 9099 70832 9141 70841
rect 9099 70792 9100 70832
rect 9140 70792 9141 70832
rect 9099 70783 9141 70792
rect 8812 70530 8852 70615
rect 8716 70036 8852 70076
rect 8626 69992 8668 70001
rect 8626 69952 8627 69992
rect 8667 69952 8756 69992
rect 8626 69943 8668 69952
rect 8716 69950 8756 69952
rect 8716 69901 8756 69910
rect 8812 69824 8852 70036
rect 8524 69187 8564 69196
rect 8716 69784 8852 69824
rect 8427 69152 8469 69161
rect 8427 69112 8428 69152
rect 8468 69112 8469 69152
rect 8427 69103 8469 69112
rect 8620 69152 8660 69161
rect 8331 69068 8373 69077
rect 8331 69028 8332 69068
rect 8372 69028 8373 69068
rect 8331 69019 8373 69028
rect 8140 64240 8276 64280
rect 8043 63944 8085 63953
rect 8043 63904 8044 63944
rect 8084 63904 8085 63944
rect 8043 63895 8085 63904
rect 8044 63104 8084 63895
rect 8044 63055 8084 63064
rect 7948 62644 8084 62684
rect 7947 62180 7989 62189
rect 7947 62140 7948 62180
rect 7988 62140 7989 62180
rect 7947 62131 7989 62140
rect 7948 62046 7988 62131
rect 7948 61424 7988 61433
rect 7851 60584 7893 60593
rect 7851 60544 7852 60584
rect 7892 60544 7893 60584
rect 7851 60535 7893 60544
rect 7948 60416 7988 61384
rect 7852 60376 7988 60416
rect 7852 59403 7892 60376
rect 8044 59660 8084 62644
rect 8140 61097 8180 64240
rect 8235 64112 8277 64121
rect 8235 64072 8236 64112
rect 8276 64072 8277 64112
rect 8235 64063 8277 64072
rect 8236 63978 8276 64063
rect 8332 63953 8372 69019
rect 8428 69018 8468 69103
rect 8620 68405 8660 69112
rect 8619 68396 8661 68405
rect 8619 68356 8620 68396
rect 8660 68356 8661 68396
rect 8619 68347 8661 68356
rect 8427 67724 8469 67733
rect 8427 67684 8428 67724
rect 8468 67684 8469 67724
rect 8427 67675 8469 67684
rect 8428 67565 8468 67675
rect 8524 67640 8564 67649
rect 8427 67556 8469 67565
rect 8427 67516 8428 67556
rect 8468 67516 8469 67556
rect 8427 67507 8469 67516
rect 8427 67052 8469 67061
rect 8427 67012 8428 67052
rect 8468 67012 8469 67052
rect 8427 67003 8469 67012
rect 8428 66968 8468 67003
rect 8428 66917 8468 66928
rect 8524 66641 8564 67600
rect 8619 67136 8661 67145
rect 8619 67096 8620 67136
rect 8660 67096 8661 67136
rect 8619 67087 8661 67096
rect 8620 67002 8660 67087
rect 8619 66800 8661 66809
rect 8619 66760 8620 66800
rect 8660 66760 8661 66800
rect 8619 66751 8661 66760
rect 8523 66632 8565 66641
rect 8523 66592 8524 66632
rect 8564 66592 8565 66632
rect 8523 66583 8565 66592
rect 8620 66473 8660 66751
rect 8619 66464 8661 66473
rect 8619 66424 8620 66464
rect 8660 66424 8661 66464
rect 8619 66415 8661 66424
rect 8716 66296 8756 69784
rect 8908 69245 8948 70624
rect 8907 69236 8949 69245
rect 8907 69196 8908 69236
rect 8948 69196 8949 69236
rect 8907 69187 8949 69196
rect 8812 69152 8852 69161
rect 8812 67817 8852 69112
rect 8908 69152 8948 69187
rect 8908 69101 8948 69112
rect 9004 69152 9044 69161
rect 8907 68060 8949 68069
rect 9004 68060 9044 69112
rect 9100 68984 9140 68993
rect 9100 68069 9140 68944
rect 8907 68020 8908 68060
rect 8948 68020 9044 68060
rect 9099 68060 9141 68069
rect 9099 68020 9100 68060
rect 9140 68020 9141 68060
rect 8907 68011 8949 68020
rect 9099 68011 9141 68020
rect 8811 67808 8853 67817
rect 8811 67768 8812 67808
rect 8852 67768 8853 67808
rect 8811 67759 8853 67768
rect 8812 67145 8852 67759
rect 8908 67472 8948 68011
rect 9292 67985 9332 71791
rect 9484 71499 9524 71968
rect 9484 71450 9524 71459
rect 9387 70916 9429 70925
rect 9387 70876 9388 70916
rect 9428 70876 9429 70916
rect 9387 70867 9429 70876
rect 9388 70664 9428 70867
rect 9388 70615 9428 70624
rect 9483 70664 9525 70673
rect 9483 70624 9484 70664
rect 9524 70624 9525 70664
rect 9483 70615 9525 70624
rect 9387 68900 9429 68909
rect 9387 68860 9388 68900
rect 9428 68860 9429 68900
rect 9387 68851 9429 68860
rect 9388 68480 9428 68851
rect 9484 68480 9524 70615
rect 9580 69152 9620 72388
rect 9676 72101 9716 72976
rect 9964 73016 10004 73060
rect 9964 72967 10004 72976
rect 10156 73016 10196 73471
rect 10252 73193 10292 74236
rect 10443 73856 10485 73865
rect 10443 73816 10444 73856
rect 10484 73816 10485 73856
rect 10443 73807 10485 73816
rect 10348 73697 10388 73782
rect 10444 73717 10484 73807
rect 10347 73688 10389 73697
rect 10347 73648 10348 73688
rect 10388 73648 10389 73688
rect 10636 73697 10676 77419
rect 10828 77225 10868 77512
rect 10827 77216 10869 77225
rect 10827 77176 10828 77216
rect 10868 77176 10869 77216
rect 10827 77167 10869 77176
rect 10827 76880 10869 76889
rect 10827 76840 10828 76880
rect 10868 76840 10869 76880
rect 10827 76831 10869 76840
rect 10828 74705 10868 76831
rect 10924 76544 10964 78007
rect 11020 77552 11060 78184
rect 11116 78308 11156 78317
rect 11212 78308 11252 79024
rect 11156 78268 11252 78308
rect 11116 77636 11156 78268
rect 11308 78065 11348 80200
rect 11403 79988 11445 79997
rect 11403 79948 11404 79988
rect 11444 79948 11445 79988
rect 11403 79939 11445 79948
rect 11404 79745 11444 79939
rect 11691 79904 11733 79913
rect 11691 79864 11692 79904
rect 11732 79864 11733 79904
rect 11691 79855 11733 79864
rect 11403 79736 11445 79745
rect 11403 79696 11404 79736
rect 11444 79696 11445 79736
rect 11403 79687 11445 79696
rect 11499 79064 11541 79073
rect 11692 79064 11732 79855
rect 11499 79024 11500 79064
rect 11540 79024 11541 79064
rect 11499 79015 11541 79024
rect 11596 79024 11692 79064
rect 11307 78056 11349 78065
rect 11307 78016 11308 78056
rect 11348 78016 11349 78056
rect 11307 78007 11349 78016
rect 11116 77596 11348 77636
rect 11308 77552 11348 77596
rect 11020 77512 11252 77552
rect 11212 77468 11252 77512
rect 11115 77132 11157 77141
rect 11115 77092 11116 77132
rect 11156 77092 11157 77132
rect 11115 77083 11157 77092
rect 11116 76712 11156 77083
rect 11116 76663 11156 76672
rect 10924 76504 11156 76544
rect 11019 75200 11061 75209
rect 11019 75160 11020 75200
rect 11060 75160 11061 75200
rect 11019 75151 11061 75160
rect 11020 75066 11060 75151
rect 10827 74696 10869 74705
rect 10827 74656 10828 74696
rect 10868 74656 10869 74696
rect 10827 74647 10869 74656
rect 10732 74453 10772 74538
rect 10828 74528 10868 74647
rect 10731 74444 10773 74453
rect 10731 74404 10732 74444
rect 10772 74404 10773 74444
rect 10731 74395 10773 74404
rect 10828 74276 10868 74488
rect 10732 74236 10868 74276
rect 11019 74276 11061 74285
rect 11019 74236 11020 74276
rect 11060 74236 11061 74276
rect 10545 73688 10585 73697
rect 10444 73668 10484 73677
rect 10347 73639 10389 73648
rect 10540 73648 10545 73688
rect 10540 73639 10585 73648
rect 10635 73688 10677 73697
rect 10635 73648 10636 73688
rect 10676 73648 10677 73688
rect 10635 73639 10677 73648
rect 10540 73361 10580 73639
rect 10539 73352 10581 73361
rect 10539 73312 10540 73352
rect 10580 73312 10581 73352
rect 10539 73303 10581 73312
rect 10443 73268 10485 73277
rect 10443 73228 10444 73268
rect 10484 73228 10485 73268
rect 10443 73219 10485 73228
rect 10251 73184 10293 73193
rect 10251 73144 10252 73184
rect 10292 73144 10293 73184
rect 10251 73135 10293 73144
rect 10444 73184 10484 73219
rect 10444 73133 10484 73144
rect 10156 72967 10196 72976
rect 10251 73016 10293 73025
rect 10251 72976 10252 73016
rect 10292 72976 10293 73016
rect 10251 72967 10293 72976
rect 10540 73016 10580 73025
rect 10252 72882 10292 72967
rect 10540 72857 10580 72976
rect 10539 72848 10581 72857
rect 10539 72808 10540 72848
rect 10580 72808 10581 72848
rect 10539 72799 10581 72808
rect 9771 72260 9813 72269
rect 9771 72220 9772 72260
rect 9812 72220 9813 72260
rect 9771 72211 9813 72220
rect 9675 72092 9717 72101
rect 9675 72052 9676 72092
rect 9716 72052 9717 72092
rect 9675 72043 9717 72052
rect 9676 71588 9716 71597
rect 9676 71429 9716 71548
rect 9675 71420 9717 71429
rect 9675 71380 9676 71420
rect 9716 71380 9717 71420
rect 9675 71371 9717 71380
rect 9772 69329 9812 72211
rect 10251 72176 10293 72185
rect 10251 72136 10252 72176
rect 10292 72136 10293 72176
rect 10251 72127 10293 72136
rect 10059 71672 10101 71681
rect 10059 71632 10060 71672
rect 10100 71632 10101 71672
rect 10059 71623 10101 71632
rect 9868 71504 9908 71513
rect 10060 71504 10100 71623
rect 9908 71464 10196 71504
rect 9868 71455 9908 71464
rect 9916 70673 9956 70682
rect 9956 70633 10004 70664
rect 9916 70624 10004 70633
rect 9964 70160 10004 70624
rect 10059 70580 10101 70589
rect 10059 70540 10060 70580
rect 10100 70540 10101 70580
rect 10059 70531 10101 70540
rect 10060 70446 10100 70531
rect 10156 70421 10196 71464
rect 10155 70412 10197 70421
rect 10155 70372 10156 70412
rect 10196 70372 10197 70412
rect 10155 70363 10197 70372
rect 10156 70160 10196 70169
rect 9964 70120 10156 70160
rect 10156 70111 10196 70120
rect 9964 69992 10004 70001
rect 9771 69320 9813 69329
rect 9771 69280 9772 69320
rect 9812 69280 9813 69320
rect 9771 69271 9813 69280
rect 9580 69103 9620 69112
rect 9964 68909 10004 69952
rect 9963 68900 10005 68909
rect 9963 68860 9964 68900
rect 10004 68860 10005 68900
rect 9963 68851 10005 68860
rect 9580 68648 9620 68657
rect 9620 68608 10004 68648
rect 9580 68599 9620 68608
rect 9772 68480 9812 68489
rect 9484 68440 9620 68480
rect 9388 68237 9428 68440
rect 9387 68228 9429 68237
rect 9387 68188 9388 68228
rect 9428 68188 9429 68228
rect 9387 68179 9429 68188
rect 9291 67976 9333 67985
rect 9291 67936 9292 67976
rect 9332 67936 9333 67976
rect 9291 67927 9333 67936
rect 9483 67808 9525 67817
rect 9483 67768 9484 67808
rect 9524 67768 9525 67808
rect 9483 67759 9525 67768
rect 9003 67724 9045 67733
rect 9003 67684 9004 67724
rect 9044 67684 9045 67724
rect 9003 67675 9045 67684
rect 9004 67640 9044 67675
rect 9484 67654 9524 67759
rect 9484 67605 9524 67614
rect 9004 67589 9044 67600
rect 9580 67565 9620 68440
rect 9676 68440 9772 68480
rect 9579 67556 9621 67565
rect 9579 67516 9580 67556
rect 9620 67516 9621 67556
rect 9579 67507 9621 67516
rect 9676 67556 9716 68440
rect 9772 68431 9812 68440
rect 9964 68480 10004 68608
rect 10155 68480 10197 68489
rect 10004 68440 10100 68480
rect 9964 68431 10004 68440
rect 9867 68396 9909 68405
rect 9867 68356 9868 68396
rect 9908 68356 9909 68396
rect 9867 68347 9909 68356
rect 9868 68262 9908 68347
rect 9771 68228 9813 68237
rect 9771 68188 9772 68228
rect 9812 68188 9813 68228
rect 9771 68179 9813 68188
rect 9676 67507 9716 67516
rect 9195 67472 9237 67481
rect 8908 67432 9140 67472
rect 8811 67136 8853 67145
rect 8811 67096 8812 67136
rect 8852 67096 8853 67136
rect 8811 67087 8853 67096
rect 8812 66968 8852 67087
rect 8908 66968 8948 66977
rect 8812 66928 8908 66968
rect 8908 66919 8948 66928
rect 8811 66800 8853 66809
rect 8811 66760 8812 66800
rect 8852 66760 8853 66800
rect 8811 66751 8853 66760
rect 8428 66256 8756 66296
rect 8428 64289 8468 66256
rect 8716 66128 8756 66137
rect 8523 64616 8565 64625
rect 8523 64576 8524 64616
rect 8564 64576 8565 64616
rect 8523 64567 8565 64576
rect 8427 64280 8469 64289
rect 8427 64240 8428 64280
rect 8468 64240 8469 64280
rect 8427 64231 8469 64240
rect 8331 63944 8373 63953
rect 8331 63904 8332 63944
rect 8372 63904 8373 63944
rect 8331 63895 8373 63904
rect 8428 63944 8468 63953
rect 8428 63869 8468 63904
rect 8524 63944 8564 64567
rect 8716 64280 8756 66088
rect 8524 63895 8564 63904
rect 8620 64240 8756 64280
rect 8812 64280 8852 66751
rect 9004 66305 9044 66390
rect 9003 66296 9045 66305
rect 9003 66256 9004 66296
rect 9044 66256 9045 66296
rect 9003 66247 9045 66256
rect 8908 66128 8948 66137
rect 8908 65708 8948 66088
rect 9004 66128 9044 66137
rect 9100 66128 9140 67432
rect 9195 67432 9196 67472
rect 9236 67432 9237 67472
rect 9195 67423 9237 67432
rect 9196 66968 9236 67423
rect 9675 67388 9717 67397
rect 9675 67348 9676 67388
rect 9716 67348 9717 67388
rect 9772 67388 9812 68179
rect 9963 68060 10005 68069
rect 9963 68020 9964 68060
rect 10004 68020 10005 68060
rect 9963 68011 10005 68020
rect 9867 67640 9909 67649
rect 9867 67600 9868 67640
rect 9908 67600 9909 67640
rect 9867 67591 9909 67600
rect 9964 67640 10004 68011
rect 9964 67591 10004 67600
rect 10060 67640 10100 68440
rect 10155 68440 10156 68480
rect 10196 68440 10197 68480
rect 10155 68431 10197 68440
rect 10156 68346 10196 68431
rect 10156 67649 10196 67734
rect 10060 67591 10100 67600
rect 10155 67640 10197 67649
rect 10155 67600 10156 67640
rect 10196 67600 10197 67640
rect 10155 67591 10197 67600
rect 9868 67506 9908 67591
rect 10252 67472 10292 72127
rect 10443 72008 10485 72017
rect 10443 71968 10444 72008
rect 10484 71968 10485 72008
rect 10443 71959 10485 71968
rect 10347 71588 10389 71597
rect 10347 71548 10348 71588
rect 10388 71548 10389 71588
rect 10347 71539 10389 71548
rect 10348 70496 10388 71539
rect 10444 70673 10484 71959
rect 10540 71345 10580 72799
rect 10636 72176 10676 72187
rect 10636 72101 10676 72136
rect 10635 72092 10677 72101
rect 10635 72052 10636 72092
rect 10676 72052 10677 72092
rect 10635 72043 10677 72052
rect 10732 71597 10772 74236
rect 11019 74227 11061 74236
rect 11020 74033 11060 74227
rect 11019 74024 11061 74033
rect 11019 73984 11020 74024
rect 11060 73984 11061 74024
rect 11019 73975 11061 73984
rect 10827 73688 10869 73697
rect 10827 73648 10828 73688
rect 10868 73648 10869 73688
rect 10827 73639 10869 73648
rect 10828 72185 10868 73639
rect 11116 73100 11156 76504
rect 11212 75461 11252 77428
rect 11308 76889 11348 77512
rect 11307 76880 11349 76889
rect 11307 76840 11308 76880
rect 11348 76840 11349 76880
rect 11307 76831 11349 76840
rect 11404 76040 11444 76049
rect 11320 75965 11360 75984
rect 11307 75956 11360 75965
rect 11404 75956 11444 76000
rect 11307 75916 11308 75956
rect 11348 75916 11444 75956
rect 11307 75907 11349 75916
rect 11500 75872 11540 79015
rect 11596 78224 11636 79024
rect 11692 79015 11732 79024
rect 11636 78184 11828 78224
rect 11596 78175 11636 78184
rect 11788 77552 11828 78184
rect 11691 76712 11733 76721
rect 11691 76672 11692 76712
rect 11732 76672 11733 76712
rect 11691 76663 11733 76672
rect 11404 75832 11540 75872
rect 11404 75629 11444 75832
rect 11596 75788 11636 75797
rect 11500 75748 11596 75788
rect 11403 75620 11445 75629
rect 11403 75580 11404 75620
rect 11444 75580 11445 75620
rect 11403 75571 11445 75580
rect 11211 75452 11253 75461
rect 11211 75412 11212 75452
rect 11252 75412 11253 75452
rect 11211 75403 11253 75412
rect 11403 75452 11445 75461
rect 11403 75412 11404 75452
rect 11444 75412 11445 75452
rect 11403 75403 11445 75412
rect 11307 75284 11349 75293
rect 11307 75244 11308 75284
rect 11348 75244 11349 75284
rect 11307 75235 11349 75244
rect 11211 75032 11253 75041
rect 11211 74992 11212 75032
rect 11252 74992 11253 75032
rect 11211 74983 11253 74992
rect 11212 74898 11252 74983
rect 11308 74528 11348 75235
rect 11308 74479 11348 74488
rect 11404 75032 11444 75403
rect 11500 75200 11540 75748
rect 11596 75739 11636 75748
rect 11500 75151 11540 75160
rect 11596 75200 11636 75209
rect 11596 75032 11636 75160
rect 11404 74992 11636 75032
rect 11404 74453 11444 74992
rect 11692 74948 11732 76663
rect 11788 75293 11828 77512
rect 11787 75284 11829 75293
rect 11787 75244 11788 75284
rect 11828 75244 11829 75284
rect 11787 75235 11829 75244
rect 11787 75032 11829 75041
rect 11787 74992 11788 75032
rect 11828 74992 11829 75032
rect 11787 74983 11829 74992
rect 11500 74908 11732 74948
rect 11403 74444 11445 74453
rect 11403 74404 11404 74444
rect 11444 74404 11445 74444
rect 11403 74395 11445 74404
rect 11211 74108 11253 74117
rect 11211 74068 11212 74108
rect 11252 74068 11253 74108
rect 11211 74059 11253 74068
rect 11403 74108 11445 74117
rect 11403 74068 11404 74108
rect 11444 74068 11445 74108
rect 11403 74059 11445 74068
rect 10924 73060 11156 73100
rect 10827 72176 10869 72185
rect 10827 72136 10828 72176
rect 10868 72136 10869 72176
rect 10827 72127 10869 72136
rect 10827 72008 10869 72017
rect 10827 71968 10828 72008
rect 10868 71968 10869 72008
rect 10827 71959 10869 71968
rect 10828 71874 10868 71959
rect 10731 71588 10773 71597
rect 10731 71548 10732 71588
rect 10772 71548 10773 71588
rect 10731 71539 10773 71548
rect 10924 71420 10964 73060
rect 11212 72176 11252 74059
rect 11404 72437 11444 74059
rect 11403 72428 11445 72437
rect 11403 72388 11404 72428
rect 11444 72388 11445 72428
rect 11403 72379 11445 72388
rect 11115 72092 11157 72101
rect 11115 72052 11116 72092
rect 11156 72052 11157 72092
rect 11115 72043 11157 72052
rect 10732 71380 10964 71420
rect 11020 72008 11060 72017
rect 10539 71336 10581 71345
rect 10539 71296 10540 71336
rect 10580 71296 10581 71336
rect 10539 71287 10581 71296
rect 10635 71252 10677 71261
rect 10635 71212 10636 71252
rect 10676 71212 10677 71252
rect 10635 71203 10677 71212
rect 10439 70664 10484 70673
rect 10479 70624 10484 70664
rect 10540 70664 10580 70675
rect 10439 70615 10479 70624
rect 10540 70589 10580 70624
rect 10636 70664 10676 71203
rect 10636 70615 10676 70624
rect 10539 70580 10581 70589
rect 10539 70540 10540 70580
rect 10580 70540 10581 70580
rect 10539 70531 10581 70540
rect 10348 70456 10484 70496
rect 10347 69152 10389 69161
rect 10347 69112 10348 69152
rect 10388 69112 10389 69152
rect 10347 69103 10389 69112
rect 10348 67892 10388 69103
rect 10348 67843 10388 67852
rect 10347 67640 10389 67649
rect 10347 67600 10348 67640
rect 10388 67600 10389 67640
rect 10347 67591 10389 67600
rect 10348 67506 10388 67591
rect 10156 67432 10292 67472
rect 9772 67348 9908 67388
rect 9675 67339 9717 67348
rect 9291 67052 9333 67061
rect 9291 67012 9292 67052
rect 9332 67012 9333 67052
rect 9291 67003 9333 67012
rect 9196 66893 9236 66928
rect 9292 66918 9332 67003
rect 9483 66968 9525 66977
rect 9483 66928 9484 66968
rect 9524 66928 9525 66968
rect 9483 66919 9525 66928
rect 9195 66884 9237 66893
rect 9195 66844 9196 66884
rect 9236 66844 9237 66884
rect 9195 66835 9237 66844
rect 9196 66804 9236 66835
rect 9291 66800 9333 66809
rect 9291 66760 9292 66800
rect 9332 66760 9333 66800
rect 9291 66751 9333 66760
rect 9196 66128 9236 66137
rect 9100 66088 9196 66128
rect 9004 65792 9044 66088
rect 9196 66079 9236 66088
rect 9292 66128 9332 66751
rect 9484 66548 9524 66919
rect 9579 66800 9621 66809
rect 9579 66760 9580 66800
rect 9620 66760 9621 66800
rect 9579 66751 9621 66760
rect 9580 66666 9620 66751
rect 9484 66508 9620 66548
rect 9483 66296 9525 66305
rect 9483 66256 9484 66296
rect 9524 66256 9525 66296
rect 9483 66247 9525 66256
rect 9292 66079 9332 66088
rect 9004 65752 9332 65792
rect 8908 65668 9236 65708
rect 8908 64709 8948 65668
rect 9196 65624 9236 65668
rect 9196 65575 9236 65584
rect 9099 65540 9141 65549
rect 9099 65500 9100 65540
rect 9140 65500 9141 65540
rect 9099 65491 9141 65500
rect 9004 65414 9044 65423
rect 9004 65372 9044 65374
rect 9100 65372 9140 65491
rect 9004 65332 9140 65372
rect 9003 65036 9045 65045
rect 9003 64996 9004 65036
rect 9044 64996 9045 65036
rect 9003 64987 9045 64996
rect 8907 64700 8949 64709
rect 8907 64660 8908 64700
rect 8948 64660 8949 64700
rect 8907 64651 8949 64660
rect 8812 64240 8948 64280
rect 8427 63860 8469 63869
rect 8427 63820 8428 63860
rect 8468 63820 8469 63860
rect 8427 63811 8469 63820
rect 8428 63029 8468 63811
rect 8523 63608 8565 63617
rect 8523 63568 8524 63608
rect 8564 63568 8565 63608
rect 8523 63559 8565 63568
rect 8427 63020 8469 63029
rect 8427 62980 8428 63020
rect 8468 62980 8469 63020
rect 8427 62971 8469 62980
rect 8236 62432 8276 62441
rect 8236 62189 8276 62392
rect 8332 62432 8372 62441
rect 8372 62392 8468 62432
rect 8332 62383 8372 62392
rect 8235 62180 8277 62189
rect 8235 62140 8236 62180
rect 8276 62140 8277 62180
rect 8235 62131 8277 62140
rect 8139 61088 8181 61097
rect 8139 61048 8140 61088
rect 8180 61048 8181 61088
rect 8139 61039 8181 61048
rect 8139 60920 8181 60929
rect 8139 60880 8140 60920
rect 8180 60880 8181 60920
rect 8139 60871 8181 60880
rect 8140 60786 8180 60871
rect 8332 60668 8372 60677
rect 8236 60628 8332 60668
rect 8236 60164 8276 60628
rect 8332 60619 8372 60628
rect 8331 60500 8373 60509
rect 8331 60460 8332 60500
rect 8372 60460 8373 60500
rect 8331 60451 8373 60460
rect 8428 60500 8468 62392
rect 8524 60929 8564 63559
rect 8620 62852 8660 64240
rect 8715 63944 8757 63953
rect 8715 63904 8716 63944
rect 8756 63904 8757 63944
rect 8715 63895 8757 63904
rect 8716 63810 8756 63895
rect 8811 63020 8853 63029
rect 8811 62980 8812 63020
rect 8852 62980 8853 63020
rect 8811 62971 8853 62980
rect 8715 62852 8757 62861
rect 8620 62812 8716 62852
rect 8756 62812 8757 62852
rect 8715 62803 8757 62812
rect 8619 62516 8661 62525
rect 8619 62476 8620 62516
rect 8660 62476 8661 62516
rect 8619 62467 8661 62476
rect 8523 60920 8565 60929
rect 8523 60880 8524 60920
rect 8564 60880 8565 60920
rect 8523 60871 8565 60880
rect 8524 60509 8564 60528
rect 8523 60500 8565 60509
rect 8428 60460 8524 60500
rect 8564 60460 8565 60500
rect 8188 60124 8276 60164
rect 8188 60122 8228 60124
rect 8188 60073 8228 60082
rect 8332 59996 8372 60451
rect 8332 59947 8372 59956
rect 8044 59620 8276 59660
rect 8044 59492 8084 59501
rect 8084 59452 8180 59492
rect 8044 59443 8084 59452
rect 7852 59354 7892 59363
rect 7756 59200 8084 59240
rect 7564 58948 7700 58988
rect 7467 58939 7509 58948
rect 7564 58568 7604 58579
rect 7564 58493 7604 58528
rect 7371 58484 7413 58493
rect 7371 58444 7372 58484
rect 7412 58444 7413 58484
rect 7371 58435 7413 58444
rect 7563 58484 7605 58493
rect 7563 58444 7564 58484
rect 7604 58444 7605 58484
rect 7563 58435 7605 58444
rect 7467 58232 7509 58241
rect 7467 58192 7468 58232
rect 7508 58192 7509 58232
rect 7660 58232 7700 58948
rect 8044 58568 8084 59200
rect 7756 58400 7796 58409
rect 7796 58360 7988 58400
rect 7756 58351 7796 58360
rect 7660 58192 7892 58232
rect 7467 58183 7509 58192
rect 7468 57896 7508 58183
rect 7275 57056 7317 57065
rect 7275 57016 7276 57056
rect 7316 57016 7317 57056
rect 7275 57007 7317 57016
rect 7276 56813 7316 57007
rect 7275 56804 7317 56813
rect 7275 56764 7276 56804
rect 7316 56764 7317 56804
rect 7275 56755 7317 56764
rect 7276 56384 7316 56393
rect 7468 56384 7508 57856
rect 7660 57644 7700 57653
rect 7700 57604 7796 57644
rect 7660 57595 7700 57604
rect 7659 57476 7701 57485
rect 7659 57436 7660 57476
rect 7700 57436 7701 57476
rect 7659 57427 7701 57436
rect 7660 56813 7700 57427
rect 7756 57070 7796 57604
rect 7756 57021 7796 57030
rect 7659 56804 7701 56813
rect 7659 56764 7660 56804
rect 7700 56764 7701 56804
rect 7659 56755 7701 56764
rect 7316 56344 7508 56384
rect 7276 56335 7316 56344
rect 7180 56176 7316 56216
rect 7084 56092 7220 56132
rect 7083 55544 7125 55553
rect 6988 55504 7084 55544
rect 7124 55504 7125 55544
rect 7083 55495 7125 55504
rect 6795 54956 6837 54965
rect 6795 54916 6796 54956
rect 6836 54916 6837 54956
rect 6795 54907 6837 54916
rect 7084 54872 7124 55495
rect 7084 54823 7124 54832
rect 6508 54664 7028 54704
rect 6891 54536 6933 54545
rect 6891 54496 6892 54536
rect 6932 54496 6933 54536
rect 6891 54487 6933 54496
rect 6604 52529 6644 52614
rect 6603 52520 6645 52529
rect 6603 52480 6604 52520
rect 6644 52480 6645 52520
rect 6603 52471 6645 52480
rect 6603 52352 6645 52361
rect 6603 52312 6604 52352
rect 6644 52312 6645 52352
rect 6603 52303 6645 52312
rect 6507 52184 6549 52193
rect 6507 52144 6508 52184
rect 6548 52144 6549 52184
rect 6507 52135 6549 52144
rect 6508 51848 6548 52135
rect 6508 51799 6548 51808
rect 6604 51848 6644 52303
rect 6411 51008 6453 51017
rect 6508 51008 6548 51017
rect 6411 50968 6412 51008
rect 6452 50968 6508 51008
rect 6411 50959 6453 50968
rect 6508 50959 6548 50968
rect 6412 50874 6452 50959
rect 6507 48824 6549 48833
rect 6507 48784 6508 48824
rect 6548 48784 6549 48824
rect 6507 48775 6549 48784
rect 6412 48740 6452 48749
rect 6412 48572 6452 48700
rect 6508 48690 6548 48775
rect 6412 48532 6548 48572
rect 6315 48404 6357 48413
rect 6315 48364 6316 48404
rect 6356 48364 6357 48404
rect 6315 48355 6357 48364
rect 6315 48236 6357 48245
rect 6315 48196 6316 48236
rect 6356 48196 6357 48236
rect 6315 48187 6357 48196
rect 6316 47909 6356 48187
rect 6411 47984 6453 47993
rect 6411 47944 6412 47984
rect 6452 47944 6453 47984
rect 6411 47935 6453 47944
rect 6315 47900 6357 47909
rect 6315 47860 6316 47900
rect 6356 47860 6357 47900
rect 6315 47851 6357 47860
rect 6220 47816 6260 47825
rect 6220 47312 6260 47776
rect 6220 47263 6260 47272
rect 6316 47312 6356 47851
rect 6412 47850 6452 47935
rect 6508 47312 6548 48532
rect 6604 48245 6644 51808
rect 6699 49664 6741 49673
rect 6699 49624 6700 49664
rect 6740 49624 6741 49664
rect 6699 49615 6741 49624
rect 6700 49496 6740 49615
rect 6700 49447 6740 49456
rect 6795 48824 6837 48833
rect 6795 48784 6796 48824
rect 6836 48784 6837 48824
rect 6795 48775 6837 48784
rect 6603 48236 6645 48245
rect 6603 48196 6604 48236
rect 6644 48196 6645 48236
rect 6603 48187 6645 48196
rect 6700 47312 6740 47321
rect 6508 47272 6700 47312
rect 6316 47263 6356 47272
rect 6604 47153 6644 47272
rect 6700 47263 6740 47272
rect 6796 47312 6836 48775
rect 6796 47263 6836 47272
rect 6603 47144 6645 47153
rect 6603 47104 6604 47144
rect 6644 47104 6645 47144
rect 6603 47095 6645 47104
rect 6411 46472 6453 46481
rect 6411 46432 6412 46472
rect 6452 46432 6453 46472
rect 6411 46423 6453 46432
rect 6412 46338 6452 46423
rect 6028 46012 6164 46052
rect 5348 44962 5588 45002
rect 5644 45800 5684 45809
rect 6028 45800 6068 46012
rect 6123 45884 6165 45893
rect 6123 45844 6124 45884
rect 6164 45844 6165 45884
rect 6123 45835 6165 45844
rect 5684 45760 6068 45800
rect 5644 44969 5684 45760
rect 5836 45548 5876 45557
rect 5740 45508 5836 45548
rect 5308 44953 5348 44962
rect 5643 44960 5685 44969
rect 4780 44911 4820 44920
rect 5643 44920 5644 44960
rect 5684 44920 5685 44960
rect 5643 44911 5685 44920
rect 5451 44876 5493 44885
rect 5451 44836 5452 44876
rect 5492 44836 5493 44876
rect 5451 44827 5493 44836
rect 5452 44742 5492 44827
rect 4928 44624 5296 44633
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 4928 44575 5296 44584
rect 5740 44540 5780 45508
rect 5836 45499 5876 45508
rect 5835 44960 5877 44969
rect 5835 44920 5836 44960
rect 5876 44920 5877 44960
rect 5835 44911 5877 44920
rect 6124 44960 6164 45835
rect 6411 45716 6453 45725
rect 6411 45676 6412 45716
rect 6452 45676 6453 45716
rect 6411 45667 6453 45676
rect 6124 44911 6164 44920
rect 5452 44500 5780 44540
rect 4875 44456 4917 44465
rect 4875 44416 4876 44456
rect 4916 44416 4917 44456
rect 4875 44407 4917 44416
rect 4436 44248 4532 44288
rect 4876 44288 4916 44407
rect 5452 44288 5492 44500
rect 5547 44372 5589 44381
rect 5547 44332 5548 44372
rect 5588 44332 5589 44372
rect 5547 44323 5589 44332
rect 4396 44239 4436 44248
rect 4876 44239 4916 44248
rect 5404 44278 5492 44288
rect 3820 44154 3860 44239
rect 5444 44248 5492 44278
rect 5548 44238 5588 44323
rect 5404 44229 5444 44238
rect 3476 44080 3764 44120
rect 3436 44071 3476 44080
rect 1612 44036 1652 44045
rect 1612 43793 1652 43996
rect 3688 43868 4056 43877
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 3688 43819 4056 43828
rect 1611 43784 1653 43793
rect 1611 43744 1612 43784
rect 1652 43744 1653 43784
rect 1611 43735 1653 43744
rect 2188 43448 2228 43459
rect 2188 43373 2228 43408
rect 2475 43448 2517 43457
rect 2475 43408 2476 43448
rect 2516 43408 2517 43448
rect 2475 43399 2517 43408
rect 3435 43448 3477 43457
rect 3435 43408 3436 43448
rect 3476 43408 3477 43448
rect 3435 43399 3477 43408
rect 3820 43448 3860 43457
rect 2187 43364 2229 43373
rect 2187 43324 2188 43364
rect 2228 43324 2229 43364
rect 2187 43315 2229 43324
rect 2091 43196 2133 43205
rect 2091 43156 2092 43196
rect 2132 43156 2133 43196
rect 2091 43147 2133 43156
rect 1803 42356 1845 42365
rect 1803 42316 1804 42356
rect 1844 42316 1845 42356
rect 1803 42307 1845 42316
rect 1611 41264 1653 41273
rect 1611 41224 1612 41264
rect 1652 41224 1653 41264
rect 1611 41215 1653 41224
rect 1612 34385 1652 41215
rect 1707 40088 1749 40097
rect 1707 40048 1708 40088
rect 1748 40048 1749 40088
rect 1707 40039 1749 40048
rect 1611 34376 1653 34385
rect 1611 34336 1612 34376
rect 1652 34336 1653 34376
rect 1611 34327 1653 34336
rect 1708 32957 1748 40039
rect 1804 38333 1844 42307
rect 1995 41180 2037 41189
rect 1995 41140 1996 41180
rect 2036 41140 2037 41180
rect 1995 41131 2037 41140
rect 1899 41096 1941 41105
rect 1899 41056 1900 41096
rect 1940 41056 1941 41096
rect 1899 41047 1941 41056
rect 1803 38324 1845 38333
rect 1803 38284 1804 38324
rect 1844 38284 1845 38324
rect 1803 38275 1845 38284
rect 1900 38249 1940 41047
rect 1996 40256 2036 41131
rect 1996 40207 2036 40216
rect 2092 40013 2132 43147
rect 2476 41936 2516 43399
rect 3436 43314 3476 43399
rect 3628 43280 3668 43289
rect 3531 43028 3573 43037
rect 3531 42988 3532 43028
rect 3572 42988 3573 43028
rect 3531 42979 3573 42988
rect 3148 42869 3188 42885
rect 3147 42860 3189 42869
rect 3147 42820 3148 42860
rect 3188 42820 3189 42860
rect 3147 42811 3189 42820
rect 2763 42776 2805 42785
rect 2763 42736 2764 42776
rect 2804 42736 2805 42776
rect 2763 42727 2805 42736
rect 2956 42776 2996 42785
rect 2764 42642 2804 42727
rect 2764 42524 2804 42533
rect 2804 42484 2900 42524
rect 2764 42475 2804 42484
rect 2763 42020 2805 42029
rect 2763 41980 2764 42020
rect 2804 41980 2805 42020
rect 2763 41971 2805 41980
rect 2283 41432 2325 41441
rect 2283 41392 2284 41432
rect 2324 41392 2325 41432
rect 2283 41383 2325 41392
rect 2284 40433 2324 41383
rect 2476 41264 2516 41896
rect 2668 41768 2708 41777
rect 2571 41348 2613 41357
rect 2571 41308 2572 41348
rect 2612 41308 2613 41348
rect 2571 41299 2613 41308
rect 2380 41224 2476 41264
rect 2188 40424 2228 40433
rect 2091 40004 2133 40013
rect 2091 39964 2092 40004
rect 2132 39964 2133 40004
rect 2091 39955 2133 39964
rect 2092 38996 2132 39955
rect 2188 39173 2228 40384
rect 2283 40424 2325 40433
rect 2283 40384 2284 40424
rect 2324 40384 2325 40424
rect 2283 40375 2325 40384
rect 2284 40290 2324 40375
rect 2380 39584 2420 41224
rect 2476 41215 2516 41224
rect 2572 41096 2612 41299
rect 2668 41273 2708 41728
rect 2667 41264 2709 41273
rect 2667 41224 2668 41264
rect 2708 41224 2709 41264
rect 2667 41215 2709 41224
rect 2668 41096 2708 41105
rect 2572 41056 2668 41096
rect 2668 41047 2708 41056
rect 2571 40424 2613 40433
rect 2571 40384 2572 40424
rect 2612 40384 2613 40424
rect 2571 40375 2613 40384
rect 2668 40424 2708 40433
rect 2572 40290 2612 40375
rect 2668 40265 2708 40384
rect 2667 40256 2709 40265
rect 2667 40216 2668 40256
rect 2708 40216 2709 40256
rect 2667 40207 2709 40216
rect 2764 40004 2804 41971
rect 2860 41936 2900 42484
rect 2956 42029 2996 42736
rect 3052 42776 3092 42785
rect 3052 42533 3092 42736
rect 3148 42761 3188 42811
rect 3244 42776 3284 42785
rect 3148 42736 3244 42761
rect 3148 42721 3284 42736
rect 3435 42776 3477 42785
rect 3435 42736 3436 42776
rect 3476 42736 3477 42776
rect 3435 42727 3477 42736
rect 3532 42776 3572 42979
rect 3628 42785 3668 43240
rect 3723 43112 3765 43121
rect 3723 43072 3724 43112
rect 3764 43072 3765 43112
rect 3723 43063 3765 43072
rect 3724 42953 3764 43063
rect 3723 42944 3765 42953
rect 3723 42904 3724 42944
rect 3764 42904 3765 42944
rect 3820 42944 3860 43408
rect 3916 43448 3956 43457
rect 3916 43205 3956 43408
rect 4108 43448 4148 43457
rect 4148 43408 4820 43448
rect 4108 43399 4148 43408
rect 4011 43280 4053 43289
rect 4011 43240 4012 43280
rect 4052 43240 4053 43280
rect 4011 43231 4053 43240
rect 3915 43196 3957 43205
rect 3915 43156 3916 43196
rect 3956 43156 3957 43196
rect 3915 43147 3957 43156
rect 4012 43146 4052 43231
rect 3820 42904 4628 42944
rect 3723 42895 3765 42904
rect 4204 42797 4244 42806
rect 3532 42727 3572 42736
rect 3627 42776 3669 42785
rect 3627 42736 3628 42776
rect 3668 42736 3669 42776
rect 3627 42727 3669 42736
rect 3724 42776 3764 42785
rect 3051 42524 3093 42533
rect 3051 42484 3052 42524
rect 3092 42484 3093 42524
rect 3051 42475 3093 42484
rect 2955 42020 2997 42029
rect 2955 41980 2956 42020
rect 2996 41980 2997 42020
rect 2955 41971 2997 41980
rect 2860 41887 2900 41896
rect 3051 41936 3093 41945
rect 3051 41896 3052 41936
rect 3092 41896 3093 41936
rect 3051 41887 3093 41896
rect 3148 41936 3188 42721
rect 3340 42608 3380 42617
rect 3243 42524 3285 42533
rect 3243 42484 3244 42524
rect 3284 42484 3285 42524
rect 3243 42475 3285 42484
rect 2955 41852 2997 41861
rect 2955 41812 2956 41852
rect 2996 41812 2997 41852
rect 2955 41803 2997 41812
rect 2956 41718 2996 41803
rect 3052 41802 3092 41887
rect 3148 41600 3188 41896
rect 2956 41560 3188 41600
rect 2956 41432 2996 41560
rect 2956 41383 2996 41392
rect 2859 41264 2901 41273
rect 2859 41224 2860 41264
rect 2900 41224 2901 41264
rect 2859 41215 2901 41224
rect 3148 41264 3188 41273
rect 3244 41264 3284 42475
rect 3340 41936 3380 42568
rect 3340 41887 3380 41896
rect 3436 41357 3476 42727
rect 3724 42524 3764 42736
rect 3532 42484 3764 42524
rect 3820 42776 3860 42785
rect 3820 42524 3860 42736
rect 3915 42776 3957 42785
rect 3915 42736 3916 42776
rect 3956 42736 3957 42776
rect 3915 42727 3957 42736
rect 4012 42776 4052 42785
rect 3916 42642 3956 42727
rect 4012 42608 4052 42736
rect 4107 42776 4149 42785
rect 4107 42736 4108 42776
rect 4148 42757 4204 42776
rect 4148 42736 4244 42757
rect 4300 42797 4340 42806
rect 4107 42727 4149 42736
rect 4203 42608 4245 42617
rect 4012 42568 4204 42608
rect 4244 42568 4245 42608
rect 4203 42559 4245 42568
rect 3820 42484 4148 42524
rect 3532 42104 3572 42484
rect 3688 42356 4056 42365
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 3688 42307 4056 42316
rect 3532 42055 3572 42064
rect 4108 42104 4148 42484
rect 4108 42055 4148 42064
rect 3532 41936 3572 41945
rect 3435 41348 3477 41357
rect 3435 41308 3436 41348
rect 3476 41308 3477 41348
rect 3435 41299 3477 41308
rect 3339 41264 3381 41273
rect 3244 41224 3340 41264
rect 3380 41224 3381 41264
rect 2860 40601 2900 41215
rect 3148 41021 3188 41224
rect 3339 41215 3381 41224
rect 3436 41264 3476 41299
rect 3340 41130 3380 41215
rect 3436 41213 3476 41224
rect 3436 41096 3476 41105
rect 3532 41096 3572 41896
rect 3627 41936 3669 41945
rect 3627 41896 3628 41936
rect 3668 41896 3669 41936
rect 3627 41887 3669 41896
rect 3820 41936 3860 41945
rect 3628 41802 3668 41887
rect 3820 41441 3860 41896
rect 4012 41936 4052 41947
rect 4012 41861 4052 41896
rect 4108 41936 4148 41945
rect 4148 41896 4244 41936
rect 4108 41887 4148 41896
rect 4011 41852 4053 41861
rect 4011 41812 4012 41852
rect 4052 41812 4053 41852
rect 4011 41803 4053 41812
rect 4011 41516 4053 41525
rect 4011 41476 4012 41516
rect 4052 41476 4053 41516
rect 4204 41516 4244 41896
rect 4300 41600 4340 42757
rect 4396 42776 4436 42785
rect 4396 42617 4436 42736
rect 4491 42776 4533 42785
rect 4491 42736 4492 42776
rect 4532 42736 4533 42776
rect 4491 42727 4533 42736
rect 4492 42642 4532 42727
rect 4395 42608 4437 42617
rect 4395 42568 4396 42608
rect 4436 42568 4437 42608
rect 4588 42608 4628 42904
rect 4683 42860 4725 42869
rect 4683 42820 4684 42860
rect 4724 42820 4725 42860
rect 4683 42811 4725 42820
rect 4780 42860 4820 43408
rect 4928 43112 5296 43121
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 4928 43063 5296 43072
rect 5355 43112 5397 43121
rect 5355 43072 5356 43112
rect 5396 43072 5397 43112
rect 5355 43063 5397 43072
rect 4684 42776 4724 42811
rect 4684 42725 4724 42736
rect 4588 42568 4724 42608
rect 4395 42559 4437 42568
rect 4395 42188 4437 42197
rect 4395 42148 4396 42188
rect 4436 42148 4437 42188
rect 4395 42139 4437 42148
rect 4396 42104 4436 42139
rect 4396 42053 4436 42064
rect 4587 41936 4629 41945
rect 4587 41896 4588 41936
rect 4628 41896 4629 41936
rect 4587 41887 4629 41896
rect 4684 41936 4724 42568
rect 4588 41802 4628 41887
rect 4300 41560 4628 41600
rect 4204 41476 4436 41516
rect 4011 41467 4053 41476
rect 3819 41432 3861 41441
rect 3819 41392 3820 41432
rect 3860 41392 3861 41432
rect 3819 41383 3861 41392
rect 3476 41056 3572 41096
rect 3628 41264 3668 41273
rect 3436 41047 3476 41056
rect 2956 41012 2996 41021
rect 2956 40685 2996 40972
rect 3147 41012 3189 41021
rect 3628 41012 3668 41224
rect 3723 41180 3765 41189
rect 3723 41140 3724 41180
rect 3764 41140 3765 41180
rect 3723 41131 3765 41140
rect 3724 41046 3764 41131
rect 3820 41105 3860 41190
rect 3916 41189 3956 41274
rect 4012 41264 4052 41467
rect 4396 41432 4436 41476
rect 4204 41357 4244 41388
rect 4396 41383 4436 41392
rect 4203 41348 4245 41357
rect 4203 41308 4204 41348
rect 4244 41308 4245 41348
rect 4203 41299 4245 41308
rect 4012 41215 4052 41224
rect 4204 41264 4244 41299
rect 3915 41180 3957 41189
rect 3915 41140 3916 41180
rect 3956 41140 3957 41180
rect 3915 41131 3957 41140
rect 3819 41096 3861 41105
rect 3819 41056 3820 41096
rect 3860 41056 3861 41096
rect 3819 41047 3861 41056
rect 4107 41096 4149 41105
rect 4107 41056 4108 41096
rect 4148 41056 4149 41096
rect 4107 41047 4149 41056
rect 3147 40972 3148 41012
rect 3188 40972 3189 41012
rect 3147 40963 3189 40972
rect 3532 40972 3668 41012
rect 2955 40676 2997 40685
rect 2955 40636 2956 40676
rect 2996 40636 2997 40676
rect 2955 40627 2997 40636
rect 2859 40592 2901 40601
rect 2859 40552 2860 40592
rect 2900 40552 2901 40592
rect 3148 40592 3188 40963
rect 3532 40676 3572 40972
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 4108 40676 4148 41047
rect 4204 41012 4244 41224
rect 4307 41264 4347 41272
rect 4395 41264 4437 41273
rect 4307 41263 4396 41264
rect 4347 41224 4396 41263
rect 4436 41224 4437 41264
rect 4307 41214 4347 41223
rect 4395 41215 4437 41224
rect 4492 41264 4532 41273
rect 4204 40972 4436 41012
rect 3532 40636 3860 40676
rect 4108 40636 4244 40676
rect 3148 40552 3476 40592
rect 2859 40543 2901 40552
rect 3052 40508 3092 40517
rect 2956 40468 3052 40508
rect 2859 40424 2901 40433
rect 2859 40384 2860 40424
rect 2900 40384 2901 40424
rect 2859 40375 2901 40384
rect 2572 39964 2804 40004
rect 2475 39920 2517 39929
rect 2475 39880 2476 39920
rect 2516 39880 2517 39920
rect 2475 39871 2517 39880
rect 2572 39920 2612 39964
rect 2860 39920 2900 40375
rect 2956 40181 2996 40468
rect 3052 40459 3092 40468
rect 3148 40424 3188 40433
rect 2955 40172 2997 40181
rect 2955 40132 2956 40172
rect 2996 40132 2997 40172
rect 2955 40123 2997 40132
rect 3148 40097 3188 40384
rect 3147 40088 3189 40097
rect 3147 40048 3148 40088
rect 3188 40048 3189 40088
rect 3147 40039 3189 40048
rect 2572 39871 2612 39880
rect 2668 39880 2900 39920
rect 3339 39920 3381 39929
rect 3339 39880 3340 39920
rect 3380 39880 3381 39920
rect 2476 39752 2516 39871
rect 2668 39752 2708 39880
rect 3339 39871 3381 39880
rect 2476 39703 2516 39712
rect 2572 39712 2708 39752
rect 2764 39752 2804 39761
rect 2804 39712 2900 39752
rect 2475 39584 2517 39593
rect 2380 39544 2476 39584
rect 2516 39544 2517 39584
rect 2475 39535 2517 39544
rect 2379 39416 2421 39425
rect 2379 39376 2380 39416
rect 2420 39376 2421 39416
rect 2379 39367 2421 39376
rect 2187 39164 2229 39173
rect 2187 39124 2188 39164
rect 2228 39124 2229 39164
rect 2187 39115 2229 39124
rect 2092 38956 2228 38996
rect 1899 38240 1941 38249
rect 1899 38200 1900 38240
rect 1940 38200 1941 38240
rect 1899 38191 1941 38200
rect 1803 36896 1845 36905
rect 1803 36856 1804 36896
rect 1844 36856 1845 36896
rect 1803 36847 1845 36856
rect 1804 34973 1844 36847
rect 1803 34964 1845 34973
rect 1803 34924 1804 34964
rect 1844 34924 1845 34964
rect 1803 34915 1845 34924
rect 1804 34376 1844 34385
rect 1804 34049 1844 34336
rect 1803 34040 1845 34049
rect 1803 34000 1804 34040
rect 1844 34000 1845 34040
rect 1803 33991 1845 34000
rect 1707 32948 1749 32957
rect 1707 32908 1708 32948
rect 1748 32908 1749 32948
rect 1707 32899 1749 32908
rect 1611 31436 1653 31445
rect 1611 31396 1612 31436
rect 1652 31396 1653 31436
rect 1611 31387 1653 31396
rect 1612 31352 1652 31387
rect 1612 31301 1652 31312
rect 1707 31184 1749 31193
rect 1707 31144 1708 31184
rect 1748 31144 1749 31184
rect 1707 31135 1749 31144
rect 1708 29336 1748 31135
rect 1612 29296 1748 29336
rect 1612 24632 1652 29296
rect 1708 29168 1748 29177
rect 1708 29000 1748 29128
rect 1900 29000 1940 38191
rect 1995 35216 2037 35225
rect 1995 35176 1996 35216
rect 2036 35176 2037 35216
rect 1995 35167 2037 35176
rect 2092 35216 2132 35225
rect 1996 35082 2036 35167
rect 1995 34880 2037 34889
rect 1995 34840 1996 34880
rect 2036 34840 2037 34880
rect 1995 34831 2037 34840
rect 1996 33713 2036 34831
rect 1995 33704 2037 33713
rect 1995 33664 1996 33704
rect 2036 33664 2037 33704
rect 1995 33655 2037 33664
rect 2092 32201 2132 35176
rect 2188 33872 2228 38956
rect 2380 37400 2420 39367
rect 2476 38240 2516 39535
rect 2572 38408 2612 39712
rect 2764 39703 2804 39712
rect 2763 38912 2805 38921
rect 2763 38872 2764 38912
rect 2804 38872 2805 38912
rect 2763 38863 2805 38872
rect 2667 38828 2709 38837
rect 2667 38788 2668 38828
rect 2708 38788 2709 38828
rect 2667 38779 2709 38788
rect 2668 38744 2708 38779
rect 2668 38693 2708 38704
rect 2668 38408 2708 38417
rect 2572 38368 2668 38408
rect 2668 38359 2708 38368
rect 2476 38191 2516 38200
rect 2668 37652 2708 37661
rect 2764 37652 2804 38863
rect 2860 37661 2900 39712
rect 3147 38996 3189 39005
rect 3147 38956 3148 38996
rect 3188 38956 3189 38996
rect 3147 38947 3189 38956
rect 3051 38912 3093 38921
rect 3051 38872 3052 38912
rect 3092 38872 3093 38912
rect 3051 38863 3093 38872
rect 3148 38912 3188 38947
rect 3052 38778 3092 38863
rect 3052 38408 3092 38417
rect 3148 38408 3188 38872
rect 3092 38368 3188 38408
rect 3052 38359 3092 38368
rect 2955 38072 2997 38081
rect 2955 38032 2956 38072
rect 2996 38032 2997 38072
rect 2955 38023 2997 38032
rect 2956 37938 2996 38023
rect 2708 37612 2804 37652
rect 2859 37652 2901 37661
rect 2859 37612 2860 37652
rect 2900 37612 2901 37652
rect 2668 37603 2708 37612
rect 2859 37603 2901 37612
rect 3147 37652 3189 37661
rect 3147 37612 3148 37652
rect 3188 37612 3189 37652
rect 3147 37603 3189 37612
rect 2571 37568 2613 37577
rect 2571 37528 2572 37568
rect 2612 37528 2613 37568
rect 2571 37519 2613 37528
rect 2476 37400 2516 37409
rect 2380 37360 2476 37400
rect 2476 36728 2516 37360
rect 2476 35888 2516 36688
rect 2476 35839 2516 35848
rect 2572 35216 2612 37519
rect 3004 37409 3044 37418
rect 2668 37369 3004 37400
rect 2668 37360 3044 37369
rect 2668 36896 2708 37360
rect 2859 37232 2901 37241
rect 2859 37192 2860 37232
rect 2900 37192 2901 37232
rect 2859 37183 2901 37192
rect 2860 36980 2900 37183
rect 3148 37073 3188 37603
rect 3340 37577 3380 39871
rect 3339 37568 3381 37577
rect 3339 37528 3340 37568
rect 3380 37528 3381 37568
rect 3339 37519 3381 37528
rect 3147 37064 3189 37073
rect 3147 37024 3148 37064
rect 3188 37024 3189 37064
rect 3147 37015 3189 37024
rect 2860 36940 3092 36980
rect 2668 36847 2708 36856
rect 2860 36728 2900 36737
rect 2667 36560 2709 36569
rect 2667 36520 2668 36560
rect 2708 36520 2709 36560
rect 2667 36511 2709 36520
rect 2668 36140 2708 36511
rect 2668 36091 2708 36100
rect 2476 35132 2516 35141
rect 2476 33965 2516 35092
rect 2475 33956 2517 33965
rect 2475 33916 2476 33956
rect 2516 33916 2517 33956
rect 2475 33907 2517 33916
rect 2188 33832 2420 33872
rect 1708 28960 1940 29000
rect 1996 32192 2036 32201
rect 1708 25397 1748 28960
rect 1803 26816 1845 26825
rect 1803 26776 1804 26816
rect 1844 26776 1845 26816
rect 1803 26767 1845 26776
rect 1707 25388 1749 25397
rect 1707 25348 1708 25388
rect 1748 25348 1749 25388
rect 1707 25339 1749 25348
rect 1612 22457 1652 24592
rect 1707 22532 1749 22541
rect 1707 22492 1708 22532
rect 1748 22492 1749 22532
rect 1707 22483 1749 22492
rect 1611 22448 1653 22457
rect 1611 22408 1612 22448
rect 1652 22408 1653 22448
rect 1611 22399 1653 22408
rect 1612 17921 1652 22399
rect 1708 19937 1748 22483
rect 1707 19928 1749 19937
rect 1707 19888 1708 19928
rect 1748 19888 1749 19928
rect 1707 19879 1749 19888
rect 1804 19601 1844 26767
rect 1996 26321 2036 32152
rect 2091 32192 2133 32201
rect 2091 32152 2092 32192
rect 2132 32152 2133 32192
rect 2091 32143 2133 32152
rect 2092 32058 2132 32143
rect 2188 30008 2228 33832
rect 2284 33704 2324 33713
rect 2284 31613 2324 33664
rect 2380 33704 2420 33832
rect 2475 33788 2517 33797
rect 2475 33748 2476 33788
rect 2516 33748 2517 33788
rect 2475 33739 2517 33748
rect 2380 33655 2420 33664
rect 2476 32864 2516 33739
rect 2380 32824 2476 32864
rect 2283 31604 2325 31613
rect 2283 31564 2284 31604
rect 2324 31564 2325 31604
rect 2283 31555 2325 31564
rect 2380 31277 2420 32824
rect 2476 32815 2516 32824
rect 2572 32192 2612 35176
rect 2667 35216 2709 35225
rect 2667 35176 2668 35216
rect 2708 35176 2709 35216
rect 2667 35167 2709 35176
rect 2668 33116 2708 35167
rect 2860 35057 2900 36688
rect 2955 35216 2997 35225
rect 2955 35176 2956 35216
rect 2996 35176 2997 35216
rect 2955 35167 2997 35176
rect 3052 35216 3092 36940
rect 3092 35176 3188 35216
rect 3052 35167 3092 35176
rect 2859 35048 2901 35057
rect 2859 35008 2860 35048
rect 2900 35008 2901 35048
rect 2859 34999 2901 35008
rect 2860 34217 2900 34999
rect 2859 34208 2901 34217
rect 2859 34168 2860 34208
rect 2900 34168 2901 34208
rect 2859 34159 2901 34168
rect 2668 33067 2708 33076
rect 2764 33620 2804 33629
rect 2572 32117 2612 32152
rect 2476 32108 2516 32117
rect 2476 31697 2516 32068
rect 2571 32108 2613 32117
rect 2571 32068 2572 32108
rect 2612 32068 2613 32108
rect 2571 32059 2613 32068
rect 2572 32028 2612 32059
rect 2475 31688 2517 31697
rect 2475 31648 2476 31688
rect 2516 31648 2517 31688
rect 2475 31639 2517 31648
rect 2667 31604 2709 31613
rect 2667 31564 2668 31604
rect 2708 31564 2709 31604
rect 2667 31555 2709 31564
rect 2571 31520 2613 31529
rect 2571 31480 2572 31520
rect 2612 31480 2613 31520
rect 2571 31471 2613 31480
rect 2379 31268 2421 31277
rect 2379 31228 2380 31268
rect 2420 31228 2421 31268
rect 2379 31219 2421 31228
rect 2476 30680 2516 30689
rect 2476 30521 2516 30640
rect 2475 30512 2517 30521
rect 2475 30472 2476 30512
rect 2516 30472 2517 30512
rect 2475 30463 2517 30472
rect 2572 30353 2612 31471
rect 2668 30848 2708 31555
rect 2668 30799 2708 30808
rect 2667 30596 2709 30605
rect 2667 30556 2668 30596
rect 2708 30556 2709 30596
rect 2667 30547 2709 30556
rect 2571 30344 2613 30353
rect 2571 30304 2572 30344
rect 2612 30304 2613 30344
rect 2571 30295 2613 30304
rect 2188 29968 2612 30008
rect 2380 29840 2420 29849
rect 2092 29800 2380 29840
rect 1995 26312 2037 26321
rect 1995 26272 1996 26312
rect 2036 26272 2037 26312
rect 1995 26263 2037 26272
rect 1900 24632 1940 24641
rect 1940 24592 2036 24632
rect 1900 24583 1940 24592
rect 1900 24380 1940 24389
rect 1900 23129 1940 24340
rect 1996 23885 2036 24592
rect 1995 23876 2037 23885
rect 1995 23836 1996 23876
rect 2036 23836 2037 23876
rect 1995 23827 2037 23836
rect 2092 23297 2132 29800
rect 2380 29791 2420 29800
rect 2476 29840 2516 29849
rect 2476 29672 2516 29800
rect 2380 29632 2516 29672
rect 2380 27917 2420 29632
rect 2572 29588 2612 29968
rect 2476 29548 2612 29588
rect 2379 27908 2421 27917
rect 2379 27868 2380 27908
rect 2420 27868 2421 27908
rect 2379 27859 2421 27868
rect 2476 26825 2516 29548
rect 2571 29420 2613 29429
rect 2571 29380 2572 29420
rect 2612 29380 2613 29420
rect 2571 29371 2613 29380
rect 2572 29177 2612 29371
rect 2571 29168 2613 29177
rect 2571 29128 2572 29168
rect 2612 29128 2613 29168
rect 2571 29119 2613 29128
rect 2668 28337 2708 30547
rect 2667 28328 2709 28337
rect 2667 28288 2668 28328
rect 2708 28288 2709 28328
rect 2667 28279 2709 28288
rect 2668 28194 2708 28279
rect 2764 27245 2804 33580
rect 2860 33620 2900 33629
rect 2860 31529 2900 33580
rect 2859 31520 2901 31529
rect 2859 31480 2860 31520
rect 2900 31480 2901 31520
rect 2859 31471 2901 31480
rect 2860 31352 2900 31392
rect 2956 31361 2996 35167
rect 3052 34376 3092 34385
rect 3052 33797 3092 34336
rect 3051 33788 3093 33797
rect 3051 33748 3052 33788
rect 3092 33748 3093 33788
rect 3051 33739 3093 33748
rect 3148 33690 3188 35176
rect 3243 34712 3285 34721
rect 3243 34672 3244 34712
rect 3284 34672 3285 34712
rect 3243 34663 3285 34672
rect 3244 34628 3284 34663
rect 3244 34577 3284 34588
rect 3052 33650 3188 33690
rect 3340 33704 3380 33713
rect 3052 32201 3092 33650
rect 3147 33452 3189 33461
rect 3147 33412 3148 33452
rect 3188 33412 3189 33452
rect 3147 33403 3189 33412
rect 3051 32192 3093 32201
rect 3051 32152 3052 32192
rect 3092 32152 3093 32192
rect 3051 32143 3093 32152
rect 3052 32058 3092 32143
rect 3052 31520 3092 31529
rect 3148 31520 3188 33403
rect 3340 32873 3380 33664
rect 3339 32864 3381 32873
rect 3339 32824 3340 32864
rect 3380 32824 3381 32864
rect 3339 32815 3381 32824
rect 3092 31480 3188 31520
rect 3436 31520 3476 40552
rect 3627 40508 3669 40517
rect 3627 40468 3628 40508
rect 3668 40468 3669 40508
rect 3627 40459 3669 40468
rect 3628 40424 3668 40459
rect 3628 40373 3668 40384
rect 3531 40256 3573 40265
rect 3531 40216 3532 40256
rect 3572 40216 3573 40256
rect 3531 40207 3573 40216
rect 3532 39164 3572 40207
rect 3820 39845 3860 40636
rect 3915 40592 3957 40601
rect 3915 40552 3916 40592
rect 3956 40552 3957 40592
rect 3915 40543 3957 40552
rect 3916 40088 3956 40543
rect 4107 40508 4149 40517
rect 4107 40468 4108 40508
rect 4148 40468 4149 40508
rect 4107 40459 4149 40468
rect 4108 40438 4148 40459
rect 4204 40433 4244 40636
rect 4299 40592 4341 40601
rect 4299 40552 4300 40592
rect 4340 40552 4341 40592
rect 4299 40543 4341 40552
rect 4108 40373 4148 40398
rect 4203 40424 4245 40433
rect 4203 40384 4204 40424
rect 4244 40384 4245 40424
rect 4203 40375 4245 40384
rect 4300 40340 4340 40543
rect 4396 40517 4436 40972
rect 4492 40853 4532 41224
rect 4491 40844 4533 40853
rect 4491 40804 4492 40844
rect 4532 40804 4533 40844
rect 4491 40795 4533 40804
rect 4588 40676 4628 41560
rect 4684 41441 4724 41896
rect 4780 41936 4820 42820
rect 4876 42776 4916 42787
rect 4876 42701 4916 42736
rect 5260 42776 5300 42785
rect 5356 42776 5396 43063
rect 5547 43028 5589 43037
rect 5547 42988 5548 43028
rect 5588 42988 5589 43028
rect 5547 42979 5589 42988
rect 5300 42736 5396 42776
rect 4875 42692 4917 42701
rect 4875 42652 4876 42692
rect 4916 42652 4917 42692
rect 4875 42643 4917 42652
rect 5260 42449 5300 42736
rect 5259 42440 5301 42449
rect 5259 42400 5260 42440
rect 5300 42400 5301 42440
rect 5259 42391 5301 42400
rect 5451 42440 5493 42449
rect 5451 42400 5452 42440
rect 5492 42400 5493 42440
rect 5451 42391 5493 42400
rect 5259 42272 5301 42281
rect 5259 42232 5260 42272
rect 5300 42232 5301 42272
rect 5259 42223 5301 42232
rect 4875 42188 4917 42197
rect 4875 42148 4876 42188
rect 4916 42148 4917 42188
rect 4875 42139 4917 42148
rect 4780 41887 4820 41896
rect 4876 41936 4916 42139
rect 5260 42029 5300 42223
rect 5259 42020 5301 42029
rect 5259 41980 5260 42020
rect 5300 41980 5301 42020
rect 5259 41971 5301 41980
rect 4876 41887 4916 41896
rect 5260 41936 5300 41971
rect 5260 41886 5300 41896
rect 5355 41768 5397 41777
rect 5355 41728 5356 41768
rect 5396 41728 5397 41768
rect 5355 41719 5397 41728
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 4683 41432 4725 41441
rect 4683 41392 4684 41432
rect 4724 41392 4725 41432
rect 4683 41383 4725 41392
rect 4875 41432 4917 41441
rect 4875 41392 4876 41432
rect 4916 41392 4917 41432
rect 4875 41383 4917 41392
rect 4684 41264 4724 41273
rect 4684 41105 4724 41224
rect 4779 41264 4821 41273
rect 4779 41224 4780 41264
rect 4820 41224 4821 41264
rect 4779 41215 4821 41224
rect 4876 41264 4916 41383
rect 5356 41348 5396 41719
rect 4876 41215 4916 41224
rect 5068 41308 5396 41348
rect 5068 41264 5108 41308
rect 5068 41215 5108 41224
rect 4780 41130 4820 41215
rect 4683 41096 4725 41105
rect 4683 41056 4684 41096
rect 4724 41056 4725 41096
rect 4683 41047 4725 41056
rect 4492 40636 4628 40676
rect 4779 40676 4821 40685
rect 4779 40636 4780 40676
rect 4820 40636 4821 40676
rect 4395 40508 4437 40517
rect 4395 40468 4396 40508
rect 4436 40468 4437 40508
rect 4395 40459 4437 40468
rect 4300 40291 4340 40300
rect 4396 40256 4436 40459
rect 4492 40424 4532 40636
rect 4779 40627 4821 40636
rect 4683 40592 4725 40601
rect 4683 40552 4684 40592
rect 4724 40552 4725 40592
rect 4683 40543 4725 40552
rect 4492 40375 4532 40384
rect 4587 40424 4629 40433
rect 4587 40384 4588 40424
rect 4628 40384 4629 40424
rect 4587 40375 4629 40384
rect 4684 40424 4724 40543
rect 4684 40375 4724 40384
rect 4780 40424 4820 40627
rect 4972 40592 5012 40601
rect 4780 40375 4820 40384
rect 4876 40552 4972 40592
rect 4588 40290 4628 40375
rect 4876 40256 4916 40552
rect 4972 40543 5012 40552
rect 5259 40592 5301 40601
rect 5259 40552 5260 40592
rect 5300 40552 5301 40592
rect 5259 40543 5301 40552
rect 4972 40424 5012 40435
rect 4972 40349 5012 40384
rect 5260 40424 5300 40543
rect 5356 40517 5396 41308
rect 5355 40508 5397 40517
rect 5355 40468 5356 40508
rect 5396 40468 5397 40508
rect 5355 40459 5397 40468
rect 5260 40375 5300 40384
rect 4971 40340 5013 40349
rect 4971 40300 4972 40340
rect 5012 40300 5013 40340
rect 4971 40291 5013 40300
rect 5355 40340 5397 40349
rect 5355 40300 5356 40340
rect 5396 40300 5397 40340
rect 5355 40291 5397 40300
rect 4396 40216 4532 40256
rect 4492 40172 4532 40216
rect 4684 40216 4916 40256
rect 4492 40132 4628 40172
rect 3916 40048 4244 40088
rect 3819 39836 3861 39845
rect 3819 39796 3820 39836
rect 3860 39796 3861 39836
rect 3819 39787 3861 39796
rect 4012 39752 4052 39761
rect 4204 39752 4244 40048
rect 4396 39752 4436 39761
rect 4204 39712 4396 39752
rect 4012 39509 4052 39712
rect 4396 39703 4436 39712
rect 4491 39752 4533 39761
rect 4491 39712 4492 39752
rect 4532 39712 4533 39752
rect 4491 39703 4533 39712
rect 4588 39752 4628 40132
rect 4588 39703 4628 39712
rect 4684 39752 4724 40216
rect 4779 40088 4821 40097
rect 4779 40048 4780 40088
rect 4820 40048 4821 40088
rect 4779 40039 4821 40048
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 4684 39703 4724 39712
rect 4492 39618 4532 39703
rect 4780 39584 4820 40039
rect 5356 39920 5396 40291
rect 5068 39880 5396 39920
rect 4971 39836 5013 39845
rect 4971 39796 4972 39836
rect 5012 39796 5013 39836
rect 4971 39787 5013 39796
rect 4875 39752 4917 39761
rect 4875 39712 4876 39752
rect 4916 39712 4917 39752
rect 4875 39703 4917 39712
rect 4684 39544 4820 39584
rect 4011 39500 4053 39509
rect 4011 39460 4012 39500
rect 4052 39460 4053 39500
rect 4011 39451 4053 39460
rect 4204 39500 4244 39509
rect 4244 39460 4436 39500
rect 4204 39451 4244 39460
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 4396 39248 4436 39460
rect 4396 39208 4628 39248
rect 3532 39124 3668 39164
rect 3628 38996 3668 39124
rect 3628 38921 3668 38956
rect 4107 38996 4149 39005
rect 4107 38956 4108 38996
rect 4148 38956 4149 38996
rect 4107 38947 4149 38956
rect 4395 38996 4437 39005
rect 4395 38956 4396 38996
rect 4436 38956 4437 38996
rect 4395 38947 4437 38956
rect 3532 38912 3572 38921
rect 3532 38669 3572 38872
rect 3627 38912 3669 38921
rect 3627 38872 3628 38912
rect 3668 38872 3669 38912
rect 3627 38863 3669 38872
rect 4108 38912 4148 38947
rect 3628 38832 3668 38863
rect 4108 38861 4148 38872
rect 4203 38744 4245 38753
rect 4203 38704 4204 38744
rect 4244 38704 4245 38744
rect 4203 38695 4245 38704
rect 3531 38660 3573 38669
rect 3531 38620 3532 38660
rect 3572 38620 3573 38660
rect 3531 38611 3573 38620
rect 3915 38240 3957 38249
rect 3915 38200 3916 38240
rect 3956 38200 3957 38240
rect 3915 38191 3957 38200
rect 3916 38081 3956 38191
rect 3915 38072 3957 38081
rect 3915 38032 3916 38072
rect 3956 38032 3957 38072
rect 3915 38023 3957 38032
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3531 37400 3573 37409
rect 3531 37360 3532 37400
rect 3572 37360 3573 37400
rect 3531 37351 3573 37360
rect 4011 37400 4053 37409
rect 4011 37360 4012 37400
rect 4052 37360 4053 37400
rect 4011 37351 4053 37360
rect 4108 37400 4148 37411
rect 3532 37266 3572 37351
rect 4012 36821 4052 37351
rect 4108 37325 4148 37360
rect 4107 37316 4149 37325
rect 4107 37276 4108 37316
rect 4148 37276 4149 37316
rect 4107 37267 4149 37276
rect 4011 36812 4053 36821
rect 4011 36772 4012 36812
rect 4052 36772 4053 36812
rect 4011 36763 4053 36772
rect 4107 36728 4149 36737
rect 4107 36688 4108 36728
rect 4148 36688 4149 36728
rect 4107 36679 4149 36688
rect 4108 36594 4148 36679
rect 4204 36401 4244 38695
rect 4396 37409 4436 38947
rect 4588 38926 4628 39208
rect 4588 38877 4628 38886
rect 4395 37400 4437 37409
rect 4395 37360 4396 37400
rect 4436 37360 4437 37400
rect 4395 37351 4437 37360
rect 4492 37400 4532 37411
rect 4492 37325 4532 37360
rect 4588 37400 4628 37409
rect 4491 37316 4533 37325
rect 4491 37276 4492 37316
rect 4532 37276 4533 37316
rect 4491 37267 4533 37276
rect 4299 36896 4341 36905
rect 4299 36856 4300 36896
rect 4340 36856 4341 36896
rect 4299 36847 4341 36856
rect 4300 36762 4340 36847
rect 4491 36812 4533 36821
rect 4491 36772 4492 36812
rect 4532 36772 4533 36812
rect 4491 36763 4533 36772
rect 4492 36728 4532 36763
rect 4203 36392 4245 36401
rect 4203 36352 4204 36392
rect 4244 36352 4245 36392
rect 4203 36343 4245 36352
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 4012 35888 4052 35897
rect 4012 35477 4052 35848
rect 4492 35729 4532 36688
rect 4588 36569 4628 37360
rect 4587 36560 4629 36569
rect 4587 36520 4588 36560
rect 4628 36520 4629 36560
rect 4587 36511 4629 36520
rect 4491 35720 4533 35729
rect 4491 35680 4492 35720
rect 4532 35680 4533 35720
rect 4491 35671 4533 35680
rect 4011 35468 4053 35477
rect 4011 35428 4012 35468
rect 4052 35428 4053 35468
rect 4011 35419 4053 35428
rect 3723 35300 3765 35309
rect 3723 35260 3724 35300
rect 3764 35260 3765 35300
rect 3723 35251 3765 35260
rect 3532 35202 3572 35211
rect 3724 35166 3764 35251
rect 3532 34721 3572 35162
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 3531 34712 3573 34721
rect 3531 34672 3532 34712
rect 3572 34672 3573 34712
rect 3531 34663 3573 34672
rect 4491 34628 4533 34637
rect 4491 34588 4492 34628
rect 4532 34588 4533 34628
rect 4491 34579 4533 34588
rect 4011 34460 4053 34469
rect 4011 34420 4012 34460
rect 4052 34420 4053 34460
rect 4011 34411 4053 34420
rect 4012 34376 4052 34411
rect 4012 34133 4052 34336
rect 4203 34376 4245 34385
rect 4203 34336 4204 34376
rect 4244 34336 4245 34376
rect 4203 34327 4245 34336
rect 4011 34124 4053 34133
rect 4011 34084 4012 34124
rect 4052 34084 4053 34124
rect 4011 34075 4053 34084
rect 4011 33872 4053 33881
rect 4011 33832 4012 33872
rect 4052 33832 4053 33872
rect 4011 33823 4053 33832
rect 4012 33738 4052 33823
rect 3820 33690 3860 33699
rect 3820 33461 3860 33650
rect 3819 33452 3861 33461
rect 3819 33412 3820 33452
rect 3860 33412 3861 33452
rect 3819 33403 3861 33412
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 4204 32864 4244 34327
rect 4299 33704 4341 33713
rect 4299 33664 4300 33704
rect 4340 33664 4341 33704
rect 4299 33655 4341 33664
rect 4300 33570 4340 33655
rect 4204 32815 4244 32824
rect 4492 32789 4532 34579
rect 4587 33368 4629 33377
rect 4587 33328 4588 33368
rect 4628 33328 4629 33368
rect 4587 33319 4629 33328
rect 4491 32780 4533 32789
rect 4491 32740 4492 32780
rect 4532 32740 4533 32780
rect 4491 32731 4533 32740
rect 3723 32276 3765 32285
rect 3723 32236 3724 32276
rect 3764 32236 3765 32276
rect 3723 32227 3765 32236
rect 3532 32178 3572 32187
rect 3724 32142 3764 32227
rect 3532 31604 3572 32138
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 3532 31564 3668 31604
rect 3436 31480 3572 31520
rect 3052 31471 3092 31480
rect 2860 31277 2900 31312
rect 2955 31352 2997 31361
rect 2955 31312 2956 31352
rect 2996 31312 2997 31352
rect 2955 31303 2997 31312
rect 3340 31352 3380 31361
rect 2859 31268 2901 31277
rect 2859 31228 2860 31268
rect 2900 31228 2901 31268
rect 2859 31219 2901 31228
rect 2860 30521 2900 31219
rect 2956 31109 2996 31303
rect 2955 31100 2997 31109
rect 2955 31060 2956 31100
rect 2996 31060 2997 31100
rect 2955 31051 2997 31060
rect 3147 31100 3189 31109
rect 3147 31060 3148 31100
rect 3188 31060 3189 31100
rect 3147 31051 3189 31060
rect 3051 30764 3093 30773
rect 3051 30724 3052 30764
rect 3092 30724 3093 30764
rect 3051 30715 3093 30724
rect 2859 30512 2901 30521
rect 2859 30472 2860 30512
rect 2900 30472 2901 30512
rect 2859 30463 2901 30472
rect 2955 29924 2997 29933
rect 2955 29884 2956 29924
rect 2996 29884 2997 29924
rect 2955 29875 2997 29884
rect 2860 29840 2900 29849
rect 2860 29765 2900 29800
rect 2956 29790 2996 29875
rect 2859 29756 2901 29765
rect 2859 29716 2860 29756
rect 2900 29716 2901 29756
rect 2859 29707 2901 29716
rect 2860 29093 2900 29707
rect 2956 29168 2996 29177
rect 2859 29084 2901 29093
rect 2859 29044 2860 29084
rect 2900 29044 2901 29084
rect 2859 29035 2901 29044
rect 2956 28001 2996 29128
rect 2955 27992 2997 28001
rect 2955 27952 2956 27992
rect 2996 27952 2997 27992
rect 2955 27943 2997 27952
rect 2860 27656 2900 27665
rect 2763 27236 2805 27245
rect 2763 27196 2764 27236
rect 2804 27196 2805 27236
rect 2763 27187 2805 27196
rect 2860 27068 2900 27616
rect 2955 27656 2997 27665
rect 2955 27616 2956 27656
rect 2996 27616 2997 27656
rect 2955 27607 2997 27616
rect 2956 27522 2996 27607
rect 2955 27320 2997 27329
rect 2955 27280 2956 27320
rect 2996 27280 2997 27320
rect 2955 27271 2997 27280
rect 2764 27028 2900 27068
rect 2380 26816 2420 26825
rect 2380 25565 2420 26776
rect 2475 26816 2517 26825
rect 2475 26776 2476 26816
rect 2516 26776 2517 26816
rect 2475 26767 2517 26776
rect 2476 26682 2516 26767
rect 2764 26732 2804 27028
rect 2860 26825 2900 26910
rect 2956 26900 2996 27271
rect 2956 26851 2996 26860
rect 2859 26816 2901 26825
rect 2859 26776 2860 26816
rect 2900 26776 2901 26816
rect 2859 26767 2901 26776
rect 2572 26692 2804 26732
rect 2475 26480 2517 26489
rect 2475 26440 2476 26480
rect 2516 26440 2517 26480
rect 2475 26431 2517 26440
rect 2476 26144 2516 26431
rect 2379 25556 2421 25565
rect 2379 25516 2380 25556
rect 2420 25516 2421 25556
rect 2379 25507 2421 25516
rect 2476 25481 2516 26104
rect 2475 25472 2517 25481
rect 2475 25432 2476 25472
rect 2516 25432 2517 25472
rect 2475 25423 2517 25432
rect 2476 25304 2516 25315
rect 2476 25229 2516 25264
rect 2475 25220 2517 25229
rect 2475 25180 2476 25220
rect 2516 25180 2517 25220
rect 2475 25171 2517 25180
rect 2187 24632 2229 24641
rect 2187 24592 2188 24632
rect 2228 24592 2229 24632
rect 2187 24583 2229 24592
rect 2284 24632 2324 24641
rect 2188 24498 2228 24583
rect 2187 23960 2229 23969
rect 2187 23920 2188 23960
rect 2228 23920 2229 23960
rect 2284 23960 2324 24592
rect 2284 23920 2420 23960
rect 2187 23911 2229 23920
rect 2091 23288 2133 23297
rect 2091 23248 2092 23288
rect 2132 23248 2133 23288
rect 2091 23239 2133 23248
rect 1899 23120 1941 23129
rect 1899 23080 1900 23120
rect 1940 23080 1941 23120
rect 1899 23071 1941 23080
rect 2188 22625 2228 23911
rect 2284 23792 2324 23801
rect 2187 22616 2229 22625
rect 2187 22576 2188 22616
rect 2228 22576 2229 22616
rect 2187 22567 2229 22576
rect 2284 21776 2324 23752
rect 2380 23792 2420 23920
rect 2380 22541 2420 23752
rect 2476 23120 2516 25171
rect 2379 22532 2421 22541
rect 2379 22492 2380 22532
rect 2420 22492 2421 22532
rect 2379 22483 2421 22492
rect 2476 22280 2516 23080
rect 2572 22532 2612 26692
rect 3052 26480 3092 30715
rect 3148 30017 3188 31051
rect 3340 30773 3380 31312
rect 3435 31352 3477 31361
rect 3435 31312 3436 31352
rect 3476 31312 3477 31352
rect 3435 31303 3477 31312
rect 3436 31218 3476 31303
rect 3339 30764 3381 30773
rect 3339 30724 3340 30764
rect 3380 30724 3381 30764
rect 3339 30715 3381 30724
rect 3532 30605 3572 31480
rect 3339 30596 3381 30605
rect 3339 30556 3340 30596
rect 3380 30556 3381 30596
rect 3339 30547 3381 30556
rect 3531 30596 3573 30605
rect 3531 30556 3532 30596
rect 3572 30556 3573 30596
rect 3531 30547 3573 30556
rect 3147 30008 3189 30017
rect 3147 29968 3148 30008
rect 3188 29968 3189 30008
rect 3147 29959 3189 29968
rect 3147 29336 3189 29345
rect 3147 29296 3148 29336
rect 3188 29296 3189 29336
rect 3147 29287 3189 29296
rect 3148 29202 3188 29287
rect 3147 29084 3189 29093
rect 3147 29044 3148 29084
rect 3188 29044 3189 29084
rect 3147 29035 3189 29044
rect 3148 28505 3188 29035
rect 3340 28916 3380 30547
rect 3628 30428 3668 31564
rect 3820 31352 3860 31361
rect 3820 31025 3860 31312
rect 3915 31352 3957 31361
rect 3915 31312 3916 31352
rect 3956 31312 3957 31352
rect 3915 31303 3957 31312
rect 4395 31352 4437 31361
rect 4395 31312 4396 31352
rect 4436 31312 4437 31352
rect 4395 31303 4437 31312
rect 3916 31218 3956 31303
rect 4396 31218 4436 31303
rect 3819 31016 3861 31025
rect 3819 30976 3820 31016
rect 3860 30976 3861 31016
rect 3819 30967 3861 30976
rect 4492 30932 4532 32731
rect 4396 30892 4532 30932
rect 3820 30680 3860 30691
rect 3820 30605 3860 30640
rect 3819 30596 3861 30605
rect 3819 30556 3820 30596
rect 3860 30556 3861 30596
rect 3819 30547 3861 30556
rect 3532 30388 3668 30428
rect 3436 29840 3476 29849
rect 3436 29597 3476 29800
rect 3435 29588 3477 29597
rect 3435 29548 3436 29588
rect 3476 29548 3477 29588
rect 3435 29539 3477 29548
rect 3436 29093 3476 29539
rect 3532 29345 3572 30388
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 3627 30008 3669 30017
rect 3627 29968 3628 30008
rect 3668 29968 3669 30008
rect 3627 29959 3669 29968
rect 3531 29336 3573 29345
rect 3531 29296 3532 29336
rect 3572 29296 3573 29336
rect 3531 29287 3573 29296
rect 3435 29084 3477 29093
rect 3435 29044 3436 29084
rect 3476 29044 3477 29084
rect 3435 29035 3477 29044
rect 3628 29000 3668 29959
rect 3964 29849 4004 29858
rect 4299 29840 4341 29849
rect 4004 29809 4244 29840
rect 3964 29800 4244 29809
rect 4107 29672 4149 29681
rect 4107 29632 4108 29672
rect 4148 29632 4149 29672
rect 4107 29623 4149 29632
rect 4108 29538 4148 29623
rect 4204 29336 4244 29800
rect 4299 29800 4300 29840
rect 4340 29800 4341 29840
rect 4299 29791 4341 29800
rect 4300 29706 4340 29791
rect 4300 29336 4340 29345
rect 4204 29296 4300 29336
rect 4300 29287 4340 29296
rect 3532 28960 3668 29000
rect 3340 28876 3476 28916
rect 3147 28496 3189 28505
rect 3147 28456 3148 28496
rect 3188 28456 3189 28496
rect 3147 28447 3189 28456
rect 3147 28328 3189 28337
rect 3147 28288 3148 28328
rect 3188 28288 3189 28328
rect 3147 28279 3189 28288
rect 3148 26489 3188 28279
rect 3339 27740 3381 27749
rect 3339 27700 3340 27740
rect 3380 27700 3381 27740
rect 3339 27691 3381 27700
rect 3243 27656 3285 27665
rect 3243 27616 3244 27656
rect 3284 27616 3285 27656
rect 3243 27607 3285 27616
rect 2764 26440 3092 26480
rect 3147 26480 3189 26489
rect 3147 26440 3148 26480
rect 3188 26440 3189 26480
rect 2667 26312 2709 26321
rect 2667 26272 2668 26312
rect 2708 26272 2709 26312
rect 2667 26263 2709 26272
rect 2668 26178 2708 26263
rect 2668 25556 2708 25565
rect 2764 25556 2804 26440
rect 3147 26431 3189 26440
rect 3244 26237 3284 27607
rect 3340 27572 3380 27691
rect 3340 27161 3380 27532
rect 3436 27656 3476 28876
rect 3532 28580 3572 28960
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 3532 28540 3668 28580
rect 3339 27152 3381 27161
rect 3339 27112 3340 27152
rect 3380 27112 3381 27152
rect 3339 27103 3381 27112
rect 3436 27077 3476 27616
rect 3628 27413 3668 28540
rect 4011 28496 4053 28505
rect 4011 28456 4012 28496
rect 4052 28456 4053 28496
rect 4011 28447 4053 28456
rect 3916 28328 3956 28339
rect 3916 28253 3956 28288
rect 3915 28244 3957 28253
rect 3915 28204 3916 28244
rect 3956 28204 3957 28244
rect 3915 28195 3957 28204
rect 4012 28076 4052 28447
rect 4107 28328 4149 28337
rect 4107 28288 4108 28328
rect 4148 28288 4149 28328
rect 4107 28279 4149 28288
rect 4300 28328 4340 28337
rect 4396 28328 4436 30892
rect 4491 30512 4533 30521
rect 4491 30472 4492 30512
rect 4532 30472 4533 30512
rect 4491 30463 4533 30472
rect 4492 29168 4532 30463
rect 4492 28505 4532 29128
rect 4491 28496 4533 28505
rect 4491 28456 4492 28496
rect 4532 28456 4533 28496
rect 4491 28447 4533 28456
rect 4340 28288 4532 28328
rect 4300 28279 4340 28288
rect 4108 28244 4148 28279
rect 4108 28193 4148 28204
rect 4012 28036 4148 28076
rect 3916 27656 3956 27665
rect 3916 27497 3956 27616
rect 3915 27488 3957 27497
rect 3915 27448 3916 27488
rect 3956 27448 3957 27488
rect 3915 27439 3957 27448
rect 3627 27404 3669 27413
rect 3627 27364 3628 27404
rect 3668 27364 3669 27404
rect 3627 27355 3669 27364
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 3435 27068 3477 27077
rect 3435 27028 3436 27068
rect 3476 27028 3477 27068
rect 3435 27019 3477 27028
rect 3627 27068 3669 27077
rect 4108 27068 4148 28036
rect 3627 27028 3628 27068
rect 3668 27028 3669 27068
rect 3627 27019 3669 27028
rect 3820 27028 4148 27068
rect 4396 27642 4436 27651
rect 3339 26984 3381 26993
rect 3339 26944 3340 26984
rect 3380 26944 3381 26984
rect 3339 26935 3381 26944
rect 3243 26228 3285 26237
rect 3243 26188 3244 26228
rect 3284 26188 3285 26228
rect 3243 26179 3285 26188
rect 3051 26144 3093 26153
rect 3051 26104 3052 26144
rect 3092 26104 3093 26144
rect 3051 26095 3093 26104
rect 2955 26060 2997 26069
rect 2955 26020 2956 26060
rect 2996 26020 2997 26060
rect 2955 26011 2997 26020
rect 2708 25516 2804 25556
rect 2859 25556 2901 25565
rect 2859 25516 2860 25556
rect 2900 25516 2901 25556
rect 2668 25507 2708 25516
rect 2859 25507 2901 25516
rect 2860 25422 2900 25507
rect 2956 25229 2996 26011
rect 3052 26010 3092 26095
rect 3244 25733 3284 26179
rect 3243 25724 3285 25733
rect 3243 25684 3244 25724
rect 3284 25684 3285 25724
rect 3243 25675 3285 25684
rect 3051 25472 3093 25481
rect 3051 25432 3052 25472
rect 3092 25432 3093 25472
rect 3051 25423 3093 25432
rect 3052 25304 3092 25423
rect 3052 25255 3092 25264
rect 2955 25220 2997 25229
rect 2955 25180 2956 25220
rect 2996 25180 2997 25220
rect 2955 25171 2997 25180
rect 2763 24632 2805 24641
rect 2763 24592 2764 24632
rect 2804 24592 2805 24632
rect 2763 24583 2805 24592
rect 3243 24632 3285 24641
rect 3243 24592 3244 24632
rect 3284 24592 3285 24632
rect 3243 24583 3285 24592
rect 2668 24548 2708 24557
rect 2668 23960 2708 24508
rect 2764 24498 2804 24583
rect 3051 24548 3093 24557
rect 3051 24508 3052 24548
rect 3092 24508 3093 24548
rect 3051 24499 3093 24508
rect 2955 24380 2997 24389
rect 2955 24340 2956 24380
rect 2996 24340 2997 24380
rect 2955 24331 2997 24340
rect 2763 23960 2805 23969
rect 2668 23920 2764 23960
rect 2804 23920 2805 23960
rect 2763 23911 2805 23920
rect 2764 23876 2804 23911
rect 2764 23825 2804 23836
rect 2860 23792 2900 23803
rect 2860 23717 2900 23752
rect 2859 23708 2901 23717
rect 2859 23668 2860 23708
rect 2900 23668 2901 23708
rect 2859 23659 2901 23668
rect 2667 23288 2709 23297
rect 2667 23248 2668 23288
rect 2708 23248 2709 23288
rect 2667 23239 2709 23248
rect 2668 23154 2708 23239
rect 2668 22532 2708 22541
rect 2572 22492 2668 22532
rect 2668 22483 2708 22492
rect 2860 22280 2900 22291
rect 2516 22240 2612 22280
rect 2476 22231 2516 22240
rect 1996 21736 2324 21776
rect 2380 21736 2516 21776
rect 1900 21356 1940 21365
rect 1803 19592 1845 19601
rect 1803 19552 1804 19592
rect 1844 19552 1845 19592
rect 1803 19543 1845 19552
rect 1611 17912 1653 17921
rect 1611 17872 1612 17912
rect 1652 17872 1653 17912
rect 1611 17863 1653 17872
rect 1611 15476 1653 15485
rect 1611 15436 1612 15476
rect 1652 15436 1653 15476
rect 1611 15427 1653 15436
rect 1515 15392 1557 15401
rect 1515 15352 1516 15392
rect 1556 15352 1557 15392
rect 1515 15343 1557 15352
rect 1516 14552 1556 14561
rect 1268 14008 1364 14048
rect 1228 13999 1268 14008
rect 1228 11696 1268 11705
rect 1324 11696 1364 14008
rect 1420 14512 1516 14552
rect 1420 13217 1460 14512
rect 1516 14503 1556 14512
rect 1612 14384 1652 15427
rect 1900 15317 1940 21316
rect 1996 20189 2036 21736
rect 2380 21692 2420 21736
rect 2092 21652 2420 21692
rect 2476 21692 2516 21736
rect 2092 21524 2132 21652
rect 2476 21643 2516 21652
rect 2572 21594 2612 22240
rect 2860 22205 2900 22240
rect 2859 22196 2901 22205
rect 2859 22156 2860 22196
rect 2900 22156 2901 22196
rect 2859 22147 2901 22156
rect 2476 21554 2612 21594
rect 2668 21594 2708 21603
rect 2092 21475 2132 21484
rect 2283 21524 2325 21533
rect 2283 21484 2284 21524
rect 2324 21484 2325 21524
rect 2283 21475 2325 21484
rect 1995 20180 2037 20189
rect 1995 20140 1996 20180
rect 2036 20140 2037 20180
rect 1995 20131 2037 20140
rect 1995 19760 2037 19769
rect 1995 19720 1996 19760
rect 2036 19720 2037 19760
rect 1995 19711 2037 19720
rect 1996 15737 2036 19711
rect 2091 19592 2133 19601
rect 2091 19552 2092 19592
rect 2132 19552 2133 19592
rect 2091 19543 2133 19552
rect 1995 15728 2037 15737
rect 1995 15688 1996 15728
rect 2036 15688 2037 15728
rect 1995 15679 2037 15688
rect 1899 15308 1941 15317
rect 1899 15268 1900 15308
rect 1940 15268 1941 15308
rect 1899 15259 1941 15268
rect 1708 14804 1748 14813
rect 1708 14477 1748 14764
rect 1996 14720 2036 15679
rect 2092 15653 2132 19543
rect 2284 19256 2324 21475
rect 2476 20768 2516 21554
rect 2668 20852 2708 21554
rect 2476 20096 2516 20728
rect 2476 20047 2516 20056
rect 2572 20812 2708 20852
rect 2476 19256 2516 19265
rect 2284 19216 2476 19256
rect 2476 19207 2516 19216
rect 2475 18668 2517 18677
rect 2475 18628 2476 18668
rect 2516 18628 2517 18668
rect 2475 18619 2517 18628
rect 2476 18534 2516 18619
rect 2572 17996 2612 20812
rect 2956 20768 2996 24331
rect 2668 20728 2996 20768
rect 2668 20684 2708 20728
rect 2668 20635 2708 20644
rect 3052 20516 3092 24499
rect 3244 24498 3284 24583
rect 3340 24128 3380 26935
rect 3435 26816 3477 26825
rect 3435 26776 3436 26816
rect 3476 26776 3477 26816
rect 3435 26767 3477 26776
rect 3436 24977 3476 26767
rect 3628 26480 3668 27019
rect 3532 26440 3668 26480
rect 3532 25817 3572 26440
rect 3820 26153 3860 27028
rect 4300 26984 4340 26993
rect 4012 26944 4300 26984
rect 4012 26900 4052 26944
rect 4300 26935 4340 26944
rect 3964 26860 4052 26900
rect 3964 26858 4004 26860
rect 3964 26809 4004 26818
rect 4203 26816 4245 26825
rect 4203 26776 4204 26816
rect 4244 26776 4245 26816
rect 4203 26767 4245 26776
rect 4107 26648 4149 26657
rect 4107 26608 4108 26648
rect 4148 26608 4149 26648
rect 4107 26599 4149 26608
rect 4108 26514 4148 26599
rect 4204 26228 4244 26767
rect 4396 26312 4436 27602
rect 4492 27488 4532 28288
rect 4588 27908 4628 33319
rect 4684 31445 4724 39544
rect 4876 39005 4916 39703
rect 4972 39702 5012 39787
rect 5068 39752 5108 39880
rect 5068 39703 5108 39712
rect 5260 39752 5300 39763
rect 5260 39677 5300 39712
rect 5259 39668 5301 39677
rect 5259 39628 5260 39668
rect 5300 39628 5301 39668
rect 5259 39619 5301 39628
rect 5355 39080 5397 39089
rect 5355 39040 5356 39080
rect 5396 39040 5397 39080
rect 5355 39031 5397 39040
rect 4875 38996 4917 39005
rect 4875 38956 4876 38996
rect 4916 38956 4917 38996
rect 4875 38947 4917 38956
rect 5260 38912 5300 38921
rect 4780 38744 4820 38753
rect 5260 38744 5300 38872
rect 5356 38912 5396 39031
rect 5356 38863 5396 38872
rect 5260 38704 5396 38744
rect 4780 38333 4820 38704
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5356 38408 5396 38704
rect 5356 38359 5396 38368
rect 4779 38324 4821 38333
rect 4779 38284 4780 38324
rect 4820 38284 4821 38324
rect 4779 38275 4821 38284
rect 5163 38240 5205 38249
rect 5163 38200 5164 38240
rect 5204 38200 5205 38240
rect 5163 38191 5205 38200
rect 5164 38106 5204 38191
rect 5452 37745 5492 42391
rect 5548 42029 5588 42979
rect 5643 42860 5685 42869
rect 5643 42820 5644 42860
rect 5684 42820 5685 42860
rect 5643 42811 5685 42820
rect 5547 42020 5589 42029
rect 5547 41980 5548 42020
rect 5588 41980 5589 42020
rect 5547 41971 5589 41980
rect 5547 41348 5589 41357
rect 5547 41308 5548 41348
rect 5588 41308 5589 41348
rect 5547 41299 5589 41308
rect 5548 38417 5588 41299
rect 5547 38408 5589 38417
rect 5547 38368 5548 38408
rect 5588 38368 5589 38408
rect 5547 38359 5589 38368
rect 5548 38240 5588 38251
rect 5548 38165 5588 38200
rect 5547 38156 5589 38165
rect 5547 38116 5548 38156
rect 5588 38116 5589 38156
rect 5547 38107 5589 38116
rect 5644 37820 5684 42811
rect 5836 41600 5876 44911
rect 6412 44288 6452 45667
rect 6892 45137 6932 54487
rect 6988 51848 7028 54664
rect 7083 53780 7125 53789
rect 7083 53740 7084 53780
rect 7124 53740 7125 53780
rect 7083 53731 7125 53740
rect 6988 51799 7028 51808
rect 7084 51848 7124 53731
rect 7180 52529 7220 56092
rect 7179 52520 7221 52529
rect 7179 52480 7180 52520
rect 7220 52480 7221 52520
rect 7179 52471 7221 52480
rect 7084 51799 7124 51808
rect 7180 51680 7220 52471
rect 7084 51640 7220 51680
rect 6988 48824 7028 48833
rect 6988 47825 7028 48784
rect 6987 47816 7029 47825
rect 6987 47776 6988 47816
rect 7028 47776 7029 47816
rect 6987 47767 7029 47776
rect 6988 47405 7028 47767
rect 6987 47396 7029 47405
rect 6987 47356 6988 47396
rect 7028 47356 7029 47396
rect 6987 47347 7029 47356
rect 7084 45389 7124 51640
rect 7179 50336 7221 50345
rect 7179 50296 7180 50336
rect 7220 50296 7221 50336
rect 7179 50287 7221 50296
rect 7180 50202 7220 50287
rect 7276 49916 7316 56176
rect 7468 56132 7508 56141
rect 7468 55460 7508 56092
rect 7468 55420 7604 55460
rect 7564 54867 7604 55420
rect 7564 54818 7604 54827
rect 7660 54704 7700 56755
rect 7755 56636 7797 56645
rect 7755 56596 7756 56636
rect 7796 56596 7797 56636
rect 7755 56587 7797 56596
rect 7756 55553 7796 56587
rect 7755 55544 7797 55553
rect 7755 55504 7756 55544
rect 7796 55504 7797 55544
rect 7755 55495 7797 55504
rect 7756 55410 7796 55495
rect 7755 54956 7797 54965
rect 7755 54916 7756 54956
rect 7796 54916 7797 54956
rect 7755 54907 7797 54916
rect 7756 54822 7796 54907
rect 7564 54664 7700 54704
rect 7564 54200 7604 54664
rect 7659 54536 7701 54545
rect 7659 54496 7660 54536
rect 7700 54496 7701 54536
rect 7659 54487 7701 54496
rect 7468 54160 7604 54200
rect 7468 51680 7508 54160
rect 7563 54032 7605 54041
rect 7563 53992 7564 54032
rect 7604 53992 7605 54032
rect 7563 53983 7605 53992
rect 7564 53898 7604 53983
rect 7563 52940 7605 52949
rect 7563 52900 7564 52940
rect 7604 52900 7605 52940
rect 7563 52891 7605 52900
rect 7564 51848 7604 52891
rect 7564 51799 7604 51808
rect 7468 51640 7604 51680
rect 7372 50084 7412 50093
rect 7412 50044 7508 50084
rect 7372 50035 7412 50044
rect 7276 49876 7412 49916
rect 7179 49076 7221 49085
rect 7179 49036 7180 49076
rect 7220 49036 7221 49076
rect 7179 49027 7221 49036
rect 7180 48161 7220 49027
rect 7179 48152 7221 48161
rect 7179 48112 7180 48152
rect 7220 48112 7221 48152
rect 7179 48103 7221 48112
rect 7180 47993 7220 48103
rect 7179 47984 7221 47993
rect 7179 47944 7180 47984
rect 7220 47944 7221 47984
rect 7179 47935 7221 47944
rect 7275 47396 7317 47405
rect 7275 47356 7276 47396
rect 7316 47356 7317 47396
rect 7275 47347 7317 47356
rect 7276 47312 7316 47347
rect 7276 47261 7316 47272
rect 7275 45464 7317 45473
rect 7275 45424 7276 45464
rect 7316 45424 7317 45464
rect 7275 45415 7317 45424
rect 7083 45380 7125 45389
rect 7083 45340 7084 45380
rect 7124 45340 7125 45380
rect 7083 45331 7125 45340
rect 6891 45128 6933 45137
rect 6891 45088 6892 45128
rect 6932 45088 6933 45128
rect 6891 45079 6933 45088
rect 7276 44960 7316 45415
rect 7372 45389 7412 49876
rect 7468 48819 7508 50044
rect 7564 49085 7604 51640
rect 7660 51185 7700 54487
rect 7756 53864 7796 53873
rect 7756 53528 7796 53824
rect 7852 53705 7892 58192
rect 7948 57896 7988 58360
rect 8044 58073 8084 58528
rect 8043 58064 8085 58073
rect 8043 58024 8044 58064
rect 8084 58024 8085 58064
rect 8043 58015 8085 58024
rect 7948 57847 7988 57856
rect 8043 57896 8085 57905
rect 8043 57856 8044 57896
rect 8084 57856 8085 57896
rect 8043 57847 8085 57856
rect 8044 57762 8084 57847
rect 8140 57476 8180 59452
rect 8044 57436 8180 57476
rect 7947 57140 7989 57149
rect 7947 57100 7948 57140
rect 7988 57100 7989 57140
rect 7947 57091 7989 57100
rect 7948 56972 7988 57091
rect 7948 56923 7988 56932
rect 7948 55469 7988 55554
rect 7947 55460 7989 55469
rect 7947 55420 7948 55460
rect 7988 55420 7989 55460
rect 7947 55411 7989 55420
rect 8044 55133 8084 57436
rect 8139 57056 8181 57065
rect 8139 57016 8140 57056
rect 8180 57016 8181 57056
rect 8139 57007 8181 57016
rect 8140 56922 8180 57007
rect 8139 56720 8181 56729
rect 8139 56680 8140 56720
rect 8180 56680 8181 56720
rect 8139 56671 8181 56680
rect 8043 55124 8085 55133
rect 8043 55084 8044 55124
rect 8084 55084 8085 55124
rect 8043 55075 8085 55084
rect 8140 54545 8180 56671
rect 8236 56057 8276 59620
rect 8428 59585 8468 60460
rect 8523 60451 8565 60460
rect 8523 59660 8565 59669
rect 8523 59620 8524 59660
rect 8564 59620 8565 59660
rect 8523 59611 8565 59620
rect 8427 59576 8469 59585
rect 8427 59536 8428 59576
rect 8468 59536 8469 59576
rect 8427 59527 8469 59536
rect 8331 59408 8373 59417
rect 8331 59368 8332 59408
rect 8372 59368 8373 59408
rect 8331 59359 8373 59368
rect 8332 57065 8372 59359
rect 8427 57896 8469 57905
rect 8427 57856 8428 57896
rect 8468 57856 8469 57896
rect 8427 57847 8469 57856
rect 8524 57896 8564 59611
rect 8620 59585 8660 62467
rect 8716 62432 8756 62803
rect 8716 62383 8756 62392
rect 8812 62432 8852 62971
rect 8812 62383 8852 62392
rect 8908 61760 8948 64240
rect 9004 62525 9044 64987
rect 9100 64616 9140 65332
rect 9195 65120 9237 65129
rect 9195 65080 9196 65120
rect 9236 65080 9237 65120
rect 9195 65071 9237 65080
rect 9100 64541 9140 64576
rect 9099 64532 9141 64541
rect 9099 64492 9100 64532
rect 9140 64492 9141 64532
rect 9099 64483 9141 64492
rect 9099 64364 9141 64373
rect 9099 64324 9100 64364
rect 9140 64324 9141 64364
rect 9099 64315 9141 64324
rect 9003 62516 9045 62525
rect 9003 62476 9004 62516
rect 9044 62476 9045 62516
rect 9003 62467 9045 62476
rect 8908 61720 9044 61760
rect 8811 61592 8853 61601
rect 8811 61552 8812 61592
rect 8852 61552 8853 61592
rect 8811 61543 8853 61552
rect 8908 61592 8948 61603
rect 8812 60920 8852 61543
rect 8908 61517 8948 61552
rect 8907 61508 8949 61517
rect 8907 61468 8908 61508
rect 8948 61468 8949 61508
rect 8907 61459 8949 61468
rect 8812 60871 8852 60880
rect 8907 60920 8949 60929
rect 8907 60880 8908 60920
rect 8948 60880 8949 60920
rect 8907 60871 8949 60880
rect 8908 60752 8948 60871
rect 8812 60712 8948 60752
rect 8619 59576 8661 59585
rect 8619 59536 8620 59576
rect 8660 59536 8661 59576
rect 8619 59527 8661 59536
rect 8620 59417 8660 59527
rect 8619 59408 8661 59417
rect 8619 59368 8620 59408
rect 8660 59368 8661 59408
rect 8619 59359 8661 59368
rect 8715 58064 8757 58073
rect 8715 58024 8716 58064
rect 8756 58024 8757 58064
rect 8715 58015 8757 58024
rect 8564 57856 8660 57896
rect 8524 57847 8564 57856
rect 8428 57485 8468 57847
rect 8427 57476 8469 57485
rect 8427 57436 8428 57476
rect 8468 57436 8469 57476
rect 8427 57427 8469 57436
rect 8331 57056 8373 57065
rect 8331 57016 8332 57056
rect 8372 57016 8373 57056
rect 8331 57007 8373 57016
rect 8427 56804 8469 56813
rect 8427 56764 8428 56804
rect 8468 56764 8469 56804
rect 8427 56755 8469 56764
rect 8235 56048 8277 56057
rect 8235 56008 8236 56048
rect 8276 56008 8277 56048
rect 8235 55999 8277 56008
rect 8332 55553 8372 55638
rect 8236 55544 8276 55553
rect 8236 55385 8276 55504
rect 8331 55544 8373 55553
rect 8331 55504 8332 55544
rect 8372 55504 8373 55544
rect 8331 55495 8373 55504
rect 8235 55376 8277 55385
rect 8235 55336 8236 55376
rect 8276 55336 8277 55376
rect 8235 55327 8277 55336
rect 8331 55292 8373 55301
rect 8331 55252 8332 55292
rect 8372 55252 8373 55292
rect 8331 55243 8373 55252
rect 8139 54536 8181 54545
rect 8139 54496 8140 54536
rect 8180 54496 8181 54536
rect 8139 54487 8181 54496
rect 8139 54368 8181 54377
rect 8139 54328 8140 54368
rect 8180 54328 8181 54368
rect 8139 54319 8181 54328
rect 8044 54032 8084 54041
rect 7851 53696 7893 53705
rect 7851 53656 7852 53696
rect 7892 53656 7893 53696
rect 7851 53647 7893 53656
rect 8044 53528 8084 53992
rect 7756 53488 8084 53528
rect 8140 54032 8180 54319
rect 8140 53444 8180 53992
rect 8332 53780 8372 55243
rect 8428 54872 8468 56755
rect 8523 56720 8565 56729
rect 8523 56680 8524 56720
rect 8564 56680 8565 56720
rect 8523 56671 8565 56680
rect 8524 56384 8564 56671
rect 8524 56335 8564 56344
rect 8620 55460 8660 57856
rect 8716 55721 8756 58015
rect 8812 57644 8852 60712
rect 8907 58904 8949 58913
rect 8907 58864 8908 58904
rect 8948 58864 8949 58904
rect 8907 58855 8949 58864
rect 8908 58241 8948 58855
rect 8907 58232 8949 58241
rect 8907 58192 8908 58232
rect 8948 58192 8949 58232
rect 8907 58183 8949 58192
rect 9004 58064 9044 61720
rect 8908 58024 9044 58064
rect 8908 57905 8948 58024
rect 8907 57896 8949 57905
rect 8907 57856 8908 57896
rect 8948 57856 8949 57896
rect 8907 57847 8949 57856
rect 9004 57896 9044 57907
rect 9004 57821 9044 57856
rect 9003 57812 9045 57821
rect 9003 57772 9004 57812
rect 9044 57772 9045 57812
rect 9003 57763 9045 57772
rect 8812 57604 9044 57644
rect 8811 57476 8853 57485
rect 8811 57436 8812 57476
rect 8852 57436 8853 57476
rect 8811 57427 8853 57436
rect 8715 55712 8757 55721
rect 8715 55672 8716 55712
rect 8756 55672 8757 55712
rect 8715 55663 8757 55672
rect 8812 55628 8852 57427
rect 8716 55544 8756 55553
rect 8620 55420 8663 55460
rect 8623 55376 8663 55420
rect 8615 55336 8663 55376
rect 8615 55292 8655 55336
rect 8615 55252 8660 55292
rect 8523 55208 8565 55217
rect 8523 55168 8524 55208
rect 8564 55168 8565 55208
rect 8523 55159 8565 55168
rect 8428 54823 8468 54832
rect 8524 54368 8564 55159
rect 7756 53404 8180 53444
rect 8236 53740 8372 53780
rect 8428 54328 8564 54368
rect 7756 51689 7796 53404
rect 8236 53360 8276 53740
rect 7948 53320 8236 53360
rect 7851 52856 7893 52865
rect 7851 52816 7852 52856
rect 7892 52816 7893 52856
rect 7851 52807 7893 52816
rect 7852 52520 7892 52807
rect 7755 51680 7797 51689
rect 7755 51640 7756 51680
rect 7796 51640 7797 51680
rect 7755 51631 7797 51640
rect 7852 51428 7892 52480
rect 7948 51605 7988 53320
rect 8236 53311 8276 53320
rect 8332 52520 8372 52529
rect 8044 52436 8084 52445
rect 8332 52436 8372 52480
rect 8084 52396 8372 52436
rect 8428 52520 8468 54328
rect 8523 54032 8565 54041
rect 8523 53992 8524 54032
rect 8564 53992 8565 54032
rect 8523 53983 8565 53992
rect 8620 54032 8660 55252
rect 8716 54041 8756 55504
rect 8812 55460 8852 55588
rect 8811 55420 8852 55460
rect 8811 55376 8851 55420
rect 8811 55336 8852 55376
rect 8524 53898 8564 53983
rect 8620 53873 8660 53992
rect 8715 54032 8757 54041
rect 8715 53992 8716 54032
rect 8756 53992 8757 54032
rect 8715 53983 8757 53992
rect 8619 53864 8661 53873
rect 8619 53824 8620 53864
rect 8660 53824 8661 53864
rect 8619 53815 8661 53824
rect 8716 53789 8756 53983
rect 8715 53780 8757 53789
rect 8715 53740 8716 53780
rect 8756 53740 8757 53780
rect 8715 53731 8757 53740
rect 8523 53696 8565 53705
rect 8523 53656 8524 53696
rect 8564 53656 8565 53696
rect 8812 53696 8852 55336
rect 8812 53656 8948 53696
rect 8523 53647 8565 53656
rect 8044 52387 8084 52396
rect 8428 52361 8468 52480
rect 8427 52352 8469 52361
rect 8427 52312 8428 52352
rect 8468 52312 8469 52352
rect 8427 52303 8469 52312
rect 8235 51932 8277 51941
rect 8235 51892 8236 51932
rect 8276 51892 8277 51932
rect 8235 51883 8277 51892
rect 8044 51834 8084 51843
rect 8236 51798 8276 51883
rect 7947 51596 7989 51605
rect 7947 51556 7948 51596
rect 7988 51556 7989 51596
rect 7947 51547 7989 51556
rect 7756 51388 7892 51428
rect 7659 51176 7701 51185
rect 7659 51136 7660 51176
rect 7700 51136 7701 51176
rect 7659 51127 7701 51136
rect 7659 51008 7701 51017
rect 7659 50968 7660 51008
rect 7700 50968 7701 51008
rect 7659 50959 7701 50968
rect 7756 51008 7796 51388
rect 7851 51260 7893 51269
rect 7851 51220 7852 51260
rect 7892 51220 7893 51260
rect 7851 51211 7893 51220
rect 7948 51260 7988 51269
rect 8044 51260 8084 51794
rect 8524 51764 8564 53647
rect 8715 53528 8757 53537
rect 8715 53488 8716 53528
rect 8756 53488 8757 53528
rect 8715 53479 8757 53488
rect 8619 53108 8661 53117
rect 8619 53068 8620 53108
rect 8660 53068 8661 53108
rect 8619 53059 8661 53068
rect 8620 51932 8660 53059
rect 8716 52445 8756 53479
rect 8812 52520 8852 52529
rect 8715 52436 8757 52445
rect 8715 52396 8716 52436
rect 8756 52396 8757 52436
rect 8715 52387 8757 52396
rect 8620 51892 8756 51932
rect 8620 51764 8660 51773
rect 8524 51724 8620 51764
rect 8620 51715 8660 51724
rect 8235 51680 8277 51689
rect 8235 51640 8236 51680
rect 8276 51640 8277 51680
rect 8235 51631 8277 51640
rect 7988 51220 8084 51260
rect 7948 51211 7988 51220
rect 7660 50336 7700 50959
rect 7756 50765 7796 50968
rect 7755 50756 7797 50765
rect 7755 50716 7756 50756
rect 7796 50716 7797 50756
rect 7755 50707 7797 50716
rect 7756 50336 7796 50345
rect 7660 50296 7756 50336
rect 7756 50287 7796 50296
rect 7852 50168 7892 51211
rect 7947 50336 7989 50345
rect 7947 50296 7948 50336
rect 7988 50296 7989 50336
rect 7947 50287 7989 50296
rect 7756 50128 7892 50168
rect 7563 49076 7605 49085
rect 7563 49036 7564 49076
rect 7604 49036 7605 49076
rect 7563 49027 7605 49036
rect 7660 48908 7700 48917
rect 7468 48770 7508 48779
rect 7564 48868 7660 48908
rect 7564 47237 7604 48868
rect 7660 48859 7700 48868
rect 7659 48320 7701 48329
rect 7659 48280 7660 48320
rect 7700 48280 7701 48320
rect 7659 48271 7701 48280
rect 7660 47984 7700 48271
rect 7660 47657 7700 47944
rect 7659 47648 7701 47657
rect 7659 47608 7660 47648
rect 7700 47608 7701 47648
rect 7659 47599 7701 47608
rect 7756 47396 7796 50128
rect 7948 49496 7988 50287
rect 8139 49832 8181 49841
rect 8139 49792 8140 49832
rect 8180 49792 8181 49832
rect 8139 49783 8181 49792
rect 8140 49748 8180 49783
rect 8140 49697 8180 49708
rect 8236 49580 8276 51631
rect 8428 51596 8468 51605
rect 8428 50849 8468 51556
rect 8619 51596 8661 51605
rect 8619 51556 8620 51596
rect 8660 51556 8661 51596
rect 8619 51547 8661 51556
rect 8523 51260 8565 51269
rect 8523 51220 8524 51260
rect 8564 51220 8565 51260
rect 8523 51211 8565 51220
rect 8524 51008 8564 51211
rect 8524 50959 8564 50968
rect 8427 50840 8469 50849
rect 8427 50800 8428 50840
rect 8468 50800 8469 50840
rect 8427 50791 8469 50800
rect 8620 50765 8660 51547
rect 8716 51269 8756 51892
rect 8715 51260 8757 51269
rect 8715 51220 8716 51260
rect 8756 51220 8757 51260
rect 8715 51211 8757 51220
rect 8619 50756 8661 50765
rect 8619 50716 8620 50756
rect 8660 50716 8661 50756
rect 8619 50707 8661 50716
rect 8331 50000 8373 50009
rect 8331 49960 8332 50000
rect 8372 49960 8373 50000
rect 8331 49951 8373 49960
rect 7948 49447 7988 49456
rect 8140 49540 8276 49580
rect 7947 49076 7989 49085
rect 7947 49036 7948 49076
rect 7988 49036 7989 49076
rect 7947 49027 7989 49036
rect 7948 48824 7988 49027
rect 7948 48775 7988 48784
rect 8043 48824 8085 48833
rect 8043 48784 8044 48824
rect 8084 48784 8085 48824
rect 8043 48775 8085 48784
rect 8044 48690 8084 48775
rect 7947 48068 7989 48077
rect 7947 48028 7948 48068
rect 7988 48028 7989 48068
rect 7947 48019 7989 48028
rect 7660 47356 7796 47396
rect 7852 47816 7892 47825
rect 7563 47228 7605 47237
rect 7563 47188 7564 47228
rect 7604 47188 7605 47228
rect 7563 47179 7605 47188
rect 7660 47144 7700 47356
rect 7852 47312 7892 47776
rect 7948 47480 7988 48019
rect 7948 47431 7988 47440
rect 7804 47302 7892 47312
rect 7844 47272 7892 47302
rect 7804 47253 7844 47262
rect 7660 47104 7796 47144
rect 7659 46640 7701 46649
rect 7659 46600 7660 46640
rect 7700 46600 7701 46640
rect 7659 46591 7701 46600
rect 7660 46472 7700 46591
rect 7660 45473 7700 46432
rect 7756 45893 7796 47104
rect 8140 46640 8180 49540
rect 8235 48992 8277 49001
rect 8235 48952 8236 48992
rect 8276 48952 8277 48992
rect 8235 48943 8277 48952
rect 8236 48824 8276 48943
rect 8236 48775 8276 48784
rect 8236 48572 8276 48581
rect 8236 47993 8276 48532
rect 8235 47984 8277 47993
rect 8235 47944 8236 47984
rect 8276 47944 8277 47984
rect 8235 47935 8277 47944
rect 8332 47144 8372 49951
rect 8427 49832 8469 49841
rect 8427 49792 8428 49832
rect 8468 49792 8469 49832
rect 8427 49783 8469 49792
rect 8428 49496 8468 49783
rect 8523 49748 8565 49757
rect 8523 49708 8524 49748
rect 8564 49708 8565 49748
rect 8523 49699 8565 49708
rect 8428 49447 8468 49456
rect 8524 49496 8564 49699
rect 8524 49447 8564 49456
rect 8620 49328 8660 50707
rect 8524 49288 8660 49328
rect 8428 48824 8468 48835
rect 8428 48749 8468 48784
rect 8427 48740 8469 48749
rect 8427 48700 8428 48740
rect 8468 48700 8469 48740
rect 8427 48691 8469 48700
rect 8524 47312 8564 49288
rect 8812 48152 8852 52480
rect 8908 52520 8948 53656
rect 8908 52361 8948 52480
rect 8907 52352 8949 52361
rect 8907 52312 8908 52352
rect 8948 52312 8949 52352
rect 8907 52303 8949 52312
rect 9004 50345 9044 57604
rect 9100 54032 9140 64315
rect 9196 55460 9236 65071
rect 9292 64868 9332 65752
rect 9387 65456 9429 65465
rect 9387 65416 9388 65456
rect 9428 65416 9429 65456
rect 9387 65407 9429 65416
rect 9292 64625 9332 64828
rect 9291 64616 9333 64625
rect 9291 64576 9292 64616
rect 9332 64576 9333 64616
rect 9291 64567 9333 64576
rect 9388 64205 9428 65407
rect 9484 64639 9524 66247
rect 9580 65129 9620 66508
rect 9676 65297 9716 67339
rect 9771 67220 9813 67229
rect 9771 67180 9772 67220
rect 9812 67180 9813 67220
rect 9771 67171 9813 67180
rect 9772 66968 9812 67171
rect 9868 67145 9908 67348
rect 9867 67136 9909 67145
rect 9867 67096 9868 67136
rect 9908 67096 9909 67136
rect 9867 67087 9909 67096
rect 9772 66919 9812 66928
rect 9675 65288 9717 65297
rect 9675 65248 9676 65288
rect 9716 65248 9717 65288
rect 9675 65239 9717 65248
rect 9579 65120 9621 65129
rect 9868 65120 9908 67087
rect 9579 65080 9580 65120
rect 9620 65080 9621 65120
rect 9579 65071 9621 65080
rect 9676 65080 9908 65120
rect 9579 64700 9621 64709
rect 9579 64660 9580 64700
rect 9620 64660 9621 64700
rect 9579 64651 9621 64660
rect 9484 64590 9524 64599
rect 9580 64616 9620 64651
rect 9580 64565 9620 64576
rect 9484 64532 9524 64541
rect 9387 64196 9429 64205
rect 9387 64156 9388 64196
rect 9428 64156 9429 64196
rect 9387 64147 9429 64156
rect 9387 63944 9429 63953
rect 9387 63904 9388 63944
rect 9428 63904 9429 63944
rect 9387 63895 9429 63904
rect 9291 63104 9333 63113
rect 9291 63064 9292 63104
rect 9332 63064 9333 63104
rect 9291 63055 9333 63064
rect 9292 62970 9332 63055
rect 9291 62516 9333 62525
rect 9291 62476 9292 62516
rect 9332 62476 9333 62516
rect 9291 62467 9333 62476
rect 9292 62432 9332 62467
rect 9292 58736 9332 62392
rect 9388 61517 9428 63895
rect 9484 63281 9524 64492
rect 9676 63356 9716 65080
rect 9772 64616 9812 64625
rect 9772 64448 9812 64576
rect 9867 64616 9909 64625
rect 9867 64576 9868 64616
rect 9908 64576 9909 64616
rect 9867 64567 9909 64576
rect 10022 64616 10064 64625
rect 10022 64576 10023 64616
rect 10063 64576 10064 64616
rect 10022 64567 10064 64576
rect 9868 64482 9908 64567
rect 10023 64482 10063 64567
rect 9772 64408 9813 64448
rect 9773 64364 9813 64408
rect 9772 64324 9813 64364
rect 9772 64121 9812 64324
rect 10059 64280 10101 64289
rect 10059 64240 10060 64280
rect 10100 64240 10101 64280
rect 10059 64231 10101 64240
rect 9771 64112 9813 64121
rect 9771 64072 9772 64112
rect 9812 64072 9813 64112
rect 9771 64063 9813 64072
rect 9964 63944 10004 63953
rect 9964 63701 10004 63904
rect 9963 63692 10005 63701
rect 9963 63652 9964 63692
rect 10004 63652 10005 63692
rect 9963 63643 10005 63652
rect 9676 63316 10004 63356
rect 9483 63272 9525 63281
rect 9483 63232 9484 63272
rect 9524 63232 9525 63272
rect 9483 63223 9525 63232
rect 9772 63113 9812 63198
rect 9867 63188 9909 63197
rect 9867 63148 9868 63188
rect 9908 63148 9909 63188
rect 9867 63139 9909 63148
rect 9771 63104 9813 63113
rect 9771 63064 9772 63104
rect 9812 63064 9813 63104
rect 9771 63055 9813 63064
rect 9868 63104 9908 63139
rect 9868 63053 9908 63064
rect 9484 62936 9524 62945
rect 9964 62936 10004 63316
rect 9524 62896 9812 62936
rect 9484 62887 9524 62896
rect 9483 62684 9525 62693
rect 9483 62644 9484 62684
rect 9524 62644 9525 62684
rect 9483 62635 9525 62644
rect 9387 61508 9429 61517
rect 9387 61468 9388 61508
rect 9428 61468 9429 61508
rect 9387 61459 9429 61468
rect 9484 59249 9524 62635
rect 9772 62427 9812 62896
rect 9772 62378 9812 62387
rect 9868 62896 10004 62936
rect 9675 62012 9717 62021
rect 9675 61972 9676 62012
rect 9716 61972 9717 62012
rect 9675 61963 9717 61972
rect 9579 61676 9621 61685
rect 9579 61636 9580 61676
rect 9620 61636 9621 61676
rect 9579 61627 9621 61636
rect 9580 59408 9620 61627
rect 9483 59240 9525 59249
rect 9483 59200 9484 59240
rect 9524 59200 9525 59240
rect 9483 59191 9525 59200
rect 9580 58913 9620 59368
rect 9579 58904 9621 58913
rect 9579 58864 9580 58904
rect 9620 58864 9621 58904
rect 9579 58855 9621 58864
rect 9292 58696 9428 58736
rect 9292 58568 9332 58579
rect 9292 58493 9332 58528
rect 9291 58484 9333 58493
rect 9291 58444 9292 58484
rect 9332 58444 9333 58484
rect 9291 58435 9333 58444
rect 9292 57905 9332 58435
rect 9291 57896 9333 57905
rect 9291 57856 9292 57896
rect 9332 57856 9333 57896
rect 9291 57847 9333 57856
rect 9388 57821 9428 58696
rect 9676 58568 9716 61963
rect 9771 61088 9813 61097
rect 9771 61048 9772 61088
rect 9812 61048 9813 61088
rect 9771 61039 9813 61048
rect 9772 60593 9812 61039
rect 9868 60845 9908 62896
rect 9963 62516 10005 62525
rect 9963 62476 9964 62516
rect 10004 62476 10005 62516
rect 9963 62467 10005 62476
rect 9964 62382 10004 62467
rect 10060 61088 10100 64231
rect 10156 63953 10196 67432
rect 10444 65297 10484 70456
rect 10635 70412 10677 70421
rect 10635 70372 10636 70412
rect 10676 70372 10677 70412
rect 10635 70363 10677 70372
rect 10636 68909 10676 70363
rect 10635 68900 10677 68909
rect 10635 68860 10636 68900
rect 10676 68860 10677 68900
rect 10635 68851 10677 68860
rect 10540 67640 10580 67649
rect 10540 66893 10580 67600
rect 10636 67640 10676 67649
rect 10539 66884 10581 66893
rect 10539 66844 10540 66884
rect 10580 66844 10581 66884
rect 10539 66835 10581 66844
rect 10636 66809 10676 67600
rect 10635 66800 10677 66809
rect 10635 66760 10636 66800
rect 10676 66760 10677 66800
rect 10635 66751 10677 66760
rect 10539 66632 10581 66641
rect 10539 66592 10540 66632
rect 10580 66592 10581 66632
rect 10539 66583 10581 66592
rect 10251 65288 10293 65297
rect 10251 65248 10252 65288
rect 10292 65248 10293 65288
rect 10251 65239 10293 65248
rect 10443 65288 10485 65297
rect 10443 65248 10444 65288
rect 10484 65248 10485 65288
rect 10443 65239 10485 65248
rect 10252 64616 10292 65239
rect 10540 65120 10580 66583
rect 10635 66548 10677 66557
rect 10635 66508 10636 66548
rect 10676 66508 10677 66548
rect 10635 66499 10677 66508
rect 10636 65456 10676 66499
rect 10636 65129 10676 65416
rect 10444 65080 10580 65120
rect 10635 65120 10677 65129
rect 10635 65080 10636 65120
rect 10676 65080 10677 65120
rect 10252 64373 10292 64576
rect 10347 64616 10389 64625
rect 10347 64576 10348 64616
rect 10388 64576 10389 64616
rect 10347 64567 10389 64576
rect 10348 64482 10388 64567
rect 10251 64364 10293 64373
rect 10251 64324 10252 64364
rect 10292 64324 10293 64364
rect 10251 64315 10293 64324
rect 10444 64280 10484 65080
rect 10635 65071 10677 65080
rect 10539 64952 10581 64961
rect 10539 64912 10540 64952
rect 10580 64912 10581 64952
rect 10539 64903 10581 64912
rect 10348 64240 10484 64280
rect 10155 63944 10197 63953
rect 10155 63904 10156 63944
rect 10196 63904 10197 63944
rect 10155 63895 10197 63904
rect 10348 63944 10388 64240
rect 10156 63692 10196 63701
rect 10156 63113 10196 63652
rect 10348 63365 10388 63904
rect 10443 63944 10485 63953
rect 10443 63904 10444 63944
rect 10484 63904 10485 63944
rect 10443 63895 10485 63904
rect 10347 63356 10389 63365
rect 10347 63316 10348 63356
rect 10388 63316 10389 63356
rect 10347 63307 10389 63316
rect 10251 63272 10293 63281
rect 10251 63232 10252 63272
rect 10292 63232 10293 63272
rect 10251 63223 10293 63232
rect 10252 63188 10292 63223
rect 10252 63137 10292 63148
rect 10347 63188 10389 63197
rect 10347 63148 10348 63188
rect 10388 63148 10389 63188
rect 10347 63139 10389 63148
rect 10155 63104 10197 63113
rect 10155 63064 10156 63104
rect 10196 63064 10197 63104
rect 10155 63055 10197 63064
rect 10348 63054 10388 63139
rect 10251 63020 10293 63029
rect 10251 62980 10252 63020
rect 10292 62980 10293 63020
rect 10251 62971 10293 62980
rect 10252 62357 10292 62971
rect 10444 62852 10484 63895
rect 10348 62812 10484 62852
rect 10251 62348 10293 62357
rect 10251 62308 10252 62348
rect 10292 62308 10293 62348
rect 10251 62299 10293 62308
rect 10348 62180 10388 62812
rect 10443 62348 10485 62357
rect 10443 62308 10444 62348
rect 10484 62308 10485 62348
rect 10443 62299 10485 62308
rect 10252 62140 10388 62180
rect 10155 61676 10197 61685
rect 10155 61636 10156 61676
rect 10196 61636 10197 61676
rect 10155 61627 10197 61636
rect 10156 61592 10196 61627
rect 10156 61541 10196 61552
rect 10155 61340 10197 61349
rect 10252 61340 10292 62140
rect 10155 61300 10156 61340
rect 10196 61300 10292 61340
rect 10348 61424 10388 61433
rect 10155 61291 10197 61300
rect 9964 61048 10100 61088
rect 9867 60836 9909 60845
rect 9867 60796 9868 60836
rect 9908 60796 9909 60836
rect 9867 60787 9909 60796
rect 9771 60584 9813 60593
rect 9771 60544 9772 60584
rect 9812 60544 9813 60584
rect 9771 60535 9813 60544
rect 9964 59669 10004 61048
rect 10059 60920 10101 60929
rect 10059 60880 10060 60920
rect 10100 60880 10101 60920
rect 10059 60871 10101 60880
rect 10060 60786 10100 60871
rect 10156 60332 10196 61291
rect 10252 61013 10292 61098
rect 10251 61004 10293 61013
rect 10251 60964 10252 61004
rect 10292 60964 10293 61004
rect 10348 61004 10388 61384
rect 10444 61181 10484 62299
rect 10540 61592 10580 64903
rect 10636 64448 10676 64457
rect 10636 63113 10676 64408
rect 10732 63197 10772 71380
rect 11020 71336 11060 71968
rect 10828 71296 11060 71336
rect 11116 71504 11156 72043
rect 10828 70664 10868 71296
rect 11116 71252 11156 71464
rect 11020 71212 11156 71252
rect 10924 70925 10964 71010
rect 10923 70916 10965 70925
rect 10923 70876 10924 70916
rect 10964 70876 10965 70916
rect 10923 70867 10965 70876
rect 10828 70615 10868 70624
rect 10923 70664 10965 70673
rect 10923 70624 10924 70664
rect 10964 70624 10965 70664
rect 10923 70615 10965 70624
rect 10924 70530 10964 70615
rect 11020 70412 11060 71212
rect 11212 71000 11252 72136
rect 11308 72176 11348 72185
rect 11308 72017 11348 72136
rect 11307 72008 11349 72017
rect 11307 71968 11308 72008
rect 11348 71968 11349 72008
rect 11307 71959 11349 71968
rect 11500 71672 11540 74908
rect 11788 74523 11828 74983
rect 11788 74474 11828 74483
rect 11884 73100 11924 80368
rect 11979 79400 12021 79409
rect 11979 79360 11980 79400
rect 12020 79360 12021 79400
rect 11979 79351 12021 79360
rect 11980 76712 12020 79351
rect 12076 79241 12116 80536
rect 12267 80240 12309 80249
rect 12267 80200 12268 80240
rect 12308 80200 12309 80240
rect 12267 80191 12309 80200
rect 12268 79997 12308 80191
rect 12267 79988 12309 79997
rect 12172 79948 12268 79988
rect 12308 79948 12309 79988
rect 12172 79325 12212 79948
rect 12267 79939 12309 79948
rect 12364 79913 12404 81367
rect 12460 80249 12500 81544
rect 12556 81341 12596 82720
rect 12652 82760 12692 82771
rect 12652 82685 12692 82720
rect 12651 82676 12693 82685
rect 12651 82636 12652 82676
rect 12692 82636 12693 82676
rect 12651 82627 12693 82636
rect 12652 82265 12692 82627
rect 12748 82592 12788 82601
rect 12651 82256 12693 82265
rect 12651 82216 12652 82256
rect 12692 82216 12693 82256
rect 12651 82207 12693 82216
rect 12652 82088 12692 82097
rect 12652 81929 12692 82048
rect 12651 81920 12693 81929
rect 12651 81880 12652 81920
rect 12692 81880 12693 81920
rect 12651 81871 12693 81880
rect 12555 81332 12597 81341
rect 12555 81292 12556 81332
rect 12596 81292 12597 81332
rect 12555 81283 12597 81292
rect 12459 80240 12501 80249
rect 12459 80200 12460 80240
rect 12500 80200 12501 80240
rect 12459 80191 12501 80200
rect 12363 79904 12405 79913
rect 12363 79864 12364 79904
rect 12404 79864 12405 79904
rect 12363 79855 12405 79864
rect 12267 79820 12309 79829
rect 12267 79780 12268 79820
rect 12308 79780 12309 79820
rect 12267 79771 12309 79780
rect 12268 79652 12308 79771
rect 12364 79757 12404 79766
rect 12364 79652 12404 79717
rect 12268 79612 12404 79652
rect 12556 79568 12596 79577
rect 12268 79528 12556 79568
rect 12171 79316 12213 79325
rect 12171 79276 12172 79316
rect 12212 79276 12213 79316
rect 12171 79267 12213 79276
rect 12075 79232 12117 79241
rect 12075 79192 12076 79232
rect 12116 79192 12117 79232
rect 12075 79183 12117 79192
rect 12076 78653 12116 79183
rect 12268 79064 12308 79528
rect 12556 79519 12596 79528
rect 12220 79054 12308 79064
rect 12260 79024 12308 79054
rect 12364 79148 12404 79157
rect 12220 79005 12260 79014
rect 12364 78821 12404 79108
rect 12555 79064 12597 79073
rect 12555 79024 12556 79064
rect 12596 79024 12597 79064
rect 12555 79015 12597 79024
rect 12556 78930 12596 79015
rect 12363 78812 12405 78821
rect 12363 78772 12364 78812
rect 12404 78772 12405 78812
rect 12363 78763 12405 78772
rect 12075 78644 12117 78653
rect 12075 78604 12076 78644
rect 12116 78604 12117 78644
rect 12075 78595 12117 78604
rect 12076 78233 12116 78238
rect 12075 78229 12117 78233
rect 12075 78184 12076 78229
rect 12116 78184 12117 78229
rect 12075 78175 12117 78184
rect 12076 78094 12116 78175
rect 12364 78149 12404 78763
rect 12171 78140 12213 78149
rect 12268 78140 12308 78149
rect 12171 78100 12172 78140
rect 12212 78100 12268 78140
rect 12171 78091 12213 78100
rect 12268 78091 12308 78100
rect 12363 78140 12405 78149
rect 12363 78100 12364 78140
rect 12404 78100 12405 78140
rect 12363 78091 12405 78100
rect 11980 76672 12116 76712
rect 11979 75620 12021 75629
rect 11979 75580 11980 75620
rect 12020 75580 12021 75620
rect 11979 75571 12021 75580
rect 11980 75461 12020 75571
rect 11979 75452 12021 75461
rect 11979 75412 11980 75452
rect 12020 75412 12021 75452
rect 11979 75403 12021 75412
rect 11979 75284 12021 75293
rect 11979 75244 11980 75284
rect 12020 75244 12021 75284
rect 11979 75235 12021 75244
rect 12076 75284 12116 76672
rect 12172 76385 12212 78091
rect 12460 77678 12500 77687
rect 12363 77636 12405 77645
rect 12460 77636 12500 77638
rect 12363 77596 12364 77636
rect 12404 77596 12500 77636
rect 12363 77587 12405 77596
rect 12316 77510 12356 77519
rect 12356 77470 12500 77510
rect 12316 77461 12356 77470
rect 12267 77300 12309 77309
rect 12267 77260 12268 77300
rect 12308 77260 12309 77300
rect 12267 77251 12309 77260
rect 12268 76973 12308 77251
rect 12267 76964 12309 76973
rect 12267 76924 12268 76964
rect 12308 76924 12309 76964
rect 12267 76915 12309 76924
rect 12171 76376 12213 76385
rect 12171 76336 12172 76376
rect 12212 76336 12213 76376
rect 12171 76327 12213 76336
rect 12172 76040 12212 76049
rect 12268 76040 12308 76915
rect 12460 76880 12500 77470
rect 12556 76880 12596 76889
rect 12460 76840 12556 76880
rect 12556 76831 12596 76840
rect 12363 76712 12405 76721
rect 12363 76672 12364 76712
rect 12404 76672 12405 76712
rect 12363 76663 12405 76672
rect 12364 76578 12404 76663
rect 12363 76376 12405 76385
rect 12363 76336 12364 76376
rect 12404 76336 12405 76376
rect 12363 76327 12405 76336
rect 12212 76000 12308 76040
rect 12172 75991 12212 76000
rect 12171 75620 12213 75629
rect 12171 75580 12172 75620
rect 12212 75580 12213 75620
rect 12171 75571 12213 75580
rect 11980 75150 12020 75235
rect 11979 74696 12021 74705
rect 11979 74656 11980 74696
rect 12020 74656 12021 74696
rect 11979 74647 12021 74656
rect 11980 74562 12020 74647
rect 12076 74444 12116 75244
rect 11692 73060 11924 73100
rect 11980 74404 12116 74444
rect 11692 73016 11732 73060
rect 11692 72437 11732 72976
rect 11691 72428 11733 72437
rect 11691 72388 11692 72428
rect 11732 72388 11733 72428
rect 11691 72379 11733 72388
rect 11692 72185 11732 72270
rect 11883 72260 11925 72269
rect 11883 72220 11884 72260
rect 11924 72220 11925 72260
rect 11883 72211 11925 72220
rect 11691 72176 11733 72185
rect 11691 72136 11692 72176
rect 11732 72136 11733 72176
rect 11691 72127 11733 72136
rect 11884 72176 11924 72211
rect 11884 72125 11924 72136
rect 11596 72008 11636 72017
rect 11636 71968 11924 72008
rect 11596 71959 11636 71968
rect 11787 71840 11829 71849
rect 11787 71800 11788 71840
rect 11828 71800 11829 71840
rect 11787 71791 11829 71800
rect 11500 71632 11732 71672
rect 11500 71504 11540 71513
rect 11404 71464 11500 71504
rect 11307 71252 11349 71261
rect 11307 71212 11308 71252
rect 11348 71212 11349 71252
rect 11307 71203 11349 71212
rect 11308 71118 11348 71203
rect 11212 70960 11348 71000
rect 11212 70664 11252 70673
rect 11115 70580 11157 70589
rect 11115 70540 11116 70580
rect 11156 70540 11157 70580
rect 11115 70531 11157 70540
rect 11116 70446 11156 70531
rect 10924 70372 11060 70412
rect 10827 69152 10869 69161
rect 10924 69152 10964 70372
rect 11212 70169 11252 70624
rect 11308 70421 11348 70960
rect 11307 70412 11349 70421
rect 11307 70372 11308 70412
rect 11348 70372 11349 70412
rect 11307 70363 11349 70372
rect 11211 70160 11253 70169
rect 11211 70120 11212 70160
rect 11252 70120 11253 70160
rect 11211 70111 11253 70120
rect 11116 69992 11156 70001
rect 11020 69404 11060 69413
rect 11116 69404 11156 69952
rect 11212 69992 11252 70020
rect 11404 69992 11444 71464
rect 11500 71455 11540 71464
rect 11596 71504 11636 71513
rect 11500 71336 11540 71345
rect 11500 70673 11540 71296
rect 11596 71261 11636 71464
rect 11595 71252 11637 71261
rect 11595 71212 11596 71252
rect 11636 71212 11637 71252
rect 11595 71203 11637 71212
rect 11692 71084 11732 71632
rect 11788 71504 11828 71791
rect 11788 71455 11828 71464
rect 11596 71044 11732 71084
rect 11499 70664 11541 70673
rect 11499 70624 11500 70664
rect 11540 70624 11541 70664
rect 11499 70615 11541 70624
rect 11596 70076 11636 71044
rect 11884 71000 11924 71968
rect 11788 70960 11924 71000
rect 11691 70916 11733 70925
rect 11691 70876 11692 70916
rect 11732 70876 11733 70916
rect 11691 70867 11733 70876
rect 11692 70496 11732 70867
rect 11788 70673 11828 70960
rect 11980 70916 12020 74404
rect 12075 74192 12117 74201
rect 12075 74152 12076 74192
rect 12116 74152 12117 74192
rect 12075 74143 12117 74152
rect 12076 73688 12116 74143
rect 12076 73613 12116 73648
rect 12075 73604 12117 73613
rect 12075 73564 12076 73604
rect 12116 73564 12117 73604
rect 12075 73555 12117 73564
rect 12075 71252 12117 71261
rect 12075 71212 12076 71252
rect 12116 71212 12117 71252
rect 12075 71203 12117 71212
rect 12076 71009 12116 71203
rect 12075 71000 12117 71009
rect 12075 70960 12076 71000
rect 12116 70960 12117 71000
rect 12075 70951 12117 70960
rect 11884 70876 12020 70916
rect 11787 70664 11829 70673
rect 11787 70624 11788 70664
rect 11828 70624 11829 70664
rect 11787 70615 11829 70624
rect 11692 70456 11828 70496
rect 11252 69952 11444 69992
rect 11500 70036 11636 70076
rect 11212 69943 11252 69952
rect 11308 69749 11348 69952
rect 11307 69740 11349 69749
rect 11307 69700 11308 69740
rect 11348 69700 11349 69740
rect 11307 69691 11349 69700
rect 11060 69364 11156 69404
rect 11020 69355 11060 69364
rect 11211 69320 11253 69329
rect 10827 69112 10828 69152
rect 10868 69112 10964 69152
rect 11116 69280 11212 69320
rect 11252 69280 11253 69320
rect 10827 69103 10869 69112
rect 10828 69018 10868 69103
rect 10827 68900 10869 68909
rect 10827 68860 10828 68900
rect 10868 68860 10869 68900
rect 10827 68851 10869 68860
rect 10828 66053 10868 68851
rect 11020 66968 11060 66977
rect 11020 66557 11060 66928
rect 11116 66641 11156 69280
rect 11211 69271 11253 69280
rect 11212 69152 11252 69161
rect 11212 68741 11252 69112
rect 11211 68732 11253 68741
rect 11211 68692 11212 68732
rect 11252 68692 11253 68732
rect 11211 68683 11253 68692
rect 11403 68732 11445 68741
rect 11500 68732 11540 70036
rect 11692 70001 11732 70086
rect 11691 69992 11733 70001
rect 11691 69952 11692 69992
rect 11732 69952 11733 69992
rect 11691 69943 11733 69952
rect 11595 69908 11637 69917
rect 11595 69868 11596 69908
rect 11636 69868 11637 69908
rect 11595 69859 11637 69868
rect 11596 69774 11636 69859
rect 11691 69740 11733 69749
rect 11691 69700 11692 69740
rect 11732 69700 11733 69740
rect 11691 69691 11733 69700
rect 11403 68692 11404 68732
rect 11444 68692 11540 68732
rect 11403 68683 11445 68692
rect 11404 68459 11444 68683
rect 11404 68410 11444 68419
rect 11596 68228 11636 68237
rect 11500 68188 11596 68228
rect 11500 67640 11540 68188
rect 11596 68179 11636 68188
rect 11500 67591 11540 67600
rect 11596 67640 11636 67649
rect 11692 67640 11732 69691
rect 11636 67600 11732 67640
rect 11212 67052 11252 67061
rect 11252 67012 11540 67052
rect 11212 67003 11252 67012
rect 11500 66968 11540 67012
rect 11500 66919 11540 66928
rect 11596 66968 11636 67600
rect 11596 66800 11636 66928
rect 11691 66884 11733 66893
rect 11691 66844 11692 66884
rect 11732 66844 11733 66884
rect 11691 66835 11733 66844
rect 11308 66760 11636 66800
rect 11115 66632 11157 66641
rect 11115 66592 11116 66632
rect 11156 66592 11157 66632
rect 11115 66583 11157 66592
rect 11019 66548 11061 66557
rect 11019 66508 11020 66548
rect 11060 66508 11061 66548
rect 11019 66499 11061 66508
rect 11212 66128 11252 66139
rect 11212 66053 11252 66088
rect 10827 66044 10869 66053
rect 10827 66004 10828 66044
rect 10868 66004 10869 66044
rect 10827 65995 10869 66004
rect 11211 66044 11253 66053
rect 11211 66004 11212 66044
rect 11252 66004 11253 66044
rect 11211 65995 11253 66004
rect 10828 65540 10868 65549
rect 10868 65500 11156 65540
rect 10828 65491 10868 65500
rect 11116 65456 11156 65500
rect 11116 65407 11156 65416
rect 11212 65456 11252 65465
rect 11308 65456 11348 66760
rect 11692 65624 11732 66835
rect 11252 65416 11348 65456
rect 11500 65584 11732 65624
rect 10923 65120 10965 65129
rect 10923 65080 10924 65120
rect 10964 65080 10965 65120
rect 10923 65071 10965 65080
rect 10827 64616 10869 64625
rect 10827 64576 10828 64616
rect 10868 64576 10869 64616
rect 10827 64567 10869 64576
rect 10828 63701 10868 64567
rect 10924 64541 10964 65071
rect 10923 64532 10965 64541
rect 10923 64492 10924 64532
rect 10964 64492 10965 64532
rect 10923 64483 10965 64492
rect 10827 63692 10869 63701
rect 10827 63652 10828 63692
rect 10868 63652 10869 63692
rect 10827 63643 10869 63652
rect 10731 63188 10773 63197
rect 10731 63148 10732 63188
rect 10772 63148 10773 63188
rect 10731 63139 10773 63148
rect 10635 63104 10677 63113
rect 10635 63064 10636 63104
rect 10676 63064 10677 63104
rect 10635 63055 10677 63064
rect 10828 63104 10868 63113
rect 10828 62768 10868 63064
rect 10732 62728 10868 62768
rect 10732 61937 10772 62728
rect 10827 62600 10869 62609
rect 10827 62560 10828 62600
rect 10868 62560 10869 62600
rect 10827 62551 10869 62560
rect 10731 61928 10773 61937
rect 10731 61888 10732 61928
rect 10772 61888 10773 61928
rect 10731 61879 10773 61888
rect 10540 61552 10772 61592
rect 10635 61424 10677 61433
rect 10635 61384 10636 61424
rect 10676 61384 10677 61424
rect 10635 61375 10677 61384
rect 10443 61172 10485 61181
rect 10443 61132 10444 61172
rect 10484 61132 10485 61172
rect 10443 61123 10485 61132
rect 10539 61004 10581 61013
rect 10348 60964 10484 61004
rect 10251 60955 10293 60964
rect 10156 60292 10388 60332
rect 9963 59660 10005 59669
rect 9963 59620 9964 59660
rect 10004 59620 10005 59660
rect 9963 59611 10005 59620
rect 10251 59660 10293 59669
rect 10251 59620 10252 59660
rect 10292 59620 10293 59660
rect 10251 59611 10293 59620
rect 9772 59492 9812 59501
rect 9812 59452 10100 59492
rect 9772 59443 9812 59452
rect 10060 59408 10100 59452
rect 10060 59359 10100 59368
rect 10156 59408 10196 59417
rect 10156 59249 10196 59368
rect 10155 59240 10197 59249
rect 10155 59200 10156 59240
rect 10196 59200 10197 59240
rect 10155 59191 10197 59200
rect 10252 59072 10292 59611
rect 10060 59032 10292 59072
rect 9868 58652 9908 58661
rect 9580 58528 9716 58568
rect 9772 58612 9868 58652
rect 9484 58400 9524 58409
rect 9484 57891 9524 58360
rect 9484 57842 9524 57851
rect 9387 57812 9429 57821
rect 9387 57772 9388 57812
rect 9428 57772 9429 57812
rect 9387 57763 9429 57772
rect 9388 57485 9428 57763
rect 9387 57476 9429 57485
rect 9387 57436 9388 57476
rect 9428 57436 9429 57476
rect 9387 57427 9429 57436
rect 9387 57224 9429 57233
rect 9387 57184 9388 57224
rect 9428 57184 9429 57224
rect 9387 57175 9429 57184
rect 9388 57056 9428 57175
rect 9580 57056 9620 58528
rect 9675 58400 9717 58409
rect 9675 58360 9676 58400
rect 9716 58360 9717 58400
rect 9675 58351 9717 58360
rect 9676 58266 9716 58351
rect 9676 58064 9716 58073
rect 9772 58064 9812 58612
rect 9868 58603 9908 58612
rect 10060 58568 10100 59032
rect 10348 58988 10388 60292
rect 10444 60080 10484 60964
rect 10539 60964 10540 61004
rect 10580 60964 10581 61004
rect 10539 60955 10581 60964
rect 10540 60920 10580 60955
rect 10540 60869 10580 60880
rect 10636 60920 10676 61375
rect 10636 60871 10676 60880
rect 10732 60257 10772 61552
rect 10731 60248 10773 60257
rect 10731 60208 10732 60248
rect 10772 60208 10773 60248
rect 10731 60199 10773 60208
rect 10540 60080 10580 60089
rect 10444 60040 10540 60080
rect 10540 60031 10580 60040
rect 10636 60080 10676 60089
rect 10676 60040 10772 60080
rect 10636 60031 10676 60040
rect 10635 59828 10677 59837
rect 10635 59788 10636 59828
rect 10676 59788 10677 59828
rect 10635 59779 10677 59788
rect 10443 59744 10485 59753
rect 10443 59704 10444 59744
rect 10484 59704 10485 59744
rect 10443 59695 10485 59704
rect 10444 59156 10484 59695
rect 10539 59408 10581 59417
rect 10539 59368 10540 59408
rect 10580 59368 10581 59408
rect 10539 59359 10581 59368
rect 10636 59408 10676 59779
rect 10540 59274 10580 59359
rect 10444 59116 10580 59156
rect 10252 58948 10388 58988
rect 10100 58528 10196 58568
rect 10060 58519 10100 58528
rect 10059 58400 10101 58409
rect 10059 58360 10060 58400
rect 10100 58360 10101 58400
rect 10059 58351 10101 58360
rect 9716 58024 9812 58064
rect 9676 58015 9716 58024
rect 9963 57560 10005 57569
rect 9963 57520 9964 57560
rect 10004 57520 10005 57560
rect 9963 57511 10005 57520
rect 9771 57056 9813 57065
rect 9580 57016 9716 57056
rect 9292 55544 9332 55553
rect 9292 55460 9332 55504
rect 9196 55420 9332 55460
rect 9100 52949 9140 53992
rect 9099 52940 9141 52949
rect 9099 52900 9100 52940
rect 9140 52900 9141 52940
rect 9099 52891 9141 52900
rect 9292 52025 9332 55420
rect 9388 53360 9428 57016
rect 9580 56888 9620 56897
rect 9580 56393 9620 56848
rect 9579 56384 9621 56393
rect 9579 56344 9580 56384
rect 9620 56344 9621 56384
rect 9579 56335 9621 56344
rect 9579 56132 9621 56141
rect 9579 56092 9580 56132
rect 9620 56092 9621 56132
rect 9579 56083 9621 56092
rect 9483 55796 9525 55805
rect 9483 55756 9484 55796
rect 9524 55756 9525 55796
rect 9483 55747 9525 55756
rect 9484 53948 9524 55747
rect 9580 54956 9620 56083
rect 9676 55460 9716 57016
rect 9771 57016 9772 57056
rect 9812 57016 9813 57056
rect 9771 57007 9813 57016
rect 9772 56922 9812 57007
rect 9771 56636 9813 56645
rect 9771 56596 9772 56636
rect 9812 56596 9813 56636
rect 9771 56587 9813 56596
rect 9772 56384 9812 56587
rect 9964 56384 10004 57511
rect 10060 56561 10100 58351
rect 10156 57896 10196 58528
rect 10156 57065 10196 57856
rect 10155 57056 10197 57065
rect 10155 57016 10156 57056
rect 10196 57016 10197 57056
rect 10155 57007 10197 57016
rect 10059 56552 10101 56561
rect 10059 56512 10060 56552
rect 10100 56512 10101 56552
rect 10059 56503 10101 56512
rect 10156 56468 10196 56477
rect 9964 56344 10100 56384
rect 9772 56141 9812 56344
rect 9771 56132 9813 56141
rect 9771 56092 9772 56132
rect 9812 56092 9813 56132
rect 9771 56083 9813 56092
rect 9964 56132 10004 56141
rect 9820 55553 9860 55562
rect 9964 55544 10004 56092
rect 9860 55513 10004 55544
rect 9820 55504 10004 55513
rect 10060 55460 10100 56344
rect 9676 55420 9908 55460
rect 9676 54965 9716 55050
rect 9675 54956 9717 54965
rect 9580 54916 9676 54956
rect 9716 54916 9717 54956
rect 9675 54907 9717 54916
rect 9676 54872 9716 54907
rect 9676 54823 9716 54832
rect 9868 54788 9908 55420
rect 9964 55420 10100 55460
rect 9964 55376 10004 55420
rect 9964 55327 10004 55336
rect 10156 55049 10196 56428
rect 10252 56216 10292 58948
rect 10443 58484 10485 58493
rect 10443 58444 10444 58484
rect 10484 58444 10485 58484
rect 10443 58435 10485 58444
rect 10347 56468 10389 56477
rect 10347 56428 10348 56468
rect 10388 56428 10389 56468
rect 10347 56419 10389 56428
rect 10348 56379 10388 56419
rect 10348 56330 10388 56339
rect 10252 56176 10388 56216
rect 10251 56048 10293 56057
rect 10251 56008 10252 56048
rect 10292 56008 10293 56048
rect 10251 55999 10293 56008
rect 10252 55805 10292 55999
rect 10251 55796 10293 55805
rect 10251 55756 10252 55796
rect 10292 55756 10293 55796
rect 10251 55747 10293 55756
rect 10155 55040 10197 55049
rect 10155 55000 10156 55040
rect 10196 55000 10197 55040
rect 10155 54991 10197 55000
rect 10060 54872 10100 54881
rect 10252 54872 10292 55747
rect 10100 54832 10292 54872
rect 10060 54823 10100 54832
rect 9868 54748 10004 54788
rect 9868 54620 9908 54629
rect 9676 54580 9868 54620
rect 9676 54116 9716 54580
rect 9868 54571 9908 54580
rect 9628 54076 9716 54116
rect 9867 54116 9909 54125
rect 9867 54076 9868 54116
rect 9908 54076 9909 54116
rect 9628 54074 9668 54076
rect 9867 54067 9909 54076
rect 9628 54025 9668 54034
rect 9772 53948 9812 53957
rect 9484 53908 9772 53948
rect 9772 53899 9812 53908
rect 9484 53360 9524 53369
rect 9388 53320 9484 53360
rect 9484 52865 9524 53320
rect 9868 53360 9908 54067
rect 9868 53285 9908 53320
rect 9867 53276 9909 53285
rect 9867 53236 9868 53276
rect 9908 53236 9909 53276
rect 9867 53227 9909 53236
rect 9868 53196 9908 53227
rect 9676 53108 9716 53117
rect 9716 53068 9908 53108
rect 9676 53059 9716 53068
rect 9483 52856 9525 52865
rect 9483 52816 9484 52856
rect 9524 52816 9525 52856
rect 9483 52807 9525 52816
rect 9771 52856 9813 52865
rect 9771 52816 9772 52856
rect 9812 52816 9813 52856
rect 9771 52807 9813 52816
rect 9387 52520 9429 52529
rect 9387 52480 9388 52520
rect 9428 52480 9429 52520
rect 9387 52471 9429 52480
rect 9388 52386 9428 52471
rect 9291 52016 9333 52025
rect 9291 51976 9292 52016
rect 9332 51976 9333 52016
rect 9291 51967 9333 51976
rect 9292 51848 9332 51967
rect 9580 51848 9620 51857
rect 9292 51799 9332 51808
rect 9388 51808 9580 51848
rect 9291 51596 9333 51605
rect 9291 51556 9292 51596
rect 9332 51556 9333 51596
rect 9291 51547 9333 51556
rect 9292 51462 9332 51547
rect 9388 50588 9428 51808
rect 9580 51799 9620 51808
rect 9772 51008 9812 52807
rect 9868 52534 9908 53068
rect 9868 52485 9908 52494
rect 9964 52016 10004 54748
rect 10059 53948 10101 53957
rect 10059 53908 10060 53948
rect 10100 53908 10101 53948
rect 10059 53899 10101 53908
rect 10060 52436 10100 53899
rect 10060 52387 10100 52396
rect 9772 50959 9812 50968
rect 9868 51976 10004 52016
rect 9868 50840 9908 51976
rect 9964 51848 10004 51857
rect 9964 51260 10004 51808
rect 10060 51848 10100 51857
rect 10060 51689 10100 51808
rect 10059 51680 10101 51689
rect 10059 51640 10060 51680
rect 10100 51640 10101 51680
rect 10059 51631 10101 51640
rect 9964 51211 10004 51220
rect 9196 50548 9428 50588
rect 9580 50800 9908 50840
rect 9196 50420 9236 50548
rect 9196 50345 9236 50380
rect 9003 50336 9045 50345
rect 9003 50296 9004 50336
rect 9044 50296 9045 50336
rect 9003 50287 9045 50296
rect 9195 50336 9237 50345
rect 9195 50296 9196 50336
rect 9236 50296 9237 50336
rect 9195 50287 9237 50296
rect 9484 50336 9524 50345
rect 9004 50202 9044 50287
rect 9196 50256 9236 50287
rect 9388 50084 9428 50093
rect 8907 49916 8949 49925
rect 8907 49876 8908 49916
rect 8948 49876 8949 49916
rect 8907 49867 8949 49876
rect 8908 49580 8948 49867
rect 8908 49531 8948 49540
rect 9003 49580 9045 49589
rect 9003 49540 9004 49580
rect 9044 49540 9045 49580
rect 9003 49531 9045 49540
rect 9004 49446 9044 49531
rect 9003 49244 9045 49253
rect 9003 49204 9004 49244
rect 9044 49204 9045 49244
rect 9003 49195 9045 49204
rect 8812 48112 8948 48152
rect 8715 48068 8757 48077
rect 8715 48028 8716 48068
rect 8756 48028 8757 48068
rect 8715 48019 8757 48028
rect 8619 47984 8661 47993
rect 8619 47944 8620 47984
rect 8660 47944 8661 47984
rect 8619 47935 8661 47944
rect 8620 47850 8660 47935
rect 8716 47934 8756 48019
rect 8811 47984 8853 47993
rect 8811 47944 8812 47984
rect 8852 47944 8853 47984
rect 8811 47935 8853 47944
rect 8812 47850 8852 47935
rect 8908 47648 8948 48112
rect 8524 47263 8564 47272
rect 8620 47608 8948 47648
rect 9004 47984 9044 49195
rect 9388 48833 9428 50044
rect 9484 49841 9524 50296
rect 9483 49832 9525 49841
rect 9483 49792 9484 49832
rect 9524 49792 9525 49832
rect 9483 49783 9525 49792
rect 9483 49496 9525 49505
rect 9483 49456 9484 49496
rect 9524 49456 9525 49496
rect 9483 49447 9525 49456
rect 9484 49362 9524 49447
rect 9483 49160 9525 49169
rect 9483 49120 9484 49160
rect 9524 49120 9525 49160
rect 9483 49111 9525 49120
rect 9387 48824 9429 48833
rect 9387 48784 9388 48824
rect 9428 48784 9429 48824
rect 9387 48775 9429 48784
rect 8332 47104 8564 47144
rect 8427 46808 8469 46817
rect 8427 46768 8428 46808
rect 8468 46768 8469 46808
rect 8427 46759 8469 46768
rect 8140 46600 8276 46640
rect 8140 46472 8180 46481
rect 7852 46388 7892 46397
rect 8140 46388 8180 46432
rect 7892 46348 8180 46388
rect 8236 46472 8276 46600
rect 7852 46339 7892 46348
rect 7755 45884 7797 45893
rect 7755 45844 7756 45884
rect 7796 45844 7797 45884
rect 7755 45835 7797 45844
rect 8139 45884 8181 45893
rect 8139 45844 8140 45884
rect 8180 45844 8181 45884
rect 8139 45835 8181 45844
rect 7659 45464 7701 45473
rect 7659 45424 7660 45464
rect 7700 45424 7701 45464
rect 7659 45415 7701 45424
rect 7371 45380 7413 45389
rect 7371 45340 7372 45380
rect 7412 45340 7413 45380
rect 7371 45331 7413 45340
rect 7372 44960 7412 44969
rect 7276 44920 7372 44960
rect 7372 44911 7412 44920
rect 7852 44960 7892 44969
rect 7564 44876 7604 44885
rect 7852 44876 7892 44920
rect 7947 44960 7989 44969
rect 7947 44920 7948 44960
rect 7988 44920 7989 44960
rect 7947 44911 7989 44920
rect 7604 44836 7892 44876
rect 7564 44827 7604 44836
rect 7948 44826 7988 44911
rect 6412 43709 6452 44248
rect 7660 44288 7700 44297
rect 6411 43700 6453 43709
rect 6411 43660 6412 43700
rect 6452 43660 6453 43700
rect 6411 43651 6453 43660
rect 7083 43700 7125 43709
rect 7083 43660 7084 43700
rect 7124 43660 7125 43700
rect 7083 43651 7125 43660
rect 6315 43448 6357 43457
rect 6315 43408 6316 43448
rect 6356 43408 6357 43448
rect 6315 43399 6357 43408
rect 6412 43448 6452 43457
rect 6316 42104 6356 43399
rect 6220 42064 6356 42104
rect 6123 41684 6165 41693
rect 6123 41644 6124 41684
rect 6164 41644 6165 41684
rect 6123 41635 6165 41644
rect 5740 41560 5876 41600
rect 5740 40433 5780 41560
rect 5835 41432 5877 41441
rect 5835 41392 5836 41432
rect 5876 41392 5877 41432
rect 5835 41383 5877 41392
rect 5739 40424 5781 40433
rect 5739 40384 5740 40424
rect 5780 40384 5781 40424
rect 5739 40375 5781 40384
rect 5836 40424 5876 41383
rect 5931 40844 5973 40853
rect 5931 40804 5932 40844
rect 5972 40804 5973 40844
rect 5931 40795 5973 40804
rect 5836 40375 5876 40384
rect 5739 40256 5781 40265
rect 5739 40216 5740 40256
rect 5780 40216 5781 40256
rect 5739 40207 5781 40216
rect 5740 40122 5780 40207
rect 5932 40004 5972 40795
rect 6124 40676 6164 41635
rect 6220 41096 6260 42064
rect 6315 41936 6357 41945
rect 6315 41896 6316 41936
rect 6356 41896 6357 41936
rect 6315 41887 6357 41896
rect 6316 41264 6356 41887
rect 6412 41441 6452 43408
rect 6603 43448 6645 43457
rect 6603 43408 6604 43448
rect 6644 43408 6645 43448
rect 6603 43399 6645 43408
rect 6795 43448 6837 43457
rect 6795 43408 6796 43448
rect 6836 43408 6837 43448
rect 6795 43399 6837 43408
rect 6892 43448 6932 43457
rect 6508 43364 6548 43373
rect 6508 42944 6548 43324
rect 6604 43314 6644 43399
rect 6508 42904 6644 42944
rect 6508 42776 6548 42785
rect 6508 42365 6548 42736
rect 6507 42356 6549 42365
rect 6507 42316 6508 42356
rect 6548 42316 6549 42356
rect 6507 42307 6549 42316
rect 6508 41945 6548 42307
rect 6507 41936 6549 41945
rect 6507 41896 6508 41936
rect 6548 41896 6549 41936
rect 6507 41887 6549 41896
rect 6508 41802 6548 41887
rect 6604 41609 6644 42904
rect 6699 42524 6741 42533
rect 6699 42484 6700 42524
rect 6740 42484 6741 42524
rect 6699 42475 6741 42484
rect 6700 42390 6740 42475
rect 6699 41936 6741 41945
rect 6699 41896 6700 41936
rect 6740 41896 6741 41936
rect 6699 41887 6741 41896
rect 6700 41852 6740 41887
rect 6700 41801 6740 41812
rect 6603 41600 6645 41609
rect 6603 41560 6604 41600
rect 6644 41560 6645 41600
rect 6603 41551 6645 41560
rect 6411 41432 6453 41441
rect 6508 41432 6548 41441
rect 6411 41392 6412 41432
rect 6452 41392 6508 41432
rect 6548 41392 6644 41432
rect 6411 41383 6453 41392
rect 6508 41383 6548 41392
rect 6412 41298 6452 41383
rect 6604 41264 6644 41392
rect 6700 41264 6740 41273
rect 6604 41224 6700 41264
rect 6316 41215 6356 41224
rect 6700 41215 6740 41224
rect 6796 41180 6836 43399
rect 6892 43205 6932 43408
rect 7084 43448 7124 43651
rect 7084 43399 7124 43408
rect 7276 43448 7316 43457
rect 7179 43364 7221 43373
rect 7179 43324 7180 43364
rect 7220 43324 7221 43364
rect 7179 43315 7221 43324
rect 6988 43280 7028 43289
rect 7028 43240 7124 43280
rect 6988 43231 7028 43240
rect 6891 43196 6933 43205
rect 6891 43156 6892 43196
rect 6932 43156 6933 43196
rect 6891 43147 6933 43156
rect 6987 42944 7029 42953
rect 6987 42904 6988 42944
rect 7028 42904 7029 42944
rect 6987 42895 7029 42904
rect 6988 42608 7028 42895
rect 6988 42533 7028 42568
rect 6987 42524 7029 42533
rect 6987 42484 6988 42524
rect 7028 42484 7029 42524
rect 6987 42475 7029 42484
rect 6988 42197 7028 42475
rect 6987 42188 7029 42197
rect 6987 42148 6988 42188
rect 7028 42148 7029 42188
rect 6987 42139 7029 42148
rect 6892 42029 6932 42041
rect 6891 42020 6933 42029
rect 6891 41980 6892 42020
rect 6932 41980 6933 42020
rect 6891 41971 6933 41980
rect 6892 41946 6932 41971
rect 6892 41897 6932 41906
rect 6988 41936 7028 41945
rect 6988 41777 7028 41896
rect 6987 41768 7029 41777
rect 6987 41728 6988 41768
rect 7028 41728 7029 41768
rect 6987 41719 7029 41728
rect 7084 41432 7124 43240
rect 7180 42617 7220 43315
rect 7276 42785 7316 43408
rect 7372 43448 7412 43459
rect 7372 43373 7412 43408
rect 7371 43364 7413 43373
rect 7371 43324 7372 43364
rect 7412 43324 7413 43364
rect 7371 43315 7413 43324
rect 7564 43280 7604 43289
rect 7468 43240 7564 43280
rect 7371 42944 7413 42953
rect 7371 42904 7372 42944
rect 7412 42904 7413 42944
rect 7371 42895 7413 42904
rect 7275 42776 7317 42785
rect 7275 42736 7276 42776
rect 7316 42736 7317 42776
rect 7275 42727 7317 42736
rect 7372 42776 7412 42895
rect 7372 42727 7412 42736
rect 7179 42608 7221 42617
rect 7179 42568 7180 42608
rect 7220 42568 7221 42608
rect 7179 42559 7221 42568
rect 7180 42449 7220 42559
rect 7179 42440 7221 42449
rect 7179 42400 7180 42440
rect 7220 42400 7221 42440
rect 7179 42391 7221 42400
rect 7276 41945 7316 42727
rect 7372 42608 7412 42617
rect 7468 42608 7508 43240
rect 7564 43231 7604 43240
rect 7412 42568 7508 42608
rect 7372 42559 7412 42568
rect 7371 42440 7413 42449
rect 7371 42400 7372 42440
rect 7412 42400 7413 42440
rect 7371 42391 7413 42400
rect 7275 41936 7317 41945
rect 7275 41896 7276 41936
rect 7316 41896 7317 41936
rect 7275 41887 7317 41896
rect 7372 41936 7412 42391
rect 7179 41852 7221 41861
rect 7179 41812 7180 41852
rect 7220 41812 7221 41852
rect 7179 41803 7221 41812
rect 7180 41768 7220 41803
rect 7180 41717 7220 41728
rect 7275 41684 7317 41693
rect 7275 41644 7276 41684
rect 7316 41644 7317 41684
rect 7275 41635 7317 41644
rect 7008 41392 7124 41432
rect 7008 41273 7048 41392
rect 7276 41348 7316 41635
rect 7372 41441 7412 41896
rect 7468 41693 7508 42568
rect 7564 42524 7604 42533
rect 7564 42104 7604 42484
rect 7660 42365 7700 44248
rect 8140 44288 8180 45835
rect 8236 44969 8276 46432
rect 8428 45044 8468 46759
rect 8428 44995 8468 45004
rect 8235 44960 8277 44969
rect 8235 44920 8236 44960
rect 8276 44920 8277 44960
rect 8235 44911 8277 44920
rect 8332 44960 8372 44971
rect 8332 44885 8372 44920
rect 8331 44876 8373 44885
rect 8331 44836 8332 44876
rect 8372 44836 8373 44876
rect 8331 44827 8373 44836
rect 8140 44239 8180 44248
rect 7852 44036 7892 44045
rect 7756 43996 7852 44036
rect 7756 43448 7796 43996
rect 7852 43987 7892 43996
rect 7756 43399 7796 43408
rect 7852 43448 7892 43457
rect 8044 43448 8084 43457
rect 7892 43408 8044 43448
rect 7852 43196 7892 43408
rect 8044 43399 8084 43408
rect 8235 43448 8277 43457
rect 8235 43408 8236 43448
rect 8276 43408 8277 43448
rect 8235 43399 8277 43408
rect 8332 43448 8372 43457
rect 8236 43314 8276 43399
rect 8140 43280 8180 43289
rect 8044 43240 8140 43280
rect 7756 43156 7892 43196
rect 7947 43196 7989 43205
rect 7947 43156 7948 43196
rect 7988 43156 7989 43196
rect 7756 42776 7796 43156
rect 7947 43147 7989 43156
rect 7756 42727 7796 42736
rect 7852 42692 7892 42701
rect 7659 42356 7701 42365
rect 7659 42316 7660 42356
rect 7700 42316 7701 42356
rect 7659 42307 7701 42316
rect 7852 42281 7892 42652
rect 7948 42608 7988 43147
rect 8044 42692 8084 43240
rect 8140 43231 8180 43240
rect 8332 42944 8372 43408
rect 8427 43364 8469 43373
rect 8427 43324 8428 43364
rect 8468 43324 8469 43364
rect 8427 43315 8469 43324
rect 8428 43121 8468 43315
rect 8524 43205 8564 47104
rect 8620 46472 8660 47608
rect 8715 46808 8757 46817
rect 8715 46768 8716 46808
rect 8756 46768 8757 46808
rect 8715 46759 8757 46768
rect 8716 46556 8756 46759
rect 8716 46507 8756 46516
rect 8620 44885 8660 46432
rect 9004 46313 9044 47944
rect 9196 46472 9236 46481
rect 9003 46304 9045 46313
rect 9003 46264 9004 46304
rect 9044 46264 9045 46304
rect 9003 46255 9045 46264
rect 8715 45800 8757 45809
rect 8715 45760 8716 45800
rect 8756 45760 8757 45800
rect 8715 45751 8757 45760
rect 8716 45666 8756 45751
rect 9196 45305 9236 46432
rect 8907 45296 8949 45305
rect 8907 45256 8908 45296
rect 8948 45256 8949 45296
rect 8907 45247 8949 45256
rect 9195 45296 9237 45305
rect 9195 45256 9196 45296
rect 9236 45256 9237 45296
rect 9195 45247 9237 45256
rect 8908 44960 8948 45247
rect 9484 45128 9524 49111
rect 9580 45212 9620 50800
rect 10059 50588 10101 50597
rect 10059 50548 10060 50588
rect 10100 50548 10101 50588
rect 10059 50539 10101 50548
rect 9867 50336 9909 50345
rect 9867 50296 9868 50336
rect 9908 50296 9909 50336
rect 9867 50287 9909 50296
rect 9964 50336 10004 50345
rect 9771 50252 9813 50261
rect 9771 50212 9772 50252
rect 9812 50212 9813 50252
rect 9771 50203 9813 50212
rect 9676 50084 9716 50093
rect 9676 49085 9716 50044
rect 9772 49169 9812 50203
rect 9868 50000 9908 50287
rect 9964 50084 10004 50296
rect 10060 50336 10100 50539
rect 10156 50429 10196 54832
rect 10251 51596 10293 51605
rect 10251 51556 10252 51596
rect 10292 51556 10293 51596
rect 10251 51547 10293 51556
rect 10155 50420 10197 50429
rect 10155 50380 10156 50420
rect 10196 50380 10197 50420
rect 10155 50371 10197 50380
rect 10060 50287 10100 50296
rect 10059 50084 10101 50093
rect 9964 50044 10060 50084
rect 10100 50044 10101 50084
rect 10059 50035 10101 50044
rect 9868 49960 10004 50000
rect 9964 49510 10004 49960
rect 10059 49832 10101 49841
rect 10059 49792 10060 49832
rect 10100 49792 10101 49832
rect 10059 49783 10101 49792
rect 9867 49496 9909 49505
rect 9867 49456 9868 49496
rect 9908 49456 9909 49496
rect 9867 49447 9909 49456
rect 9771 49160 9813 49169
rect 9771 49120 9772 49160
rect 9812 49120 9813 49160
rect 9771 49111 9813 49120
rect 9675 49076 9717 49085
rect 9675 49036 9676 49076
rect 9716 49036 9717 49076
rect 9675 49027 9717 49036
rect 9676 48824 9716 48833
rect 9772 48824 9812 49111
rect 9868 48992 9908 49447
rect 9868 48943 9908 48952
rect 9716 48784 9812 48824
rect 9964 48824 10004 49470
rect 10060 49160 10100 49783
rect 10252 49496 10292 51547
rect 10348 51176 10388 56176
rect 10444 52184 10484 58435
rect 10540 55721 10580 59116
rect 10636 56384 10676 59368
rect 10732 59249 10772 60040
rect 10731 59240 10773 59249
rect 10731 59200 10732 59240
rect 10772 59200 10773 59240
rect 10731 59191 10773 59200
rect 10828 58493 10868 62551
rect 10827 58484 10869 58493
rect 10827 58444 10828 58484
rect 10868 58444 10869 58484
rect 10827 58435 10869 58444
rect 10828 56384 10868 56393
rect 10636 56344 10828 56384
rect 10828 56335 10868 56344
rect 10924 56216 10964 64483
rect 11212 64280 11252 65416
rect 11307 65288 11349 65297
rect 11307 65248 11308 65288
rect 11348 65248 11349 65288
rect 11307 65239 11349 65248
rect 11116 64240 11252 64280
rect 11019 64196 11061 64205
rect 11019 64156 11020 64196
rect 11060 64156 11061 64196
rect 11019 64147 11061 64156
rect 11020 63785 11060 64147
rect 11019 63776 11061 63785
rect 11019 63736 11020 63776
rect 11060 63736 11061 63776
rect 11019 63727 11061 63736
rect 11116 62609 11156 64240
rect 11308 63272 11348 65239
rect 11403 64532 11445 64541
rect 11403 64492 11404 64532
rect 11444 64492 11445 64532
rect 11403 64483 11445 64492
rect 11212 63232 11348 63272
rect 11115 62600 11157 62609
rect 11115 62560 11116 62600
rect 11156 62560 11157 62600
rect 11115 62551 11157 62560
rect 11116 62432 11156 62441
rect 11116 61769 11156 62392
rect 11115 61760 11157 61769
rect 11115 61720 11116 61760
rect 11156 61720 11157 61760
rect 11115 61711 11157 61720
rect 11019 61592 11061 61601
rect 11019 61552 11020 61592
rect 11060 61552 11061 61592
rect 11019 61543 11061 61552
rect 11020 61433 11060 61543
rect 11116 61517 11156 61711
rect 11115 61508 11157 61517
rect 11115 61468 11116 61508
rect 11156 61468 11157 61508
rect 11115 61459 11157 61468
rect 11019 61424 11061 61433
rect 11019 61384 11020 61424
rect 11060 61384 11061 61424
rect 11019 61375 11061 61384
rect 11116 60920 11156 60929
rect 11212 60920 11252 63232
rect 11308 63113 11348 63118
rect 11307 63109 11349 63113
rect 11307 63064 11308 63109
rect 11348 63064 11349 63109
rect 11307 63055 11349 63064
rect 11308 62974 11348 63055
rect 11307 61760 11349 61769
rect 11307 61720 11308 61760
rect 11348 61720 11349 61760
rect 11307 61711 11349 61720
rect 11156 60880 11252 60920
rect 11116 60871 11156 60880
rect 11020 60836 11060 60845
rect 11020 60677 11060 60796
rect 11019 60668 11061 60677
rect 11019 60628 11020 60668
rect 11060 60628 11061 60668
rect 11019 60619 11061 60628
rect 11211 60248 11253 60257
rect 11116 60173 11156 60248
rect 11211 60208 11212 60248
rect 11252 60208 11253 60248
rect 11211 60199 11253 60208
rect 11019 60164 11061 60173
rect 11019 60124 11020 60164
rect 11060 60124 11061 60164
rect 11019 60115 11061 60124
rect 11116 60164 11168 60173
rect 11167 60124 11168 60164
rect 11116 60115 11168 60124
rect 11020 59417 11060 60115
rect 11115 59912 11157 59921
rect 11115 59872 11116 59912
rect 11156 59872 11157 59912
rect 11115 59863 11157 59872
rect 11019 59408 11061 59417
rect 11019 59368 11020 59408
rect 11060 59368 11061 59408
rect 11019 59359 11061 59368
rect 11116 59408 11156 59863
rect 11212 59669 11252 60199
rect 11211 59660 11253 59669
rect 11211 59620 11212 59660
rect 11252 59620 11253 59660
rect 11211 59611 11253 59620
rect 11116 59359 11156 59368
rect 11308 59324 11348 61711
rect 11404 61265 11444 64483
rect 11500 64289 11540 65584
rect 11595 65456 11637 65465
rect 11595 65416 11596 65456
rect 11636 65416 11637 65456
rect 11595 65407 11637 65416
rect 11692 65456 11732 65584
rect 11692 65407 11732 65416
rect 11596 65322 11636 65407
rect 11788 64373 11828 70456
rect 11884 64532 11924 70876
rect 12075 70832 12117 70841
rect 11980 70792 12076 70832
rect 12116 70792 12117 70832
rect 11980 70664 12020 70792
rect 12075 70783 12117 70792
rect 11980 70615 12020 70624
rect 12075 70664 12117 70673
rect 12075 70624 12076 70664
rect 12116 70624 12117 70664
rect 12075 70615 12117 70624
rect 12076 70530 12116 70615
rect 12075 70412 12117 70421
rect 12075 70372 12076 70412
rect 12116 70372 12117 70412
rect 12075 70363 12117 70372
rect 11979 70076 12021 70085
rect 11979 70036 11980 70076
rect 12020 70036 12021 70076
rect 11979 70027 12021 70036
rect 11980 69749 12020 70027
rect 12076 70001 12116 70363
rect 12075 69992 12117 70001
rect 12075 69952 12076 69992
rect 12116 69952 12117 69992
rect 12075 69943 12117 69952
rect 12172 69992 12212 75571
rect 12268 73520 12308 73529
rect 12268 73025 12308 73480
rect 12267 73016 12309 73025
rect 12267 72976 12268 73016
rect 12308 72976 12309 73016
rect 12267 72967 12309 72976
rect 12268 71513 12308 72967
rect 12364 71849 12404 76327
rect 12652 75713 12692 81871
rect 12748 81089 12788 82552
rect 12747 81080 12789 81089
rect 12747 81040 12748 81080
rect 12788 81040 12789 81080
rect 12747 81031 12789 81040
rect 12651 75704 12693 75713
rect 12651 75664 12652 75704
rect 12692 75664 12693 75704
rect 12651 75655 12693 75664
rect 12844 75629 12884 84484
rect 13036 84449 13076 84979
rect 13132 84524 13172 85063
rect 13324 84785 13364 85936
rect 13323 84776 13365 84785
rect 13323 84736 13324 84776
rect 13364 84736 13365 84776
rect 13323 84727 13365 84736
rect 13516 84701 13556 85936
rect 13515 84692 13557 84701
rect 13515 84652 13516 84692
rect 13556 84652 13557 84692
rect 13515 84643 13557 84652
rect 13132 84475 13172 84484
rect 13708 84449 13748 85936
rect 13803 85280 13845 85289
rect 13803 85240 13804 85280
rect 13844 85240 13845 85280
rect 13803 85231 13845 85240
rect 13035 84440 13077 84449
rect 13035 84400 13036 84440
rect 13076 84400 13077 84440
rect 13035 84391 13077 84400
rect 13707 84440 13749 84449
rect 13707 84400 13708 84440
rect 13748 84400 13749 84440
rect 13707 84391 13749 84400
rect 12940 84356 12980 84365
rect 12940 84113 12980 84316
rect 13131 84356 13173 84365
rect 13131 84316 13132 84356
rect 13172 84316 13173 84356
rect 13131 84307 13173 84316
rect 13515 84356 13557 84365
rect 13515 84316 13516 84356
rect 13556 84316 13557 84356
rect 13515 84307 13557 84316
rect 12939 84104 12981 84113
rect 12939 84064 12940 84104
rect 12980 84064 12981 84104
rect 12939 84055 12981 84064
rect 12940 83432 12980 84055
rect 12940 82601 12980 83392
rect 12939 82592 12981 82601
rect 12939 82552 12940 82592
rect 12980 82552 12981 82592
rect 12939 82543 12981 82552
rect 12940 82458 12980 82543
rect 13132 79400 13172 84307
rect 13419 84272 13461 84281
rect 13419 84232 13420 84272
rect 13460 84232 13461 84272
rect 13419 84223 13461 84232
rect 13323 84104 13365 84113
rect 13323 84064 13324 84104
rect 13364 84064 13365 84104
rect 13323 84055 13365 84064
rect 13324 83970 13364 84055
rect 13323 83684 13365 83693
rect 13323 83644 13324 83684
rect 13364 83644 13365 83684
rect 13323 83635 13365 83644
rect 13036 79360 13172 79400
rect 13228 83348 13268 83357
rect 13036 77897 13076 79360
rect 13228 78317 13268 83308
rect 13324 83273 13364 83635
rect 13420 83516 13460 84223
rect 13516 84222 13556 84307
rect 13708 84272 13748 84281
rect 13804 84272 13844 85231
rect 13900 84449 13940 85936
rect 13899 84440 13941 84449
rect 13899 84400 13900 84440
rect 13940 84400 13941 84440
rect 13899 84391 13941 84400
rect 14092 84281 14132 85936
rect 13612 84232 13708 84272
rect 13748 84232 13844 84272
rect 14091 84272 14133 84281
rect 14091 84232 14092 84272
rect 14132 84232 14133 84272
rect 13515 84104 13557 84113
rect 13515 84064 13516 84104
rect 13556 84064 13557 84104
rect 13515 84055 13557 84064
rect 13516 83693 13556 84055
rect 13515 83684 13557 83693
rect 13515 83644 13516 83684
rect 13556 83644 13557 83684
rect 13515 83635 13557 83644
rect 13612 83516 13652 84232
rect 13708 84223 13748 84232
rect 14091 84223 14133 84232
rect 13707 84104 13749 84113
rect 13707 84064 13708 84104
rect 13748 84064 13749 84104
rect 13707 84055 13749 84064
rect 13420 83467 13460 83476
rect 13516 83476 13652 83516
rect 13323 83264 13365 83273
rect 13323 83224 13324 83264
rect 13364 83224 13365 83264
rect 13323 83215 13365 83224
rect 13324 80744 13364 83215
rect 13516 83021 13556 83476
rect 13611 83348 13653 83357
rect 13611 83308 13612 83348
rect 13652 83308 13653 83348
rect 13611 83299 13653 83308
rect 13612 83214 13652 83299
rect 13515 83012 13557 83021
rect 13515 82972 13516 83012
rect 13556 82972 13557 83012
rect 13515 82963 13557 82972
rect 13612 82844 13652 82853
rect 13708 82844 13748 84055
rect 13996 83600 14036 83609
rect 13803 83516 13845 83525
rect 13803 83476 13804 83516
rect 13844 83476 13845 83516
rect 13803 83467 13845 83476
rect 13804 83382 13844 83467
rect 13996 83105 14036 83560
rect 14284 83525 14324 85936
rect 14379 85364 14421 85373
rect 14379 85324 14380 85364
rect 14420 85324 14421 85364
rect 14379 85315 14421 85324
rect 14283 83516 14325 83525
rect 14283 83476 14284 83516
rect 14324 83476 14325 83516
rect 14283 83467 14325 83476
rect 14380 83105 14420 85315
rect 14476 84365 14516 85936
rect 14668 85205 14708 85936
rect 14763 85448 14805 85457
rect 14763 85408 14764 85448
rect 14804 85408 14805 85448
rect 14763 85399 14805 85408
rect 14667 85196 14709 85205
rect 14667 85156 14668 85196
rect 14708 85156 14709 85196
rect 14667 85147 14709 85156
rect 14667 84692 14709 84701
rect 14667 84652 14668 84692
rect 14708 84652 14709 84692
rect 14667 84643 14709 84652
rect 14475 84356 14517 84365
rect 14475 84316 14476 84356
rect 14516 84316 14517 84356
rect 14475 84307 14517 84316
rect 14571 84020 14613 84029
rect 14571 83980 14572 84020
rect 14612 83980 14613 84020
rect 14571 83971 14613 83980
rect 13995 83096 14037 83105
rect 13995 83056 13996 83096
rect 14036 83056 14037 83096
rect 13995 83047 14037 83056
rect 14379 83096 14421 83105
rect 14379 83056 14380 83096
rect 14420 83056 14421 83096
rect 14379 83047 14421 83056
rect 14380 82928 14420 83047
rect 14380 82888 14516 82928
rect 13652 82804 13748 82844
rect 14476 82844 14516 82888
rect 13612 82795 13652 82804
rect 14476 82795 14516 82804
rect 13900 82760 13940 82769
rect 13708 82720 13900 82760
rect 13419 82592 13461 82601
rect 13419 82552 13420 82592
rect 13460 82552 13461 82592
rect 13419 82543 13461 82552
rect 13420 82458 13460 82543
rect 13612 81500 13652 81509
rect 13708 81500 13748 82720
rect 13900 82711 13940 82720
rect 13996 82760 14036 82769
rect 14379 82760 14421 82769
rect 14036 82720 14324 82760
rect 13996 82711 14036 82720
rect 14284 82256 14324 82720
rect 14379 82720 14380 82760
rect 14420 82720 14421 82760
rect 14379 82711 14421 82720
rect 14380 82626 14420 82711
rect 14572 82601 14612 83971
rect 14571 82592 14613 82601
rect 14571 82552 14572 82592
rect 14612 82552 14613 82592
rect 14571 82543 14613 82552
rect 14284 82216 14612 82256
rect 14092 82172 14132 82181
rect 14132 82132 14516 82172
rect 14092 82123 14132 82132
rect 13652 81460 13748 81500
rect 13900 82088 13940 82097
rect 13612 81451 13652 81460
rect 13900 81257 13940 82048
rect 14476 82088 14516 82132
rect 14476 82039 14516 82048
rect 14572 82088 14612 82216
rect 14379 82004 14421 82013
rect 14379 81964 14380 82004
rect 14420 81964 14421 82004
rect 14379 81955 14421 81964
rect 14283 81920 14325 81929
rect 14283 81880 14284 81920
rect 14324 81880 14325 81920
rect 14283 81871 14325 81880
rect 13420 81248 13460 81257
rect 13804 81248 13844 81257
rect 13420 80921 13460 81208
rect 13708 81208 13804 81248
rect 13419 80912 13461 80921
rect 13419 80872 13420 80912
rect 13460 80872 13461 80912
rect 13419 80863 13461 80872
rect 13324 80704 13460 80744
rect 13323 80576 13365 80585
rect 13323 80536 13324 80576
rect 13364 80536 13365 80576
rect 13323 80527 13365 80536
rect 13324 79829 13364 80527
rect 13323 79820 13365 79829
rect 13323 79780 13324 79820
rect 13364 79780 13365 79820
rect 13323 79771 13365 79780
rect 13420 79736 13460 80704
rect 13515 80660 13557 80669
rect 13515 80620 13516 80660
rect 13556 80620 13557 80660
rect 13515 80611 13557 80620
rect 13516 80526 13556 80611
rect 13708 80408 13748 81208
rect 13804 81199 13844 81208
rect 13899 81248 13941 81257
rect 13899 81208 13900 81248
rect 13940 81208 13941 81248
rect 13899 81199 13941 81208
rect 13900 80921 13940 81199
rect 13899 80912 13941 80921
rect 13899 80872 13900 80912
rect 13940 80872 13941 80912
rect 13899 80863 13941 80872
rect 13803 80660 13845 80669
rect 13803 80620 13804 80660
rect 13844 80620 13845 80660
rect 13803 80611 13845 80620
rect 13804 80576 13844 80611
rect 13804 80525 13844 80536
rect 13900 80576 13940 80585
rect 13708 80368 13844 80408
rect 13708 79736 13748 79745
rect 13420 79696 13708 79736
rect 13419 78560 13461 78569
rect 13419 78520 13420 78560
rect 13460 78520 13461 78560
rect 13419 78511 13461 78520
rect 13227 78308 13269 78317
rect 13227 78268 13228 78308
rect 13268 78268 13269 78308
rect 13227 78259 13269 78268
rect 13323 78224 13365 78233
rect 13323 78184 13324 78224
rect 13364 78184 13365 78224
rect 13323 78175 13365 78184
rect 13420 78224 13460 78511
rect 13420 78175 13460 78184
rect 13324 78090 13364 78175
rect 13035 77888 13077 77897
rect 13035 77848 13036 77888
rect 13076 77848 13077 77888
rect 13035 77839 13077 77848
rect 13420 77552 13460 77561
rect 13460 77512 13556 77552
rect 13420 77503 13460 77512
rect 13419 76712 13461 76721
rect 13419 76672 13420 76712
rect 13460 76672 13461 76712
rect 13419 76663 13461 76672
rect 13323 76628 13365 76637
rect 13323 76588 13324 76628
rect 13364 76588 13365 76628
rect 13323 76579 13365 76588
rect 12843 75620 12885 75629
rect 12843 75580 12844 75620
rect 12884 75580 12885 75620
rect 12843 75571 12885 75580
rect 13035 75284 13077 75293
rect 13035 75244 13036 75284
rect 13076 75244 13077 75284
rect 13035 75235 13077 75244
rect 13036 75214 13076 75235
rect 12555 75200 12597 75209
rect 12555 75160 12556 75200
rect 12596 75160 12597 75200
rect 12555 75151 12597 75160
rect 12556 75066 12596 75151
rect 13036 75149 13076 75174
rect 13228 75032 13268 75041
rect 12652 74992 13228 75032
rect 12459 74864 12501 74873
rect 12459 74824 12460 74864
rect 12500 74824 12501 74864
rect 12459 74815 12501 74824
rect 12460 74696 12500 74815
rect 12460 74647 12500 74656
rect 12555 74528 12597 74537
rect 12555 74488 12556 74528
rect 12596 74488 12597 74528
rect 12555 74479 12597 74488
rect 12460 73688 12500 73697
rect 12460 73193 12500 73648
rect 12459 73184 12501 73193
rect 12459 73144 12460 73184
rect 12500 73144 12501 73184
rect 12459 73135 12501 73144
rect 12363 71840 12405 71849
rect 12363 71800 12364 71840
rect 12404 71800 12405 71840
rect 12363 71791 12405 71800
rect 12364 71597 12404 71628
rect 12363 71588 12405 71597
rect 12363 71548 12364 71588
rect 12404 71548 12405 71588
rect 12363 71539 12405 71548
rect 12267 71504 12309 71513
rect 12267 71464 12268 71504
rect 12308 71464 12309 71504
rect 12267 71455 12309 71464
rect 12364 71504 12404 71539
rect 12268 71370 12308 71455
rect 12364 71009 12404 71464
rect 12363 71000 12405 71009
rect 12363 70960 12364 71000
rect 12404 70960 12405 71000
rect 12363 70951 12405 70960
rect 12267 70916 12309 70925
rect 12267 70876 12268 70916
rect 12308 70876 12309 70916
rect 12267 70867 12309 70876
rect 12268 70782 12308 70867
rect 12460 70841 12500 70926
rect 12459 70832 12501 70841
rect 12459 70792 12460 70832
rect 12500 70792 12501 70832
rect 12459 70783 12501 70792
rect 12268 70664 12308 70673
rect 12556 70664 12596 74479
rect 12652 74444 12692 74992
rect 13228 74983 13268 74992
rect 13324 74780 13364 76579
rect 13420 76049 13460 76663
rect 13516 76469 13556 77512
rect 13515 76460 13557 76469
rect 13515 76420 13516 76460
rect 13556 76420 13557 76460
rect 13515 76411 13557 76420
rect 13419 76040 13461 76049
rect 13419 76000 13420 76040
rect 13460 76000 13461 76040
rect 13419 75991 13461 76000
rect 13420 75906 13460 75991
rect 13516 75965 13556 76411
rect 13515 75956 13557 75965
rect 13515 75916 13516 75956
rect 13556 75916 13557 75956
rect 13515 75907 13557 75916
rect 13612 75788 13652 75797
rect 13515 75368 13557 75377
rect 13515 75328 13516 75368
rect 13556 75328 13557 75368
rect 13515 75319 13557 75328
rect 13516 75200 13556 75319
rect 13612 75293 13652 75748
rect 13611 75284 13653 75293
rect 13611 75244 13612 75284
rect 13652 75244 13653 75284
rect 13611 75235 13653 75244
rect 13516 75151 13556 75160
rect 13324 74740 13556 74780
rect 12843 74528 12885 74537
rect 12843 74488 12844 74528
rect 12884 74488 12885 74528
rect 12843 74479 12885 74488
rect 12940 74528 12980 74537
rect 12652 74395 12692 74404
rect 12844 74394 12884 74479
rect 12940 73772 12980 74488
rect 13036 74528 13076 74537
rect 13036 73856 13076 74488
rect 13131 74528 13173 74537
rect 13131 74488 13132 74528
rect 13172 74488 13173 74528
rect 13131 74479 13173 74488
rect 13420 74528 13460 74537
rect 13132 74394 13172 74479
rect 13420 73949 13460 74488
rect 13516 74528 13556 74740
rect 13419 73940 13461 73949
rect 13419 73900 13420 73940
rect 13460 73900 13461 73940
rect 13419 73891 13461 73900
rect 13036 73816 13364 73856
rect 12940 73732 13076 73772
rect 12939 73604 12981 73613
rect 12939 73564 12940 73604
rect 12980 73564 12981 73604
rect 12939 73555 12981 73564
rect 12940 73016 12980 73555
rect 12651 72932 12693 72941
rect 12651 72892 12652 72932
rect 12692 72892 12693 72932
rect 12651 72883 12693 72892
rect 12652 71597 12692 72883
rect 12843 72680 12885 72689
rect 12843 72640 12844 72680
rect 12884 72640 12885 72680
rect 12843 72631 12885 72640
rect 12844 71672 12884 72631
rect 12940 72176 12980 72976
rect 13036 72512 13076 73732
rect 13131 73688 13173 73697
rect 13131 73648 13132 73688
rect 13172 73648 13173 73688
rect 13131 73639 13173 73648
rect 13132 72941 13172 73639
rect 13324 73100 13364 73816
rect 13516 73697 13556 74488
rect 13611 74528 13653 74537
rect 13611 74488 13612 74528
rect 13652 74488 13653 74528
rect 13611 74479 13653 74488
rect 13515 73688 13557 73697
rect 13515 73648 13516 73688
rect 13556 73648 13557 73688
rect 13515 73639 13557 73648
rect 13612 73520 13652 74479
rect 13708 74117 13748 79696
rect 13804 79232 13844 80368
rect 13900 79409 13940 80536
rect 14284 80501 14324 81871
rect 14380 80576 14420 81955
rect 14572 81920 14612 82048
rect 14283 80492 14325 80501
rect 14283 80452 14284 80492
rect 14324 80452 14325 80492
rect 14283 80443 14325 80452
rect 14284 80358 14324 80443
rect 14380 79493 14420 80536
rect 14476 81880 14612 81920
rect 14379 79484 14421 79493
rect 14379 79444 14380 79484
rect 14420 79444 14421 79484
rect 14379 79435 14421 79444
rect 13899 79400 13941 79409
rect 13899 79360 13900 79400
rect 13940 79360 13941 79400
rect 13899 79351 13941 79360
rect 14476 79325 14516 81880
rect 14571 81752 14613 81761
rect 14571 81712 14572 81752
rect 14612 81712 14613 81752
rect 14571 81703 14613 81712
rect 14475 79316 14517 79325
rect 14475 79276 14476 79316
rect 14516 79276 14517 79316
rect 14475 79267 14517 79276
rect 13804 79192 13940 79232
rect 13803 79064 13845 79073
rect 13803 79024 13804 79064
rect 13844 79024 13845 79064
rect 13803 79015 13845 79024
rect 13804 78930 13844 79015
rect 13900 78737 13940 79192
rect 14379 79064 14421 79073
rect 14379 79024 14380 79064
rect 14420 79024 14516 79064
rect 14379 79015 14421 79024
rect 14091 78980 14133 78989
rect 14091 78940 14092 78980
rect 14132 78940 14133 78980
rect 14091 78931 14133 78940
rect 13996 78812 14036 78821
rect 13899 78728 13941 78737
rect 13899 78688 13900 78728
rect 13940 78688 13941 78728
rect 13899 78679 13941 78688
rect 13803 78392 13845 78401
rect 13803 78352 13804 78392
rect 13844 78352 13845 78392
rect 13803 78343 13845 78352
rect 13804 78308 13844 78343
rect 13804 78257 13844 78268
rect 13900 78224 13940 78235
rect 13996 78233 14036 78772
rect 13900 78149 13940 78184
rect 13995 78224 14037 78233
rect 13995 78184 13996 78224
rect 14036 78184 14037 78224
rect 13995 78175 14037 78184
rect 13899 78140 13941 78149
rect 13899 78100 13900 78140
rect 13940 78100 13941 78140
rect 13899 78091 13941 78100
rect 13996 76040 14036 76049
rect 13899 75704 13941 75713
rect 13899 75664 13900 75704
rect 13940 75664 13941 75704
rect 13899 75655 13941 75664
rect 13803 75116 13845 75125
rect 13803 75076 13804 75116
rect 13844 75076 13845 75116
rect 13803 75067 13845 75076
rect 13707 74108 13749 74117
rect 13707 74068 13708 74108
rect 13748 74068 13749 74108
rect 13707 74059 13749 74068
rect 13707 73772 13749 73781
rect 13707 73732 13708 73772
rect 13748 73732 13749 73772
rect 13707 73723 13749 73732
rect 13708 73688 13748 73723
rect 13708 73637 13748 73648
rect 13612 73480 13748 73520
rect 13516 73109 13556 73140
rect 13324 73051 13364 73060
rect 13515 73100 13557 73109
rect 13515 73060 13516 73100
rect 13556 73060 13557 73100
rect 13515 73051 13557 73060
rect 13420 73016 13460 73025
rect 13131 72932 13173 72941
rect 13131 72892 13132 72932
rect 13172 72892 13173 72932
rect 13131 72883 13173 72892
rect 13132 72764 13172 72773
rect 13420 72764 13460 72976
rect 13516 73016 13556 73051
rect 13516 72965 13556 72976
rect 13611 73016 13653 73025
rect 13611 72976 13612 73016
rect 13652 72976 13653 73016
rect 13611 72967 13653 72976
rect 13612 72882 13652 72967
rect 13515 72848 13557 72857
rect 13515 72808 13516 72848
rect 13556 72808 13557 72848
rect 13515 72799 13557 72808
rect 13172 72724 13460 72764
rect 13132 72715 13172 72724
rect 13036 72472 13364 72512
rect 13324 72428 13364 72472
rect 13324 72379 13364 72388
rect 13420 72185 13460 72724
rect 13132 72176 13172 72185
rect 12940 72136 13132 72176
rect 13132 72127 13172 72136
rect 13419 72176 13461 72185
rect 13419 72136 13420 72176
rect 13460 72136 13461 72176
rect 13419 72127 13461 72136
rect 13516 72176 13556 72799
rect 13612 72260 13652 72269
rect 13708 72260 13748 73480
rect 13804 73193 13844 75067
rect 13900 74705 13940 75655
rect 13996 75629 14036 76000
rect 13995 75620 14037 75629
rect 13995 75580 13996 75620
rect 14036 75580 14037 75620
rect 13995 75571 14037 75580
rect 13995 74948 14037 74957
rect 13995 74908 13996 74948
rect 14036 74908 14037 74948
rect 13995 74899 14037 74908
rect 13899 74696 13941 74705
rect 13899 74656 13900 74696
rect 13940 74656 13941 74696
rect 13899 74647 13941 74656
rect 13900 74528 13940 74647
rect 13900 74108 13940 74488
rect 13996 74528 14036 74899
rect 13996 74369 14036 74488
rect 13995 74360 14037 74369
rect 13995 74320 13996 74360
rect 14036 74320 14037 74360
rect 13995 74311 14037 74320
rect 13900 74068 14036 74108
rect 13899 73940 13941 73949
rect 13899 73900 13900 73940
rect 13940 73900 13941 73940
rect 13899 73891 13941 73900
rect 13900 73806 13940 73891
rect 13996 73688 14036 74068
rect 13900 73648 14036 73688
rect 13803 73184 13845 73193
rect 13803 73144 13804 73184
rect 13844 73144 13845 73184
rect 13803 73135 13845 73144
rect 13900 73109 13940 73648
rect 13995 73520 14037 73529
rect 13995 73480 13996 73520
rect 14036 73480 14037 73520
rect 13995 73471 14037 73480
rect 13899 73100 13941 73109
rect 13899 73060 13900 73100
rect 13940 73060 13941 73100
rect 13899 73051 13941 73060
rect 13803 73016 13845 73025
rect 13803 72976 13804 73016
rect 13844 72976 13845 73016
rect 13803 72967 13845 72976
rect 13996 73016 14036 73471
rect 13652 72220 13748 72260
rect 13612 72211 13652 72220
rect 13420 72017 13460 72127
rect 13324 72008 13364 72017
rect 13035 71924 13077 71933
rect 13035 71884 13036 71924
rect 13076 71884 13077 71924
rect 13035 71875 13077 71884
rect 12844 71632 12980 71672
rect 12651 71588 12693 71597
rect 12651 71548 12652 71588
rect 12692 71548 12693 71588
rect 12651 71539 12693 71548
rect 12844 71504 12884 71513
rect 12940 71504 12980 71632
rect 12748 71462 12788 71471
rect 12884 71464 12980 71504
rect 12844 71455 12884 71464
rect 12748 71420 12788 71422
rect 12308 70624 12596 70664
rect 12652 71380 12788 71420
rect 12268 70615 12308 70624
rect 12652 70505 12692 71380
rect 12747 70832 12789 70841
rect 12747 70792 12748 70832
rect 12788 70792 12789 70832
rect 12747 70783 12789 70792
rect 12748 70706 12788 70783
rect 12748 70657 12788 70666
rect 12843 70664 12885 70673
rect 12843 70624 12844 70664
rect 12884 70624 12885 70664
rect 12843 70615 12885 70624
rect 12651 70496 12693 70505
rect 12651 70456 12652 70496
rect 12692 70456 12693 70496
rect 12651 70447 12693 70456
rect 12844 70244 12884 70615
rect 12748 70204 12884 70244
rect 12212 69952 12308 69992
rect 12172 69943 12212 69952
rect 11979 69740 12021 69749
rect 11979 69700 11980 69740
rect 12020 69700 12021 69740
rect 11979 69691 12021 69700
rect 11979 67724 12021 67733
rect 11979 67684 11980 67724
rect 12020 67684 12021 67724
rect 11979 67675 12021 67684
rect 11980 66968 12020 67675
rect 11980 66919 12020 66928
rect 12076 67640 12116 69943
rect 12171 69740 12213 69749
rect 12171 69700 12172 69740
rect 12212 69700 12213 69740
rect 12171 69691 12213 69700
rect 12076 66893 12116 67600
rect 12075 66884 12117 66893
rect 12075 66844 12076 66884
rect 12116 66844 12117 66884
rect 12075 66835 12117 66844
rect 12076 66750 12116 66835
rect 12172 66632 12212 69691
rect 12268 66977 12308 69952
rect 12652 69978 12692 69987
rect 12652 69404 12692 69938
rect 12652 69355 12692 69364
rect 12459 69152 12501 69161
rect 12459 69112 12460 69152
rect 12500 69112 12501 69152
rect 12459 69103 12501 69112
rect 12363 68228 12405 68237
rect 12363 68188 12364 68228
rect 12404 68188 12405 68228
rect 12363 68179 12405 68188
rect 12364 68094 12404 68179
rect 12363 67976 12405 67985
rect 12363 67936 12364 67976
rect 12404 67936 12405 67976
rect 12363 67927 12405 67936
rect 12364 67733 12404 67927
rect 12363 67724 12405 67733
rect 12363 67684 12364 67724
rect 12404 67684 12405 67724
rect 12363 67675 12405 67684
rect 12267 66968 12309 66977
rect 12267 66928 12268 66968
rect 12308 66928 12309 66968
rect 12267 66919 12309 66928
rect 12076 66592 12212 66632
rect 12076 64616 12116 66592
rect 12171 65456 12213 65465
rect 12268 65456 12308 66919
rect 12364 66548 12404 67675
rect 12460 66800 12500 69103
rect 12555 68732 12597 68741
rect 12555 68692 12556 68732
rect 12596 68692 12597 68732
rect 12555 68683 12597 68692
rect 12556 68480 12596 68683
rect 12556 67985 12596 68440
rect 12555 67976 12597 67985
rect 12555 67936 12556 67976
rect 12596 67936 12597 67976
rect 12555 67927 12597 67936
rect 12556 67640 12596 67649
rect 12556 66977 12596 67600
rect 12748 67388 12788 70204
rect 12844 70076 12884 70085
rect 12844 69245 12884 70036
rect 12843 69236 12885 69245
rect 12843 69196 12844 69236
rect 12884 69196 12885 69236
rect 12843 69187 12885 69196
rect 12652 67348 12788 67388
rect 12555 66968 12597 66977
rect 12555 66928 12556 66968
rect 12596 66928 12597 66968
rect 12555 66919 12597 66928
rect 12460 66760 12596 66800
rect 12459 66548 12501 66557
rect 12364 66508 12460 66548
rect 12500 66508 12501 66548
rect 12459 66499 12501 66508
rect 12363 66380 12405 66389
rect 12363 66340 12364 66380
rect 12404 66340 12405 66380
rect 12363 66331 12405 66340
rect 12364 65717 12404 66331
rect 12460 66128 12500 66499
rect 12460 66079 12500 66088
rect 12363 65708 12405 65717
rect 12363 65668 12364 65708
rect 12404 65668 12405 65708
rect 12363 65659 12405 65668
rect 12171 65416 12172 65456
rect 12212 65416 12308 65456
rect 12171 65407 12213 65416
rect 12172 65322 12212 65407
rect 11884 64492 12020 64532
rect 11787 64364 11829 64373
rect 11787 64324 11788 64364
rect 11828 64324 11829 64364
rect 11787 64315 11829 64324
rect 11499 64280 11541 64289
rect 11499 64240 11500 64280
rect 11540 64240 11541 64280
rect 11499 64231 11541 64240
rect 11499 64112 11541 64121
rect 11499 64072 11500 64112
rect 11540 64072 11541 64112
rect 11499 64063 11541 64072
rect 11500 63356 11540 64063
rect 11595 63944 11637 63953
rect 11595 63904 11596 63944
rect 11636 63904 11637 63944
rect 11980 63944 12020 64492
rect 12076 64121 12116 64576
rect 12364 64280 12404 65659
rect 12268 64240 12404 64280
rect 12459 64280 12501 64289
rect 12459 64240 12460 64280
rect 12500 64240 12501 64280
rect 12075 64112 12117 64121
rect 12075 64072 12076 64112
rect 12116 64072 12117 64112
rect 12075 64063 12117 64072
rect 12268 63944 12308 64240
rect 12459 64231 12501 64240
rect 12363 64112 12405 64121
rect 12363 64072 12364 64112
rect 12404 64072 12405 64112
rect 12363 64063 12405 64072
rect 11980 63904 12116 63944
rect 11595 63895 11637 63904
rect 11596 63533 11636 63895
rect 11788 63692 11828 63701
rect 11595 63524 11637 63533
rect 11595 63484 11596 63524
rect 11636 63484 11637 63524
rect 11595 63475 11637 63484
rect 11500 63316 11732 63356
rect 11692 63020 11732 63316
rect 11788 63123 11828 63652
rect 11883 63356 11925 63365
rect 11883 63316 11884 63356
rect 11924 63316 11925 63356
rect 11883 63307 11925 63316
rect 11884 63113 11924 63307
rect 11788 63074 11828 63083
rect 11883 63104 11925 63113
rect 11883 63064 11884 63104
rect 11924 63064 11925 63104
rect 11883 63055 11925 63064
rect 11692 62980 11828 63020
rect 11500 62936 11540 62945
rect 11540 62896 11732 62936
rect 11500 62887 11540 62896
rect 11499 62768 11541 62777
rect 11499 62728 11500 62768
rect 11540 62728 11541 62768
rect 11499 62719 11541 62728
rect 11403 61256 11445 61265
rect 11403 61216 11404 61256
rect 11444 61216 11445 61256
rect 11403 61207 11445 61216
rect 11212 59284 11348 59324
rect 11019 59240 11061 59249
rect 11212 59240 11252 59284
rect 11500 59240 11540 62719
rect 11596 60920 11636 60929
rect 11596 60257 11636 60880
rect 11595 60248 11637 60257
rect 11595 60208 11596 60248
rect 11636 60208 11637 60248
rect 11595 60199 11637 60208
rect 11596 60080 11636 60091
rect 11596 60005 11636 60040
rect 11595 59996 11637 60005
rect 11595 59956 11596 59996
rect 11636 59956 11637 59996
rect 11595 59947 11637 59956
rect 11019 59200 11020 59240
rect 11060 59200 11061 59240
rect 11019 59191 11061 59200
rect 11116 59200 11252 59240
rect 11308 59200 11540 59240
rect 11596 59394 11636 59403
rect 11020 58829 11060 59191
rect 11019 58820 11061 58829
rect 11019 58780 11020 58820
rect 11060 58780 11061 58820
rect 11019 58771 11061 58780
rect 11019 57224 11061 57233
rect 11019 57184 11020 57224
rect 11060 57184 11061 57224
rect 11019 57175 11061 57184
rect 11020 57065 11060 57175
rect 11019 57056 11061 57065
rect 11019 57016 11020 57056
rect 11060 57016 11061 57056
rect 11019 57007 11061 57016
rect 11020 56922 11060 57007
rect 10828 56176 10964 56216
rect 10539 55712 10581 55721
rect 10539 55672 10540 55712
rect 10580 55672 10581 55712
rect 10539 55663 10581 55672
rect 10444 52144 10772 52184
rect 10539 52016 10581 52025
rect 10539 51976 10540 52016
rect 10580 51976 10581 52016
rect 10539 51967 10581 51976
rect 10540 51848 10580 51967
rect 10540 51799 10580 51808
rect 10635 51848 10677 51857
rect 10635 51808 10636 51848
rect 10676 51808 10677 51848
rect 10635 51799 10677 51808
rect 10443 51764 10485 51773
rect 10443 51724 10444 51764
rect 10484 51724 10485 51764
rect 10443 51715 10485 51724
rect 10444 51630 10484 51715
rect 10348 51136 10484 51176
rect 10348 51008 10388 51019
rect 10348 50933 10388 50968
rect 10347 50924 10389 50933
rect 10347 50884 10348 50924
rect 10388 50884 10389 50924
rect 10347 50875 10389 50884
rect 10347 50336 10389 50345
rect 10347 50296 10348 50336
rect 10388 50296 10389 50336
rect 10347 50287 10389 50296
rect 10348 50202 10388 50287
rect 10444 49673 10484 51136
rect 10636 50597 10676 51799
rect 10635 50588 10677 50597
rect 10635 50548 10636 50588
rect 10676 50548 10677 50588
rect 10635 50539 10677 50548
rect 10443 49664 10485 49673
rect 10443 49624 10444 49664
rect 10484 49624 10485 49664
rect 10443 49615 10485 49624
rect 10540 49505 10580 49591
rect 10348 49496 10388 49505
rect 10252 49456 10348 49496
rect 10348 49447 10388 49456
rect 10444 49496 10484 49505
rect 10155 49412 10197 49421
rect 10155 49372 10156 49412
rect 10196 49372 10197 49412
rect 10155 49363 10197 49372
rect 10156 49278 10196 49363
rect 10060 49120 10292 49160
rect 10060 48824 10100 48833
rect 9964 48784 10060 48824
rect 9676 48775 9716 48784
rect 10060 48775 10100 48784
rect 10156 48824 10196 48833
rect 9867 47732 9909 47741
rect 9867 47692 9868 47732
rect 9908 47692 9909 47732
rect 9867 47683 9909 47692
rect 9772 47312 9812 47321
rect 9676 47272 9772 47312
rect 9676 46733 9716 47272
rect 9772 47263 9812 47272
rect 9771 46892 9813 46901
rect 9771 46852 9772 46892
rect 9812 46852 9813 46892
rect 9771 46843 9813 46852
rect 9675 46724 9717 46733
rect 9675 46684 9676 46724
rect 9716 46684 9717 46724
rect 9675 46675 9717 46684
rect 9772 46556 9812 46843
rect 9724 46516 9812 46556
rect 9724 46514 9764 46516
rect 9724 46465 9764 46474
rect 9868 46388 9908 47683
rect 10156 47321 10196 48784
rect 10252 48824 10292 49120
rect 10348 48992 10388 49001
rect 10444 48992 10484 49456
rect 10539 49504 10581 49505
rect 10539 49456 10540 49504
rect 10580 49456 10581 49504
rect 10539 49447 10581 49456
rect 10636 49328 10676 49337
rect 10636 49085 10676 49288
rect 10635 49076 10677 49085
rect 10635 49036 10636 49076
rect 10676 49036 10677 49076
rect 10635 49027 10677 49036
rect 10388 48952 10484 48992
rect 10348 48943 10388 48952
rect 10636 48833 10676 48918
rect 10252 48775 10292 48784
rect 10347 48824 10389 48833
rect 10347 48784 10348 48824
rect 10388 48784 10389 48824
rect 10347 48775 10389 48784
rect 10635 48824 10677 48833
rect 10635 48784 10636 48824
rect 10676 48784 10677 48824
rect 10635 48775 10677 48784
rect 10251 48320 10293 48329
rect 10251 48280 10252 48320
rect 10292 48280 10293 48320
rect 10251 48271 10293 48280
rect 10252 48026 10292 48271
rect 10252 47977 10292 47986
rect 10348 47900 10388 48775
rect 10732 48656 10772 52144
rect 10828 51689 10868 56176
rect 11116 56132 11156 59200
rect 11308 59156 11348 59200
rect 11212 59116 11348 59156
rect 11212 58577 11252 59116
rect 11307 58904 11349 58913
rect 11307 58864 11308 58904
rect 11348 58864 11349 58904
rect 11307 58855 11349 58864
rect 11211 58568 11253 58577
rect 11211 58528 11212 58568
rect 11252 58528 11253 58568
rect 11211 58519 11253 58528
rect 11308 58568 11348 58855
rect 11403 58820 11445 58829
rect 11403 58780 11404 58820
rect 11444 58780 11445 58820
rect 11403 58771 11445 58780
rect 11500 58820 11540 58829
rect 11596 58820 11636 59354
rect 11540 58780 11636 58820
rect 11500 58771 11540 58780
rect 11404 58652 11444 58771
rect 11404 58612 11540 58652
rect 11308 58519 11348 58528
rect 11403 57980 11445 57989
rect 11403 57940 11404 57980
rect 11444 57940 11445 57980
rect 11403 57931 11445 57940
rect 11404 57896 11444 57931
rect 11404 57845 11444 57856
rect 11500 57728 11540 58612
rect 11404 57688 11540 57728
rect 11307 57476 11349 57485
rect 11307 57436 11308 57476
rect 11348 57436 11349 57476
rect 11307 57427 11349 57436
rect 11212 56888 11252 56897
rect 11212 56477 11252 56848
rect 11308 56729 11348 57427
rect 11404 56972 11444 57688
rect 11596 57644 11636 57653
rect 11500 57604 11596 57644
rect 11500 57075 11540 57604
rect 11596 57595 11636 57604
rect 11500 57026 11540 57035
rect 11596 57056 11636 57065
rect 11596 56972 11636 57016
rect 11404 56932 11636 56972
rect 11500 56813 11540 56932
rect 11499 56804 11541 56813
rect 11499 56764 11500 56804
rect 11540 56764 11541 56804
rect 11499 56755 11541 56764
rect 11307 56720 11349 56729
rect 11307 56680 11308 56720
rect 11348 56680 11349 56720
rect 11307 56671 11349 56680
rect 11595 56720 11637 56729
rect 11595 56680 11596 56720
rect 11636 56680 11637 56720
rect 11595 56671 11637 56680
rect 11403 56636 11445 56645
rect 11403 56596 11404 56636
rect 11444 56596 11445 56636
rect 11403 56587 11445 56596
rect 11307 56552 11349 56561
rect 11307 56512 11308 56552
rect 11348 56512 11349 56552
rect 11307 56503 11349 56512
rect 11211 56468 11253 56477
rect 11211 56428 11212 56468
rect 11252 56428 11253 56468
rect 11211 56419 11253 56428
rect 11308 56384 11348 56503
rect 11308 56335 11348 56344
rect 11404 56384 11444 56587
rect 11308 56225 11348 56244
rect 11307 56216 11349 56225
rect 11404 56216 11444 56344
rect 11307 56176 11308 56216
rect 11348 56176 11444 56216
rect 11499 56216 11541 56225
rect 11499 56176 11500 56216
rect 11540 56176 11541 56216
rect 11307 56167 11349 56176
rect 11499 56167 11541 56176
rect 10924 56092 11156 56132
rect 10827 51680 10869 51689
rect 10827 51640 10828 51680
rect 10868 51640 10869 51680
rect 10827 51631 10869 51640
rect 10827 50336 10869 50345
rect 10827 50296 10828 50336
rect 10868 50296 10869 50336
rect 10827 50287 10869 50296
rect 10828 50202 10868 50287
rect 10924 49664 10964 56092
rect 11500 56048 11540 56167
rect 11404 56008 11540 56048
rect 11596 56048 11636 56671
rect 11692 56225 11732 62896
rect 11788 61433 11828 62980
rect 11884 62970 11924 63055
rect 12076 62861 12116 63904
rect 12172 63904 12268 63944
rect 11883 62852 11925 62861
rect 11883 62812 11884 62852
rect 11924 62812 11925 62852
rect 11883 62803 11925 62812
rect 12075 62852 12117 62861
rect 12075 62812 12076 62852
rect 12116 62812 12117 62852
rect 12075 62803 12117 62812
rect 11787 61424 11829 61433
rect 11787 61384 11788 61424
rect 11828 61384 11829 61424
rect 11787 61375 11829 61384
rect 11787 61172 11829 61181
rect 11787 61132 11788 61172
rect 11828 61132 11829 61172
rect 11787 61123 11829 61132
rect 11788 60005 11828 61123
rect 11787 59996 11829 60005
rect 11787 59956 11788 59996
rect 11828 59956 11829 59996
rect 11787 59947 11829 59956
rect 11787 59492 11829 59501
rect 11787 59452 11788 59492
rect 11828 59452 11829 59492
rect 11787 59443 11829 59452
rect 11788 59358 11828 59443
rect 11884 58064 11924 62803
rect 12172 62777 12212 63904
rect 12268 63895 12308 63904
rect 12364 63440 12404 64063
rect 12268 63400 12404 63440
rect 12268 63188 12308 63400
rect 12363 63272 12405 63281
rect 12363 63232 12364 63272
rect 12404 63232 12405 63272
rect 12363 63223 12405 63232
rect 12171 62768 12213 62777
rect 12171 62728 12172 62768
rect 12212 62728 12213 62768
rect 12171 62719 12213 62728
rect 12171 62180 12213 62189
rect 12076 62140 12172 62180
rect 12212 62140 12213 62180
rect 11979 61760 12021 61769
rect 11979 61720 11980 61760
rect 12020 61720 12021 61760
rect 11979 61711 12021 61720
rect 11980 59744 12020 61711
rect 12076 60915 12116 62140
rect 12171 62131 12213 62140
rect 12268 61844 12308 63148
rect 12364 63188 12404 63223
rect 12364 63137 12404 63148
rect 12460 63029 12500 64231
rect 12459 63020 12501 63029
rect 12459 62980 12460 63020
rect 12500 62980 12501 63020
rect 12459 62971 12501 62980
rect 12364 62432 12404 62443
rect 12556 62432 12596 66760
rect 12652 66641 12692 67348
rect 12747 67052 12789 67061
rect 12747 67012 12748 67052
rect 12788 67012 12789 67052
rect 12747 67003 12789 67012
rect 12651 66632 12693 66641
rect 12651 66592 12652 66632
rect 12692 66592 12693 66632
rect 12651 66583 12693 66592
rect 12652 65960 12692 65969
rect 12652 65451 12692 65920
rect 12748 65540 12788 67003
rect 12844 66800 12884 69187
rect 12940 67145 12980 71464
rect 13036 70841 13076 71875
rect 13227 71840 13269 71849
rect 13227 71800 13228 71840
rect 13268 71800 13269 71840
rect 13324 71840 13364 71968
rect 13419 72008 13461 72017
rect 13419 71968 13420 72008
rect 13460 71968 13461 72008
rect 13419 71959 13461 71968
rect 13419 71840 13461 71849
rect 13324 71800 13420 71840
rect 13460 71800 13461 71840
rect 13227 71791 13269 71800
rect 13419 71791 13461 71800
rect 13131 71504 13173 71513
rect 13131 71464 13132 71504
rect 13172 71464 13173 71504
rect 13131 71455 13173 71464
rect 13035 70832 13077 70841
rect 13035 70792 13036 70832
rect 13076 70792 13077 70832
rect 13035 70783 13077 70792
rect 13036 70496 13076 70783
rect 13132 70664 13172 71455
rect 13132 70615 13172 70624
rect 13036 70456 13172 70496
rect 13035 68228 13077 68237
rect 13035 68188 13036 68228
rect 13076 68188 13077 68228
rect 13035 68179 13077 68188
rect 13036 67654 13076 68179
rect 13132 68144 13172 70456
rect 13228 70160 13268 71791
rect 13419 71672 13461 71681
rect 13419 71632 13420 71672
rect 13460 71632 13461 71672
rect 13419 71623 13461 71632
rect 13323 71504 13365 71513
rect 13323 71464 13324 71504
rect 13364 71464 13365 71504
rect 13323 71455 13365 71464
rect 13324 71009 13364 71455
rect 13323 71000 13365 71009
rect 13323 70960 13324 71000
rect 13364 70960 13365 71000
rect 13323 70951 13365 70960
rect 13420 70664 13460 71623
rect 13228 70120 13364 70160
rect 13227 69992 13269 70001
rect 13227 69952 13228 69992
rect 13268 69952 13269 69992
rect 13227 69943 13269 69952
rect 13228 69858 13268 69943
rect 13227 69320 13269 69329
rect 13227 69280 13228 69320
rect 13268 69280 13269 69320
rect 13227 69271 13269 69280
rect 13228 69152 13268 69271
rect 13228 68573 13268 69112
rect 13227 68564 13269 68573
rect 13227 68524 13228 68564
rect 13268 68524 13269 68564
rect 13227 68515 13269 68524
rect 13324 68321 13364 70120
rect 13420 70001 13460 70624
rect 13419 69992 13461 70001
rect 13419 69952 13420 69992
rect 13460 69952 13461 69992
rect 13419 69943 13461 69952
rect 13420 69077 13460 69943
rect 13516 69824 13556 72136
rect 13804 72176 13844 72967
rect 13996 72344 14036 72976
rect 13804 72127 13844 72136
rect 13900 72304 14036 72344
rect 13803 72008 13845 72017
rect 13803 71968 13804 72008
rect 13844 71968 13845 72008
rect 13803 71959 13845 71968
rect 13804 71499 13844 71959
rect 13804 71450 13844 71459
rect 13516 69784 13748 69824
rect 13419 69068 13461 69077
rect 13419 69028 13420 69068
rect 13460 69028 13461 69068
rect 13419 69019 13461 69028
rect 13323 68312 13365 68321
rect 13323 68272 13324 68312
rect 13364 68272 13365 68312
rect 13323 68263 13365 68272
rect 13132 68104 13556 68144
rect 13036 67605 13076 67614
rect 13227 67472 13269 67481
rect 13420 67472 13460 67481
rect 13227 67432 13228 67472
rect 13268 67432 13269 67472
rect 13227 67423 13269 67432
rect 13324 67432 13420 67472
rect 13228 67338 13268 67423
rect 13324 67220 13364 67432
rect 13420 67423 13460 67432
rect 13132 67180 13364 67220
rect 12939 67136 12981 67145
rect 12939 67096 12940 67136
rect 12980 67096 12981 67136
rect 12939 67087 12981 67096
rect 13132 66968 13172 67180
rect 13084 66958 13172 66968
rect 13124 66928 13172 66958
rect 13228 67052 13268 67061
rect 13084 66909 13124 66918
rect 12844 66760 13172 66800
rect 13035 66632 13077 66641
rect 13035 66592 13036 66632
rect 13076 66592 13077 66632
rect 13035 66583 13077 66592
rect 12844 66128 12884 66137
rect 12844 65717 12884 66088
rect 12843 65708 12885 65717
rect 12843 65668 12844 65708
rect 12884 65668 12885 65708
rect 12843 65659 12885 65668
rect 12844 65540 12884 65549
rect 12748 65500 12844 65540
rect 12652 65402 12692 65411
rect 12652 64616 12692 64625
rect 12692 64576 12788 64616
rect 12652 64567 12692 64576
rect 12748 64373 12788 64576
rect 12747 64364 12789 64373
rect 12747 64324 12748 64364
rect 12788 64324 12789 64364
rect 12747 64315 12789 64324
rect 12844 64289 12884 65500
rect 13036 65045 13076 66583
rect 13035 65036 13077 65045
rect 13035 64996 13036 65036
rect 13076 64996 13077 65036
rect 13035 64987 13077 64996
rect 12651 64280 12693 64289
rect 12651 64240 12652 64280
rect 12692 64240 12693 64280
rect 12651 64231 12693 64240
rect 12843 64280 12885 64289
rect 13036 64280 13076 64987
rect 12843 64240 12844 64280
rect 12884 64240 12885 64280
rect 12843 64231 12885 64240
rect 12940 64240 13076 64280
rect 12364 62357 12404 62392
rect 12460 62392 12596 62432
rect 12363 62348 12405 62357
rect 12363 62308 12364 62348
rect 12404 62308 12405 62348
rect 12363 62299 12405 62308
rect 12268 61804 12404 61844
rect 12268 61601 12308 61686
rect 12267 61592 12309 61601
rect 12267 61552 12268 61592
rect 12308 61552 12309 61592
rect 12267 61543 12309 61552
rect 12171 61256 12213 61265
rect 12171 61216 12172 61256
rect 12212 61216 12213 61256
rect 12171 61207 12213 61216
rect 12076 60866 12116 60875
rect 12172 60164 12212 61207
rect 12364 61088 12404 61804
rect 12460 61592 12500 62392
rect 12556 62189 12596 62274
rect 12555 62180 12597 62189
rect 12555 62140 12556 62180
rect 12596 62140 12597 62180
rect 12555 62131 12597 62140
rect 12460 61552 12596 61592
rect 12460 61424 12500 61433
rect 12460 61265 12500 61384
rect 12459 61256 12501 61265
rect 12459 61216 12460 61256
rect 12500 61216 12501 61256
rect 12459 61207 12501 61216
rect 12364 61048 12500 61088
rect 12268 61004 12308 61013
rect 12308 60964 12404 61004
rect 12268 60955 12308 60964
rect 12267 60416 12309 60425
rect 12267 60376 12268 60416
rect 12308 60376 12309 60416
rect 12267 60367 12309 60376
rect 12124 60124 12212 60164
rect 12124 60122 12164 60124
rect 12124 60073 12164 60082
rect 12268 59996 12308 60367
rect 12268 59947 12308 59956
rect 12364 59753 12404 60964
rect 12363 59744 12405 59753
rect 11980 59704 12212 59744
rect 11979 59576 12021 59585
rect 11979 59536 11980 59576
rect 12020 59536 12021 59576
rect 11979 59527 12021 59536
rect 11980 59249 12020 59527
rect 11979 59240 12021 59249
rect 11979 59200 11980 59240
rect 12020 59200 12021 59240
rect 11979 59191 12021 59200
rect 11788 58024 11924 58064
rect 11788 57140 11828 58024
rect 11884 57896 11924 57905
rect 11980 57896 12020 59191
rect 11924 57856 12020 57896
rect 11884 57847 11924 57856
rect 11980 57140 12020 57149
rect 11788 57100 11980 57140
rect 11788 56561 11828 57100
rect 11980 57091 12020 57100
rect 12076 57056 12116 57067
rect 12076 56981 12116 57016
rect 12075 56972 12117 56981
rect 12075 56932 12076 56972
rect 12116 56932 12117 56972
rect 12075 56923 12117 56932
rect 11979 56804 12021 56813
rect 11979 56764 11980 56804
rect 12020 56764 12021 56804
rect 11979 56755 12021 56764
rect 11787 56552 11829 56561
rect 11787 56512 11788 56552
rect 11828 56512 11829 56552
rect 11787 56503 11829 56512
rect 11788 56384 11828 56393
rect 11691 56216 11733 56225
rect 11691 56176 11692 56216
rect 11732 56176 11733 56216
rect 11691 56167 11733 56176
rect 11788 56132 11828 56344
rect 11883 56384 11925 56393
rect 11883 56344 11884 56384
rect 11924 56344 11925 56384
rect 11883 56335 11925 56344
rect 11884 56250 11924 56335
rect 11980 56132 12020 56755
rect 11788 56092 12020 56132
rect 12172 56048 12212 59704
rect 12363 59704 12364 59744
rect 12404 59704 12405 59744
rect 12363 59695 12405 59704
rect 12460 59492 12500 61048
rect 12556 60089 12596 61552
rect 12652 60341 12692 64231
rect 12843 64028 12885 64037
rect 12843 63988 12844 64028
rect 12884 63988 12885 64028
rect 12843 63979 12885 63988
rect 12747 63776 12789 63785
rect 12747 63736 12748 63776
rect 12788 63736 12789 63776
rect 12747 63727 12789 63736
rect 12748 61097 12788 63727
rect 12844 63104 12884 63979
rect 12844 61181 12884 63064
rect 12940 62105 12980 64240
rect 13036 62180 13076 62189
rect 12939 62096 12981 62105
rect 12939 62056 12940 62096
rect 12980 62056 12981 62096
rect 12939 62047 12981 62056
rect 13036 61853 13076 62140
rect 13035 61844 13077 61853
rect 13035 61804 13036 61844
rect 13076 61804 13077 61844
rect 13035 61795 13077 61804
rect 12843 61172 12885 61181
rect 12843 61132 12844 61172
rect 12884 61132 12885 61172
rect 12843 61123 12885 61132
rect 12747 61088 12789 61097
rect 12747 61048 12748 61088
rect 12788 61048 12789 61088
rect 12747 61039 12789 61048
rect 12748 60920 12788 61039
rect 12844 60920 12884 60929
rect 12748 60880 12844 60920
rect 12837 60875 12884 60880
rect 12844 60871 12884 60875
rect 13035 60836 13077 60845
rect 12940 60796 13036 60836
rect 13076 60796 13077 60836
rect 12940 60752 12980 60796
rect 13035 60787 13077 60796
rect 12748 60712 12980 60752
rect 12651 60332 12693 60341
rect 12651 60292 12652 60332
rect 12692 60292 12693 60332
rect 12651 60283 12693 60292
rect 12652 60173 12692 60204
rect 12651 60164 12693 60173
rect 12651 60124 12652 60164
rect 12692 60124 12693 60164
rect 12651 60115 12693 60124
rect 12555 60080 12597 60089
rect 12555 60040 12556 60080
rect 12596 60040 12597 60080
rect 12555 60031 12597 60040
rect 12652 60080 12692 60115
rect 12652 59921 12692 60040
rect 12651 59912 12693 59921
rect 12651 59872 12652 59912
rect 12692 59872 12693 59912
rect 12651 59863 12693 59872
rect 12748 59576 12788 60712
rect 13035 60668 13077 60677
rect 13035 60628 13036 60668
rect 13076 60628 13077 60668
rect 13035 60619 13077 60628
rect 13036 59585 13076 60619
rect 12748 59527 12788 59536
rect 12843 59576 12885 59585
rect 12843 59536 12844 59576
rect 12884 59536 12885 59576
rect 12843 59527 12885 59536
rect 13035 59576 13077 59585
rect 13035 59536 13036 59576
rect 13076 59536 13077 59576
rect 13035 59527 13077 59536
rect 12268 59452 12500 59492
rect 12268 57233 12308 59452
rect 12556 59408 12596 59417
rect 12460 59368 12556 59408
rect 12363 58568 12405 58577
rect 12363 58528 12364 58568
rect 12404 58528 12405 58568
rect 12363 58519 12405 58528
rect 12364 57821 12404 58519
rect 12363 57812 12405 57821
rect 12363 57772 12364 57812
rect 12404 57772 12405 57812
rect 12363 57763 12405 57772
rect 12267 57224 12309 57233
rect 12267 57184 12268 57224
rect 12308 57184 12309 57224
rect 12267 57175 12309 57184
rect 12268 56981 12308 57175
rect 12267 56972 12309 56981
rect 12267 56932 12268 56972
rect 12308 56932 12309 56972
rect 12267 56923 12309 56932
rect 12267 56720 12309 56729
rect 12267 56680 12268 56720
rect 12308 56680 12309 56720
rect 12267 56671 12309 56680
rect 11596 56008 11732 56048
rect 11115 55964 11157 55973
rect 11115 55924 11116 55964
rect 11156 55924 11157 55964
rect 11115 55915 11157 55924
rect 11019 55712 11061 55721
rect 11019 55672 11020 55712
rect 11060 55672 11061 55712
rect 11019 55663 11061 55672
rect 11020 52949 11060 55663
rect 11116 53957 11156 55915
rect 11307 54956 11349 54965
rect 11307 54916 11308 54956
rect 11348 54916 11349 54956
rect 11307 54907 11349 54916
rect 11308 54872 11348 54907
rect 11308 54209 11348 54832
rect 11307 54200 11349 54209
rect 11307 54160 11308 54200
rect 11348 54160 11349 54200
rect 11307 54151 11349 54160
rect 11115 53948 11157 53957
rect 11115 53908 11116 53948
rect 11156 53908 11157 53948
rect 11115 53899 11157 53908
rect 11212 53864 11252 53873
rect 11115 53696 11157 53705
rect 11115 53656 11116 53696
rect 11156 53656 11157 53696
rect 11115 53647 11157 53656
rect 11116 53360 11156 53647
rect 11212 53537 11252 53824
rect 11308 53705 11348 54151
rect 11404 54116 11444 56008
rect 11596 55553 11636 55638
rect 11500 55544 11540 55553
rect 11500 55040 11540 55504
rect 11595 55544 11637 55553
rect 11595 55504 11596 55544
rect 11636 55504 11637 55544
rect 11595 55495 11637 55504
rect 11500 54991 11540 55000
rect 11404 54067 11444 54076
rect 11595 54116 11637 54125
rect 11595 54076 11596 54116
rect 11636 54076 11637 54116
rect 11595 54067 11637 54076
rect 11596 54032 11636 54067
rect 11596 53981 11636 53992
rect 11403 53948 11445 53957
rect 11403 53908 11404 53948
rect 11444 53908 11445 53948
rect 11403 53899 11445 53908
rect 11404 53789 11444 53899
rect 11403 53780 11445 53789
rect 11403 53740 11404 53780
rect 11444 53740 11445 53780
rect 11403 53731 11445 53740
rect 11307 53696 11349 53705
rect 11307 53656 11308 53696
rect 11348 53656 11349 53696
rect 11307 53647 11349 53656
rect 11211 53528 11253 53537
rect 11211 53488 11212 53528
rect 11252 53488 11253 53528
rect 11692 53528 11732 56008
rect 11980 56008 12212 56048
rect 11787 55964 11829 55973
rect 11787 55924 11788 55964
rect 11828 55924 11829 55964
rect 11787 55915 11829 55924
rect 11788 55553 11828 55915
rect 11787 55544 11829 55553
rect 11787 55504 11788 55544
rect 11828 55504 11829 55544
rect 11787 55495 11829 55504
rect 11980 55544 12020 56008
rect 12171 55628 12213 55637
rect 12171 55588 12172 55628
rect 12212 55588 12213 55628
rect 12171 55579 12213 55588
rect 11980 55495 12020 55504
rect 12076 55544 12116 55553
rect 11788 54872 11828 55495
rect 11788 54823 11828 54832
rect 12076 54452 12116 55504
rect 11884 54412 12116 54452
rect 11692 53488 11828 53528
rect 11211 53479 11253 53488
rect 11320 53453 11360 53472
rect 11308 53444 11360 53453
rect 11348 53404 11444 53444
rect 11308 53395 11348 53404
rect 11404 53360 11444 53404
rect 11596 53360 11636 53369
rect 11404 53320 11596 53360
rect 11116 53311 11156 53320
rect 11596 53311 11636 53320
rect 11692 53360 11732 53369
rect 11211 53276 11253 53285
rect 11211 53236 11212 53276
rect 11252 53236 11253 53276
rect 11211 53227 11253 53236
rect 11019 52940 11061 52949
rect 11019 52900 11020 52940
rect 11060 52900 11061 52940
rect 11019 52891 11061 52900
rect 11115 52688 11157 52697
rect 11115 52648 11116 52688
rect 11156 52648 11157 52688
rect 11115 52639 11157 52648
rect 11019 52520 11061 52529
rect 11019 52480 11020 52520
rect 11060 52480 11061 52520
rect 11019 52471 11061 52480
rect 11020 51857 11060 52471
rect 11116 51941 11156 52639
rect 11115 51932 11157 51941
rect 11115 51892 11116 51932
rect 11156 51892 11157 51932
rect 11115 51883 11157 51892
rect 11019 51848 11061 51857
rect 11019 51808 11020 51848
rect 11060 51808 11061 51848
rect 11019 51799 11061 51808
rect 11020 51714 11060 51799
rect 11116 50345 11156 51883
rect 11212 50933 11252 53227
rect 11307 53192 11349 53201
rect 11307 53152 11308 53192
rect 11348 53152 11349 53192
rect 11307 53143 11349 53152
rect 11211 50924 11253 50933
rect 11211 50884 11212 50924
rect 11252 50884 11253 50924
rect 11211 50875 11253 50884
rect 11211 50420 11253 50429
rect 11211 50380 11212 50420
rect 11252 50380 11253 50420
rect 11211 50371 11253 50380
rect 11115 50336 11157 50345
rect 11115 50296 11116 50336
rect 11156 50296 11157 50336
rect 11115 50287 11157 50296
rect 10924 49624 11156 49664
rect 10828 49496 10868 49507
rect 10828 49421 10868 49456
rect 11019 49496 11061 49505
rect 11019 49456 11020 49496
rect 11060 49456 11061 49496
rect 11019 49447 11061 49456
rect 10827 49412 10869 49421
rect 10827 49372 10828 49412
rect 10868 49372 10869 49412
rect 10827 49363 10869 49372
rect 11020 49362 11060 49447
rect 10252 47860 10388 47900
rect 10540 48616 10772 48656
rect 10924 49328 10964 49337
rect 10155 47312 10197 47321
rect 10155 47272 10156 47312
rect 10196 47272 10197 47312
rect 10155 47263 10197 47272
rect 10059 47144 10101 47153
rect 10059 47104 10060 47144
rect 10100 47104 10101 47144
rect 10059 47095 10101 47104
rect 9964 47060 10004 47069
rect 9964 46901 10004 47020
rect 9963 46892 10005 46901
rect 9963 46852 9964 46892
rect 10004 46852 10005 46892
rect 9963 46843 10005 46852
rect 9963 46724 10005 46733
rect 9963 46684 9964 46724
rect 10004 46684 10005 46724
rect 9963 46675 10005 46684
rect 9868 46339 9908 46348
rect 9964 45800 10004 46675
rect 9964 45305 10004 45760
rect 9963 45296 10005 45305
rect 9963 45256 9964 45296
rect 10004 45256 10005 45296
rect 9963 45247 10005 45256
rect 9580 45172 9716 45212
rect 8908 44911 8948 44920
rect 9004 45088 9524 45128
rect 8619 44876 8661 44885
rect 8619 44836 8620 44876
rect 8660 44836 8661 44876
rect 8619 44827 8661 44836
rect 8523 43196 8565 43205
rect 8523 43156 8524 43196
rect 8564 43156 8565 43196
rect 8523 43147 8565 43156
rect 8427 43112 8469 43121
rect 8427 43072 8428 43112
rect 8468 43072 8469 43112
rect 8427 43063 8469 43072
rect 8524 42944 8564 42953
rect 8332 42904 8524 42944
rect 8524 42895 8564 42904
rect 8044 42643 8084 42652
rect 8140 42776 8180 42785
rect 7948 42559 7988 42568
rect 7851 42272 7893 42281
rect 8140 42272 8180 42736
rect 8332 42776 8372 42785
rect 8235 42440 8277 42449
rect 8235 42400 8236 42440
rect 8276 42400 8277 42440
rect 8332 42440 8372 42736
rect 8427 42776 8469 42785
rect 8427 42736 8428 42776
rect 8468 42736 8469 42776
rect 8427 42727 8469 42736
rect 8620 42776 8660 42785
rect 8428 42642 8468 42727
rect 8332 42400 8564 42440
rect 8235 42391 8277 42400
rect 7851 42232 7852 42272
rect 7892 42232 7893 42272
rect 7851 42223 7893 42232
rect 7948 42232 8180 42272
rect 7564 42064 7796 42104
rect 7756 41945 7796 42064
rect 7563 41936 7605 41945
rect 7563 41896 7564 41936
rect 7604 41896 7605 41936
rect 7563 41887 7605 41896
rect 7660 41936 7700 41945
rect 7467 41684 7509 41693
rect 7467 41644 7468 41684
rect 7508 41644 7509 41684
rect 7467 41635 7509 41644
rect 7564 41441 7604 41887
rect 7660 41777 7700 41896
rect 7755 41936 7797 41945
rect 7755 41896 7756 41936
rect 7796 41896 7797 41936
rect 7755 41887 7797 41896
rect 7659 41768 7701 41777
rect 7659 41728 7660 41768
rect 7700 41728 7701 41768
rect 7659 41719 7701 41728
rect 7851 41768 7893 41777
rect 7851 41728 7852 41768
rect 7892 41728 7893 41768
rect 7851 41719 7893 41728
rect 7852 41634 7892 41719
rect 7755 41600 7797 41609
rect 7755 41560 7756 41600
rect 7796 41560 7797 41600
rect 7948 41600 7988 42232
rect 8236 42197 8276 42391
rect 8427 42272 8469 42281
rect 8427 42232 8428 42272
rect 8468 42232 8469 42272
rect 8427 42223 8469 42232
rect 8235 42188 8277 42197
rect 8235 42148 8236 42188
rect 8276 42148 8277 42188
rect 8235 42139 8277 42148
rect 8043 41936 8085 41945
rect 8043 41896 8044 41936
rect 8084 41896 8085 41936
rect 8043 41887 8085 41896
rect 8140 41936 8180 41945
rect 8044 41802 8084 41887
rect 8140 41777 8180 41896
rect 8235 41852 8277 41861
rect 8235 41812 8236 41852
rect 8276 41812 8277 41852
rect 8235 41803 8277 41812
rect 8139 41768 8181 41777
rect 8139 41728 8140 41768
rect 8180 41728 8181 41768
rect 8139 41719 8181 41728
rect 8236 41718 8276 41803
rect 8332 41768 8372 41777
rect 8235 41600 8277 41609
rect 7948 41560 8180 41600
rect 7755 41551 7797 41560
rect 7371 41432 7413 41441
rect 7371 41392 7372 41432
rect 7412 41392 7413 41432
rect 7371 41383 7413 41392
rect 7563 41432 7605 41441
rect 7563 41392 7564 41432
rect 7604 41392 7605 41432
rect 7563 41383 7605 41392
rect 6988 41264 7048 41273
rect 7028 41224 7048 41264
rect 7274 41308 7316 41348
rect 6988 41215 7028 41224
rect 7274 41222 7314 41308
rect 6786 41140 6796 41170
rect 6786 41130 6836 41140
rect 7084 41180 7124 41189
rect 7274 41173 7314 41182
rect 7372 41264 7412 41273
rect 6699 41096 6741 41105
rect 6220 41056 6356 41096
rect 6316 40769 6356 41056
rect 6699 41056 6700 41096
rect 6740 41056 6741 41096
rect 6699 41047 6741 41056
rect 6507 40844 6549 40853
rect 6507 40804 6508 40844
rect 6548 40804 6549 40844
rect 6507 40795 6549 40804
rect 6315 40760 6357 40769
rect 6315 40720 6316 40760
rect 6356 40720 6357 40760
rect 6315 40711 6357 40720
rect 6220 40676 6260 40685
rect 6124 40636 6220 40676
rect 6220 40627 6260 40636
rect 6028 40592 6068 40601
rect 6068 40552 6164 40592
rect 6028 40543 6068 40552
rect 6124 40424 6164 40552
rect 6220 40424 6260 40433
rect 6124 40384 6220 40424
rect 6220 40375 6260 40384
rect 6412 40424 6452 40433
rect 6027 40340 6069 40349
rect 6027 40300 6028 40340
rect 6068 40300 6069 40340
rect 6027 40291 6069 40300
rect 5740 39964 5972 40004
rect 5740 38996 5780 39964
rect 5740 38947 5780 38956
rect 5836 38912 5876 38921
rect 5836 37820 5876 38872
rect 6028 38585 6068 40291
rect 6412 38921 6452 40384
rect 6508 40424 6548 40795
rect 6700 40592 6740 41047
rect 6786 41012 6826 41130
rect 6786 40972 6932 41012
rect 6892 40853 6932 40972
rect 6891 40844 6933 40853
rect 6891 40804 6892 40844
rect 6932 40804 6933 40844
rect 6891 40795 6933 40804
rect 6987 40676 7029 40685
rect 6987 40636 6988 40676
rect 7028 40636 7029 40676
rect 7084 40676 7124 41140
rect 7372 41105 7412 41224
rect 7371 41096 7413 41105
rect 7180 41054 7220 41063
rect 7371 41056 7372 41096
rect 7412 41056 7413 41096
rect 7371 41047 7413 41056
rect 7180 40844 7220 41014
rect 7180 40804 7508 40844
rect 7468 40685 7508 40804
rect 7180 40676 7220 40685
rect 7084 40636 7180 40676
rect 6987 40627 7029 40636
rect 7180 40627 7220 40636
rect 7467 40676 7509 40685
rect 7467 40636 7468 40676
rect 7508 40636 7509 40676
rect 7467 40627 7509 40636
rect 6796 40592 6836 40601
rect 6700 40552 6796 40592
rect 6836 40552 6932 40592
rect 6796 40543 6836 40552
rect 6892 40438 6932 40552
rect 6988 40542 7028 40627
rect 7276 40517 7316 40602
rect 7371 40592 7413 40601
rect 7371 40552 7372 40592
rect 7412 40552 7413 40592
rect 7371 40543 7413 40552
rect 7275 40508 7317 40517
rect 7275 40468 7276 40508
rect 7316 40468 7317 40508
rect 7275 40459 7317 40468
rect 7173 40441 7213 40450
rect 6508 40375 6548 40384
rect 6795 40424 6837 40433
rect 6795 40384 6796 40424
rect 6836 40384 6837 40424
rect 6892 40401 7173 40438
rect 6892 40398 7213 40401
rect 7173 40392 7213 40398
rect 6795 40375 6837 40384
rect 6796 40290 6836 40375
rect 7275 40340 7317 40349
rect 7275 40300 7276 40340
rect 7316 40300 7317 40340
rect 7275 40291 7317 40300
rect 7276 39929 7316 40291
rect 6699 39920 6741 39929
rect 6699 39880 6700 39920
rect 6740 39880 6741 39920
rect 6699 39871 6741 39880
rect 7275 39920 7317 39929
rect 7275 39880 7276 39920
rect 7316 39880 7317 39920
rect 7372 39920 7412 40543
rect 7467 40424 7509 40433
rect 7564 40424 7604 41383
rect 7756 41264 7796 41551
rect 8043 41432 8085 41441
rect 8043 41392 8044 41432
rect 8084 41392 8085 41432
rect 8043 41383 8085 41392
rect 7947 41348 7989 41357
rect 7947 41308 7948 41348
rect 7988 41308 7989 41348
rect 7947 41299 7989 41308
rect 7756 41215 7796 41224
rect 7852 41264 7892 41273
rect 7852 41096 7892 41224
rect 7948 41214 7988 41299
rect 8044 41298 8084 41383
rect 7756 41056 7892 41096
rect 7659 40508 7701 40517
rect 7659 40468 7660 40508
rect 7700 40468 7701 40508
rect 7659 40459 7701 40468
rect 7467 40384 7468 40424
rect 7508 40384 7604 40424
rect 7467 40375 7509 40384
rect 7468 40290 7508 40375
rect 7660 39929 7700 40459
rect 7756 40013 7796 41056
rect 8044 41012 8084 41021
rect 7851 40592 7893 40601
rect 7851 40552 7852 40592
rect 7892 40552 7893 40592
rect 7851 40543 7893 40552
rect 7852 40424 7892 40543
rect 7852 40375 7892 40384
rect 7947 40424 7989 40433
rect 7947 40384 7948 40424
rect 7988 40384 7989 40424
rect 8044 40424 8084 40972
rect 8140 40676 8180 41560
rect 8235 41560 8236 41600
rect 8276 41560 8277 41600
rect 8235 41551 8277 41560
rect 8140 40627 8180 40636
rect 8140 40424 8180 40433
rect 8044 40384 8140 40424
rect 8236 40424 8276 41551
rect 8332 41525 8372 41728
rect 8428 41768 8468 42223
rect 8428 41719 8468 41728
rect 8331 41516 8373 41525
rect 8331 41476 8332 41516
rect 8372 41476 8373 41516
rect 8331 41467 8373 41476
rect 8427 41432 8469 41441
rect 8427 41392 8428 41432
rect 8468 41392 8469 41432
rect 8427 41383 8469 41392
rect 8524 41432 8564 42400
rect 8620 41768 8660 42736
rect 8715 42776 8757 42785
rect 8715 42736 8716 42776
rect 8756 42736 8757 42776
rect 8715 42727 8757 42736
rect 8873 42761 8913 42770
rect 8716 42642 8756 42727
rect 8873 42440 8913 42721
rect 8873 42400 8948 42440
rect 8800 41945 8840 41964
rect 8800 41936 8852 41945
rect 8716 41896 8812 41936
rect 8716 41777 8756 41896
rect 8812 41887 8852 41896
rect 8908 41936 8948 42400
rect 8620 41719 8660 41728
rect 8715 41768 8757 41777
rect 8715 41728 8716 41768
rect 8756 41728 8757 41768
rect 8715 41719 8757 41728
rect 8715 41600 8757 41609
rect 8715 41560 8716 41600
rect 8756 41560 8757 41600
rect 8715 41551 8757 41560
rect 8524 41383 8564 41392
rect 8619 41432 8661 41441
rect 8619 41392 8620 41432
rect 8660 41392 8661 41432
rect 8619 41383 8661 41392
rect 8331 41348 8373 41357
rect 8331 41308 8332 41348
rect 8372 41308 8373 41348
rect 8331 41299 8373 41308
rect 8332 41264 8372 41299
rect 8332 41213 8372 41224
rect 8428 41264 8468 41383
rect 8428 41215 8468 41224
rect 8620 41264 8660 41383
rect 8716 41273 8756 41551
rect 8908 41525 8948 41896
rect 9004 41609 9044 45088
rect 9579 45044 9621 45053
rect 9579 45004 9580 45044
rect 9620 45004 9621 45044
rect 9579 44995 9621 45004
rect 9436 44969 9476 44978
rect 9476 44929 9524 44960
rect 9436 44920 9524 44929
rect 9484 44456 9524 44920
rect 9580 44876 9620 44995
rect 9580 44827 9620 44836
rect 9580 44456 9620 44465
rect 9484 44416 9580 44456
rect 9580 44407 9620 44416
rect 9387 44288 9429 44297
rect 9387 44248 9388 44288
rect 9428 44248 9429 44288
rect 9387 44239 9429 44248
rect 9388 44154 9428 44239
rect 9387 43532 9429 43541
rect 9387 43492 9388 43532
rect 9428 43492 9429 43532
rect 9387 43483 9429 43492
rect 9388 43448 9428 43483
rect 9388 43397 9428 43408
rect 9292 43280 9332 43289
rect 9100 43240 9292 43280
rect 9100 42785 9140 43240
rect 9292 43231 9332 43240
rect 9676 42944 9716 45172
rect 9964 44297 10004 45247
rect 9963 44288 10005 44297
rect 9963 44248 9964 44288
rect 10004 44248 10005 44288
rect 9963 44239 10005 44248
rect 9580 42904 9716 42944
rect 9484 42860 9524 42869
rect 9099 42776 9141 42785
rect 9099 42736 9100 42776
rect 9140 42736 9141 42776
rect 9099 42727 9141 42736
rect 9292 42776 9332 42785
rect 9484 42776 9524 42820
rect 9332 42736 9524 42776
rect 9100 42642 9140 42727
rect 9195 42608 9237 42617
rect 9195 42568 9196 42608
rect 9236 42568 9237 42608
rect 9195 42559 9237 42568
rect 9099 42524 9141 42533
rect 9099 42484 9100 42524
rect 9140 42484 9141 42524
rect 9099 42475 9141 42484
rect 9100 41777 9140 42475
rect 9196 42474 9236 42559
rect 9292 42104 9332 42736
rect 9387 42608 9429 42617
rect 9387 42568 9388 42608
rect 9428 42568 9429 42608
rect 9387 42559 9429 42568
rect 9196 42064 9332 42104
rect 9196 41936 9236 42064
rect 9099 41768 9141 41777
rect 9099 41728 9100 41768
rect 9140 41728 9141 41768
rect 9099 41719 9141 41728
rect 9003 41600 9045 41609
rect 9003 41560 9004 41600
rect 9044 41560 9045 41600
rect 9003 41551 9045 41560
rect 8907 41516 8949 41525
rect 8907 41476 8908 41516
rect 8948 41476 8949 41516
rect 8907 41467 8949 41476
rect 9196 41273 9236 41896
rect 9292 41936 9332 41945
rect 9292 41693 9332 41896
rect 9388 41936 9428 42559
rect 9388 41887 9428 41896
rect 9483 41768 9525 41777
rect 9483 41728 9484 41768
rect 9524 41728 9525 41768
rect 9483 41719 9525 41728
rect 9291 41684 9333 41693
rect 9291 41644 9292 41684
rect 9332 41644 9333 41684
rect 9291 41635 9333 41644
rect 9484 41634 9524 41719
rect 9292 41441 9332 41526
rect 9291 41432 9333 41441
rect 9580 41432 9620 42904
rect 9676 42776 9716 42785
rect 9716 42736 9908 42776
rect 9676 42727 9716 42736
rect 9868 41936 9908 42736
rect 9868 41861 9908 41896
rect 9867 41852 9909 41861
rect 9867 41812 9868 41852
rect 9908 41812 9909 41852
rect 9867 41803 9909 41812
rect 9676 41768 9716 41777
rect 9716 41728 9812 41768
rect 9676 41719 9716 41728
rect 9675 41600 9717 41609
rect 9675 41560 9676 41600
rect 9716 41560 9717 41600
rect 9675 41551 9717 41560
rect 9291 41392 9292 41432
rect 9332 41392 9333 41432
rect 9291 41383 9333 41392
rect 9388 41392 9620 41432
rect 8620 40937 8660 41224
rect 8715 41264 8757 41273
rect 8715 41224 8716 41264
rect 8756 41224 8757 41264
rect 8715 41215 8757 41224
rect 8812 41264 8852 41273
rect 8427 40928 8469 40937
rect 8427 40888 8428 40928
rect 8468 40888 8469 40928
rect 8427 40879 8469 40888
rect 8619 40928 8661 40937
rect 8619 40888 8620 40928
rect 8660 40888 8661 40928
rect 8619 40879 8661 40888
rect 8331 40676 8373 40685
rect 8331 40636 8332 40676
rect 8372 40636 8373 40676
rect 8331 40627 8373 40636
rect 8332 40542 8372 40627
rect 8332 40424 8372 40433
rect 8236 40384 8332 40424
rect 7947 40375 7989 40384
rect 8140 40375 8180 40384
rect 8332 40375 8372 40384
rect 7948 40290 7988 40375
rect 8235 40256 8277 40265
rect 8235 40216 8236 40256
rect 8276 40216 8277 40256
rect 8235 40207 8277 40216
rect 7851 40172 7893 40181
rect 7851 40132 7852 40172
rect 7892 40132 7893 40172
rect 7851 40123 7893 40132
rect 7755 40004 7797 40013
rect 7755 39964 7756 40004
rect 7796 39964 7797 40004
rect 7755 39955 7797 39964
rect 7659 39920 7701 39929
rect 7372 39880 7508 39920
rect 7275 39871 7317 39880
rect 6700 39786 6740 39871
rect 6507 39752 6549 39761
rect 6507 39712 6508 39752
rect 6548 39712 6549 39752
rect 6507 39703 6549 39712
rect 6891 39752 6933 39761
rect 6891 39712 6892 39752
rect 6932 39712 6933 39752
rect 6891 39703 6933 39712
rect 7276 39752 7316 39871
rect 6508 39341 6548 39703
rect 6507 39332 6549 39341
rect 6507 39292 6508 39332
rect 6548 39292 6549 39332
rect 6507 39283 6549 39292
rect 6892 39089 6932 39703
rect 6987 39584 7029 39593
rect 6987 39544 6988 39584
rect 7028 39544 7029 39584
rect 6987 39535 7029 39544
rect 6988 39450 7028 39535
rect 6891 39080 6933 39089
rect 6891 39040 6892 39080
rect 6932 39040 6933 39080
rect 6891 39031 6933 39040
rect 6844 38921 6884 38930
rect 6316 38912 6356 38921
rect 6027 38576 6069 38585
rect 6027 38536 6028 38576
rect 6068 38536 6069 38576
rect 6027 38527 6069 38536
rect 6219 38156 6261 38165
rect 6219 38116 6220 38156
rect 6260 38116 6261 38156
rect 6219 38107 6261 38116
rect 6220 37829 6260 38107
rect 5548 37780 5684 37820
rect 5740 37780 5876 37820
rect 6219 37820 6261 37829
rect 6219 37780 6220 37820
rect 6260 37780 6261 37820
rect 5451 37736 5493 37745
rect 5451 37696 5452 37736
rect 5492 37696 5493 37736
rect 5451 37687 5493 37696
rect 5548 37568 5588 37780
rect 5740 37577 5780 37780
rect 6219 37771 6261 37780
rect 5835 37652 5877 37661
rect 5835 37612 5836 37652
rect 5876 37612 5877 37652
rect 5835 37603 5877 37612
rect 5356 37528 5588 37568
rect 5739 37568 5781 37577
rect 5739 37528 5740 37568
rect 5780 37528 5781 37568
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 5259 36728 5301 36737
rect 5259 36688 5260 36728
rect 5300 36688 5301 36728
rect 5259 36679 5301 36688
rect 5260 35888 5300 36679
rect 5260 35729 5300 35848
rect 5259 35720 5301 35729
rect 5259 35680 5260 35720
rect 5300 35680 5301 35720
rect 5259 35671 5301 35680
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 5356 35384 5396 37528
rect 5739 37519 5781 37528
rect 5452 37400 5492 37409
rect 5740 37400 5780 37409
rect 5492 37360 5740 37400
rect 5452 36905 5492 37360
rect 5740 37351 5780 37360
rect 5836 37400 5876 37603
rect 6316 37568 6356 38872
rect 6411 38912 6453 38921
rect 6411 38872 6412 38912
rect 6452 38872 6453 38912
rect 7276 38912 7316 39712
rect 7371 39752 7413 39761
rect 7371 39712 7372 39752
rect 7412 39712 7413 39752
rect 7371 39703 7413 39712
rect 7372 39618 7412 39703
rect 6884 38881 6932 38912
rect 6844 38872 6932 38881
rect 6411 38863 6453 38872
rect 6892 38408 6932 38872
rect 7276 38863 7316 38872
rect 7372 38912 7412 38921
rect 7468 38912 7508 39880
rect 7659 39880 7660 39920
rect 7700 39880 7701 39920
rect 7659 39871 7701 39880
rect 7660 39752 7700 39871
rect 7756 39752 7796 39761
rect 7660 39712 7756 39752
rect 7756 39703 7796 39712
rect 7852 39752 7892 40123
rect 8043 40088 8085 40097
rect 8043 40048 8044 40088
rect 8084 40048 8085 40088
rect 8043 40039 8085 40048
rect 7947 39920 7989 39929
rect 7947 39880 7948 39920
rect 7988 39880 7989 39920
rect 7947 39871 7989 39880
rect 7852 39703 7892 39712
rect 7563 39332 7605 39341
rect 7563 39292 7564 39332
rect 7604 39292 7605 39332
rect 7563 39283 7605 39292
rect 7412 38872 7508 38912
rect 6987 38828 7029 38837
rect 6987 38788 6988 38828
rect 7028 38788 7029 38828
rect 6987 38779 7029 38788
rect 6988 38694 7028 38779
rect 6988 38408 7028 38417
rect 6892 38368 6988 38408
rect 6988 38359 7028 38368
rect 6795 38240 6837 38249
rect 6795 38200 6796 38240
rect 6836 38200 6837 38240
rect 6795 38191 6837 38200
rect 6796 37577 6836 38191
rect 7372 37820 7412 38872
rect 7467 38660 7509 38669
rect 7467 38620 7468 38660
rect 7508 38620 7509 38660
rect 7467 38611 7509 38620
rect 7180 37780 7412 37820
rect 6795 37568 6837 37577
rect 6316 37528 6644 37568
rect 5836 37351 5876 37360
rect 5932 37400 5972 37409
rect 5548 37232 5588 37241
rect 5588 37192 5684 37232
rect 5548 37183 5588 37192
rect 5451 36896 5493 36905
rect 5451 36856 5452 36896
rect 5492 36856 5493 36896
rect 5451 36847 5493 36856
rect 5452 36569 5492 36847
rect 5644 36653 5684 37192
rect 5932 37064 5972 37360
rect 6027 37400 6069 37409
rect 6316 37400 6356 37409
rect 6027 37360 6028 37400
rect 6068 37360 6069 37400
rect 6027 37351 6069 37360
rect 6124 37360 6316 37400
rect 6028 37266 6068 37351
rect 5836 37024 5972 37064
rect 5739 36728 5781 36737
rect 5739 36688 5740 36728
rect 5780 36688 5781 36728
rect 5739 36679 5781 36688
rect 5643 36644 5685 36653
rect 5643 36604 5644 36644
rect 5684 36604 5685 36644
rect 5643 36595 5685 36604
rect 5451 36560 5493 36569
rect 5451 36520 5452 36560
rect 5492 36520 5493 36560
rect 5451 36511 5493 36520
rect 5451 36140 5493 36149
rect 5451 36100 5452 36140
rect 5492 36100 5493 36140
rect 5451 36091 5493 36100
rect 5452 36006 5492 36091
rect 5644 35888 5684 36595
rect 5740 36594 5780 36679
rect 5836 36149 5876 37024
rect 5932 36896 5972 36905
rect 6124 36896 6164 37360
rect 6316 37351 6356 37360
rect 6411 37400 6453 37409
rect 6411 37360 6412 37400
rect 6452 37360 6453 37400
rect 6411 37351 6453 37360
rect 6508 37400 6548 37409
rect 6412 37266 6452 37351
rect 6219 37232 6261 37241
rect 6219 37192 6220 37232
rect 6260 37192 6261 37232
rect 6219 37183 6261 37192
rect 6220 37098 6260 37183
rect 6411 37064 6453 37073
rect 6508 37064 6548 37360
rect 6411 37024 6412 37064
rect 6452 37024 6548 37064
rect 6411 37015 6453 37024
rect 6604 36980 6644 37528
rect 6795 37528 6796 37568
rect 6836 37528 6837 37568
rect 6795 37519 6837 37528
rect 6700 37400 6740 37409
rect 6700 37073 6740 37360
rect 7083 37232 7125 37241
rect 7083 37192 7084 37232
rect 7124 37192 7125 37232
rect 7083 37183 7125 37192
rect 6699 37064 6741 37073
rect 6699 37024 6700 37064
rect 6740 37024 6741 37064
rect 6699 37015 6741 37024
rect 5972 36856 6164 36896
rect 6507 36940 6644 36980
rect 6507 36896 6547 36940
rect 6795 36896 6837 36905
rect 6507 36856 6548 36896
rect 5932 36847 5972 36856
rect 6124 36728 6164 36856
rect 6219 36812 6261 36821
rect 6219 36772 6220 36812
rect 6260 36772 6261 36812
rect 6219 36763 6261 36772
rect 6124 36679 6164 36688
rect 6220 36678 6260 36763
rect 6315 36728 6357 36737
rect 6315 36688 6316 36728
rect 6356 36688 6357 36728
rect 6315 36679 6357 36688
rect 6412 36709 6452 36718
rect 6316 36594 6356 36679
rect 6315 36476 6357 36485
rect 6315 36436 6316 36476
rect 6356 36436 6357 36476
rect 6315 36427 6357 36436
rect 6027 36308 6069 36317
rect 6027 36268 6028 36308
rect 6068 36268 6069 36308
rect 6027 36259 6069 36268
rect 5835 36140 5877 36149
rect 5835 36100 5836 36140
rect 5876 36100 5877 36140
rect 5835 36091 5877 36100
rect 5740 35888 5780 35897
rect 5644 35848 5740 35888
rect 5740 35839 5780 35848
rect 5836 35888 5876 35897
rect 5452 35720 5492 35729
rect 5452 35393 5492 35680
rect 5643 35720 5685 35729
rect 5643 35680 5644 35720
rect 5684 35680 5685 35720
rect 5643 35671 5685 35680
rect 5164 35344 5396 35384
rect 5451 35384 5493 35393
rect 5451 35344 5452 35384
rect 5492 35344 5493 35384
rect 4971 34964 5013 34973
rect 4971 34924 4972 34964
rect 5012 34924 5013 34964
rect 4971 34915 5013 34924
rect 4972 34385 5012 34915
rect 4971 34376 5013 34385
rect 4971 34336 4972 34376
rect 5012 34336 5013 34376
rect 4971 34327 5013 34336
rect 5164 34208 5204 35344
rect 5451 35335 5493 35344
rect 5259 35216 5301 35225
rect 5259 35176 5260 35216
rect 5300 35176 5301 35216
rect 5259 35167 5301 35176
rect 5356 35216 5396 35225
rect 5260 35082 5300 35167
rect 5259 34880 5301 34889
rect 5259 34840 5260 34880
rect 5300 34840 5301 34880
rect 5259 34831 5301 34840
rect 5260 34376 5300 34831
rect 5356 34544 5396 35176
rect 5451 35216 5493 35225
rect 5451 35176 5452 35216
rect 5492 35176 5493 35216
rect 5451 35167 5493 35176
rect 5548 35216 5588 35225
rect 5452 35082 5492 35167
rect 5548 34721 5588 35176
rect 5644 34889 5684 35671
rect 5836 35552 5876 35848
rect 5931 35888 5973 35897
rect 5931 35848 5932 35888
rect 5972 35848 5973 35888
rect 5931 35839 5973 35848
rect 6028 35888 6068 36259
rect 6028 35839 6068 35848
rect 6316 35888 6356 36427
rect 6412 36149 6452 36669
rect 6411 36140 6453 36149
rect 6411 36100 6412 36140
rect 6452 36100 6453 36140
rect 6411 36091 6453 36100
rect 5932 35754 5972 35839
rect 5836 35512 6260 35552
rect 5931 35384 5973 35393
rect 5931 35344 5932 35384
rect 5972 35344 5973 35384
rect 5931 35335 5973 35344
rect 5740 35216 5780 35225
rect 5643 34880 5685 34889
rect 5643 34840 5644 34880
rect 5684 34840 5685 34880
rect 5643 34831 5685 34840
rect 5547 34712 5589 34721
rect 5740 34712 5780 35176
rect 5836 35216 5876 35227
rect 5836 35141 5876 35176
rect 5932 35216 5972 35335
rect 6027 35300 6069 35309
rect 6027 35260 6028 35300
rect 6068 35260 6069 35300
rect 6027 35251 6069 35260
rect 5932 35167 5972 35176
rect 6028 35166 6068 35251
rect 6123 35216 6165 35225
rect 6123 35176 6124 35216
rect 6164 35176 6165 35216
rect 6123 35167 6165 35176
rect 5835 35132 5877 35141
rect 5835 35092 5836 35132
rect 5876 35092 5877 35132
rect 5835 35083 5877 35092
rect 5547 34672 5548 34712
rect 5588 34672 5589 34712
rect 5547 34663 5589 34672
rect 5644 34672 5780 34712
rect 5835 34712 5877 34721
rect 5835 34672 5836 34712
rect 5876 34672 5877 34712
rect 5451 34544 5493 34553
rect 5356 34504 5452 34544
rect 5492 34504 5493 34544
rect 5451 34495 5493 34504
rect 5452 34410 5492 34495
rect 5260 34292 5300 34336
rect 5260 34252 5492 34292
rect 5164 34168 5396 34208
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 5356 32360 5396 34168
rect 5452 33704 5492 34252
rect 5548 33704 5588 33713
rect 5452 33664 5548 33704
rect 5452 32864 5492 33664
rect 5548 33655 5588 33664
rect 5644 33536 5684 34672
rect 5835 34663 5877 34672
rect 5836 34544 5876 34663
rect 5740 34504 5876 34544
rect 5740 34376 5780 34504
rect 5740 34327 5780 34336
rect 5835 34376 5877 34385
rect 6124 34376 6164 35167
rect 6220 35057 6260 35512
rect 6316 35216 6356 35848
rect 6316 35141 6356 35176
rect 6411 35216 6453 35225
rect 6411 35176 6412 35216
rect 6452 35176 6453 35216
rect 6411 35167 6453 35176
rect 6315 35132 6357 35141
rect 6315 35092 6316 35132
rect 6356 35092 6357 35132
rect 6315 35083 6357 35092
rect 6219 35048 6261 35057
rect 6316 35052 6356 35083
rect 6219 35008 6220 35048
rect 6260 35008 6261 35048
rect 6219 34999 6261 35008
rect 6219 34796 6261 34805
rect 6219 34756 6220 34796
rect 6260 34756 6261 34796
rect 6219 34747 6261 34756
rect 5835 34336 5836 34376
rect 5876 34336 5877 34376
rect 5835 34327 5877 34336
rect 5932 34336 6124 34376
rect 5836 34242 5876 34327
rect 5739 33788 5781 33797
rect 5739 33748 5740 33788
rect 5780 33748 5781 33788
rect 5739 33739 5781 33748
rect 5740 33654 5780 33739
rect 5932 33704 5972 34336
rect 6124 34327 6164 34336
rect 6220 34376 6260 34747
rect 6315 34544 6357 34553
rect 6315 34504 6316 34544
rect 6356 34504 6357 34544
rect 6315 34495 6357 34504
rect 6220 34327 6260 34336
rect 6316 34376 6356 34495
rect 6027 34208 6069 34217
rect 6027 34168 6028 34208
rect 6068 34168 6069 34208
rect 6027 34159 6069 34168
rect 6028 34074 6068 34159
rect 6219 34124 6261 34133
rect 6219 34084 6220 34124
rect 6260 34084 6261 34124
rect 6219 34075 6261 34084
rect 6123 33872 6165 33881
rect 6123 33832 6124 33872
rect 6164 33832 6165 33872
rect 6123 33823 6165 33832
rect 5548 33496 5684 33536
rect 5548 32948 5588 33496
rect 5644 33116 5684 33125
rect 5932 33116 5972 33664
rect 6027 33704 6069 33713
rect 6027 33664 6028 33704
rect 6068 33664 6069 33704
rect 6027 33655 6069 33664
rect 6028 33570 6068 33655
rect 5684 33076 5972 33116
rect 5644 33067 5684 33076
rect 5931 32948 5973 32957
rect 5548 32908 5684 32948
rect 5492 32824 5588 32864
rect 5452 32815 5492 32824
rect 5452 32360 5492 32369
rect 5356 32320 5452 32360
rect 5452 31529 5492 32320
rect 5548 31613 5588 32824
rect 5644 31697 5684 32908
rect 5931 32908 5932 32948
rect 5972 32908 5973 32948
rect 5931 32899 5973 32908
rect 5835 32864 5877 32873
rect 5835 32824 5836 32864
rect 5876 32824 5877 32864
rect 5835 32815 5877 32824
rect 5836 32730 5876 32815
rect 5932 32814 5972 32899
rect 6028 32864 6068 32873
rect 6124 32864 6164 33823
rect 6068 32824 6164 32864
rect 6028 32815 6068 32824
rect 5931 32696 5973 32705
rect 5931 32656 5932 32696
rect 5972 32656 5973 32696
rect 5931 32647 5973 32656
rect 5740 32192 5780 32201
rect 5740 31865 5780 32152
rect 5739 31856 5781 31865
rect 5739 31816 5740 31856
rect 5780 31816 5781 31856
rect 5739 31807 5781 31816
rect 5643 31688 5685 31697
rect 5643 31648 5644 31688
rect 5684 31648 5685 31688
rect 5643 31639 5685 31648
rect 5547 31604 5589 31613
rect 5547 31564 5548 31604
rect 5588 31564 5589 31604
rect 5547 31555 5589 31564
rect 5451 31520 5493 31529
rect 5451 31480 5452 31520
rect 5492 31480 5493 31520
rect 5451 31471 5493 31480
rect 4683 31436 4725 31445
rect 4683 31396 4684 31436
rect 4724 31396 4725 31436
rect 4683 31387 4725 31396
rect 4876 31357 4916 31366
rect 4876 31184 4916 31317
rect 5067 31268 5109 31277
rect 5067 31228 5068 31268
rect 5108 31228 5109 31268
rect 5067 31219 5109 31228
rect 4780 31144 4916 31184
rect 4683 31016 4725 31025
rect 4683 30976 4684 31016
rect 4724 30976 4725 31016
rect 4683 30967 4725 30976
rect 4684 28673 4724 30967
rect 4780 30857 4820 31144
rect 5068 31134 5108 31219
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4779 30848 4821 30857
rect 4779 30808 4780 30848
rect 4820 30808 4821 30848
rect 4779 30799 4821 30808
rect 5259 30848 5301 30857
rect 5259 30808 5260 30848
rect 5300 30808 5301 30848
rect 5259 30799 5301 30808
rect 5452 30848 5492 31471
rect 5643 31436 5685 31445
rect 5643 31396 5644 31436
rect 5684 31396 5685 31436
rect 5643 31387 5685 31396
rect 5452 30799 5492 30808
rect 5548 31352 5588 31361
rect 5260 30714 5300 30799
rect 5548 30689 5588 31312
rect 5644 31352 5684 31387
rect 5068 30680 5108 30689
rect 5068 30521 5108 30640
rect 5547 30680 5589 30689
rect 5547 30640 5548 30680
rect 5588 30640 5589 30680
rect 5547 30631 5589 30640
rect 5067 30512 5109 30521
rect 5644 30512 5684 31312
rect 5835 31016 5877 31025
rect 5835 30976 5836 31016
rect 5876 30976 5877 31016
rect 5835 30967 5877 30976
rect 5739 30680 5781 30689
rect 5739 30640 5740 30680
rect 5780 30640 5781 30680
rect 5739 30631 5781 30640
rect 5067 30472 5068 30512
rect 5108 30472 5109 30512
rect 5067 30463 5109 30472
rect 5452 30472 5684 30512
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 4683 28664 4725 28673
rect 4683 28624 4684 28664
rect 4724 28624 4725 28664
rect 4683 28615 4725 28624
rect 4684 28085 4724 28615
rect 4683 28076 4725 28085
rect 4683 28036 4684 28076
rect 4724 28036 4725 28076
rect 4683 28027 4725 28036
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4588 27868 4820 27908
rect 4587 27740 4629 27749
rect 4587 27700 4588 27740
rect 4628 27700 4629 27740
rect 4587 27691 4629 27700
rect 4588 27606 4628 27691
rect 4492 27448 4628 27488
rect 4492 26816 4532 26825
rect 4492 26489 4532 26776
rect 4491 26480 4533 26489
rect 4491 26440 4492 26480
rect 4532 26440 4533 26480
rect 4491 26431 4533 26440
rect 4492 26312 4532 26321
rect 4396 26272 4492 26312
rect 4492 26263 4532 26272
rect 4108 26188 4244 26228
rect 3819 26144 3861 26153
rect 3819 26104 3820 26144
rect 3860 26104 3861 26144
rect 3819 26095 3861 26104
rect 3531 25808 3573 25817
rect 3531 25768 3532 25808
rect 3572 25768 3573 25808
rect 3531 25759 3573 25768
rect 3532 25061 3572 25759
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 3531 25052 3573 25061
rect 3531 25012 3532 25052
rect 3572 25012 3573 25052
rect 3531 25003 3573 25012
rect 3435 24968 3477 24977
rect 3435 24928 3436 24968
rect 3476 24928 3477 24968
rect 3435 24919 3477 24928
rect 3148 24088 3380 24128
rect 3148 21608 3188 24088
rect 3436 23876 3476 24919
rect 3915 24800 3957 24809
rect 3915 24760 3916 24800
rect 3956 24760 3957 24800
rect 3915 24751 3957 24760
rect 3916 24666 3956 24751
rect 3531 24632 3573 24641
rect 3531 24592 3532 24632
rect 3572 24592 3573 24632
rect 4108 24632 4148 26188
rect 4299 26144 4341 26153
rect 4299 26104 4300 26144
rect 4340 26104 4341 26144
rect 4299 26095 4341 26104
rect 4300 26010 4340 26095
rect 4299 25472 4341 25481
rect 4299 25432 4300 25472
rect 4340 25432 4341 25472
rect 4299 25423 4341 25432
rect 4300 25304 4340 25423
rect 4300 25255 4340 25264
rect 4491 25304 4533 25313
rect 4491 25264 4492 25304
rect 4532 25264 4533 25304
rect 4491 25255 4533 25264
rect 4492 25170 4532 25255
rect 4300 24632 4340 24641
rect 3531 24583 3573 24592
rect 3724 24618 3764 24627
rect 3532 24053 3572 24583
rect 4108 24592 4300 24632
rect 3724 24389 3764 24578
rect 4300 24473 4340 24592
rect 4299 24464 4341 24473
rect 4299 24424 4300 24464
rect 4340 24424 4341 24464
rect 4299 24415 4341 24424
rect 3723 24380 3765 24389
rect 3723 24340 3724 24380
rect 3764 24340 3765 24380
rect 3723 24331 3765 24340
rect 4203 24380 4245 24389
rect 4203 24340 4204 24380
rect 4244 24340 4245 24380
rect 4203 24331 4245 24340
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 3531 24044 3573 24053
rect 3531 24004 3532 24044
rect 3572 24004 3573 24044
rect 3531 23995 3573 24004
rect 3435 23836 3476 23876
rect 3340 23792 3380 23801
rect 3340 23633 3380 23752
rect 3435 23708 3475 23836
rect 3435 23668 3476 23708
rect 3339 23624 3381 23633
rect 3339 23584 3340 23624
rect 3380 23584 3381 23624
rect 3339 23575 3381 23584
rect 3148 20777 3188 21568
rect 3243 21608 3285 21617
rect 3243 21568 3244 21608
rect 3284 21568 3285 21608
rect 3243 21559 3285 21568
rect 3147 20768 3189 20777
rect 3147 20728 3148 20768
rect 3188 20728 3189 20768
rect 3147 20719 3189 20728
rect 2668 20476 3092 20516
rect 2668 20264 2708 20476
rect 3148 20432 3188 20719
rect 2668 20215 2708 20224
rect 2860 20392 3188 20432
rect 2667 20096 2709 20105
rect 2667 20056 2668 20096
rect 2708 20056 2709 20096
rect 2667 20047 2709 20056
rect 2668 19508 2708 20047
rect 2668 19459 2708 19468
rect 2763 19256 2805 19265
rect 2763 19216 2764 19256
rect 2804 19216 2805 19256
rect 2763 19207 2805 19216
rect 2668 18570 2708 18579
rect 2668 18173 2708 18530
rect 2667 18164 2709 18173
rect 2667 18124 2668 18164
rect 2708 18124 2709 18164
rect 2667 18115 2709 18124
rect 2668 17996 2708 18005
rect 2572 17956 2668 17996
rect 2668 17947 2708 17956
rect 2475 17744 2517 17753
rect 2475 17704 2476 17744
rect 2516 17704 2517 17744
rect 2475 17695 2517 17704
rect 2188 17156 2228 17165
rect 2091 15644 2133 15653
rect 2091 15604 2092 15644
rect 2132 15604 2133 15644
rect 2091 15595 2133 15604
rect 1996 14671 2036 14680
rect 1707 14468 1749 14477
rect 1707 14428 1708 14468
rect 1748 14428 1749 14468
rect 1707 14419 1749 14428
rect 1516 14344 1652 14384
rect 1419 13208 1461 13217
rect 1419 13168 1420 13208
rect 1460 13168 1461 13208
rect 1419 13159 1461 13168
rect 1419 13040 1461 13049
rect 1419 13000 1420 13040
rect 1460 13000 1461 13040
rect 1419 12991 1461 13000
rect 1420 12906 1460 12991
rect 1516 12788 1556 14344
rect 1803 14216 1845 14225
rect 1803 14176 1804 14216
rect 1844 14176 1845 14216
rect 1803 14167 1845 14176
rect 1804 13460 1844 14167
rect 2091 13628 2133 13637
rect 2091 13588 2092 13628
rect 2132 13588 2133 13628
rect 2091 13579 2133 13588
rect 1804 13411 1844 13420
rect 1611 13292 1653 13301
rect 1611 13252 1612 13292
rect 1652 13252 1653 13292
rect 1611 13243 1653 13252
rect 1996 13292 2036 13301
rect 1612 13158 1652 13243
rect 1996 13133 2036 13252
rect 1995 13124 2037 13133
rect 1995 13084 1996 13124
rect 2036 13084 2037 13124
rect 1995 13075 2037 13084
rect 1268 11656 1364 11696
rect 1420 12748 1556 12788
rect 1228 11647 1268 11656
rect 1420 10436 1460 12748
rect 2092 12620 2132 13579
rect 1996 12580 2132 12620
rect 1707 12452 1749 12461
rect 1707 12412 1708 12452
rect 1748 12412 1749 12452
rect 1707 12403 1749 12412
rect 1708 12318 1748 12403
rect 1516 12284 1556 12293
rect 1516 10940 1556 12244
rect 1803 12284 1845 12293
rect 1803 12244 1804 12284
rect 1844 12244 1845 12284
rect 1803 12235 1845 12244
rect 1900 12284 1940 12293
rect 1707 11108 1749 11117
rect 1707 11068 1708 11108
rect 1748 11068 1749 11108
rect 1707 11059 1749 11068
rect 1708 10940 1748 11059
rect 1516 10900 1652 10940
rect 1516 10772 1556 10781
rect 1420 10396 1470 10436
rect 1430 10268 1470 10396
rect 1420 10228 1470 10268
rect 1228 10184 1268 10193
rect 1420 10184 1460 10228
rect 1516 10193 1556 10732
rect 1268 10144 1460 10184
rect 1515 10184 1557 10193
rect 1515 10144 1516 10184
rect 1556 10144 1557 10184
rect 1228 10135 1268 10144
rect 1515 10135 1557 10144
rect 1515 10016 1557 10025
rect 1515 9976 1516 10016
rect 1556 9976 1557 10016
rect 1515 9967 1557 9976
rect 1323 9932 1365 9941
rect 1323 9892 1324 9932
rect 1364 9892 1365 9932
rect 1323 9883 1365 9892
rect 1131 8756 1173 8765
rect 1131 8716 1132 8756
rect 1172 8716 1173 8756
rect 1131 8707 1173 8716
rect 1228 8672 1268 8681
rect 1324 8672 1364 9883
rect 1419 9848 1461 9857
rect 1419 9808 1420 9848
rect 1460 9808 1461 9848
rect 1419 9799 1461 9808
rect 1420 9680 1460 9799
rect 1420 9631 1460 9640
rect 1268 8632 1364 8672
rect 1228 8623 1268 8632
rect 1419 8504 1461 8513
rect 1419 8464 1420 8504
rect 1460 8464 1461 8504
rect 1419 8455 1461 8464
rect 1227 8000 1269 8009
rect 1227 7960 1228 8000
rect 1268 7960 1269 8000
rect 1227 7951 1269 7960
rect 1228 7866 1268 7951
rect 1323 7916 1365 7925
rect 1323 7876 1324 7916
rect 1364 7876 1365 7916
rect 1323 7867 1365 7876
rect 1131 7832 1173 7841
rect 1131 7792 1132 7832
rect 1172 7792 1173 7832
rect 1131 7783 1173 7792
rect 1035 7160 1077 7169
rect 1035 7120 1036 7160
rect 1076 7120 1077 7160
rect 1035 7111 1077 7120
rect 843 6824 885 6833
rect 843 6784 844 6824
rect 884 6784 885 6824
rect 843 6775 885 6784
rect 171 1784 213 1793
rect 171 1744 172 1784
rect 212 1744 213 1784
rect 171 1735 213 1744
rect 1036 953 1076 7111
rect 1132 2213 1172 7783
rect 1227 6488 1269 6497
rect 1227 6448 1228 6488
rect 1268 6448 1269 6488
rect 1227 6439 1269 6448
rect 1228 4976 1268 6439
rect 1228 4927 1268 4936
rect 1228 4136 1268 4145
rect 1324 4136 1364 7867
rect 1420 5900 1460 8455
rect 1516 7160 1556 9967
rect 1612 9532 1652 10900
rect 1708 10891 1748 10900
rect 1612 9492 1748 9532
rect 1611 9428 1653 9437
rect 1611 9388 1612 9428
rect 1652 9388 1653 9428
rect 1611 9379 1653 9388
rect 1612 9294 1652 9379
rect 1611 7496 1653 7505
rect 1611 7456 1612 7496
rect 1652 7456 1653 7496
rect 1611 7447 1653 7456
rect 1516 7111 1556 7120
rect 1516 5900 1556 5909
rect 1420 5860 1516 5900
rect 1516 5851 1556 5860
rect 1419 5228 1461 5237
rect 1419 5188 1420 5228
rect 1460 5188 1461 5228
rect 1419 5179 1461 5188
rect 1268 4096 1364 4136
rect 1228 4087 1268 4096
rect 1420 3884 1460 5179
rect 1324 3844 1460 3884
rect 1324 3716 1364 3844
rect 1228 3676 1364 3716
rect 1419 3716 1461 3725
rect 1419 3676 1420 3716
rect 1460 3676 1461 3716
rect 1131 2204 1173 2213
rect 1131 2164 1132 2204
rect 1172 2164 1173 2204
rect 1131 2155 1173 2164
rect 1228 1952 1268 3676
rect 1419 3667 1461 3676
rect 1323 3548 1365 3557
rect 1323 3508 1324 3548
rect 1364 3508 1365 3548
rect 1323 3499 1365 3508
rect 1324 3414 1364 3499
rect 1420 3128 1460 3667
rect 1516 3632 1556 3641
rect 1612 3632 1652 7447
rect 1708 6404 1748 9492
rect 1804 9437 1844 12235
rect 1900 11873 1940 12244
rect 1899 11864 1941 11873
rect 1899 11824 1900 11864
rect 1940 11824 1941 11864
rect 1899 11815 1941 11824
rect 1899 11192 1941 11201
rect 1899 11152 1900 11192
rect 1940 11152 1941 11192
rect 1899 11143 1941 11152
rect 1900 11058 1940 11143
rect 1996 10445 2036 12580
rect 2091 12452 2133 12461
rect 2091 12412 2092 12452
rect 2132 12412 2133 12452
rect 2091 12403 2133 12412
rect 2092 12318 2132 12403
rect 2091 12116 2133 12125
rect 2091 12076 2092 12116
rect 2132 12076 2133 12116
rect 2091 12067 2133 12076
rect 2092 10940 2132 12067
rect 2188 12041 2228 17116
rect 2380 17058 2420 17067
rect 2283 14552 2325 14561
rect 2283 14512 2284 14552
rect 2324 14512 2325 14552
rect 2283 14503 2325 14512
rect 2284 13460 2324 14503
rect 2380 13637 2420 17018
rect 2476 15560 2516 17695
rect 2667 17660 2709 17669
rect 2667 17620 2668 17660
rect 2708 17620 2709 17660
rect 2667 17611 2709 17620
rect 2668 16829 2708 17611
rect 2667 16820 2709 16829
rect 2667 16780 2668 16820
rect 2708 16780 2709 16820
rect 2667 16771 2709 16780
rect 2764 16400 2804 19207
rect 2860 17072 2900 20392
rect 3244 19265 3284 21559
rect 3436 19517 3476 23668
rect 3532 23633 3572 23995
rect 3868 23801 3908 23810
rect 4204 23792 4244 24331
rect 3908 23761 4148 23792
rect 3868 23752 4148 23761
rect 3531 23624 3573 23633
rect 3531 23584 3532 23624
rect 3572 23584 3573 23624
rect 3531 23575 3573 23584
rect 4011 23624 4053 23633
rect 4011 23584 4012 23624
rect 4052 23584 4053 23624
rect 4011 23575 4053 23584
rect 4012 23490 4052 23575
rect 3724 23213 3764 23244
rect 3723 23204 3765 23213
rect 3723 23164 3724 23204
rect 3764 23164 3765 23204
rect 3723 23155 3765 23164
rect 3724 23120 3764 23155
rect 3724 23045 3764 23080
rect 3723 23036 3765 23045
rect 3723 22996 3724 23036
rect 3764 22996 3765 23036
rect 3723 22987 3765 22996
rect 4108 22952 4148 23752
rect 4244 23752 4436 23792
rect 4204 23743 4244 23752
rect 4108 22912 4340 22952
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 4011 22532 4053 22541
rect 4011 22492 4012 22532
rect 4052 22492 4053 22532
rect 4011 22483 4053 22492
rect 4300 22532 4340 22912
rect 4300 22483 4340 22492
rect 4012 22280 4052 22483
rect 4108 22280 4148 22289
rect 4012 22240 4108 22280
rect 4012 21701 4052 22240
rect 4108 22231 4148 22240
rect 4299 22112 4341 22121
rect 4299 22072 4300 22112
rect 4340 22072 4341 22112
rect 4299 22063 4341 22072
rect 4011 21692 4053 21701
rect 4011 21652 4012 21692
rect 4052 21652 4053 21692
rect 4011 21643 4053 21652
rect 3628 21533 3668 21618
rect 4108 21608 4148 21617
rect 3627 21524 3669 21533
rect 3627 21484 3628 21524
rect 3668 21484 3669 21524
rect 3627 21475 3669 21484
rect 3724 21524 3764 21533
rect 3724 21356 3764 21484
rect 3532 21316 3764 21356
rect 3435 19508 3477 19517
rect 3435 19468 3436 19508
rect 3476 19468 3477 19508
rect 3435 19459 3477 19468
rect 2860 16661 2900 17032
rect 2956 19256 2996 19265
rect 2859 16652 2901 16661
rect 2859 16612 2860 16652
rect 2900 16612 2901 16652
rect 2859 16603 2901 16612
rect 2764 16360 2900 16400
rect 2668 16232 2708 16241
rect 2476 15511 2516 15520
rect 2572 16192 2668 16232
rect 2475 15392 2517 15401
rect 2475 15352 2476 15392
rect 2516 15352 2517 15392
rect 2475 15343 2517 15352
rect 2476 14645 2516 15343
rect 2475 14636 2517 14645
rect 2475 14596 2476 14636
rect 2516 14596 2517 14636
rect 2475 14587 2517 14596
rect 2476 14048 2516 14587
rect 2379 13628 2421 13637
rect 2379 13588 2380 13628
rect 2420 13588 2421 13628
rect 2379 13579 2421 13588
rect 2284 13420 2420 13460
rect 2284 13208 2324 13217
rect 2284 12536 2324 13168
rect 2380 13208 2420 13420
rect 2380 13159 2420 13168
rect 2476 12629 2516 14008
rect 2475 12620 2517 12629
rect 2475 12580 2476 12620
rect 2516 12580 2517 12620
rect 2475 12571 2517 12580
rect 2284 12496 2420 12536
rect 2284 12284 2324 12293
rect 2187 12032 2229 12041
rect 2187 11992 2188 12032
rect 2228 11992 2229 12032
rect 2187 11983 2229 11992
rect 2187 11192 2229 11201
rect 2187 11152 2188 11192
rect 2228 11152 2229 11192
rect 2187 11143 2229 11152
rect 2092 10891 2132 10900
rect 2188 10772 2228 11143
rect 2092 10732 2228 10772
rect 1995 10436 2037 10445
rect 1995 10396 1996 10436
rect 2036 10396 2037 10436
rect 1995 10387 2037 10396
rect 1803 9428 1845 9437
rect 1803 9388 1804 9428
rect 1844 9388 1845 9428
rect 1803 9379 1845 9388
rect 1995 9428 2037 9437
rect 1995 9388 1996 9428
rect 2036 9388 2037 9428
rect 1995 9379 2037 9388
rect 1996 9294 2036 9379
rect 1804 9260 1844 9269
rect 1804 8177 1844 9220
rect 1899 9176 1941 9185
rect 1899 9136 1900 9176
rect 1940 9136 1941 9176
rect 1899 9127 1941 9136
rect 1803 8168 1845 8177
rect 1803 8128 1804 8168
rect 1844 8128 1845 8168
rect 1803 8119 1845 8128
rect 1708 6364 1844 6404
rect 1707 6236 1749 6245
rect 1707 6196 1708 6236
rect 1748 6196 1749 6236
rect 1707 6187 1749 6196
rect 1708 5732 1748 6187
rect 1708 5683 1748 5692
rect 1707 4472 1749 4481
rect 1707 4432 1708 4472
rect 1748 4432 1749 4472
rect 1707 4423 1749 4432
rect 1556 3592 1652 3632
rect 1516 3583 1556 3592
rect 1708 3380 1748 4423
rect 1804 4136 1844 6364
rect 1900 5900 1940 9127
rect 1995 8084 2037 8093
rect 1995 8044 1996 8084
rect 2036 8044 2037 8084
rect 1995 8035 2037 8044
rect 1900 5851 1940 5860
rect 1996 5732 2036 8035
rect 2092 8009 2132 10732
rect 2187 10520 2229 10529
rect 2187 10480 2188 10520
rect 2228 10480 2229 10520
rect 2187 10471 2229 10480
rect 2188 9680 2228 10471
rect 2284 9689 2324 12244
rect 2188 9631 2228 9640
rect 2283 9680 2325 9689
rect 2283 9640 2284 9680
rect 2324 9640 2325 9680
rect 2283 9631 2325 9640
rect 2380 9532 2420 12496
rect 2476 12452 2516 12461
rect 2476 12041 2516 12412
rect 2475 12032 2517 12041
rect 2475 11992 2476 12032
rect 2516 11992 2517 12032
rect 2475 11983 2517 11992
rect 2475 11864 2517 11873
rect 2475 11824 2476 11864
rect 2516 11824 2517 11864
rect 2475 11815 2517 11824
rect 2476 11696 2516 11815
rect 2476 11647 2516 11656
rect 2572 11621 2612 16192
rect 2668 16183 2708 16192
rect 2764 16232 2804 16241
rect 2764 15989 2804 16192
rect 2763 15980 2805 15989
rect 2763 15940 2764 15980
rect 2804 15940 2805 15980
rect 2763 15931 2805 15940
rect 2668 15728 2708 15737
rect 2860 15728 2900 16360
rect 2708 15688 2900 15728
rect 2668 15679 2708 15688
rect 2859 15560 2901 15569
rect 2859 15520 2860 15560
rect 2900 15520 2901 15560
rect 2859 15511 2901 15520
rect 2860 15392 2900 15511
rect 2860 15343 2900 15352
rect 2956 14468 2996 19216
rect 3052 19256 3092 19265
rect 3052 19004 3092 19216
rect 3243 19256 3285 19265
rect 3243 19216 3244 19256
rect 3284 19216 3285 19256
rect 3243 19207 3285 19216
rect 3436 19256 3476 19265
rect 3052 18964 3284 19004
rect 3147 18836 3189 18845
rect 3147 18796 3148 18836
rect 3188 18796 3189 18836
rect 3147 18787 3189 18796
rect 3148 18584 3188 18787
rect 3052 18544 3148 18584
rect 3052 16904 3092 18544
rect 3148 18535 3188 18544
rect 3147 17408 3189 17417
rect 3147 17368 3148 17408
rect 3188 17368 3189 17408
rect 3147 17359 3189 17368
rect 3148 16988 3188 17359
rect 3244 17249 3284 18964
rect 3339 18500 3381 18509
rect 3339 18460 3340 18500
rect 3380 18460 3381 18500
rect 3339 18451 3381 18460
rect 3340 17417 3380 18451
rect 3436 18332 3476 19216
rect 3532 19256 3572 21316
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 4011 20852 4053 20861
rect 4011 20812 4012 20852
rect 4052 20812 4053 20852
rect 4011 20803 4053 20812
rect 4012 20768 4052 20803
rect 4012 20717 4052 20728
rect 3724 20096 3764 20107
rect 3724 20021 3764 20056
rect 3723 20012 3765 20021
rect 3723 19972 3724 20012
rect 3764 19972 3765 20012
rect 3723 19963 3765 19972
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 3627 19508 3669 19517
rect 3627 19468 3628 19508
rect 3668 19468 3669 19508
rect 3627 19459 3669 19468
rect 3532 19097 3572 19216
rect 3531 19088 3573 19097
rect 3531 19048 3532 19088
rect 3572 19048 3573 19088
rect 3531 19039 3573 19048
rect 3628 18584 3668 19459
rect 4011 19256 4053 19265
rect 4011 19216 4012 19256
rect 4052 19216 4053 19256
rect 4011 19207 4053 19216
rect 4012 18845 4052 19207
rect 4011 18836 4053 18845
rect 4011 18796 4012 18836
rect 4052 18796 4053 18836
rect 4011 18787 4053 18796
rect 3628 18509 3668 18544
rect 4108 18752 4148 21568
rect 4203 21608 4245 21617
rect 4203 21568 4204 21608
rect 4244 21568 4245 21608
rect 4203 21559 4245 21568
rect 4204 21474 4244 21559
rect 4300 19265 4340 22063
rect 4396 19349 4436 23752
rect 4588 20180 4628 27448
rect 4683 26144 4725 26153
rect 4683 26104 4684 26144
rect 4724 26104 4725 26144
rect 4683 26095 4725 26104
rect 4684 22205 4724 26095
rect 4780 23120 4820 27868
rect 5355 27740 5397 27749
rect 5355 27700 5356 27740
rect 5396 27700 5397 27740
rect 5355 27691 5397 27700
rect 4875 27656 4917 27665
rect 4875 27616 4876 27656
rect 4916 27616 4917 27656
rect 4875 27607 4917 27616
rect 4876 27522 4916 27607
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 5163 24632 5205 24641
rect 5163 24592 5164 24632
rect 5204 24592 5205 24632
rect 5163 24583 5205 24592
rect 5164 23801 5204 24583
rect 5259 24548 5301 24557
rect 5259 24508 5260 24548
rect 5300 24508 5301 24548
rect 5259 24499 5301 24508
rect 5163 23792 5205 23801
rect 5163 23752 5164 23792
rect 5204 23752 5205 23792
rect 5163 23743 5205 23752
rect 5260 23717 5300 24499
rect 5259 23708 5301 23717
rect 5259 23668 5260 23708
rect 5300 23668 5301 23708
rect 5259 23659 5301 23668
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 5356 23381 5396 27691
rect 5452 25397 5492 30472
rect 5547 30260 5589 30269
rect 5547 30220 5548 30260
rect 5588 30220 5589 30260
rect 5547 30211 5589 30220
rect 5548 29840 5588 30211
rect 5740 30092 5780 30631
rect 5740 30043 5780 30052
rect 5548 29791 5588 29800
rect 5739 29672 5781 29681
rect 5739 29632 5740 29672
rect 5780 29632 5781 29672
rect 5739 29623 5781 29632
rect 5740 29168 5780 29623
rect 5740 29119 5780 29128
rect 5739 29000 5781 29009
rect 5739 28960 5740 29000
rect 5780 28960 5781 29000
rect 5739 28951 5781 28960
rect 5740 28589 5780 28951
rect 5739 28580 5781 28589
rect 5739 28540 5740 28580
rect 5780 28540 5781 28580
rect 5739 28531 5781 28540
rect 5836 28421 5876 30967
rect 5932 30680 5972 32647
rect 6028 31352 6068 31361
rect 6028 31025 6068 31312
rect 6124 31352 6164 31363
rect 6124 31277 6164 31312
rect 6123 31268 6165 31277
rect 6123 31228 6124 31268
rect 6164 31228 6165 31268
rect 6123 31219 6165 31228
rect 6027 31016 6069 31025
rect 6027 30976 6028 31016
rect 6068 30976 6069 31016
rect 6027 30967 6069 30976
rect 6028 30680 6068 30689
rect 5932 30640 6028 30680
rect 5835 28412 5877 28421
rect 5835 28372 5836 28412
rect 5876 28372 5877 28412
rect 5835 28363 5877 28372
rect 5548 28328 5588 28337
rect 5548 28253 5588 28288
rect 5643 28328 5685 28337
rect 5643 28288 5644 28328
rect 5684 28288 5685 28328
rect 5643 28279 5685 28288
rect 5547 28244 5589 28253
rect 5547 28204 5548 28244
rect 5588 28204 5589 28244
rect 5547 28195 5589 28204
rect 5548 27749 5588 28195
rect 5547 27740 5589 27749
rect 5547 27700 5548 27740
rect 5588 27700 5589 27740
rect 5547 27691 5589 27700
rect 5547 27404 5589 27413
rect 5547 27364 5548 27404
rect 5588 27364 5589 27404
rect 5547 27355 5589 27364
rect 5451 25388 5493 25397
rect 5451 25348 5452 25388
rect 5492 25348 5493 25388
rect 5451 25339 5493 25348
rect 5548 24800 5588 27355
rect 5644 25472 5684 28279
rect 5740 28160 5780 28169
rect 5835 28160 5877 28169
rect 5780 28120 5836 28160
rect 5876 28120 5877 28160
rect 5740 28111 5780 28120
rect 5835 28111 5877 28120
rect 5739 27320 5781 27329
rect 5739 27280 5740 27320
rect 5780 27280 5781 27320
rect 5739 27271 5781 27280
rect 5740 26816 5780 27271
rect 5740 26573 5780 26776
rect 5739 26564 5781 26573
rect 5739 26524 5740 26564
rect 5780 26524 5781 26564
rect 5739 26515 5781 26524
rect 5836 25817 5876 28111
rect 5932 28085 5972 30640
rect 6028 30631 6068 30640
rect 6123 30680 6165 30689
rect 6123 30640 6124 30680
rect 6164 30640 6165 30680
rect 6123 30631 6165 30640
rect 6124 30521 6164 30631
rect 6220 30605 6260 34075
rect 6316 33704 6356 34336
rect 6316 32864 6356 33664
rect 6316 32815 6356 32824
rect 6412 31445 6452 35167
rect 6508 34637 6548 36856
rect 6795 36856 6796 36896
rect 6836 36856 6837 36896
rect 6795 36847 6837 36856
rect 6603 36812 6645 36821
rect 6603 36772 6604 36812
rect 6644 36772 6645 36812
rect 6603 36763 6645 36772
rect 6604 36728 6644 36763
rect 6796 36762 6836 36847
rect 6604 36677 6644 36688
rect 6700 36728 6740 36737
rect 6603 36476 6645 36485
rect 6603 36436 6604 36476
rect 6644 36436 6645 36476
rect 6603 36427 6645 36436
rect 6604 36065 6644 36427
rect 6700 36317 6740 36688
rect 6892 36728 6932 36737
rect 6892 36560 6932 36688
rect 7084 36728 7124 37183
rect 7084 36679 7124 36688
rect 7084 36560 7124 36569
rect 6892 36520 7084 36560
rect 7084 36511 7124 36520
rect 6699 36308 6741 36317
rect 6699 36268 6700 36308
rect 6740 36268 6741 36308
rect 6699 36259 6741 36268
rect 6987 36140 7029 36149
rect 6987 36100 6988 36140
rect 7028 36100 7029 36140
rect 6987 36091 7029 36100
rect 6603 36056 6645 36065
rect 6603 36016 6604 36056
rect 6644 36016 6645 36056
rect 6603 36007 6645 36016
rect 6988 36006 7028 36091
rect 7180 36056 7220 37780
rect 7468 37325 7508 38611
rect 7467 37316 7509 37325
rect 7467 37276 7468 37316
rect 7508 37276 7509 37316
rect 7467 37267 7509 37276
rect 7467 37148 7509 37157
rect 7467 37108 7468 37148
rect 7508 37108 7509 37148
rect 7467 37099 7509 37108
rect 7275 36728 7317 36737
rect 7275 36688 7276 36728
rect 7316 36688 7317 36728
rect 7275 36679 7317 36688
rect 7372 36728 7412 36737
rect 7468 36728 7508 37099
rect 7564 36905 7604 39283
rect 7659 39164 7701 39173
rect 7659 39124 7660 39164
rect 7700 39124 7701 39164
rect 7659 39115 7701 39124
rect 7660 38081 7700 39115
rect 7755 38996 7797 39005
rect 7755 38956 7756 38996
rect 7796 38956 7797 38996
rect 7755 38947 7797 38956
rect 7756 38862 7796 38947
rect 7851 38912 7893 38921
rect 7851 38872 7852 38912
rect 7892 38872 7893 38912
rect 7851 38863 7893 38872
rect 7852 38778 7892 38863
rect 7659 38072 7701 38081
rect 7659 38032 7660 38072
rect 7700 38032 7701 38072
rect 7659 38023 7701 38032
rect 7948 37820 7988 39871
rect 7756 37780 7988 37820
rect 7659 36980 7701 36989
rect 7659 36940 7660 36980
rect 7700 36940 7701 36980
rect 7659 36931 7701 36940
rect 7563 36896 7605 36905
rect 7563 36856 7564 36896
rect 7604 36856 7605 36896
rect 7563 36847 7605 36856
rect 7660 36896 7700 36931
rect 7756 36896 7796 37780
rect 7947 37568 7989 37577
rect 7947 37528 7948 37568
rect 7988 37528 7989 37568
rect 7947 37519 7989 37528
rect 7948 37400 7988 37519
rect 7948 37351 7988 37360
rect 7756 36856 7892 36896
rect 7660 36845 7700 36856
rect 7564 36728 7604 36737
rect 7468 36688 7564 36728
rect 7084 36016 7220 36056
rect 6604 35888 6644 35897
rect 6604 35729 6644 35848
rect 6699 35804 6741 35813
rect 6699 35764 6700 35804
rect 6740 35764 6741 35804
rect 6699 35755 6741 35764
rect 6603 35720 6645 35729
rect 6603 35680 6604 35720
rect 6644 35680 6645 35720
rect 6603 35671 6645 35680
rect 6700 35670 6740 35755
rect 6987 35636 7029 35645
rect 6987 35596 6988 35636
rect 7028 35596 7029 35636
rect 6987 35587 7029 35596
rect 6604 35216 6644 35225
rect 6604 34889 6644 35176
rect 6700 35216 6740 35225
rect 6603 34880 6645 34889
rect 6603 34840 6604 34880
rect 6644 34840 6645 34880
rect 6603 34831 6645 34840
rect 6700 34721 6740 35176
rect 6988 35048 7028 35587
rect 7084 35225 7124 36016
rect 7180 35888 7220 35897
rect 7180 35393 7220 35848
rect 7276 35888 7316 36679
rect 7276 35839 7316 35848
rect 7372 35645 7412 36688
rect 7564 36679 7604 36688
rect 7756 36728 7796 36739
rect 7756 36653 7796 36688
rect 7755 36644 7797 36653
rect 7755 36604 7756 36644
rect 7796 36604 7797 36644
rect 7755 36595 7797 36604
rect 7468 35888 7508 35897
rect 7371 35636 7413 35645
rect 7371 35596 7372 35636
rect 7412 35596 7413 35636
rect 7371 35587 7413 35596
rect 7179 35384 7221 35393
rect 7179 35344 7180 35384
rect 7220 35344 7221 35384
rect 7179 35335 7221 35344
rect 7468 35309 7508 35848
rect 7563 35888 7605 35897
rect 7563 35848 7564 35888
rect 7604 35848 7605 35888
rect 7563 35839 7605 35848
rect 7755 35888 7797 35897
rect 7755 35848 7756 35888
rect 7796 35848 7797 35888
rect 7755 35839 7797 35848
rect 7564 35754 7604 35839
rect 7756 35754 7796 35839
rect 7467 35300 7509 35309
rect 7467 35260 7468 35300
rect 7508 35260 7509 35300
rect 7467 35251 7509 35260
rect 7083 35216 7125 35225
rect 7083 35176 7084 35216
rect 7124 35176 7125 35216
rect 7083 35167 7125 35176
rect 7180 35216 7220 35225
rect 6988 34999 7028 35008
rect 6699 34712 6741 34721
rect 6699 34672 6700 34712
rect 6740 34672 6741 34712
rect 6699 34663 6741 34672
rect 6507 34628 6549 34637
rect 6507 34588 6508 34628
rect 6548 34588 6549 34628
rect 6507 34579 6549 34588
rect 7180 34553 7220 35176
rect 7276 34964 7316 34973
rect 7179 34544 7221 34553
rect 6604 34504 7028 34544
rect 6508 34376 6548 34385
rect 6508 34049 6548 34336
rect 6604 34376 6644 34504
rect 6604 34327 6644 34336
rect 6796 34376 6836 34385
rect 6988 34376 7028 34504
rect 7179 34504 7180 34544
rect 7220 34504 7221 34544
rect 7179 34495 7221 34504
rect 6836 34336 6932 34376
rect 6796 34327 6836 34336
rect 6699 34292 6741 34301
rect 6699 34252 6700 34292
rect 6740 34252 6741 34292
rect 6699 34243 6741 34252
rect 6700 34158 6740 34243
rect 6795 34208 6837 34217
rect 6795 34168 6796 34208
rect 6836 34168 6837 34208
rect 6795 34159 6837 34168
rect 6507 34040 6549 34049
rect 6507 34000 6508 34040
rect 6548 34000 6549 34040
rect 6507 33991 6549 34000
rect 6507 33788 6549 33797
rect 6507 33748 6508 33788
rect 6548 33748 6549 33788
rect 6507 33739 6549 33748
rect 6508 32873 6548 33739
rect 6604 33704 6644 33713
rect 6604 33545 6644 33664
rect 6700 33704 6740 33713
rect 6603 33536 6645 33545
rect 6603 33496 6604 33536
rect 6644 33496 6645 33536
rect 6603 33487 6645 33496
rect 6603 33284 6645 33293
rect 6603 33244 6604 33284
rect 6644 33244 6645 33284
rect 6603 33235 6645 33244
rect 6507 32864 6549 32873
rect 6507 32824 6508 32864
rect 6548 32824 6549 32864
rect 6507 32815 6549 32824
rect 6604 32864 6644 33235
rect 6700 32948 6740 33664
rect 6796 33368 6836 34159
rect 6892 33956 6932 34336
rect 6988 34327 7028 34336
rect 7083 34376 7125 34385
rect 7083 34336 7084 34376
rect 7124 34336 7125 34376
rect 7083 34327 7125 34336
rect 7180 34376 7220 34385
rect 7084 34242 7124 34327
rect 7180 34133 7220 34336
rect 7276 34376 7316 34924
rect 7659 34880 7701 34889
rect 7659 34840 7660 34880
rect 7700 34840 7701 34880
rect 7659 34831 7701 34840
rect 7563 34376 7605 34385
rect 7316 34336 7508 34376
rect 7276 34327 7316 34336
rect 7179 34124 7221 34133
rect 7179 34084 7180 34124
rect 7220 34084 7221 34124
rect 7179 34075 7221 34084
rect 6892 33916 7412 33956
rect 7372 33872 7412 33916
rect 7468 33881 7508 34336
rect 7563 34336 7564 34376
rect 7604 34336 7605 34376
rect 7563 34327 7605 34336
rect 7564 34242 7604 34327
rect 7660 34301 7700 34831
rect 7659 34292 7701 34301
rect 7659 34252 7660 34292
rect 7700 34252 7701 34292
rect 7659 34243 7701 34252
rect 7563 34040 7605 34049
rect 7563 34000 7564 34040
rect 7604 34000 7605 34040
rect 7563 33991 7605 34000
rect 7372 33823 7412 33832
rect 7467 33872 7509 33881
rect 7467 33832 7468 33872
rect 7508 33832 7509 33872
rect 7467 33823 7509 33832
rect 7180 33704 7220 33713
rect 6988 33536 7028 33545
rect 7180 33536 7220 33664
rect 7275 33704 7317 33713
rect 7468 33704 7508 33713
rect 7275 33664 7276 33704
rect 7316 33664 7317 33704
rect 7275 33655 7317 33664
rect 7372 33664 7468 33704
rect 7276 33570 7316 33655
rect 7028 33496 7220 33536
rect 6988 33487 7028 33496
rect 6796 33328 7316 33368
rect 6987 33116 7029 33125
rect 6987 33076 6988 33116
rect 7028 33076 7029 33116
rect 6987 33067 7029 33076
rect 6988 32982 7028 33067
rect 7179 32948 7221 32957
rect 6700 32908 6836 32948
rect 6604 32815 6644 32824
rect 6700 32780 6740 32789
rect 6603 31520 6645 31529
rect 6603 31480 6604 31520
rect 6644 31480 6645 31520
rect 6603 31471 6645 31480
rect 6411 31436 6453 31445
rect 6411 31396 6412 31436
rect 6452 31396 6453 31436
rect 6411 31387 6453 31396
rect 6507 31352 6549 31361
rect 6507 31312 6508 31352
rect 6548 31312 6549 31352
rect 6507 31303 6549 31312
rect 6604 31352 6644 31471
rect 6604 31303 6644 31312
rect 6219 30596 6261 30605
rect 6219 30556 6220 30596
rect 6260 30556 6261 30596
rect 6219 30547 6261 30556
rect 6123 30512 6165 30521
rect 6123 30472 6124 30512
rect 6164 30472 6165 30512
rect 6123 30463 6165 30472
rect 6508 30269 6548 31303
rect 6603 31016 6645 31025
rect 6603 30976 6604 31016
rect 6644 30976 6645 31016
rect 6603 30967 6645 30976
rect 6604 30353 6644 30967
rect 6603 30344 6645 30353
rect 6603 30304 6604 30344
rect 6644 30304 6645 30344
rect 6603 30295 6645 30304
rect 6507 30260 6549 30269
rect 6507 30220 6508 30260
rect 6548 30220 6549 30260
rect 6507 30211 6549 30220
rect 6316 29840 6356 29849
rect 6220 29672 6260 29681
rect 6124 29632 6220 29672
rect 6027 29168 6069 29177
rect 6027 29128 6028 29168
rect 6068 29128 6069 29168
rect 6027 29119 6069 29128
rect 6124 29168 6164 29632
rect 6220 29623 6260 29632
rect 6316 29168 6356 29800
rect 6412 29840 6452 29849
rect 6412 29672 6452 29800
rect 6508 29840 6548 29849
rect 6604 29840 6644 30295
rect 6700 30185 6740 32740
rect 6796 31865 6836 32908
rect 7179 32908 7180 32948
rect 7220 32908 7221 32948
rect 7179 32899 7221 32908
rect 7180 32864 7220 32899
rect 7180 32813 7220 32824
rect 7276 32864 7316 33328
rect 7372 33200 7412 33664
rect 7468 33655 7508 33664
rect 7564 33536 7604 33991
rect 7852 33872 7892 36856
rect 7756 33832 7892 33872
rect 7659 33788 7701 33797
rect 7659 33748 7660 33788
rect 7700 33748 7701 33788
rect 7659 33739 7701 33748
rect 7660 33704 7700 33739
rect 7660 33653 7700 33664
rect 7660 33536 7700 33545
rect 7564 33496 7660 33536
rect 7660 33487 7700 33496
rect 7372 33160 7508 33200
rect 7276 32815 7316 32824
rect 7371 32864 7413 32873
rect 7371 32824 7372 32864
rect 7412 32824 7413 32864
rect 7371 32815 7413 32824
rect 7468 32864 7508 33160
rect 7756 33032 7796 33832
rect 7851 33704 7893 33713
rect 7851 33664 7852 33704
rect 7892 33664 7893 33704
rect 7851 33655 7893 33664
rect 7948 33704 7988 33713
rect 7852 33570 7892 33655
rect 7851 33452 7893 33461
rect 7851 33412 7852 33452
rect 7892 33412 7893 33452
rect 7851 33403 7893 33412
rect 7468 32815 7508 32824
rect 7660 32992 7796 33032
rect 7083 32780 7125 32789
rect 7083 32740 7084 32780
rect 7124 32740 7125 32780
rect 7083 32731 7125 32740
rect 6988 32192 7028 32201
rect 6891 32024 6933 32033
rect 6891 31984 6892 32024
rect 6932 31984 6933 32024
rect 6891 31975 6933 31984
rect 6795 31856 6837 31865
rect 6795 31816 6796 31856
rect 6836 31816 6837 31856
rect 6795 31807 6837 31816
rect 6795 31520 6837 31529
rect 6795 31480 6796 31520
rect 6836 31480 6837 31520
rect 6795 31471 6837 31480
rect 6796 30269 6836 31471
rect 6795 30260 6837 30269
rect 6795 30220 6796 30260
rect 6836 30220 6837 30260
rect 6795 30211 6837 30220
rect 6699 30176 6741 30185
rect 6699 30136 6700 30176
rect 6740 30136 6741 30176
rect 6699 30127 6741 30136
rect 6548 29800 6644 29840
rect 6700 29840 6740 29849
rect 6508 29791 6548 29800
rect 6700 29672 6740 29800
rect 6412 29632 6740 29672
rect 6796 29672 6836 29681
rect 6412 29252 6452 29632
rect 6603 29504 6645 29513
rect 6603 29464 6604 29504
rect 6644 29464 6645 29504
rect 6603 29455 6645 29464
rect 6604 29252 6644 29455
rect 6699 29336 6741 29345
rect 6699 29296 6700 29336
rect 6740 29296 6741 29336
rect 6699 29287 6741 29296
rect 6412 29212 6548 29252
rect 6124 29119 6164 29128
rect 6220 29128 6356 29168
rect 6028 29034 6068 29119
rect 6220 28916 6260 29128
rect 6411 29084 6453 29093
rect 6028 28876 6260 28916
rect 6316 29044 6412 29084
rect 6452 29044 6453 29084
rect 6316 28916 6356 29044
rect 6411 29035 6453 29044
rect 6508 29009 6548 29212
rect 6604 29203 6644 29212
rect 6700 29168 6740 29287
rect 6700 29119 6740 29128
rect 6507 29000 6549 29009
rect 6796 29000 6836 29632
rect 6892 29513 6932 31975
rect 6988 31949 7028 32152
rect 6987 31940 7029 31949
rect 6987 31900 6988 31940
rect 7028 31900 7029 31940
rect 6987 31891 7029 31900
rect 6987 31604 7029 31613
rect 7084 31604 7124 32731
rect 7372 32730 7412 32815
rect 7467 32696 7509 32705
rect 7467 32656 7468 32696
rect 7508 32656 7509 32696
rect 7467 32647 7509 32656
rect 6987 31564 6988 31604
rect 7028 31564 7124 31604
rect 7180 31940 7220 31949
rect 6987 31555 7029 31564
rect 6891 29504 6933 29513
rect 6891 29464 6892 29504
rect 6932 29464 6933 29504
rect 6891 29455 6933 29464
rect 6988 29429 7028 31555
rect 7180 31520 7220 31900
rect 7084 31480 7220 31520
rect 7468 31520 7508 32647
rect 7660 32192 7700 32992
rect 7756 32864 7796 32873
rect 7852 32864 7892 33403
rect 7948 33125 7988 33664
rect 8044 33209 8084 40039
rect 8139 39416 8181 39425
rect 8139 39376 8140 39416
rect 8180 39376 8181 39416
rect 8139 39367 8181 39376
rect 8140 37820 8180 39367
rect 8236 38912 8276 40207
rect 8428 40097 8468 40879
rect 8523 40508 8565 40517
rect 8523 40468 8524 40508
rect 8564 40468 8565 40508
rect 8523 40459 8565 40468
rect 8524 40424 8564 40459
rect 8524 40373 8564 40384
rect 8620 40424 8660 40433
rect 8716 40424 8756 41215
rect 8812 40433 8852 41224
rect 8908 41264 8948 41273
rect 8908 40685 8948 41224
rect 9003 41264 9045 41273
rect 9003 41224 9004 41264
rect 9044 41224 9045 41264
rect 9003 41215 9045 41224
rect 9100 41264 9140 41273
rect 9004 41130 9044 41215
rect 9100 40844 9140 41224
rect 9195 41264 9237 41273
rect 9195 41224 9196 41264
rect 9236 41224 9237 41264
rect 9195 41215 9237 41224
rect 9292 41264 9332 41273
rect 9004 40804 9140 40844
rect 8907 40676 8949 40685
rect 8907 40636 8908 40676
rect 8948 40636 8949 40676
rect 8907 40627 8949 40636
rect 8908 40517 8948 40548
rect 8907 40508 8949 40517
rect 8907 40468 8908 40508
rect 8948 40468 8949 40508
rect 8907 40459 8949 40468
rect 8660 40384 8756 40424
rect 8811 40424 8853 40433
rect 8811 40384 8812 40424
rect 8852 40384 8853 40424
rect 8620 40375 8660 40384
rect 8811 40375 8853 40384
rect 8908 40424 8948 40459
rect 8908 40256 8948 40384
rect 9004 40265 9044 40804
rect 9100 40601 9140 40686
rect 9099 40592 9141 40601
rect 9099 40552 9100 40592
rect 9140 40552 9141 40592
rect 9099 40543 9141 40552
rect 9100 40424 9140 40433
rect 9196 40424 9236 41215
rect 9292 41189 9332 41224
rect 9291 41180 9333 41189
rect 9291 41140 9292 41180
rect 9332 41140 9333 41180
rect 9291 41131 9333 41140
rect 9292 40433 9332 41131
rect 9140 40384 9236 40424
rect 9100 40375 9140 40384
rect 8812 40216 8948 40256
rect 9003 40256 9045 40265
rect 9003 40216 9004 40256
rect 9044 40216 9045 40256
rect 8427 40088 8469 40097
rect 8427 40048 8428 40088
rect 8468 40048 8469 40088
rect 8427 40039 8469 40048
rect 8331 39920 8373 39929
rect 8331 39880 8332 39920
rect 8372 39880 8373 39920
rect 8331 39871 8373 39880
rect 8332 39752 8372 39871
rect 8428 39845 8468 40039
rect 8523 39920 8565 39929
rect 8523 39880 8524 39920
rect 8564 39880 8565 39920
rect 8523 39871 8565 39880
rect 8427 39836 8469 39845
rect 8427 39796 8428 39836
rect 8468 39796 8469 39836
rect 8427 39787 8469 39796
rect 8332 39703 8372 39712
rect 8524 39677 8564 39871
rect 8812 39738 8852 40216
rect 9003 40207 9045 40216
rect 8907 40088 8949 40097
rect 8907 40048 8908 40088
rect 8948 40048 8949 40088
rect 8907 40039 8949 40048
rect 8523 39668 8565 39677
rect 8523 39628 8524 39668
rect 8564 39628 8565 39668
rect 8523 39619 8565 39628
rect 8331 38912 8373 38921
rect 8236 38872 8332 38912
rect 8372 38872 8373 38912
rect 8331 38863 8373 38872
rect 8332 38778 8372 38863
rect 8140 37780 8276 37820
rect 8139 37232 8181 37241
rect 8139 37192 8140 37232
rect 8180 37192 8181 37232
rect 8139 37183 8181 37192
rect 8140 37098 8180 37183
rect 8139 36896 8181 36905
rect 8139 36856 8140 36896
rect 8180 36856 8181 36896
rect 8139 36847 8181 36856
rect 8043 33200 8085 33209
rect 8043 33160 8044 33200
rect 8084 33160 8085 33200
rect 8043 33151 8085 33160
rect 7947 33116 7989 33125
rect 7947 33076 7948 33116
rect 7988 33076 7989 33116
rect 7947 33067 7989 33076
rect 8140 32948 8180 36847
rect 8236 33881 8276 37780
rect 8331 37484 8373 37493
rect 8331 37444 8332 37484
rect 8372 37444 8373 37484
rect 8331 37435 8373 37444
rect 8332 37400 8372 37435
rect 8332 37349 8372 37360
rect 8331 37232 8373 37241
rect 8331 37192 8332 37232
rect 8372 37192 8373 37232
rect 8331 37183 8373 37192
rect 8332 36728 8372 37183
rect 8332 36679 8372 36688
rect 8428 36728 8468 36737
rect 8428 36149 8468 36688
rect 8427 36140 8469 36149
rect 8427 36100 8428 36140
rect 8468 36100 8469 36140
rect 8427 36091 8469 36100
rect 8428 35729 8468 36091
rect 8427 35720 8469 35729
rect 8427 35680 8428 35720
rect 8468 35680 8469 35720
rect 8427 35671 8469 35680
rect 8524 34385 8564 39619
rect 8812 38926 8852 39698
rect 8619 38912 8661 38921
rect 8619 38872 8620 38912
rect 8660 38872 8661 38912
rect 8812 38877 8852 38886
rect 8619 38863 8661 38872
rect 8620 35309 8660 38863
rect 8908 37820 8948 40039
rect 9196 40004 9236 40384
rect 9291 40424 9333 40433
rect 9291 40384 9292 40424
rect 9332 40384 9333 40424
rect 9291 40375 9333 40384
rect 9291 40256 9333 40265
rect 9291 40216 9292 40256
rect 9332 40216 9333 40256
rect 9291 40207 9333 40216
rect 9292 40122 9332 40207
rect 9388 40088 9428 41392
rect 9484 41264 9524 41273
rect 9484 40433 9524 41224
rect 9580 41264 9620 41273
rect 9580 41021 9620 41224
rect 9579 41012 9621 41021
rect 9579 40972 9580 41012
rect 9620 40972 9621 41012
rect 9579 40963 9621 40972
rect 9676 40844 9716 41551
rect 9772 41357 9812 41728
rect 10060 41693 10100 47095
rect 10252 46397 10292 47860
rect 10444 47816 10484 47825
rect 10348 47776 10444 47816
rect 10348 47312 10388 47776
rect 10444 47767 10484 47776
rect 10348 47263 10388 47272
rect 10444 47312 10484 47321
rect 10444 46985 10484 47272
rect 10443 46976 10485 46985
rect 10443 46936 10444 46976
rect 10484 46936 10485 46976
rect 10443 46927 10485 46936
rect 10251 46388 10293 46397
rect 10251 46348 10252 46388
rect 10292 46348 10293 46388
rect 10251 46339 10293 46348
rect 10252 45893 10292 46339
rect 10251 45884 10293 45893
rect 10251 45844 10252 45884
rect 10292 45844 10293 45884
rect 10251 45835 10293 45844
rect 10348 45800 10388 45809
rect 10348 45641 10388 45760
rect 10347 45632 10389 45641
rect 10347 45592 10348 45632
rect 10388 45592 10389 45632
rect 10347 45583 10389 45592
rect 10156 45548 10196 45557
rect 10156 44960 10196 45508
rect 10444 45137 10484 46927
rect 10443 45128 10485 45137
rect 10443 45088 10444 45128
rect 10484 45088 10485 45128
rect 10443 45079 10485 45088
rect 10156 44911 10196 44920
rect 10252 44960 10292 44969
rect 10540 44960 10580 48616
rect 10924 47993 10964 49288
rect 11019 49160 11061 49169
rect 11019 49120 11020 49160
rect 11060 49120 11061 49160
rect 11019 49111 11061 49120
rect 10923 47984 10965 47993
rect 10923 47944 10924 47984
rect 10964 47944 10965 47984
rect 10923 47935 10965 47944
rect 11020 47984 11060 49111
rect 11020 47935 11060 47944
rect 11116 47816 11156 49624
rect 11212 49496 11252 50371
rect 11212 49253 11252 49456
rect 11211 49244 11253 49253
rect 11211 49204 11212 49244
rect 11252 49204 11253 49244
rect 11211 49195 11253 49204
rect 11211 48908 11253 48917
rect 11211 48868 11212 48908
rect 11252 48868 11253 48908
rect 11211 48859 11253 48868
rect 11212 48749 11252 48859
rect 11211 48740 11253 48749
rect 11211 48700 11212 48740
rect 11252 48700 11253 48740
rect 11211 48691 11253 48700
rect 11211 47900 11253 47909
rect 11211 47860 11212 47900
rect 11252 47860 11253 47900
rect 11211 47851 11253 47860
rect 10732 47776 11156 47816
rect 10732 45044 10772 47776
rect 11019 47648 11061 47657
rect 11019 47608 11020 47648
rect 11060 47608 11061 47648
rect 11019 47599 11061 47608
rect 10923 47312 10965 47321
rect 10923 47272 10924 47312
rect 10964 47272 10965 47312
rect 10923 47263 10965 47272
rect 10827 47228 10869 47237
rect 10827 47188 10828 47228
rect 10868 47188 10869 47228
rect 10827 47179 10869 47188
rect 10828 47094 10868 47179
rect 10924 47178 10964 47263
rect 10923 46472 10965 46481
rect 10923 46432 10924 46472
rect 10964 46432 10965 46472
rect 10923 46423 10965 46432
rect 10924 45641 10964 46423
rect 10923 45632 10965 45641
rect 10923 45592 10924 45632
rect 10964 45592 10965 45632
rect 10923 45583 10965 45592
rect 10732 44995 10772 45004
rect 10292 44920 10580 44960
rect 10635 44960 10677 44969
rect 10635 44920 10636 44960
rect 10676 44920 10677 44960
rect 10252 44456 10292 44920
rect 10635 44911 10677 44920
rect 10636 44826 10676 44911
rect 10156 44416 10292 44456
rect 10156 44120 10196 44416
rect 10252 44288 10292 44297
rect 11020 44288 11060 47599
rect 10292 44248 11060 44288
rect 11212 44960 11252 47851
rect 10252 44239 10292 44248
rect 10156 44080 10388 44120
rect 10059 41684 10101 41693
rect 10059 41644 10060 41684
rect 10100 41644 10101 41684
rect 10059 41635 10101 41644
rect 10251 41600 10293 41609
rect 10251 41560 10252 41600
rect 10292 41560 10293 41600
rect 10251 41551 10293 41560
rect 10252 41432 10292 41551
rect 10252 41383 10292 41392
rect 9771 41348 9813 41357
rect 9771 41308 9772 41348
rect 9812 41308 9813 41348
rect 9771 41299 9813 41308
rect 9963 41348 10005 41357
rect 9963 41308 9964 41348
rect 10004 41308 10005 41348
rect 9963 41299 10005 41308
rect 9867 41264 9909 41273
rect 9867 41224 9868 41264
rect 9908 41224 9909 41264
rect 9867 41215 9909 41224
rect 9964 41264 10004 41299
rect 9868 41096 9908 41215
rect 9964 41213 10004 41224
rect 10060 41264 10100 41273
rect 9868 41056 10004 41096
rect 9771 41012 9813 41021
rect 9771 40972 9772 41012
rect 9812 40972 9813 41012
rect 9771 40963 9813 40972
rect 9580 40804 9716 40844
rect 9483 40424 9525 40433
rect 9483 40384 9484 40424
rect 9524 40384 9525 40424
rect 9483 40375 9525 40384
rect 9580 40424 9620 40804
rect 9675 40676 9717 40685
rect 9675 40636 9676 40676
rect 9716 40636 9717 40676
rect 9675 40627 9717 40636
rect 9676 40508 9716 40627
rect 9772 40592 9812 40963
rect 9964 40685 10004 41056
rect 10060 40769 10100 41224
rect 10251 41264 10293 41273
rect 10251 41224 10252 41264
rect 10292 41224 10293 41264
rect 10251 41215 10293 41224
rect 10059 40760 10101 40769
rect 10059 40720 10060 40760
rect 10100 40720 10101 40760
rect 10059 40711 10101 40720
rect 9963 40676 10005 40685
rect 9963 40636 9964 40676
rect 10004 40636 10005 40676
rect 9963 40627 10005 40636
rect 9772 40543 9812 40552
rect 9867 40592 9909 40601
rect 9867 40552 9868 40592
rect 9908 40552 9909 40592
rect 9867 40543 9909 40552
rect 9676 40459 9716 40468
rect 9868 40508 9908 40543
rect 9868 40457 9908 40468
rect 9580 40265 9620 40384
rect 9964 40424 10004 40627
rect 10059 40592 10101 40601
rect 10059 40552 10060 40592
rect 10100 40552 10101 40592
rect 10059 40543 10101 40552
rect 9964 40375 10004 40384
rect 9579 40256 9621 40265
rect 9579 40216 9580 40256
rect 9620 40216 9621 40256
rect 9579 40207 9621 40216
rect 9483 40088 9525 40097
rect 9388 40048 9484 40088
rect 9524 40048 9525 40088
rect 9483 40039 9525 40048
rect 9196 39964 9427 40004
rect 9004 39920 9044 39929
rect 9387 39920 9427 39964
rect 9044 39880 9236 39920
rect 9387 39880 9428 39920
rect 9004 39871 9044 39880
rect 9196 39677 9236 39880
rect 9388 39752 9428 39880
rect 9772 39836 9812 39845
rect 9812 39796 9908 39836
rect 9772 39787 9812 39796
rect 9676 39752 9716 39761
rect 9388 39703 9428 39712
rect 9484 39712 9676 39752
rect 9195 39668 9237 39677
rect 9195 39628 9196 39668
rect 9236 39628 9237 39668
rect 9195 39619 9237 39628
rect 9004 38828 9044 38837
rect 9484 38828 9524 39712
rect 9676 39703 9716 39712
rect 9771 39668 9813 39677
rect 9771 39628 9772 39668
rect 9812 39628 9813 39668
rect 9771 39619 9813 39628
rect 9579 39584 9621 39593
rect 9579 39544 9580 39584
rect 9620 39544 9621 39584
rect 9579 39535 9621 39544
rect 9580 38912 9620 39535
rect 9675 39332 9717 39341
rect 9675 39292 9676 39332
rect 9716 39292 9717 39332
rect 9675 39283 9717 39292
rect 9580 38863 9620 38872
rect 9044 38788 9524 38828
rect 9004 38779 9044 38788
rect 9291 38492 9333 38501
rect 9291 38452 9292 38492
rect 9332 38452 9333 38492
rect 9291 38443 9333 38452
rect 9292 38240 9332 38443
rect 9292 38191 9332 38200
rect 8908 37780 9044 37820
rect 8715 37652 8757 37661
rect 8715 37612 8716 37652
rect 8756 37612 8757 37652
rect 8715 37603 8757 37612
rect 8716 37409 8756 37603
rect 8715 37400 8757 37409
rect 8715 37360 8716 37400
rect 8756 37360 8757 37400
rect 8715 37351 8757 37360
rect 8716 36644 8756 37351
rect 8812 36644 8852 36653
rect 8716 36604 8812 36644
rect 8619 35300 8661 35309
rect 8619 35260 8620 35300
rect 8660 35260 8661 35300
rect 8619 35251 8661 35260
rect 8523 34376 8565 34385
rect 8523 34336 8524 34376
rect 8564 34336 8565 34376
rect 8523 34327 8565 34336
rect 8716 34049 8756 36604
rect 8812 36595 8852 36604
rect 8907 36644 8949 36653
rect 8907 36604 8908 36644
rect 8948 36604 8949 36644
rect 8907 36595 8949 36604
rect 8908 36510 8948 36595
rect 9004 36140 9044 37780
rect 9579 37568 9621 37577
rect 9579 37528 9580 37568
rect 9620 37528 9621 37568
rect 9579 37519 9621 37528
rect 9580 37400 9620 37519
rect 9580 37351 9620 37360
rect 9388 36728 9428 36737
rect 9676 36728 9716 39283
rect 9772 39080 9812 39619
rect 9868 39593 9908 39796
rect 10060 39738 10100 40543
rect 10252 40517 10292 41215
rect 10348 40601 10388 44080
rect 10923 43532 10965 43541
rect 10923 43492 10924 43532
rect 10964 43492 10965 43532
rect 10923 43483 10965 43492
rect 10924 42776 10964 43483
rect 10924 42727 10964 42736
rect 11115 42188 11157 42197
rect 11115 42148 11116 42188
rect 11156 42148 11157 42188
rect 11115 42139 11157 42148
rect 11116 41945 11156 42139
rect 11115 41936 11157 41945
rect 11115 41896 11116 41936
rect 11156 41896 11157 41936
rect 11115 41887 11157 41896
rect 11116 41802 11156 41887
rect 11212 41861 11252 44920
rect 11308 42701 11348 53143
rect 11692 52109 11732 53320
rect 11691 52100 11733 52109
rect 11691 52060 11692 52100
rect 11732 52060 11733 52100
rect 11691 52051 11733 52060
rect 11692 51932 11732 51941
rect 11404 51892 11692 51932
rect 11404 51101 11444 51892
rect 11692 51883 11732 51892
rect 11500 51834 11540 51843
rect 11500 51353 11540 51794
rect 11788 51596 11828 53488
rect 11884 53033 11924 54412
rect 11979 54284 12021 54293
rect 11979 54244 11980 54284
rect 12020 54244 12021 54284
rect 11979 54235 12021 54244
rect 11883 53024 11925 53033
rect 11883 52984 11884 53024
rect 11924 52984 11925 53024
rect 11883 52975 11925 52984
rect 11596 51556 11828 51596
rect 11499 51344 11541 51353
rect 11499 51304 11500 51344
rect 11540 51304 11541 51344
rect 11499 51295 11541 51304
rect 11596 51176 11636 51556
rect 11788 51269 11828 51354
rect 11787 51260 11829 51269
rect 11787 51220 11788 51260
rect 11828 51220 11829 51260
rect 11787 51211 11829 51220
rect 11500 51136 11636 51176
rect 11403 51092 11445 51101
rect 11403 51052 11404 51092
rect 11444 51052 11445 51092
rect 11403 51043 11445 51052
rect 11403 50588 11445 50597
rect 11403 50548 11404 50588
rect 11444 50548 11445 50588
rect 11403 50539 11445 50548
rect 11404 49169 11444 50539
rect 11403 49160 11445 49169
rect 11403 49120 11404 49160
rect 11444 49120 11445 49160
rect 11403 49111 11445 49120
rect 11500 48992 11540 51136
rect 11787 51092 11829 51101
rect 11787 51052 11788 51092
rect 11828 51052 11829 51092
rect 11787 51043 11829 51052
rect 11404 48952 11540 48992
rect 11596 51008 11636 51017
rect 11404 47405 11444 48952
rect 11596 48833 11636 50968
rect 11691 50672 11733 50681
rect 11691 50632 11692 50672
rect 11732 50632 11733 50672
rect 11691 50623 11733 50632
rect 11595 48824 11637 48833
rect 11595 48784 11596 48824
rect 11636 48784 11637 48824
rect 11595 48775 11637 48784
rect 11596 48245 11636 48775
rect 11595 48236 11637 48245
rect 11595 48196 11596 48236
rect 11636 48196 11637 48236
rect 11595 48187 11637 48196
rect 11403 47396 11445 47405
rect 11403 47356 11404 47396
rect 11444 47356 11445 47396
rect 11403 47347 11445 47356
rect 11404 47312 11444 47347
rect 11404 47262 11444 47272
rect 11692 47153 11732 50623
rect 11788 48572 11828 51043
rect 11884 50093 11924 52975
rect 11980 52277 12020 54235
rect 12172 54116 12212 55579
rect 12268 54293 12308 56671
rect 12364 56384 12404 57763
rect 12364 56335 12404 56344
rect 12363 56216 12405 56225
rect 12363 56176 12364 56216
rect 12404 56176 12405 56216
rect 12363 56167 12405 56176
rect 12364 55637 12404 56167
rect 12363 55628 12405 55637
rect 12363 55588 12364 55628
rect 12404 55588 12405 55628
rect 12363 55579 12405 55588
rect 12363 55460 12405 55469
rect 12363 55420 12364 55460
rect 12404 55420 12405 55460
rect 12363 55411 12405 55420
rect 12267 54284 12309 54293
rect 12267 54244 12268 54284
rect 12308 54244 12309 54284
rect 12267 54235 12309 54244
rect 12172 54076 12308 54116
rect 12075 53528 12117 53537
rect 12075 53488 12076 53528
rect 12116 53488 12117 53528
rect 12075 53479 12117 53488
rect 12076 53360 12116 53479
rect 12076 53311 12116 53320
rect 12171 53276 12213 53285
rect 12171 53236 12172 53276
rect 12212 53236 12213 53276
rect 12171 53227 12213 53236
rect 12172 53142 12212 53227
rect 12268 53024 12308 54076
rect 12172 52984 12308 53024
rect 11979 52268 12021 52277
rect 11979 52228 11980 52268
rect 12020 52228 12021 52268
rect 11979 52219 12021 52228
rect 12075 51680 12117 51689
rect 12075 51640 12076 51680
rect 12116 51640 12117 51680
rect 12075 51631 12117 51640
rect 12076 51017 12116 51631
rect 12172 51101 12212 52984
rect 12268 51848 12308 51857
rect 12268 51605 12308 51808
rect 12267 51596 12309 51605
rect 12267 51556 12268 51596
rect 12308 51556 12309 51596
rect 12267 51547 12309 51556
rect 12171 51092 12213 51101
rect 12171 51052 12172 51092
rect 12212 51052 12213 51092
rect 12171 51043 12213 51052
rect 12075 51008 12117 51017
rect 12075 50968 12076 51008
rect 12116 50968 12117 51008
rect 12075 50959 12117 50968
rect 11979 50588 12021 50597
rect 11979 50548 11980 50588
rect 12020 50548 12021 50588
rect 11979 50539 12021 50548
rect 11883 50084 11925 50093
rect 11883 50044 11884 50084
rect 11924 50044 11925 50084
rect 11883 50035 11925 50044
rect 11980 49673 12020 50539
rect 12076 50336 12116 50959
rect 12268 50765 12308 51547
rect 12267 50756 12309 50765
rect 12267 50716 12268 50756
rect 12308 50716 12309 50756
rect 12267 50707 12309 50716
rect 12364 50597 12404 55411
rect 12363 50588 12405 50597
rect 12363 50548 12364 50588
rect 12404 50548 12405 50588
rect 12363 50539 12405 50548
rect 12460 50504 12500 59368
rect 12556 59359 12596 59368
rect 12651 59408 12693 59417
rect 12651 59368 12652 59408
rect 12692 59368 12693 59408
rect 12651 59359 12693 59368
rect 12844 59408 12884 59527
rect 13036 59442 13076 59527
rect 12844 59359 12884 59368
rect 12652 59274 12692 59359
rect 12940 58652 12980 58661
rect 12747 58400 12789 58409
rect 12747 58360 12748 58400
rect 12788 58360 12789 58400
rect 12747 58351 12789 58360
rect 12748 58266 12788 58351
rect 12651 58064 12693 58073
rect 12651 58024 12652 58064
rect 12692 58024 12693 58064
rect 12651 58015 12693 58024
rect 12555 57392 12597 57401
rect 12555 57352 12556 57392
rect 12596 57352 12597 57392
rect 12555 57343 12597 57352
rect 12556 57056 12596 57343
rect 12556 57007 12596 57016
rect 12555 56468 12597 56477
rect 12555 56428 12556 56468
rect 12596 56428 12597 56468
rect 12555 56419 12597 56428
rect 12556 56225 12596 56419
rect 12555 56216 12597 56225
rect 12555 56176 12556 56216
rect 12596 56176 12597 56216
rect 12555 56167 12597 56176
rect 12555 55964 12597 55973
rect 12555 55924 12556 55964
rect 12596 55924 12597 55964
rect 12555 55915 12597 55924
rect 12556 55544 12596 55915
rect 12556 55495 12596 55504
rect 12652 53705 12692 58015
rect 12747 57980 12789 57989
rect 12747 57940 12748 57980
rect 12788 57940 12789 57980
rect 12747 57931 12789 57940
rect 12651 53696 12693 53705
rect 12651 53656 12652 53696
rect 12692 53656 12693 53696
rect 12651 53647 12693 53656
rect 12652 53360 12692 53647
rect 12652 53311 12692 53320
rect 12651 53192 12693 53201
rect 12651 53152 12652 53192
rect 12692 53152 12693 53192
rect 12651 53143 12693 53152
rect 12652 51008 12692 53143
rect 12748 51185 12788 57931
rect 12940 56972 12980 58612
rect 13132 58073 13172 66760
rect 13228 66725 13268 67012
rect 13227 66716 13269 66725
rect 13227 66676 13228 66716
rect 13268 66676 13269 66716
rect 13227 66667 13269 66676
rect 13228 66389 13268 66667
rect 13227 66380 13269 66389
rect 13227 66340 13228 66380
rect 13268 66340 13269 66380
rect 13227 66331 13269 66340
rect 13516 64280 13556 68104
rect 13611 67724 13653 67733
rect 13611 67684 13612 67724
rect 13652 67684 13653 67724
rect 13611 67675 13653 67684
rect 13612 67640 13652 67675
rect 13612 67589 13652 67600
rect 13516 64240 13652 64280
rect 13515 63944 13557 63953
rect 13515 63904 13516 63944
rect 13556 63904 13557 63944
rect 13515 63895 13557 63904
rect 13516 63810 13556 63895
rect 13323 63692 13365 63701
rect 13323 63652 13324 63692
rect 13364 63652 13365 63692
rect 13323 63643 13365 63652
rect 13324 63118 13364 63643
rect 13324 63069 13364 63078
rect 13516 62936 13556 62945
rect 13228 62896 13516 62936
rect 13228 62348 13268 62896
rect 13516 62887 13556 62896
rect 13228 62299 13268 62308
rect 13515 62180 13557 62189
rect 13515 62140 13516 62180
rect 13556 62140 13557 62180
rect 13515 62131 13557 62140
rect 13323 61928 13365 61937
rect 13323 61888 13324 61928
rect 13364 61888 13365 61928
rect 13323 61879 13365 61888
rect 13228 61592 13268 61601
rect 13228 60593 13268 61552
rect 13227 60584 13269 60593
rect 13227 60544 13228 60584
rect 13268 60544 13269 60584
rect 13227 60535 13269 60544
rect 13227 60080 13269 60089
rect 13227 60040 13228 60080
rect 13268 60040 13269 60080
rect 13227 60031 13269 60040
rect 13228 59408 13268 60031
rect 13228 59359 13268 59368
rect 13131 58064 13173 58073
rect 13131 58024 13132 58064
rect 13172 58024 13173 58064
rect 13131 58015 13173 58024
rect 13324 57989 13364 61879
rect 13419 61256 13461 61265
rect 13419 61216 13420 61256
rect 13460 61216 13461 61256
rect 13419 61207 13461 61216
rect 13323 57980 13365 57989
rect 13323 57940 13324 57980
rect 13364 57940 13365 57980
rect 13323 57931 13365 57940
rect 13131 57896 13173 57905
rect 13131 57856 13132 57896
rect 13172 57856 13173 57896
rect 13131 57847 13173 57856
rect 13132 57762 13172 57847
rect 13324 57644 13364 57653
rect 13132 57604 13324 57644
rect 13132 57140 13172 57604
rect 13324 57595 13364 57604
rect 13420 57224 13460 61207
rect 13516 59081 13556 62131
rect 13612 60761 13652 64240
rect 13708 64037 13748 69784
rect 13803 68984 13845 68993
rect 13803 68944 13804 68984
rect 13844 68944 13845 68984
rect 13803 68935 13845 68944
rect 13804 68480 13844 68935
rect 13804 68431 13844 68440
rect 13803 68312 13845 68321
rect 13803 68272 13804 68312
rect 13844 68272 13845 68312
rect 13803 68263 13845 68272
rect 13707 64028 13749 64037
rect 13707 63988 13708 64028
rect 13748 63988 13749 64028
rect 13707 63979 13749 63988
rect 13707 63692 13749 63701
rect 13707 63652 13708 63692
rect 13748 63652 13749 63692
rect 13707 63643 13749 63652
rect 13708 63558 13748 63643
rect 13707 62096 13749 62105
rect 13707 62056 13708 62096
rect 13748 62056 13749 62096
rect 13707 62047 13749 62056
rect 13611 60752 13653 60761
rect 13611 60712 13612 60752
rect 13652 60712 13653 60752
rect 13611 60703 13653 60712
rect 13515 59072 13557 59081
rect 13515 59032 13516 59072
rect 13556 59032 13557 59072
rect 13515 59023 13557 59032
rect 13708 58913 13748 62047
rect 13804 60509 13844 68263
rect 13900 65288 13940 72304
rect 13996 72176 14036 72187
rect 13996 72101 14036 72136
rect 13995 72092 14037 72101
rect 13995 72052 13996 72092
rect 14036 72052 14037 72092
rect 13995 72043 14037 72052
rect 13995 71588 14037 71597
rect 13995 71548 13996 71588
rect 14036 71548 14037 71588
rect 13995 71539 14037 71548
rect 13996 71454 14036 71539
rect 14092 69329 14132 78931
rect 14380 78930 14420 79015
rect 14187 78812 14229 78821
rect 14187 78772 14188 78812
rect 14228 78772 14229 78812
rect 14187 78763 14229 78772
rect 14188 78678 14228 78763
rect 14283 78644 14325 78653
rect 14283 78604 14284 78644
rect 14324 78604 14325 78644
rect 14283 78595 14325 78604
rect 14187 78140 14229 78149
rect 14187 78100 14188 78140
rect 14228 78100 14229 78140
rect 14187 78091 14229 78100
rect 14188 71933 14228 78091
rect 14284 73688 14324 78595
rect 14380 78224 14420 78233
rect 14380 76553 14420 78184
rect 14476 76721 14516 79024
rect 14475 76712 14517 76721
rect 14475 76672 14476 76712
rect 14516 76672 14517 76712
rect 14475 76663 14517 76672
rect 14572 76712 14612 81703
rect 14668 78989 14708 84643
rect 14764 83264 14804 85399
rect 14860 84113 14900 85936
rect 14956 84272 14996 84281
rect 14859 84104 14901 84113
rect 14859 84064 14860 84104
rect 14900 84064 14901 84104
rect 14859 84055 14901 84064
rect 14956 83609 14996 84232
rect 14955 83600 14997 83609
rect 14955 83560 14956 83600
rect 14996 83560 14997 83600
rect 14955 83551 14997 83560
rect 15052 83525 15092 85936
rect 15244 84785 15284 85936
rect 15243 84776 15285 84785
rect 15243 84736 15244 84776
rect 15284 84736 15285 84776
rect 15243 84727 15285 84736
rect 15340 84281 15380 84366
rect 15339 84272 15381 84281
rect 15339 84232 15340 84272
rect 15380 84232 15381 84272
rect 15339 84223 15381 84232
rect 15148 84104 15188 84113
rect 15188 84064 15380 84104
rect 15148 84055 15188 84064
rect 15147 83852 15189 83861
rect 15147 83812 15148 83852
rect 15188 83812 15189 83852
rect 15147 83803 15189 83812
rect 15051 83516 15093 83525
rect 15051 83476 15052 83516
rect 15092 83476 15093 83516
rect 15051 83467 15093 83476
rect 14764 83224 14996 83264
rect 14763 83096 14805 83105
rect 14763 83056 14764 83096
rect 14804 83056 14805 83096
rect 14763 83047 14805 83056
rect 14764 82013 14804 83047
rect 14956 82769 14996 83224
rect 14955 82760 14997 82769
rect 14955 82720 14956 82760
rect 14996 82720 14997 82760
rect 14955 82711 14997 82720
rect 14956 82626 14996 82711
rect 14763 82004 14805 82013
rect 14763 81964 14764 82004
rect 14804 81964 14805 82004
rect 14763 81955 14805 81964
rect 14956 82004 14996 82015
rect 15052 82013 15092 82098
rect 14956 81929 14996 81964
rect 15051 82004 15093 82013
rect 15051 81964 15052 82004
rect 15092 81964 15093 82004
rect 15051 81955 15093 81964
rect 14955 81920 14997 81929
rect 14955 81880 14956 81920
rect 14996 81880 14997 81920
rect 14955 81871 14997 81880
rect 15051 81668 15093 81677
rect 15051 81628 15052 81668
rect 15092 81628 15093 81668
rect 15051 81619 15093 81628
rect 15052 81257 15092 81619
rect 15051 81248 15093 81257
rect 15051 81208 15052 81248
rect 15092 81208 15093 81248
rect 15051 81199 15093 81208
rect 15052 81114 15092 81199
rect 14859 80744 14901 80753
rect 14859 80704 14860 80744
rect 14900 80704 14901 80744
rect 14859 80695 14901 80704
rect 14860 80576 14900 80695
rect 14763 80240 14805 80249
rect 14763 80200 14764 80240
rect 14804 80200 14805 80240
rect 14763 80191 14805 80200
rect 14667 78980 14709 78989
rect 14667 78940 14668 78980
rect 14708 78940 14709 78980
rect 14667 78931 14709 78940
rect 14667 77720 14709 77729
rect 14667 77680 14668 77720
rect 14708 77680 14709 77720
rect 14667 77671 14709 77680
rect 14668 77552 14708 77671
rect 14764 77552 14804 80191
rect 14860 79400 14900 80536
rect 15148 79988 15188 83803
rect 15243 83600 15285 83609
rect 15243 83560 15244 83600
rect 15284 83560 15285 83600
rect 15243 83551 15285 83560
rect 15244 81677 15284 83551
rect 15340 81920 15380 84064
rect 15436 83945 15476 85936
rect 15435 83936 15477 83945
rect 15435 83896 15436 83936
rect 15476 83896 15477 83936
rect 15628 83936 15668 85936
rect 15820 84617 15860 85936
rect 16012 84869 16052 85936
rect 16204 84944 16244 85936
rect 16108 84904 16244 84944
rect 16011 84860 16053 84869
rect 16011 84820 16012 84860
rect 16052 84820 16053 84860
rect 16011 84811 16053 84820
rect 15819 84608 15861 84617
rect 15819 84568 15820 84608
rect 15860 84568 15861 84608
rect 15819 84559 15861 84568
rect 15628 83896 15764 83936
rect 15435 83887 15477 83896
rect 15436 83348 15476 83357
rect 15436 82774 15476 83308
rect 15627 83348 15669 83357
rect 15627 83308 15628 83348
rect 15668 83308 15669 83348
rect 15627 83299 15669 83308
rect 15628 83214 15668 83299
rect 15436 82725 15476 82734
rect 15531 82760 15573 82769
rect 15531 82720 15532 82760
rect 15572 82720 15573 82760
rect 15531 82711 15573 82720
rect 15532 82088 15572 82711
rect 15628 82592 15668 82603
rect 15628 82517 15668 82552
rect 15627 82508 15669 82517
rect 15627 82468 15628 82508
rect 15668 82468 15669 82508
rect 15627 82459 15669 82468
rect 15572 82048 15668 82088
rect 15532 82039 15572 82048
rect 15340 81880 15572 81920
rect 15243 81668 15285 81677
rect 15243 81628 15244 81668
rect 15284 81628 15285 81668
rect 15243 81619 15285 81628
rect 15436 81089 15476 81174
rect 15244 81080 15284 81089
rect 15435 81080 15477 81089
rect 15284 81040 15380 81080
rect 15244 81031 15284 81040
rect 15340 80571 15380 81040
rect 15435 81040 15436 81080
rect 15476 81040 15477 81080
rect 15435 81031 15477 81040
rect 15532 80912 15572 81880
rect 15340 80522 15380 80531
rect 15436 80872 15572 80912
rect 15148 79948 15284 79988
rect 14955 79820 14997 79829
rect 14955 79780 14956 79820
rect 14996 79780 14997 79820
rect 14955 79771 14997 79780
rect 14956 79736 14996 79771
rect 14956 79685 14996 79696
rect 15147 79652 15189 79661
rect 15147 79612 15148 79652
rect 15188 79612 15189 79652
rect 15147 79603 15189 79612
rect 15148 79518 15188 79603
rect 14860 79360 14996 79400
rect 14859 78812 14901 78821
rect 14859 78772 14860 78812
rect 14900 78772 14901 78812
rect 14859 78763 14901 78772
rect 14860 78238 14900 78763
rect 14956 78401 14996 79360
rect 14955 78392 14997 78401
rect 14955 78352 14956 78392
rect 14996 78352 14997 78392
rect 14955 78343 14997 78352
rect 15244 78317 15284 79948
rect 15340 79736 15380 79745
rect 15436 79736 15476 80872
rect 15628 80753 15668 82048
rect 15724 81500 15764 83896
rect 16108 83861 16148 84904
rect 16203 84776 16245 84785
rect 16203 84736 16204 84776
rect 16244 84736 16245 84776
rect 16203 84727 16245 84736
rect 16107 83852 16149 83861
rect 16107 83812 16108 83852
rect 16148 83812 16149 83852
rect 16107 83803 16149 83812
rect 15819 83516 15861 83525
rect 15819 83476 15820 83516
rect 15860 83476 15861 83516
rect 15819 83467 15861 83476
rect 16204 83516 16244 84727
rect 16204 83467 16244 83476
rect 15820 83382 15860 83467
rect 15915 83432 15957 83441
rect 15915 83392 15916 83432
rect 15956 83392 15957 83432
rect 15915 83383 15957 83392
rect 15819 83012 15861 83021
rect 15819 82972 15820 83012
rect 15860 82972 15861 83012
rect 15819 82963 15861 82972
rect 15820 82760 15860 82963
rect 15820 82711 15860 82720
rect 15916 81920 15956 83383
rect 16012 83357 16052 83442
rect 16011 83348 16053 83357
rect 16011 83308 16012 83348
rect 16052 83308 16053 83348
rect 16011 83299 16053 83308
rect 16299 83348 16341 83357
rect 16299 83308 16300 83348
rect 16340 83308 16341 83348
rect 16299 83299 16341 83308
rect 16011 83180 16053 83189
rect 16011 83140 16012 83180
rect 16052 83140 16053 83180
rect 16011 83131 16053 83140
rect 16012 82083 16052 83131
rect 16107 82508 16149 82517
rect 16107 82468 16108 82508
rect 16148 82468 16149 82508
rect 16107 82459 16149 82468
rect 16012 82034 16052 82043
rect 16108 81920 16148 82459
rect 16203 82340 16245 82349
rect 16203 82300 16204 82340
rect 16244 82300 16245 82340
rect 16203 82291 16245 82300
rect 16204 82172 16244 82291
rect 16204 82097 16244 82132
rect 16203 82088 16245 82097
rect 16203 82048 16204 82088
rect 16244 82048 16245 82088
rect 16203 82039 16245 82048
rect 15916 81880 16052 81920
rect 16108 81880 16244 81920
rect 15724 81451 15764 81460
rect 15916 81332 15956 81341
rect 15724 81292 15916 81332
rect 15627 80744 15669 80753
rect 15627 80704 15628 80744
rect 15668 80704 15669 80744
rect 15627 80695 15669 80704
rect 15532 80660 15572 80669
rect 15532 80333 15572 80620
rect 15627 80576 15669 80585
rect 15627 80536 15628 80576
rect 15668 80536 15669 80576
rect 15627 80527 15669 80536
rect 15531 80324 15573 80333
rect 15531 80284 15532 80324
rect 15572 80284 15573 80324
rect 15531 80275 15573 80284
rect 15532 79988 15572 79997
rect 15628 79988 15668 80527
rect 15572 79948 15668 79988
rect 15532 79939 15572 79948
rect 15380 79696 15476 79736
rect 15531 79736 15573 79745
rect 15531 79696 15532 79736
rect 15572 79696 15573 79736
rect 15340 79157 15380 79696
rect 15531 79687 15573 79696
rect 15532 79602 15572 79687
rect 15435 79316 15477 79325
rect 15435 79276 15436 79316
rect 15476 79276 15477 79316
rect 15435 79267 15477 79276
rect 15339 79148 15381 79157
rect 15339 79108 15340 79148
rect 15380 79108 15381 79148
rect 15339 79099 15381 79108
rect 15243 78308 15285 78317
rect 15243 78268 15244 78308
rect 15284 78268 15285 78308
rect 15243 78259 15285 78268
rect 14860 78189 14900 78198
rect 14955 78224 14997 78233
rect 14955 78184 14956 78224
rect 14996 78184 14997 78224
rect 14955 78175 14997 78184
rect 15339 78224 15381 78233
rect 15339 78184 15340 78224
rect 15380 78184 15381 78224
rect 15339 78175 15381 78184
rect 15436 78224 15476 79267
rect 15627 79232 15669 79241
rect 15627 79192 15628 79232
rect 15668 79192 15669 79232
rect 15627 79183 15669 79192
rect 15531 79064 15573 79073
rect 15531 79024 15532 79064
rect 15572 79024 15573 79064
rect 15531 79015 15573 79024
rect 15628 79064 15668 79183
rect 14860 77720 14900 77729
rect 14956 77720 14996 78175
rect 15052 78140 15092 78149
rect 15092 78100 15284 78140
rect 15052 78091 15092 78100
rect 14900 77680 14996 77720
rect 14860 77671 14900 77680
rect 14764 77512 14900 77552
rect 14668 77057 14708 77512
rect 14667 77048 14709 77057
rect 14667 77008 14668 77048
rect 14708 77008 14709 77048
rect 14667 76999 14709 77008
rect 14763 76796 14805 76805
rect 14763 76756 14764 76796
rect 14804 76756 14805 76796
rect 14763 76747 14805 76756
rect 14379 76544 14421 76553
rect 14379 76504 14380 76544
rect 14420 76504 14421 76544
rect 14379 76495 14421 76504
rect 14380 75713 14420 76495
rect 14379 75704 14421 75713
rect 14379 75664 14380 75704
rect 14420 75664 14421 75704
rect 14379 75655 14421 75664
rect 14475 74528 14517 74537
rect 14475 74488 14476 74528
rect 14516 74488 14517 74528
rect 14475 74479 14517 74488
rect 14476 74394 14516 74479
rect 14284 73529 14324 73648
rect 14283 73520 14325 73529
rect 14283 73480 14284 73520
rect 14324 73480 14325 73520
rect 14283 73471 14325 73480
rect 14283 73016 14325 73025
rect 14283 72976 14284 73016
rect 14324 72976 14325 73016
rect 14283 72967 14325 72976
rect 14187 71924 14229 71933
rect 14187 71884 14188 71924
rect 14228 71884 14229 71924
rect 14187 71875 14229 71884
rect 14187 71756 14229 71765
rect 14187 71716 14188 71756
rect 14228 71716 14229 71756
rect 14187 71707 14229 71716
rect 14188 71504 14228 71707
rect 14188 71455 14228 71464
rect 14187 70496 14229 70505
rect 14187 70456 14188 70496
rect 14228 70456 14229 70496
rect 14187 70447 14229 70456
rect 14091 69320 14133 69329
rect 14091 69280 14092 69320
rect 14132 69280 14133 69320
rect 14188 69320 14228 70447
rect 14284 70001 14324 72967
rect 14572 72101 14612 76672
rect 14667 76712 14709 76721
rect 14667 76672 14668 76712
rect 14708 76672 14709 76712
rect 14667 76663 14709 76672
rect 14668 74789 14708 76663
rect 14764 75200 14804 76747
rect 14667 74780 14709 74789
rect 14667 74740 14668 74780
rect 14708 74740 14709 74780
rect 14667 74731 14709 74740
rect 14764 73781 14804 75160
rect 14763 73772 14805 73781
rect 14763 73732 14764 73772
rect 14804 73732 14805 73772
rect 14763 73723 14805 73732
rect 14860 73100 14900 77512
rect 15244 77468 15284 78100
rect 15340 78090 15380 78175
rect 15436 78149 15476 78184
rect 15435 78140 15477 78149
rect 15435 78100 15436 78140
rect 15476 78100 15477 78140
rect 15435 78091 15477 78100
rect 15532 77720 15572 79015
rect 15628 78653 15668 79024
rect 15627 78644 15669 78653
rect 15627 78604 15628 78644
rect 15668 78604 15669 78644
rect 15627 78595 15669 78604
rect 15244 77419 15284 77428
rect 15340 77680 15572 77720
rect 15051 77300 15093 77309
rect 15051 77260 15052 77300
rect 15092 77260 15093 77300
rect 15051 77251 15093 77260
rect 15052 77166 15092 77251
rect 15243 76880 15285 76889
rect 15243 76840 15244 76880
rect 15284 76840 15285 76880
rect 15243 76831 15285 76840
rect 15244 76040 15284 76831
rect 15244 75991 15284 76000
rect 15051 75956 15093 75965
rect 15051 75916 15052 75956
rect 15092 75916 15093 75956
rect 15051 75907 15093 75916
rect 14956 75032 14996 75041
rect 14956 74523 14996 74992
rect 15052 74948 15092 75907
rect 15340 75545 15380 77680
rect 15532 77552 15572 77561
rect 15436 77512 15532 77552
rect 15436 76301 15476 77512
rect 15532 77503 15572 77512
rect 15724 76964 15764 81292
rect 15916 81283 15956 81292
rect 15819 80576 15861 80585
rect 15819 80536 15820 80576
rect 15860 80536 15861 80576
rect 15819 80527 15861 80536
rect 16012 80576 16052 81880
rect 16108 81089 16148 81174
rect 16107 81080 16149 81089
rect 16107 81040 16108 81080
rect 16148 81040 16149 81080
rect 16107 81031 16149 81040
rect 16204 80912 16244 81880
rect 16012 80527 16052 80536
rect 16108 80872 16244 80912
rect 15820 80442 15860 80527
rect 15819 80324 15861 80333
rect 15819 80284 15820 80324
rect 15860 80284 15861 80324
rect 15819 80275 15861 80284
rect 15820 80190 15860 80275
rect 15915 80156 15957 80165
rect 15915 80116 15916 80156
rect 15956 80116 15957 80156
rect 15915 80107 15957 80116
rect 15820 79736 15860 79747
rect 15820 79661 15860 79696
rect 15916 79736 15956 80107
rect 15819 79652 15861 79661
rect 15819 79612 15820 79652
rect 15860 79612 15861 79652
rect 15819 79603 15861 79612
rect 15819 79484 15861 79493
rect 15819 79444 15820 79484
rect 15860 79444 15861 79484
rect 15819 79435 15861 79444
rect 15820 78728 15860 79435
rect 15916 79409 15956 79696
rect 15915 79400 15957 79409
rect 15915 79360 15916 79400
rect 15956 79360 15957 79400
rect 15915 79351 15957 79360
rect 15915 79064 15957 79073
rect 15915 79024 15916 79064
rect 15956 79024 15957 79064
rect 15915 79015 15957 79024
rect 15916 78930 15956 79015
rect 16011 78728 16053 78737
rect 15820 78688 15956 78728
rect 15819 78560 15861 78569
rect 15819 78520 15820 78560
rect 15860 78520 15861 78560
rect 15819 78511 15861 78520
rect 15820 78308 15860 78511
rect 15820 78259 15860 78268
rect 15916 78233 15956 78688
rect 16011 78688 16012 78728
rect 16052 78688 16053 78728
rect 16011 78679 16053 78688
rect 15915 78224 15957 78233
rect 15915 78184 15916 78224
rect 15956 78184 15957 78224
rect 15915 78175 15957 78184
rect 15916 78090 15956 78175
rect 15915 77720 15957 77729
rect 15915 77680 15916 77720
rect 15956 77680 15957 77720
rect 15915 77671 15957 77680
rect 15532 76924 15764 76964
rect 15435 76292 15477 76301
rect 15435 76252 15436 76292
rect 15476 76252 15477 76292
rect 15435 76243 15477 76252
rect 15435 76124 15477 76133
rect 15435 76084 15436 76124
rect 15476 76084 15477 76124
rect 15435 76075 15477 76084
rect 15339 75536 15381 75545
rect 15339 75496 15340 75536
rect 15380 75496 15381 75536
rect 15339 75487 15381 75496
rect 15436 75368 15476 76075
rect 15244 75328 15476 75368
rect 15244 75200 15284 75328
rect 15532 75284 15572 76924
rect 15916 76889 15956 77671
rect 15915 76880 15957 76889
rect 15915 76840 15916 76880
rect 15956 76840 15957 76880
rect 15915 76831 15957 76840
rect 15820 76712 15860 76721
rect 15916 76712 15956 76831
rect 15860 76672 15956 76712
rect 16012 76712 16052 78679
rect 16108 77552 16148 80872
rect 16300 80669 16340 83299
rect 16396 81500 16436 85936
rect 16588 84440 16628 85936
rect 16588 84400 16724 84440
rect 16588 84272 16628 84281
rect 16588 83609 16628 84232
rect 16492 83600 16532 83609
rect 16492 83273 16532 83560
rect 16587 83600 16629 83609
rect 16587 83560 16588 83600
rect 16628 83560 16629 83600
rect 16587 83551 16629 83560
rect 16491 83264 16533 83273
rect 16491 83224 16492 83264
rect 16532 83224 16533 83264
rect 16491 83215 16533 83224
rect 16492 81920 16532 81929
rect 16492 81845 16532 81880
rect 16491 81836 16533 81845
rect 16491 81796 16492 81836
rect 16532 81796 16533 81836
rect 16491 81787 16533 81796
rect 16492 81785 16532 81787
rect 16587 81500 16629 81509
rect 16396 81460 16532 81500
rect 16396 81332 16436 81341
rect 16396 81089 16436 81292
rect 16395 81080 16437 81089
rect 16395 81040 16396 81080
rect 16436 81040 16437 81080
rect 16395 81031 16437 81040
rect 16492 80744 16532 81460
rect 16587 81460 16588 81500
rect 16628 81460 16629 81500
rect 16587 81451 16629 81460
rect 16588 81366 16628 81451
rect 16684 80744 16724 84400
rect 16780 84281 16820 85936
rect 16972 84449 17012 85936
rect 16971 84440 17013 84449
rect 16971 84400 16972 84440
rect 17012 84400 17013 84440
rect 16971 84391 17013 84400
rect 16779 84272 16821 84281
rect 16779 84232 16780 84272
rect 16820 84232 16821 84272
rect 16779 84223 16821 84232
rect 16780 84104 16820 84113
rect 16780 83189 16820 84064
rect 17067 84104 17109 84113
rect 17067 84064 17068 84104
rect 17108 84064 17109 84104
rect 17067 84055 17109 84064
rect 17068 83970 17108 84055
rect 16971 83684 17013 83693
rect 16971 83644 16972 83684
rect 17012 83644 17013 83684
rect 16971 83635 17013 83644
rect 16779 83180 16821 83189
rect 16779 83140 16780 83180
rect 16820 83140 16821 83180
rect 16779 83131 16821 83140
rect 16779 82424 16821 82433
rect 16779 82384 16780 82424
rect 16820 82384 16821 82424
rect 16779 82375 16821 82384
rect 16780 82088 16820 82375
rect 16780 81248 16820 82048
rect 16780 81199 16820 81208
rect 16972 80921 17012 83635
rect 17068 82760 17108 82769
rect 16971 80912 17013 80921
rect 16971 80872 16972 80912
rect 17012 80872 17013 80912
rect 16971 80863 17013 80872
rect 16492 80704 16628 80744
rect 16684 80704 17012 80744
rect 16299 80660 16341 80669
rect 16299 80620 16300 80660
rect 16340 80620 16341 80660
rect 16299 80611 16341 80620
rect 16204 80576 16244 80585
rect 16204 80492 16244 80536
rect 16492 80576 16532 80585
rect 16204 80452 16340 80492
rect 16204 80324 16244 80333
rect 16204 79073 16244 80284
rect 16300 80249 16340 80452
rect 16395 80324 16437 80333
rect 16395 80284 16396 80324
rect 16436 80284 16437 80324
rect 16395 80275 16437 80284
rect 16299 80240 16341 80249
rect 16299 80200 16300 80240
rect 16340 80200 16341 80240
rect 16299 80191 16341 80200
rect 16299 80072 16341 80081
rect 16299 80032 16300 80072
rect 16340 80032 16341 80072
rect 16299 80023 16341 80032
rect 16300 79820 16340 80023
rect 16396 79997 16436 80275
rect 16395 79988 16437 79997
rect 16395 79948 16396 79988
rect 16436 79948 16437 79988
rect 16395 79939 16437 79948
rect 16300 79771 16340 79780
rect 16396 79820 16436 79939
rect 16492 79913 16532 80536
rect 16491 79904 16533 79913
rect 16491 79864 16492 79904
rect 16532 79864 16533 79904
rect 16491 79855 16533 79864
rect 16299 79652 16341 79661
rect 16299 79612 16300 79652
rect 16340 79612 16341 79652
rect 16299 79603 16341 79612
rect 16203 79064 16245 79073
rect 16203 79024 16204 79064
rect 16244 79024 16245 79064
rect 16203 79015 16245 79024
rect 16300 77729 16340 79603
rect 16396 78569 16436 79780
rect 16491 79232 16533 79241
rect 16491 79192 16492 79232
rect 16532 79192 16533 79232
rect 16491 79183 16533 79192
rect 16395 78560 16437 78569
rect 16395 78520 16396 78560
rect 16436 78520 16437 78560
rect 16395 78511 16437 78520
rect 16395 78392 16437 78401
rect 16395 78352 16396 78392
rect 16436 78352 16437 78392
rect 16395 78343 16437 78352
rect 16396 78224 16436 78343
rect 16396 78175 16436 78184
rect 16299 77720 16341 77729
rect 16299 77680 16300 77720
rect 16340 77680 16341 77720
rect 16299 77671 16341 77680
rect 16395 77552 16437 77561
rect 16108 77512 16340 77552
rect 16204 76712 16244 76721
rect 16012 76672 16204 76712
rect 15820 76663 15860 76672
rect 16012 76544 16052 76553
rect 15724 76504 16012 76544
rect 15627 76040 15669 76049
rect 15627 76000 15628 76040
rect 15668 76000 15669 76040
rect 15627 75991 15669 76000
rect 15724 76040 15764 76504
rect 15915 76124 15957 76133
rect 15915 76084 15916 76124
rect 15956 76084 15957 76124
rect 15915 76075 15957 76084
rect 15724 75991 15764 76000
rect 15916 76040 15956 76075
rect 15628 75906 15668 75991
rect 15916 75989 15956 76000
rect 15724 75872 15764 75881
rect 15532 75244 15668 75284
rect 15244 75151 15284 75160
rect 15339 75200 15381 75209
rect 15339 75160 15340 75200
rect 15380 75160 15381 75200
rect 15339 75151 15381 75160
rect 15052 74908 15284 74948
rect 15051 74780 15093 74789
rect 15051 74740 15052 74780
rect 15092 74740 15093 74780
rect 15051 74731 15093 74740
rect 14956 74474 14996 74483
rect 14764 73060 14900 73100
rect 14667 72176 14709 72185
rect 14667 72136 14668 72176
rect 14708 72136 14709 72176
rect 14667 72127 14709 72136
rect 14571 72092 14613 72101
rect 14571 72052 14572 72092
rect 14612 72052 14613 72092
rect 14571 72043 14613 72052
rect 14379 71588 14421 71597
rect 14379 71548 14380 71588
rect 14420 71548 14421 71588
rect 14379 71539 14421 71548
rect 14380 71504 14420 71539
rect 14572 71513 14612 72043
rect 14380 71453 14420 71464
rect 14571 71504 14613 71513
rect 14571 71464 14572 71504
rect 14612 71464 14613 71504
rect 14571 71455 14613 71464
rect 14572 71370 14612 71455
rect 14380 71252 14420 71261
rect 14420 71212 14612 71252
rect 14380 71203 14420 71212
rect 14572 70925 14612 71212
rect 14379 70916 14421 70925
rect 14379 70876 14380 70916
rect 14420 70876 14421 70916
rect 14379 70867 14421 70876
rect 14571 70916 14613 70925
rect 14571 70876 14572 70916
rect 14612 70876 14613 70916
rect 14571 70867 14613 70876
rect 14283 69992 14325 70001
rect 14283 69952 14284 69992
rect 14324 69952 14325 69992
rect 14283 69943 14325 69952
rect 14188 69280 14324 69320
rect 14091 69271 14133 69280
rect 14187 69152 14229 69161
rect 14187 69112 14188 69152
rect 14228 69112 14229 69152
rect 14187 69103 14229 69112
rect 14188 68489 14228 69103
rect 14187 68480 14229 68489
rect 14187 68440 14188 68480
rect 14228 68440 14229 68480
rect 14187 68431 14229 68440
rect 14188 68346 14228 68431
rect 14284 68405 14324 69280
rect 14380 68984 14420 70867
rect 14668 70664 14708 72127
rect 14572 70624 14668 70664
rect 14476 69992 14516 70001
rect 14476 69161 14516 69952
rect 14475 69152 14517 69161
rect 14475 69112 14476 69152
rect 14516 69112 14517 69152
rect 14475 69103 14517 69112
rect 14380 68944 14516 68984
rect 14283 68396 14325 68405
rect 14283 68356 14284 68396
rect 14324 68356 14325 68396
rect 14283 68347 14325 68356
rect 13996 68228 14036 68237
rect 14036 68188 14420 68228
rect 13996 68179 14036 68188
rect 14380 66968 14420 68188
rect 14380 66919 14420 66928
rect 14476 66968 14516 68944
rect 14572 68732 14612 70624
rect 14668 70615 14708 70624
rect 14667 70076 14709 70085
rect 14667 70036 14668 70076
rect 14708 70036 14709 70076
rect 14667 70027 14709 70036
rect 14668 69942 14708 70027
rect 14764 69413 14804 73060
rect 15052 72185 15092 74731
rect 15147 74612 15189 74621
rect 15147 74572 15148 74612
rect 15188 74572 15189 74612
rect 15147 74563 15189 74572
rect 15148 74478 15188 74563
rect 15244 74360 15284 74908
rect 15148 74320 15284 74360
rect 15051 72176 15093 72185
rect 15051 72136 15052 72176
rect 15092 72136 15093 72176
rect 15051 72127 15093 72136
rect 15148 71588 15188 74320
rect 15340 73865 15380 75151
rect 15531 75032 15573 75041
rect 15531 74992 15532 75032
rect 15572 74992 15573 75032
rect 15531 74983 15573 74992
rect 15532 74898 15572 74983
rect 15628 74612 15668 75244
rect 15724 75200 15764 75832
rect 15724 75151 15764 75160
rect 15820 75200 15860 75209
rect 15820 75041 15860 75160
rect 15915 75200 15957 75209
rect 15915 75160 15916 75200
rect 15956 75160 15957 75200
rect 15915 75151 15957 75160
rect 16012 75200 16052 76504
rect 16107 76124 16149 76133
rect 16107 76084 16108 76124
rect 16148 76084 16149 76124
rect 16107 76075 16149 76084
rect 16108 75536 16148 76075
rect 16204 76040 16244 76672
rect 16204 75991 16244 76000
rect 16108 75496 16249 75536
rect 16012 75151 16052 75160
rect 16108 75200 16148 75209
rect 15819 75032 15861 75041
rect 15819 74992 15820 75032
rect 15860 74992 15861 75032
rect 15819 74983 15861 74992
rect 15916 75032 15956 75151
rect 15916 74983 15956 74992
rect 15628 74563 15668 74572
rect 16011 74276 16053 74285
rect 16011 74236 16012 74276
rect 16052 74236 16053 74276
rect 16011 74227 16053 74236
rect 15339 73856 15381 73865
rect 15339 73816 15340 73856
rect 15380 73816 15381 73856
rect 15339 73807 15381 73816
rect 15532 73688 15572 73697
rect 15243 73184 15285 73193
rect 15243 73144 15244 73184
rect 15284 73144 15285 73184
rect 15243 73135 15285 73144
rect 15244 73016 15284 73135
rect 15244 72353 15284 72976
rect 15435 72848 15477 72857
rect 15435 72808 15436 72848
rect 15476 72808 15477 72848
rect 15435 72799 15477 72808
rect 15436 72714 15476 72799
rect 15532 72512 15572 73648
rect 16012 73688 16052 74227
rect 16108 73940 16148 75160
rect 16209 75200 16249 75496
rect 16209 75151 16249 75160
rect 16203 74360 16245 74369
rect 16203 74320 16204 74360
rect 16244 74320 16245 74360
rect 16203 74311 16245 74320
rect 16108 73891 16148 73900
rect 16107 73772 16149 73781
rect 16107 73732 16108 73772
rect 16148 73732 16149 73772
rect 16107 73723 16149 73732
rect 16012 73639 16052 73648
rect 15724 73520 15764 73529
rect 15724 73100 15764 73480
rect 15628 73060 15764 73100
rect 15628 72680 15668 73060
rect 15820 73016 15860 73025
rect 15724 72997 15764 73006
rect 15724 72857 15764 72957
rect 15723 72848 15765 72857
rect 15723 72808 15724 72848
rect 15764 72808 15765 72848
rect 15723 72799 15765 72808
rect 15628 72640 15764 72680
rect 15532 72472 15668 72512
rect 15339 72428 15381 72437
rect 15339 72388 15340 72428
rect 15380 72388 15381 72428
rect 15339 72379 15381 72388
rect 15243 72344 15285 72353
rect 15243 72304 15244 72344
rect 15284 72304 15285 72344
rect 15243 72295 15285 72304
rect 15243 72176 15285 72185
rect 15243 72136 15244 72176
rect 15284 72136 15285 72176
rect 15243 72127 15285 72136
rect 15244 72042 15284 72127
rect 15148 71548 15284 71588
rect 15147 71420 15189 71429
rect 15147 71380 15148 71420
rect 15188 71380 15189 71420
rect 15147 71371 15189 71380
rect 15051 70916 15093 70925
rect 15051 70876 15052 70916
rect 15092 70876 15093 70916
rect 15051 70867 15093 70876
rect 14955 70748 14997 70757
rect 14955 70708 14956 70748
rect 14996 70708 14997 70748
rect 14955 70699 14997 70708
rect 14860 70496 14900 70505
rect 14956 70496 14996 70699
rect 15052 70664 15092 70867
rect 15148 70757 15188 71371
rect 15244 70925 15284 71548
rect 15243 70916 15285 70925
rect 15243 70876 15244 70916
rect 15284 70876 15285 70916
rect 15243 70867 15285 70876
rect 15147 70748 15189 70757
rect 15147 70708 15148 70748
rect 15188 70708 15189 70748
rect 15147 70699 15189 70708
rect 15052 70615 15092 70624
rect 15243 70664 15285 70673
rect 15243 70624 15244 70664
rect 15284 70624 15285 70664
rect 15243 70615 15285 70624
rect 15147 70580 15189 70589
rect 15147 70540 15148 70580
rect 15188 70540 15189 70580
rect 15147 70531 15189 70540
rect 14956 70456 15092 70496
rect 14763 69404 14805 69413
rect 14763 69364 14764 69404
rect 14804 69364 14805 69404
rect 14860 69404 14900 70456
rect 14955 70076 14997 70085
rect 14955 70036 14956 70076
rect 14996 70036 14997 70076
rect 14955 70027 14997 70036
rect 14956 69992 14996 70027
rect 14956 69941 14996 69952
rect 15052 69992 15092 70456
rect 15148 70446 15188 70531
rect 15244 70530 15284 70615
rect 15340 70160 15380 72379
rect 15435 72008 15477 72017
rect 15435 71968 15436 72008
rect 15476 71968 15477 72008
rect 15435 71959 15477 71968
rect 15436 71874 15476 71959
rect 15628 71513 15668 72472
rect 15724 72176 15764 72640
rect 15724 72127 15764 72136
rect 15820 72176 15860 72976
rect 15915 72932 15957 72941
rect 15915 72892 15916 72932
rect 15956 72892 15957 72932
rect 15915 72883 15957 72892
rect 15820 71672 15860 72136
rect 15724 71632 15860 71672
rect 15627 71504 15669 71513
rect 15627 71464 15628 71504
rect 15668 71464 15669 71504
rect 15627 71455 15669 71464
rect 15724 71429 15764 71632
rect 15819 71504 15861 71513
rect 15819 71464 15820 71504
rect 15860 71464 15861 71504
rect 15819 71455 15861 71464
rect 15723 71420 15765 71429
rect 15723 71380 15724 71420
rect 15764 71380 15765 71420
rect 15723 71371 15765 71380
rect 15820 71370 15860 71455
rect 15435 71336 15477 71345
rect 15435 71296 15436 71336
rect 15476 71296 15477 71336
rect 15435 71287 15477 71296
rect 15436 70169 15476 71287
rect 15819 70916 15861 70925
rect 15819 70876 15820 70916
rect 15860 70876 15861 70916
rect 15819 70867 15861 70876
rect 15531 70580 15573 70589
rect 15531 70540 15532 70580
rect 15572 70540 15573 70580
rect 15531 70531 15573 70540
rect 14860 69364 14996 69404
rect 14763 69355 14805 69364
rect 14667 68984 14709 68993
rect 14667 68944 14668 68984
rect 14708 68944 14709 68984
rect 14667 68935 14709 68944
rect 14668 68850 14708 68935
rect 14764 68900 14804 69355
rect 14956 69152 14996 69364
rect 14956 69103 14996 69112
rect 15052 69152 15092 69952
rect 15052 69103 15092 69112
rect 15148 70120 15380 70160
rect 15435 70160 15477 70169
rect 15435 70120 15436 70160
rect 15476 70120 15477 70160
rect 14764 68860 15092 68900
rect 14572 68692 14708 68732
rect 14571 68564 14613 68573
rect 14571 68524 14572 68564
rect 14612 68524 14613 68564
rect 14571 68515 14613 68524
rect 14476 66800 14516 66928
rect 14380 66760 14516 66800
rect 14091 66128 14133 66137
rect 14091 66088 14092 66128
rect 14132 66088 14133 66128
rect 14091 66079 14133 66088
rect 14092 65994 14132 66079
rect 14284 65960 14324 65969
rect 14284 65456 14324 65920
rect 14284 65407 14324 65416
rect 14380 65456 14420 66760
rect 14476 66128 14516 66137
rect 14572 66128 14612 68515
rect 14516 66088 14612 66128
rect 14476 66079 14516 66088
rect 14571 65876 14613 65885
rect 14571 65836 14572 65876
rect 14612 65836 14613 65876
rect 14571 65827 14613 65836
rect 14380 65297 14420 65416
rect 14379 65288 14421 65297
rect 13900 65248 14324 65288
rect 14187 65120 14229 65129
rect 14187 65080 14188 65120
rect 14228 65080 14229 65120
rect 14187 65071 14229 65080
rect 13899 64616 13941 64625
rect 13899 64576 13900 64616
rect 13940 64576 13941 64616
rect 13899 64567 13941 64576
rect 13900 64482 13940 64567
rect 14092 64448 14132 64457
rect 14092 64280 14132 64408
rect 13996 64240 14132 64280
rect 13996 63944 14036 64240
rect 13996 63895 14036 63904
rect 14092 63944 14132 63953
rect 14092 63113 14132 63904
rect 14091 63104 14133 63113
rect 14091 63064 14092 63104
rect 14132 63064 14133 63104
rect 14091 63055 14133 63064
rect 13995 63020 14037 63029
rect 13995 62980 13996 63020
rect 14036 62980 14037 63020
rect 13995 62971 14037 62980
rect 13899 61844 13941 61853
rect 13899 61804 13900 61844
rect 13940 61804 13941 61844
rect 13899 61795 13941 61804
rect 13803 60500 13845 60509
rect 13803 60460 13804 60500
rect 13844 60460 13845 60500
rect 13803 60451 13845 60460
rect 13900 60425 13940 61795
rect 13996 61517 14036 62971
rect 13995 61508 14037 61517
rect 13995 61468 13996 61508
rect 14036 61468 14037 61508
rect 13995 61459 14037 61468
rect 13899 60416 13941 60425
rect 13899 60376 13900 60416
rect 13940 60376 13941 60416
rect 13899 60367 13941 60376
rect 13899 60080 13941 60089
rect 13899 60040 13900 60080
rect 13940 60040 13941 60080
rect 13899 60031 13941 60040
rect 13707 58904 13749 58913
rect 13707 58864 13708 58904
rect 13748 58864 13749 58904
rect 13707 58855 13749 58864
rect 13707 58736 13749 58745
rect 13707 58696 13708 58736
rect 13748 58696 13749 58736
rect 13707 58687 13749 58696
rect 13708 58568 13748 58687
rect 13708 57989 13748 58528
rect 13707 57980 13749 57989
rect 13707 57940 13708 57980
rect 13748 57940 13749 57980
rect 13707 57931 13749 57940
rect 13084 57100 13172 57140
rect 13324 57184 13460 57224
rect 13084 57098 13124 57100
rect 13084 57049 13124 57058
rect 13228 56972 13268 56981
rect 12940 56932 13228 56972
rect 13228 56923 13268 56932
rect 13324 56300 13364 57184
rect 13419 57056 13461 57065
rect 13419 57016 13420 57056
rect 13460 57016 13461 57056
rect 13419 57007 13461 57016
rect 13516 57056 13556 57065
rect 13420 56729 13460 57007
rect 13419 56720 13461 56729
rect 13419 56680 13420 56720
rect 13460 56680 13461 56720
rect 13419 56671 13461 56680
rect 13420 56468 13460 56671
rect 13516 56552 13556 57016
rect 13612 57056 13652 57065
rect 13612 56813 13652 57016
rect 13611 56804 13653 56813
rect 13611 56764 13612 56804
rect 13652 56764 13653 56804
rect 13611 56755 13653 56764
rect 13516 56512 13748 56552
rect 13708 56468 13748 56512
rect 13804 56468 13844 56477
rect 13420 56428 13652 56468
rect 13708 56428 13804 56468
rect 13612 56384 13652 56428
rect 13804 56419 13844 56428
rect 13612 56335 13652 56344
rect 13324 56260 13556 56300
rect 13516 56216 13556 56260
rect 13516 56176 13748 56216
rect 12939 55880 12981 55889
rect 12939 55840 12940 55880
rect 12980 55840 12981 55880
rect 12939 55831 12981 55840
rect 12940 55469 12980 55831
rect 13612 55628 13652 55637
rect 13228 55588 13612 55628
rect 13084 55553 13124 55562
rect 13124 55513 13172 55544
rect 13084 55504 13172 55513
rect 12939 55460 12981 55469
rect 12939 55420 12940 55460
rect 12980 55420 12981 55460
rect 12939 55411 12981 55420
rect 13132 55040 13172 55504
rect 13228 55460 13268 55588
rect 13612 55579 13652 55588
rect 13228 55411 13268 55420
rect 13420 55376 13460 55387
rect 13420 55301 13460 55336
rect 13515 55376 13557 55385
rect 13515 55336 13516 55376
rect 13556 55336 13557 55376
rect 13515 55327 13557 55336
rect 13419 55292 13461 55301
rect 13419 55252 13420 55292
rect 13460 55252 13461 55292
rect 13419 55243 13461 55252
rect 13228 55040 13268 55049
rect 13132 55000 13228 55040
rect 13228 54991 13268 55000
rect 13420 55040 13460 55049
rect 13516 55040 13556 55327
rect 13460 55000 13556 55040
rect 13420 54991 13460 55000
rect 13036 54872 13076 54881
rect 12843 54200 12885 54209
rect 13036 54200 13076 54832
rect 13612 54788 13652 54797
rect 12843 54160 12844 54200
rect 12884 54160 13076 54200
rect 13324 54748 13612 54788
rect 12843 54151 12885 54160
rect 12844 54032 12884 54151
rect 12844 53983 12884 53992
rect 13228 54032 13268 54043
rect 13228 53957 13268 53992
rect 13227 53948 13269 53957
rect 13227 53908 13228 53948
rect 13268 53908 13269 53948
rect 13227 53899 13269 53908
rect 13036 53864 13076 53873
rect 13076 53824 13172 53864
rect 13036 53815 13076 53824
rect 12843 53696 12885 53705
rect 12843 53656 12844 53696
rect 12884 53656 12885 53696
rect 12843 53647 12885 53656
rect 12844 52025 12884 53647
rect 13132 53355 13172 53824
rect 13228 53369 13268 53899
rect 13324 53528 13364 54748
rect 13612 54739 13652 54748
rect 13708 53528 13748 56176
rect 13324 53479 13364 53488
rect 13420 53488 13748 53528
rect 13132 53306 13172 53315
rect 13227 53360 13269 53369
rect 13227 53320 13228 53360
rect 13268 53320 13269 53360
rect 13227 53311 13269 53320
rect 13323 53276 13365 53285
rect 13323 53236 13324 53276
rect 13364 53236 13365 53276
rect 13323 53227 13365 53236
rect 13324 52529 13364 53227
rect 12939 52520 12981 52529
rect 12939 52480 12940 52520
rect 12980 52480 12981 52520
rect 12939 52471 12981 52480
rect 13323 52520 13365 52529
rect 13323 52480 13324 52520
rect 13364 52480 13365 52520
rect 13323 52471 13365 52480
rect 12843 52016 12885 52025
rect 12843 51976 12844 52016
rect 12884 51976 12885 52016
rect 12843 51967 12885 51976
rect 12747 51176 12789 51185
rect 12747 51136 12748 51176
rect 12788 51136 12789 51176
rect 12747 51127 12789 51136
rect 12748 51008 12788 51017
rect 12652 50968 12748 51008
rect 12748 50959 12788 50968
rect 12460 50464 12692 50504
rect 12556 50336 12596 50345
rect 12116 50296 12212 50336
rect 12076 50287 12116 50296
rect 11979 49664 12021 49673
rect 11979 49624 11980 49664
rect 12020 49624 12021 49664
rect 11979 49615 12021 49624
rect 11883 48824 11925 48833
rect 11883 48784 11884 48824
rect 11924 48784 11925 48824
rect 11883 48775 11925 48784
rect 11884 48690 11924 48775
rect 11980 48749 12020 49615
rect 12172 49496 12212 50296
rect 12556 50252 12596 50296
rect 12268 50212 12596 50252
rect 12652 50336 12692 50464
rect 12940 50345 12980 52471
rect 13035 52100 13077 52109
rect 13035 52060 13036 52100
rect 13076 52060 13077 52100
rect 13035 52051 13077 52060
rect 12268 50168 12308 50212
rect 12268 50119 12308 50128
rect 12652 49925 12692 50296
rect 12939 50336 12981 50345
rect 12939 50296 12940 50336
rect 12980 50296 12981 50336
rect 12939 50287 12981 50296
rect 13036 50261 13076 52051
rect 13420 50840 13460 53488
rect 13707 53360 13749 53369
rect 13707 53320 13708 53360
rect 13748 53320 13749 53360
rect 13707 53311 13749 53320
rect 13804 53360 13844 53369
rect 13611 53024 13653 53033
rect 13611 52984 13612 53024
rect 13652 52984 13653 53024
rect 13611 52975 13653 52984
rect 13515 52436 13557 52445
rect 13515 52396 13516 52436
rect 13556 52396 13557 52436
rect 13515 52387 13557 52396
rect 13516 51848 13556 52387
rect 13516 51773 13556 51808
rect 13515 51764 13557 51773
rect 13515 51724 13516 51764
rect 13556 51724 13557 51764
rect 13515 51715 13557 51724
rect 13420 50800 13556 50840
rect 13132 50294 13172 50303
rect 13035 50252 13077 50261
rect 13035 50212 13036 50252
rect 13076 50212 13077 50252
rect 13516 50261 13556 50800
rect 13612 50336 13652 52975
rect 13708 52016 13748 53311
rect 13804 52949 13844 53320
rect 13803 52940 13845 52949
rect 13803 52900 13804 52940
rect 13844 52900 13845 52940
rect 13803 52891 13845 52900
rect 13708 51967 13748 51976
rect 13803 52016 13845 52025
rect 13803 51976 13804 52016
rect 13844 51976 13845 52016
rect 13803 51967 13845 51976
rect 13804 51689 13844 51967
rect 13803 51680 13845 51689
rect 13803 51640 13804 51680
rect 13844 51640 13845 51680
rect 13803 51631 13845 51640
rect 13900 51260 13940 60031
rect 13996 57401 14036 61459
rect 14092 61013 14132 61044
rect 14091 61004 14133 61013
rect 14091 60964 14092 61004
rect 14132 60964 14133 61004
rect 14091 60955 14133 60964
rect 14092 60920 14132 60955
rect 14092 60761 14132 60880
rect 14091 60752 14133 60761
rect 14091 60712 14092 60752
rect 14132 60712 14133 60752
rect 14091 60703 14133 60712
rect 14091 60500 14133 60509
rect 14091 60460 14092 60500
rect 14132 60460 14133 60500
rect 14091 60451 14133 60460
rect 14092 60332 14132 60451
rect 14092 60283 14132 60292
rect 14092 59912 14132 59921
rect 14092 59417 14132 59872
rect 14091 59408 14133 59417
rect 14091 59368 14092 59408
rect 14132 59368 14133 59408
rect 14091 59359 14133 59368
rect 14092 57896 14132 57907
rect 14092 57821 14132 57856
rect 14091 57812 14133 57821
rect 14091 57772 14092 57812
rect 14132 57772 14133 57812
rect 14091 57763 14133 57772
rect 13995 57392 14037 57401
rect 13995 57352 13996 57392
rect 14036 57352 14037 57392
rect 13995 57343 14037 57352
rect 14091 57224 14133 57233
rect 14091 57184 14092 57224
rect 14132 57184 14133 57224
rect 14091 57175 14133 57184
rect 14092 57140 14132 57175
rect 14092 57089 14132 57100
rect 13996 57056 14036 57065
rect 13996 56804 14036 57016
rect 13996 56764 14132 56804
rect 13995 56636 14037 56645
rect 13995 56596 13996 56636
rect 14036 56596 14037 56636
rect 13995 56587 14037 56596
rect 13804 51220 13940 51260
rect 13707 51176 13749 51185
rect 13707 51136 13708 51176
rect 13748 51136 13749 51176
rect 13707 51127 13749 51136
rect 13132 50252 13172 50254
rect 13227 50252 13269 50261
rect 13132 50212 13228 50252
rect 13268 50212 13269 50252
rect 13035 50203 13077 50212
rect 13227 50203 13269 50212
rect 13515 50252 13557 50261
rect 13515 50212 13516 50252
rect 13556 50212 13557 50252
rect 13515 50203 13557 50212
rect 13419 50168 13461 50177
rect 13419 50128 13420 50168
rect 13460 50128 13461 50168
rect 13419 50119 13461 50128
rect 12651 49916 12693 49925
rect 12651 49876 12652 49916
rect 12692 49876 12693 49916
rect 12651 49867 12693 49876
rect 13035 49916 13077 49925
rect 13035 49876 13036 49916
rect 13076 49876 13077 49916
rect 13035 49867 13077 49876
rect 12460 49496 12500 49505
rect 12940 49496 12980 49505
rect 12172 49456 12460 49496
rect 11979 48740 12021 48749
rect 11979 48700 11980 48740
rect 12020 48700 12021 48740
rect 11979 48691 12021 48700
rect 12076 48572 12116 48581
rect 11788 48532 11924 48572
rect 11787 48404 11829 48413
rect 11787 48364 11788 48404
rect 11828 48364 11829 48404
rect 11787 48355 11829 48364
rect 11691 47144 11733 47153
rect 11691 47104 11692 47144
rect 11732 47104 11733 47144
rect 11691 47095 11733 47104
rect 11403 46136 11445 46145
rect 11403 46096 11404 46136
rect 11444 46096 11445 46136
rect 11403 46087 11445 46096
rect 11307 42692 11349 42701
rect 11307 42652 11308 42692
rect 11348 42652 11349 42692
rect 11307 42643 11349 42652
rect 11307 42440 11349 42449
rect 11307 42400 11308 42440
rect 11348 42400 11349 42440
rect 11307 42391 11349 42400
rect 11308 41936 11348 42391
rect 11308 41887 11348 41896
rect 11211 41852 11253 41861
rect 11211 41812 11212 41852
rect 11252 41812 11253 41852
rect 11211 41803 11253 41812
rect 10539 41768 10581 41777
rect 10539 41728 10540 41768
rect 10580 41728 10581 41768
rect 10539 41719 10581 41728
rect 10443 41264 10485 41273
rect 10443 41224 10444 41264
rect 10484 41224 10485 41264
rect 10443 41215 10485 41224
rect 10540 41264 10580 41719
rect 11307 41684 11349 41693
rect 11307 41644 11308 41684
rect 11348 41644 11349 41684
rect 11307 41635 11349 41644
rect 10635 41600 10677 41609
rect 10635 41560 10636 41600
rect 10676 41560 10677 41600
rect 10635 41551 10677 41560
rect 10540 41215 10580 41224
rect 10636 41264 10676 41551
rect 11019 41432 11061 41441
rect 11019 41392 11020 41432
rect 11060 41392 11156 41432
rect 11019 41383 11061 41392
rect 10731 41348 10773 41357
rect 10731 41308 10732 41348
rect 10772 41308 10773 41348
rect 10731 41299 10773 41308
rect 10636 41215 10676 41224
rect 10444 41130 10484 41215
rect 10732 41214 10772 41299
rect 10924 41273 10964 41358
rect 11116 41285 11156 41392
rect 10923 41264 10965 41273
rect 10923 41224 10924 41264
rect 10964 41224 10965 41264
rect 10923 41215 10965 41224
rect 11020 41264 11060 41275
rect 11212 41273 11252 41358
rect 11116 41236 11156 41245
rect 11211 41264 11253 41273
rect 11020 41189 11060 41224
rect 11211 41224 11212 41264
rect 11252 41224 11253 41264
rect 11211 41215 11253 41224
rect 11019 41180 11061 41189
rect 11019 41140 11020 41180
rect 11060 41140 11061 41180
rect 11019 41131 11061 41140
rect 10827 40844 10869 40853
rect 10827 40804 10828 40844
rect 10868 40804 10869 40844
rect 10827 40795 10869 40804
rect 10443 40676 10485 40685
rect 10443 40636 10444 40676
rect 10484 40636 10485 40676
rect 10443 40627 10485 40636
rect 10347 40592 10389 40601
rect 10347 40552 10348 40592
rect 10388 40552 10389 40592
rect 10347 40543 10389 40552
rect 10251 40508 10293 40517
rect 10251 40468 10252 40508
rect 10292 40468 10293 40508
rect 10251 40459 10293 40468
rect 10155 40424 10197 40433
rect 10155 40384 10156 40424
rect 10196 40384 10197 40424
rect 10155 40375 10197 40384
rect 10252 40424 10292 40459
rect 10156 40290 10196 40375
rect 10252 40373 10292 40384
rect 10347 40424 10389 40433
rect 10347 40384 10348 40424
rect 10388 40384 10389 40424
rect 10347 40375 10389 40384
rect 10444 40424 10484 40627
rect 10444 40375 10484 40384
rect 10636 40424 10676 40433
rect 10348 40290 10388 40375
rect 10251 40256 10293 40265
rect 10251 40216 10252 40256
rect 10292 40216 10293 40256
rect 10251 40207 10293 40216
rect 9964 39698 10100 39738
rect 9867 39584 9909 39593
rect 9867 39544 9868 39584
rect 9908 39544 9909 39584
rect 9867 39535 9909 39544
rect 9964 39416 10004 39698
rect 10060 39584 10100 39593
rect 10252 39584 10292 40207
rect 10636 40181 10676 40384
rect 10828 40424 10868 40795
rect 10923 40676 10965 40685
rect 10923 40636 10924 40676
rect 10964 40636 10965 40676
rect 10923 40627 10965 40636
rect 10828 40375 10868 40384
rect 10732 40340 10772 40349
rect 10635 40172 10677 40181
rect 10635 40132 10636 40172
rect 10676 40132 10677 40172
rect 10635 40123 10677 40132
rect 10732 40013 10772 40300
rect 10731 40004 10773 40013
rect 10731 39964 10732 40004
rect 10772 39964 10773 40004
rect 10731 39955 10773 39964
rect 10539 39836 10581 39845
rect 10539 39796 10540 39836
rect 10580 39796 10581 39836
rect 10539 39787 10581 39796
rect 10347 39752 10389 39761
rect 10347 39712 10348 39752
rect 10388 39712 10389 39752
rect 10347 39703 10389 39712
rect 10540 39752 10580 39787
rect 10348 39618 10388 39703
rect 10540 39701 10580 39712
rect 10636 39752 10676 39761
rect 10676 39712 10772 39752
rect 10636 39703 10676 39712
rect 10100 39544 10292 39584
rect 10060 39535 10100 39544
rect 10348 39500 10388 39509
rect 9964 39376 10100 39416
rect 9772 39031 9812 39040
rect 9771 38912 9813 38921
rect 9771 38872 9772 38912
rect 9812 38872 9813 38912
rect 9771 38863 9813 38872
rect 9964 38912 10004 38923
rect 9772 38778 9812 38863
rect 9964 38837 10004 38872
rect 9963 38828 10005 38837
rect 9963 38788 9964 38828
rect 10004 38788 10005 38828
rect 9963 38779 10005 38788
rect 9964 38417 10004 38779
rect 9963 38408 10005 38417
rect 9963 38368 9964 38408
rect 10004 38368 10005 38408
rect 9963 38359 10005 38368
rect 9772 37232 9812 37241
rect 9812 37192 9908 37232
rect 9772 37183 9812 37192
rect 9676 36688 9812 36728
rect 9291 36308 9333 36317
rect 9291 36268 9292 36308
rect 9332 36268 9333 36308
rect 9291 36259 9333 36268
rect 8908 36100 9044 36140
rect 9196 36140 9236 36149
rect 9292 36140 9332 36259
rect 9236 36100 9332 36140
rect 8908 34721 8948 36100
rect 9196 36091 9236 36100
rect 9291 35972 9333 35981
rect 9291 35932 9292 35972
rect 9332 35932 9333 35972
rect 9291 35923 9333 35932
rect 9004 35888 9044 35897
rect 9004 35225 9044 35848
rect 9195 35720 9237 35729
rect 9195 35680 9196 35720
rect 9236 35680 9237 35720
rect 9195 35671 9237 35680
rect 9003 35216 9045 35225
rect 9003 35176 9004 35216
rect 9044 35176 9045 35216
rect 9003 35167 9045 35176
rect 8907 34712 8949 34721
rect 8907 34672 8908 34712
rect 8948 34672 8949 34712
rect 8907 34663 8949 34672
rect 9004 34385 9044 35167
rect 8811 34376 8853 34385
rect 8811 34336 8812 34376
rect 8852 34336 8853 34376
rect 8811 34327 8853 34336
rect 9003 34376 9045 34385
rect 9003 34336 9004 34376
rect 9044 34336 9045 34376
rect 9003 34327 9045 34336
rect 8812 34242 8852 34327
rect 9004 34208 9044 34217
rect 9004 34049 9044 34168
rect 8715 34040 8757 34049
rect 8715 34000 8716 34040
rect 8756 34000 8757 34040
rect 8715 33991 8757 34000
rect 9003 34040 9045 34049
rect 9003 34000 9004 34040
rect 9044 34000 9045 34040
rect 9003 33991 9045 34000
rect 8235 33872 8277 33881
rect 8235 33832 8236 33872
rect 8276 33832 8277 33872
rect 8235 33823 8277 33832
rect 9004 33872 9044 33881
rect 9044 33832 9140 33872
rect 8716 33797 8756 33828
rect 9004 33823 9044 33832
rect 8427 33788 8469 33797
rect 8427 33748 8428 33788
rect 8468 33748 8469 33788
rect 8427 33739 8469 33748
rect 8715 33788 8757 33797
rect 8715 33748 8716 33788
rect 8756 33748 8757 33788
rect 8715 33739 8757 33748
rect 8236 33704 8276 33713
rect 8428 33704 8468 33739
rect 8276 33664 8372 33704
rect 8236 33655 8276 33664
rect 8235 33200 8277 33209
rect 8235 33160 8236 33200
rect 8276 33160 8277 33200
rect 8235 33151 8277 33160
rect 7796 32824 7892 32864
rect 7756 32815 7796 32824
rect 7700 32152 7796 32192
rect 7660 32143 7700 32152
rect 7468 31480 7700 31520
rect 7084 31366 7124 31480
rect 7084 31317 7124 31326
rect 7275 31352 7317 31361
rect 7275 31312 7276 31352
rect 7316 31312 7317 31352
rect 7275 31303 7317 31312
rect 7276 31268 7316 31303
rect 7276 31217 7316 31228
rect 7468 31016 7508 31480
rect 7372 30976 7508 31016
rect 7564 31352 7604 31361
rect 7276 30680 7316 30689
rect 7276 30269 7316 30640
rect 7275 30260 7317 30269
rect 7275 30220 7276 30260
rect 7316 30220 7317 30260
rect 7275 30211 7317 30220
rect 7372 30092 7412 30976
rect 7468 30848 7508 30857
rect 7564 30848 7604 31312
rect 7660 31352 7700 31480
rect 7660 31303 7700 31312
rect 7659 31184 7701 31193
rect 7659 31144 7660 31184
rect 7700 31144 7701 31184
rect 7659 31135 7701 31144
rect 7508 30808 7604 30848
rect 7468 30799 7508 30808
rect 7276 30052 7412 30092
rect 6987 29420 7029 29429
rect 6987 29380 6988 29420
rect 7028 29380 7029 29420
rect 6987 29371 7029 29380
rect 7276 29345 7316 30052
rect 7563 29924 7605 29933
rect 7563 29884 7564 29924
rect 7604 29884 7605 29924
rect 7563 29875 7605 29884
rect 7564 29840 7604 29875
rect 7564 29789 7604 29800
rect 7275 29336 7317 29345
rect 7275 29296 7276 29336
rect 7316 29296 7317 29336
rect 7275 29287 7317 29296
rect 6988 29151 7028 29179
rect 6988 29093 7028 29111
rect 7276 29168 7316 29177
rect 6987 29084 7029 29093
rect 6987 29044 6988 29084
rect 7028 29044 7029 29084
rect 6987 29035 7029 29044
rect 6507 28960 6508 29000
rect 6548 28960 6549 29000
rect 6507 28951 6549 28960
rect 6604 28960 6836 29000
rect 6028 28505 6068 28876
rect 6316 28867 6356 28876
rect 6219 28748 6261 28757
rect 6219 28708 6220 28748
rect 6260 28708 6261 28748
rect 6219 28699 6261 28708
rect 6123 28580 6165 28589
rect 6123 28540 6124 28580
rect 6164 28540 6165 28580
rect 6123 28531 6165 28540
rect 6027 28496 6069 28505
rect 6027 28456 6028 28496
rect 6068 28456 6069 28496
rect 6027 28447 6069 28456
rect 6028 28169 6068 28447
rect 6027 28160 6069 28169
rect 6027 28120 6028 28160
rect 6068 28120 6069 28160
rect 6027 28111 6069 28120
rect 5931 28076 5973 28085
rect 5931 28036 5932 28076
rect 5972 28036 5973 28076
rect 5931 28027 5973 28036
rect 6124 27908 6164 28531
rect 5932 27868 6164 27908
rect 5932 26816 5972 27868
rect 6027 27740 6069 27749
rect 6027 27700 6028 27740
rect 6068 27700 6069 27740
rect 6027 27691 6069 27700
rect 5932 26767 5972 26776
rect 6028 26816 6068 27691
rect 6124 27665 6164 27750
rect 6123 27656 6165 27665
rect 6123 27616 6124 27656
rect 6164 27616 6165 27656
rect 6123 27607 6165 27616
rect 6220 27488 6260 28699
rect 6412 28337 6452 28422
rect 6411 28328 6453 28337
rect 6508 28328 6548 28951
rect 6604 28421 6644 28960
rect 7083 28748 7125 28757
rect 7083 28708 7084 28748
rect 7124 28708 7125 28748
rect 7276 28748 7316 29128
rect 7564 29168 7604 29177
rect 7660 29168 7700 31135
rect 7604 29128 7700 29168
rect 7564 29119 7604 29128
rect 7372 28916 7412 28925
rect 7412 28876 7508 28916
rect 7372 28867 7412 28876
rect 7276 28708 7412 28748
rect 7083 28699 7125 28708
rect 7084 28580 7124 28699
rect 7084 28531 7124 28540
rect 7372 28505 7412 28708
rect 7371 28496 7413 28505
rect 7371 28456 7372 28496
rect 7412 28456 7413 28496
rect 7371 28447 7413 28456
rect 6603 28412 6645 28421
rect 6603 28372 6604 28412
rect 6644 28372 6645 28412
rect 6603 28363 6645 28372
rect 6411 28288 6412 28328
rect 6452 28288 6548 28328
rect 6411 28279 6453 28288
rect 6411 28160 6453 28169
rect 6411 28120 6412 28160
rect 6452 28120 6453 28160
rect 6411 28111 6453 28120
rect 6028 26767 6068 26776
rect 6124 27448 6260 27488
rect 6124 26648 6164 27448
rect 6316 27404 6356 27413
rect 6220 27077 6260 27162
rect 6219 27068 6261 27077
rect 6219 27028 6220 27068
rect 6260 27028 6261 27068
rect 6219 27019 6261 27028
rect 6316 26825 6356 27364
rect 6220 26816 6260 26825
rect 6315 26816 6357 26825
rect 6260 26776 6316 26816
rect 6356 26776 6357 26816
rect 6220 26767 6260 26776
rect 6315 26767 6357 26776
rect 6316 26682 6356 26767
rect 6412 26648 6452 28111
rect 6507 28076 6549 28085
rect 6507 28036 6508 28076
rect 6548 28036 6549 28076
rect 6507 28027 6549 28036
rect 6508 27656 6548 28027
rect 6604 27656 6644 28363
rect 6699 28328 6741 28337
rect 7276 28328 7316 28337
rect 6699 28288 6700 28328
rect 6740 28288 6741 28328
rect 6699 28279 6741 28288
rect 6892 28288 7276 28328
rect 6700 28194 6740 28279
rect 6796 28244 6836 28255
rect 6796 28169 6836 28204
rect 6795 28160 6837 28169
rect 6795 28120 6796 28160
rect 6836 28120 6837 28160
rect 6795 28111 6837 28120
rect 6892 27824 6932 28288
rect 7276 28279 7316 28288
rect 7468 28328 7508 28876
rect 7563 28748 7605 28757
rect 7563 28708 7564 28748
rect 7604 28708 7605 28748
rect 7563 28699 7605 28708
rect 7372 28160 7412 28169
rect 6796 27784 6932 27824
rect 7180 28120 7372 28160
rect 6700 27656 6740 27665
rect 6604 27616 6700 27656
rect 6508 27572 6548 27616
rect 6700 27607 6740 27616
rect 6508 27532 6644 27572
rect 6508 27404 6548 27413
rect 6508 26816 6548 27364
rect 6604 26993 6644 27532
rect 6603 26984 6645 26993
rect 6603 26944 6604 26984
rect 6644 26944 6645 26984
rect 6603 26935 6645 26944
rect 6508 26767 6548 26776
rect 6604 26816 6644 26825
rect 6124 26608 6260 26648
rect 6412 26608 6548 26648
rect 6124 26228 6164 26237
rect 5932 26144 5972 26153
rect 5932 25901 5972 26104
rect 6027 26144 6069 26153
rect 6027 26104 6028 26144
rect 6068 26104 6069 26144
rect 6027 26095 6069 26104
rect 5931 25892 5973 25901
rect 5931 25852 5932 25892
rect 5972 25852 5973 25892
rect 5931 25843 5973 25852
rect 5835 25808 5877 25817
rect 5835 25768 5836 25808
rect 5876 25768 5877 25808
rect 5835 25759 5877 25768
rect 5932 25556 5972 25565
rect 6028 25556 6068 26095
rect 6124 26069 6164 26188
rect 6123 26060 6165 26069
rect 6123 26020 6124 26060
rect 6164 26020 6165 26060
rect 6123 26011 6165 26020
rect 6123 25892 6165 25901
rect 6123 25852 6124 25892
rect 6164 25852 6165 25892
rect 6123 25843 6165 25852
rect 5972 25516 6068 25556
rect 5932 25507 5972 25516
rect 6124 25481 6164 25843
rect 6123 25472 6165 25481
rect 5644 25432 5876 25472
rect 5739 25304 5781 25313
rect 5739 25264 5740 25304
rect 5780 25264 5781 25304
rect 5836 25304 5876 25432
rect 6123 25432 6124 25472
rect 6164 25432 6165 25472
rect 6123 25423 6165 25432
rect 6124 25304 6164 25313
rect 5836 25264 6124 25304
rect 5739 25255 5781 25264
rect 6124 25255 6164 25264
rect 6220 25304 6260 26608
rect 6315 26564 6357 26573
rect 6315 26524 6316 26564
rect 6356 26524 6357 26564
rect 6315 26515 6357 26524
rect 6316 25976 6356 26515
rect 6508 26405 6548 26608
rect 6604 26573 6644 26776
rect 6699 26816 6741 26825
rect 6699 26776 6700 26816
rect 6740 26776 6741 26816
rect 6699 26767 6741 26776
rect 6796 26816 6836 27784
rect 6892 27656 6932 27665
rect 6892 27077 6932 27616
rect 6987 27656 7029 27665
rect 6987 27616 6988 27656
rect 7028 27616 7029 27656
rect 6987 27607 7029 27616
rect 7180 27656 7220 28120
rect 7372 28111 7412 28120
rect 7275 27992 7317 28001
rect 7468 27992 7508 28288
rect 7564 28328 7604 28699
rect 7564 28279 7604 28288
rect 7275 27952 7276 27992
rect 7316 27952 7317 27992
rect 7275 27943 7317 27952
rect 7372 27952 7508 27992
rect 7180 27607 7220 27616
rect 7276 27642 7316 27943
rect 7372 27749 7412 27952
rect 7371 27740 7413 27749
rect 7371 27700 7372 27740
rect 7412 27700 7413 27740
rect 7371 27691 7413 27700
rect 7468 27656 7508 27667
rect 6988 27522 7028 27607
rect 7276 27602 7412 27642
rect 7179 27404 7221 27413
rect 7179 27364 7180 27404
rect 7220 27364 7221 27404
rect 7179 27355 7221 27364
rect 7180 27270 7220 27355
rect 6891 27068 6933 27077
rect 6891 27028 6892 27068
rect 6932 27028 6933 27068
rect 6891 27019 6933 27028
rect 7275 26984 7317 26993
rect 7275 26944 7276 26984
rect 7316 26944 7317 26984
rect 7275 26935 7317 26944
rect 6891 26900 6933 26909
rect 6891 26860 6892 26900
rect 6932 26860 6933 26900
rect 6891 26851 6933 26860
rect 6796 26767 6836 26776
rect 6700 26682 6740 26767
rect 6795 26648 6837 26657
rect 6795 26608 6796 26648
rect 6836 26608 6837 26648
rect 6795 26599 6837 26608
rect 6603 26564 6645 26573
rect 6603 26524 6604 26564
rect 6644 26524 6645 26564
rect 6603 26515 6645 26524
rect 6507 26396 6549 26405
rect 6796 26396 6836 26599
rect 6507 26356 6508 26396
rect 6548 26356 6549 26396
rect 6507 26347 6549 26356
rect 6700 26356 6836 26396
rect 6412 26153 6452 26238
rect 6411 26144 6453 26153
rect 6411 26104 6412 26144
rect 6452 26104 6453 26144
rect 6604 26129 6644 26138
rect 6411 26095 6453 26104
rect 6508 26102 6548 26111
rect 6316 25936 6452 25976
rect 6315 25808 6357 25817
rect 6315 25768 6316 25808
rect 6356 25768 6357 25808
rect 6315 25759 6357 25768
rect 5643 25220 5685 25229
rect 5643 25180 5644 25220
rect 5684 25180 5685 25220
rect 5643 25171 5685 25180
rect 5452 24760 5588 24800
rect 5452 23960 5492 24760
rect 5547 24632 5589 24641
rect 5547 24592 5548 24632
rect 5588 24592 5589 24632
rect 5547 24583 5589 24592
rect 5548 24498 5588 24583
rect 5644 24128 5684 25171
rect 5740 24641 5780 25255
rect 5931 25052 5973 25061
rect 5931 25012 5932 25052
rect 5972 25012 5973 25052
rect 5931 25003 5973 25012
rect 5739 24632 5781 24641
rect 5739 24592 5740 24632
rect 5780 24592 5781 24632
rect 5739 24583 5781 24592
rect 5740 24380 5780 24389
rect 5780 24340 5876 24380
rect 5740 24331 5780 24340
rect 5644 24088 5780 24128
rect 5644 23960 5684 23971
rect 5452 23920 5588 23960
rect 5451 23792 5493 23801
rect 5451 23752 5452 23792
rect 5492 23752 5493 23792
rect 5451 23743 5493 23752
rect 5452 23658 5492 23743
rect 5355 23372 5397 23381
rect 5355 23332 5356 23372
rect 5396 23332 5397 23372
rect 5355 23323 5397 23332
rect 4971 23288 5013 23297
rect 4971 23248 4972 23288
rect 5012 23248 5013 23288
rect 4971 23239 5013 23248
rect 5451 23288 5493 23297
rect 5451 23248 5452 23288
rect 5492 23248 5493 23288
rect 5451 23239 5493 23248
rect 4972 23120 5012 23239
rect 5356 23129 5396 23214
rect 5452 23154 5492 23239
rect 4780 23080 4916 23120
rect 4779 22616 4821 22625
rect 4779 22576 4780 22616
rect 4820 22576 4821 22616
rect 4779 22567 4821 22576
rect 4780 22299 4820 22567
rect 4876 22532 4916 23080
rect 4972 22793 5012 23080
rect 5355 23120 5397 23129
rect 5355 23080 5356 23120
rect 5396 23080 5397 23120
rect 5355 23071 5397 23080
rect 5548 23120 5588 23920
rect 5644 23885 5684 23920
rect 5643 23876 5685 23885
rect 5643 23836 5644 23876
rect 5684 23836 5685 23876
rect 5643 23827 5685 23836
rect 5548 23036 5588 23080
rect 5644 23120 5684 23827
rect 5644 23071 5684 23080
rect 5452 22996 5588 23036
rect 5164 22868 5204 22877
rect 4971 22784 5013 22793
rect 4971 22744 4972 22784
rect 5012 22744 5013 22784
rect 4971 22735 5013 22744
rect 5164 22625 5204 22828
rect 5163 22616 5205 22625
rect 5163 22576 5164 22616
rect 5204 22576 5205 22616
rect 5163 22567 5205 22576
rect 4876 22492 5012 22532
rect 4875 22364 4917 22373
rect 4875 22324 4876 22364
rect 4916 22324 4917 22364
rect 4875 22315 4917 22324
rect 4780 22250 4820 22259
rect 4876 22280 4916 22315
rect 4876 22229 4916 22240
rect 4683 22196 4725 22205
rect 4683 22156 4684 22196
rect 4724 22156 4725 22196
rect 4683 22147 4725 22156
rect 4972 22112 5012 22492
rect 5259 22448 5301 22457
rect 5259 22408 5260 22448
rect 5300 22408 5301 22448
rect 5259 22399 5301 22408
rect 5260 22364 5300 22399
rect 5260 22313 5300 22324
rect 5356 22364 5396 22373
rect 5452 22364 5492 22996
rect 5547 22868 5589 22877
rect 5547 22828 5548 22868
rect 5588 22828 5589 22868
rect 5547 22819 5589 22828
rect 5396 22324 5492 22364
rect 4780 22072 5012 22112
rect 4780 21608 4820 22072
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4780 20357 4820 21568
rect 5356 20936 5396 22324
rect 5548 21449 5588 22819
rect 5643 22784 5685 22793
rect 5643 22744 5644 22784
rect 5684 22744 5685 22784
rect 5643 22735 5685 22744
rect 5644 21608 5684 22735
rect 5740 21944 5780 24088
rect 5836 23801 5876 24340
rect 5932 24044 5972 25003
rect 6123 24968 6165 24977
rect 6123 24928 6124 24968
rect 6164 24928 6165 24968
rect 6123 24919 6165 24928
rect 6124 24632 6164 24919
rect 6220 24809 6260 25264
rect 6316 25304 6356 25759
rect 6316 25255 6356 25264
rect 6412 25304 6452 25936
rect 6508 25817 6548 26062
rect 6604 25901 6644 26089
rect 6603 25892 6645 25901
rect 6603 25852 6604 25892
rect 6644 25852 6645 25892
rect 6603 25843 6645 25852
rect 6507 25808 6549 25817
rect 6507 25768 6508 25808
rect 6548 25768 6549 25808
rect 6507 25759 6549 25768
rect 6412 25255 6452 25264
rect 6315 25136 6357 25145
rect 6315 25096 6316 25136
rect 6356 25096 6357 25136
rect 6315 25087 6357 25096
rect 6219 24800 6261 24809
rect 6219 24760 6220 24800
rect 6260 24760 6261 24800
rect 6219 24751 6261 24760
rect 6027 24548 6069 24557
rect 6124 24548 6164 24592
rect 6027 24508 6028 24548
rect 6068 24508 6164 24548
rect 6027 24499 6069 24508
rect 6316 24221 6356 25087
rect 6315 24212 6357 24221
rect 6315 24172 6316 24212
rect 6356 24172 6357 24212
rect 6315 24163 6357 24172
rect 6508 24044 6548 25759
rect 6604 25304 6644 25843
rect 6604 25255 6644 25264
rect 6700 25304 6740 26356
rect 6700 25255 6740 25264
rect 6796 25892 6836 25901
rect 6796 25304 6836 25852
rect 6892 25817 6932 26851
rect 6988 26825 7028 26910
rect 6987 26816 7029 26825
rect 6987 26776 6988 26816
rect 7028 26776 7029 26816
rect 6987 26767 7029 26776
rect 7084 26816 7124 26825
rect 7084 26573 7124 26776
rect 7276 26816 7316 26935
rect 7276 26767 7316 26776
rect 7179 26648 7221 26657
rect 7179 26608 7180 26648
rect 7220 26608 7221 26648
rect 7179 26599 7221 26608
rect 7083 26564 7125 26573
rect 7083 26524 7084 26564
rect 7124 26524 7125 26564
rect 7083 26515 7125 26524
rect 7084 26153 7124 26515
rect 7180 26514 7220 26599
rect 7372 26396 7412 27602
rect 7468 27581 7508 27616
rect 7467 27572 7509 27581
rect 7467 27532 7468 27572
rect 7508 27532 7509 27572
rect 7467 27523 7509 27532
rect 7468 26993 7508 27078
rect 7467 26984 7509 26993
rect 7467 26944 7468 26984
rect 7508 26944 7509 26984
rect 7467 26935 7509 26944
rect 7467 26816 7509 26825
rect 7467 26776 7468 26816
rect 7508 26776 7509 26816
rect 7467 26767 7509 26776
rect 7180 26356 7412 26396
rect 7083 26144 7125 26153
rect 7083 26104 7084 26144
rect 7124 26104 7125 26144
rect 7083 26095 7125 26104
rect 6891 25808 6933 25817
rect 6891 25768 6892 25808
rect 6932 25768 6933 25808
rect 6891 25759 6933 25768
rect 7083 25472 7125 25481
rect 7083 25432 7084 25472
rect 7124 25432 7125 25472
rect 7083 25423 7125 25432
rect 6796 25255 6836 25264
rect 7084 25304 7124 25423
rect 7084 25255 7124 25264
rect 6699 25136 6741 25145
rect 6699 25096 6700 25136
rect 6740 25096 6741 25136
rect 6699 25087 6741 25096
rect 6891 25136 6933 25145
rect 6891 25096 6892 25136
rect 6932 25096 6933 25136
rect 6891 25087 6933 25096
rect 5932 24004 6068 24044
rect 5932 23885 5972 23929
rect 5931 23876 5973 23885
rect 5931 23836 5932 23876
rect 5972 23836 5973 23876
rect 5931 23834 5973 23836
rect 5931 23827 5932 23834
rect 5835 23792 5877 23801
rect 5835 23752 5836 23792
rect 5876 23752 5877 23792
rect 5972 23827 5973 23834
rect 5932 23785 5972 23794
rect 6028 23792 6068 24004
rect 6412 24004 6548 24044
rect 6124 23801 6164 23886
rect 5835 23743 5877 23752
rect 6028 23743 6068 23752
rect 6123 23792 6165 23801
rect 6123 23752 6124 23792
rect 6164 23752 6165 23792
rect 6123 23743 6165 23752
rect 5836 23120 5876 23743
rect 6316 23624 6356 23633
rect 6028 23584 6316 23624
rect 5931 23288 5973 23297
rect 5931 23248 5932 23288
rect 5972 23248 5973 23288
rect 5931 23239 5973 23248
rect 5836 23071 5876 23080
rect 5932 23120 5972 23239
rect 5932 23071 5972 23080
rect 6028 23120 6068 23584
rect 6316 23575 6356 23584
rect 6123 23288 6165 23297
rect 6123 23248 6124 23288
rect 6164 23248 6165 23288
rect 6123 23239 6165 23248
rect 6124 23154 6164 23239
rect 6028 23071 6068 23080
rect 6315 23120 6357 23129
rect 6315 23080 6316 23120
rect 6356 23080 6357 23120
rect 6315 23071 6357 23080
rect 6316 22986 6356 23071
rect 5835 22280 5877 22289
rect 5835 22240 5836 22280
rect 5876 22240 5877 22280
rect 5835 22231 5877 22240
rect 6316 22285 6356 22294
rect 5836 22121 5876 22231
rect 5835 22112 5877 22121
rect 5835 22072 5836 22112
rect 5876 22072 5877 22112
rect 5835 22063 5877 22072
rect 5740 21904 5876 21944
rect 5739 21608 5781 21617
rect 5644 21568 5740 21608
rect 5780 21568 5781 21608
rect 5739 21559 5781 21568
rect 5547 21440 5589 21449
rect 5547 21400 5548 21440
rect 5588 21400 5589 21440
rect 5547 21391 5589 21400
rect 5740 21197 5780 21559
rect 5739 21188 5781 21197
rect 5739 21148 5740 21188
rect 5780 21148 5781 21188
rect 5739 21139 5781 21148
rect 5164 20896 5396 20936
rect 5164 20609 5204 20896
rect 5260 20768 5300 20777
rect 5740 20768 5780 20777
rect 5300 20728 5396 20768
rect 5260 20719 5300 20728
rect 5163 20600 5205 20609
rect 5163 20560 5164 20600
rect 5204 20560 5205 20600
rect 5163 20551 5205 20560
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5356 20432 5396 20728
rect 5452 20684 5492 20693
rect 5740 20684 5780 20728
rect 5492 20644 5780 20684
rect 5836 20768 5876 21904
rect 6028 21617 6068 21702
rect 6220 21692 6260 21701
rect 6316 21692 6356 22245
rect 6260 21652 6356 21692
rect 6220 21643 6260 21652
rect 6027 21608 6069 21617
rect 6027 21568 6028 21608
rect 6068 21568 6069 21608
rect 6027 21559 6069 21568
rect 6027 21440 6069 21449
rect 6027 21400 6028 21440
rect 6068 21400 6069 21440
rect 6027 21391 6069 21400
rect 5452 20635 5492 20644
rect 5356 20392 5492 20432
rect 4928 20383 5296 20392
rect 4779 20348 4821 20357
rect 4779 20308 4780 20348
rect 4820 20308 4821 20348
rect 4779 20299 4821 20308
rect 4492 20140 4628 20180
rect 4492 20021 4532 20140
rect 4972 20096 5012 20105
rect 4780 20056 4972 20096
rect 4491 20012 4533 20021
rect 4491 19972 4492 20012
rect 4532 19972 4533 20012
rect 4491 19963 4533 19972
rect 4491 19844 4533 19853
rect 4491 19804 4492 19844
rect 4532 19804 4533 19844
rect 4491 19795 4533 19804
rect 4395 19340 4437 19349
rect 4395 19300 4396 19340
rect 4436 19300 4437 19340
rect 4395 19291 4437 19300
rect 4492 19270 4532 19795
rect 4299 19256 4341 19265
rect 4299 19216 4300 19256
rect 4340 19216 4341 19256
rect 4492 19221 4532 19230
rect 4299 19207 4341 19216
rect 4684 19088 4724 19097
rect 4684 18929 4724 19048
rect 4683 18920 4725 18929
rect 4683 18880 4684 18920
rect 4724 18880 4725 18920
rect 4683 18871 4725 18880
rect 4108 18712 4532 18752
rect 4108 18584 4148 18712
rect 4108 18535 4148 18544
rect 4204 18584 4244 18593
rect 3627 18500 3669 18509
rect 3627 18460 3628 18500
rect 3668 18460 3669 18500
rect 3627 18451 3669 18460
rect 3724 18500 3764 18509
rect 3628 18420 3668 18451
rect 3724 18332 3764 18460
rect 3436 18292 3764 18332
rect 3435 17660 3477 17669
rect 3435 17620 3436 17660
rect 3476 17620 3477 17660
rect 3435 17611 3477 17620
rect 3339 17408 3381 17417
rect 3339 17368 3340 17408
rect 3380 17368 3381 17408
rect 3339 17359 3381 17368
rect 3243 17240 3285 17249
rect 3243 17200 3244 17240
rect 3284 17200 3285 17240
rect 3243 17191 3285 17200
rect 3340 17030 3380 17083
rect 3339 16990 3340 16997
rect 3436 17072 3476 17611
rect 3436 17023 3476 17032
rect 3380 16990 3381 16997
rect 3339 16988 3381 16990
rect 3148 16948 3284 16988
rect 3052 16864 3188 16904
rect 3051 16484 3093 16493
rect 3051 16444 3052 16484
rect 3092 16444 3093 16484
rect 3051 16435 3093 16444
rect 3052 16232 3092 16435
rect 3148 16409 3188 16864
rect 3147 16400 3189 16409
rect 3147 16360 3148 16400
rect 3188 16360 3189 16400
rect 3147 16351 3189 16360
rect 3244 16316 3284 16948
rect 3339 16948 3340 16988
rect 3380 16948 3381 16988
rect 3339 16939 3381 16948
rect 3435 16820 3477 16829
rect 3435 16780 3436 16820
rect 3476 16780 3477 16820
rect 3435 16771 3477 16780
rect 3339 16652 3381 16661
rect 3339 16612 3340 16652
rect 3380 16612 3381 16652
rect 3339 16603 3381 16612
rect 3244 16267 3284 16276
rect 3148 16232 3188 16241
rect 3052 16192 3148 16232
rect 3148 16183 3188 16192
rect 3243 15980 3285 15989
rect 3243 15940 3244 15980
rect 3284 15940 3285 15980
rect 3243 15931 3285 15940
rect 3052 15476 3092 15485
rect 3052 15233 3092 15436
rect 3147 15308 3189 15317
rect 3147 15268 3148 15308
rect 3188 15268 3189 15308
rect 3147 15259 3189 15268
rect 3051 15224 3093 15233
rect 3051 15184 3052 15224
rect 3092 15184 3093 15224
rect 3051 15175 3093 15184
rect 3051 15056 3093 15065
rect 3051 15016 3052 15056
rect 3092 15016 3093 15056
rect 3051 15007 3093 15016
rect 2764 14428 2996 14468
rect 2667 14216 2709 14225
rect 2667 14176 2668 14216
rect 2708 14176 2709 14216
rect 2667 14167 2709 14176
rect 2668 14082 2708 14167
rect 2764 13628 2804 14428
rect 2956 14048 2996 14057
rect 2859 13964 2901 13973
rect 2859 13924 2860 13964
rect 2900 13924 2901 13964
rect 2859 13915 2901 13924
rect 2668 13588 2804 13628
rect 2668 11948 2708 13588
rect 2763 13376 2805 13385
rect 2763 13336 2764 13376
rect 2804 13336 2805 13376
rect 2763 13327 2805 13336
rect 2764 13292 2804 13327
rect 2764 13241 2804 13252
rect 2860 13208 2900 13915
rect 2763 12872 2805 12881
rect 2763 12832 2764 12872
rect 2804 12832 2805 12872
rect 2763 12823 2805 12832
rect 2764 12536 2804 12823
rect 2764 12487 2804 12496
rect 2763 12116 2805 12125
rect 2763 12076 2764 12116
rect 2804 12076 2805 12116
rect 2763 12067 2805 12076
rect 2668 11899 2708 11908
rect 2571 11612 2613 11621
rect 2571 11572 2572 11612
rect 2612 11572 2613 11612
rect 2571 11563 2613 11572
rect 2475 11444 2517 11453
rect 2475 11404 2476 11444
rect 2516 11404 2517 11444
rect 2475 11395 2517 11404
rect 2284 9512 2420 9532
rect 2188 9492 2420 9512
rect 2476 10184 2516 11395
rect 2571 11024 2613 11033
rect 2571 10984 2572 11024
rect 2612 10984 2613 11024
rect 2571 10975 2613 10984
rect 2668 11024 2708 11033
rect 2572 10890 2612 10975
rect 2668 10604 2708 10984
rect 2572 10564 2708 10604
rect 2572 10184 2612 10564
rect 2667 10436 2709 10445
rect 2667 10396 2668 10436
rect 2708 10396 2709 10436
rect 2667 10387 2709 10396
rect 2668 10302 2708 10387
rect 2572 10144 2708 10184
rect 2188 9472 2324 9492
rect 2091 8000 2133 8009
rect 2091 7960 2092 8000
rect 2132 7960 2133 8000
rect 2091 7951 2133 7960
rect 2188 7757 2228 9472
rect 2380 9428 2420 9437
rect 2380 9017 2420 9388
rect 2379 9008 2421 9017
rect 2379 8968 2380 9008
rect 2420 8968 2421 9008
rect 2379 8959 2421 8968
rect 2476 8672 2516 10144
rect 2571 9848 2613 9857
rect 2571 9808 2572 9848
rect 2612 9808 2613 9848
rect 2571 9799 2613 9808
rect 2572 8840 2612 9799
rect 2668 9680 2708 10144
rect 2764 9857 2804 12067
rect 2860 11948 2900 13168
rect 2956 12965 2996 14008
rect 3052 14048 3092 15007
rect 3052 13999 3092 14008
rect 2955 12956 2997 12965
rect 2955 12916 2956 12956
rect 2996 12916 2997 12956
rect 2955 12907 2997 12916
rect 3148 12125 3188 15259
rect 3244 15149 3284 15931
rect 3243 15140 3285 15149
rect 3243 15100 3244 15140
rect 3284 15100 3285 15140
rect 3243 15091 3285 15100
rect 3243 14720 3285 14729
rect 3243 14680 3244 14720
rect 3284 14680 3285 14720
rect 3243 14671 3285 14680
rect 3244 14586 3284 14671
rect 3243 14132 3285 14141
rect 3243 14092 3244 14132
rect 3284 14092 3285 14132
rect 3243 14083 3285 14092
rect 3244 12881 3284 14083
rect 3340 13208 3380 16603
rect 3436 14972 3476 16771
rect 3532 16493 3572 18292
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 3819 17072 3861 17081
rect 3819 17032 3820 17072
rect 3860 17032 3861 17072
rect 3819 17023 3861 17032
rect 3916 17072 3956 17081
rect 3956 17032 4148 17072
rect 3916 17023 3956 17032
rect 3820 16938 3860 17023
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3531 16484 3573 16493
rect 4108 16484 4148 17032
rect 3531 16444 3532 16484
rect 3572 16444 3573 16484
rect 3531 16435 3573 16444
rect 4012 16444 4148 16484
rect 3723 16400 3765 16409
rect 3723 16360 3724 16400
rect 3764 16360 3765 16400
rect 3723 16351 3765 16360
rect 3531 16316 3573 16325
rect 3531 16276 3532 16316
rect 3572 16276 3573 16316
rect 3531 16267 3573 16276
rect 3436 14923 3476 14932
rect 3532 14804 3572 16267
rect 3724 16232 3764 16351
rect 3764 16192 3860 16232
rect 3724 16183 3764 16192
rect 3723 15644 3765 15653
rect 3723 15604 3724 15644
rect 3764 15604 3765 15644
rect 3723 15595 3765 15604
rect 3724 15560 3764 15595
rect 3724 15509 3764 15520
rect 3820 15401 3860 16192
rect 3819 15392 3861 15401
rect 3819 15352 3820 15392
rect 3860 15352 3861 15392
rect 3819 15343 3861 15352
rect 4012 15317 4052 16444
rect 4204 16400 4244 18544
rect 4396 17744 4436 17753
rect 4396 16409 4436 17704
rect 4108 16360 4244 16400
rect 4395 16400 4437 16409
rect 4395 16360 4396 16400
rect 4436 16360 4437 16400
rect 4011 15308 4053 15317
rect 4011 15268 4012 15308
rect 4052 15268 4053 15308
rect 4011 15259 4053 15268
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3436 14764 3572 14804
rect 3819 14804 3861 14813
rect 3819 14764 3820 14804
rect 3860 14764 3861 14804
rect 3436 14048 3476 14764
rect 3819 14755 3861 14764
rect 3820 14670 3860 14755
rect 3628 14552 3668 14561
rect 3436 13385 3476 14008
rect 3531 14048 3573 14057
rect 3531 14008 3532 14048
rect 3572 14008 3573 14048
rect 3531 13999 3573 14008
rect 3532 13914 3572 13999
rect 3628 13889 3668 14512
rect 4108 14225 4148 16360
rect 4395 16351 4437 16360
rect 4252 16241 4292 16250
rect 4292 16201 4340 16232
rect 4252 16192 4340 16201
rect 4203 14888 4245 14897
rect 4203 14848 4204 14888
rect 4244 14848 4245 14888
rect 4203 14839 4245 14848
rect 4204 14720 4244 14839
rect 4107 14216 4149 14225
rect 4107 14176 4108 14216
rect 4148 14176 4149 14216
rect 4107 14167 4149 14176
rect 4012 14048 4052 14059
rect 4012 13973 4052 14008
rect 4011 13964 4053 13973
rect 4011 13924 4012 13964
rect 4052 13924 4053 13964
rect 4011 13915 4053 13924
rect 3627 13880 3669 13889
rect 3627 13840 3628 13880
rect 3668 13840 3669 13880
rect 3627 13831 3669 13840
rect 3688 13628 4056 13637
rect 4204 13628 4244 14680
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 4108 13588 4244 13628
rect 3435 13376 3477 13385
rect 3435 13336 3436 13376
rect 3476 13336 3477 13376
rect 3435 13327 3477 13336
rect 3820 13213 3860 13222
rect 3380 13168 3572 13208
rect 3340 13159 3380 13168
rect 3243 12872 3285 12881
rect 3243 12832 3244 12872
rect 3284 12832 3285 12872
rect 3243 12823 3285 12832
rect 3339 12284 3381 12293
rect 3339 12244 3340 12284
rect 3380 12244 3381 12284
rect 3339 12235 3381 12244
rect 3147 12116 3189 12125
rect 3147 12076 3148 12116
rect 3188 12076 3189 12116
rect 3147 12067 3189 12076
rect 2860 11908 3188 11948
rect 3051 11780 3093 11789
rect 3051 11740 3052 11780
rect 3092 11740 3093 11780
rect 3051 11731 3093 11740
rect 3052 11646 3092 11731
rect 2859 11528 2901 11537
rect 2859 11488 2860 11528
rect 2900 11488 2901 11528
rect 2859 11479 2901 11488
rect 2860 11394 2900 11479
rect 2955 11024 2997 11033
rect 2955 10984 2956 11024
rect 2996 10984 2997 11024
rect 2955 10975 2997 10984
rect 2859 10352 2901 10361
rect 2859 10312 2860 10352
rect 2900 10312 2901 10352
rect 2859 10303 2901 10312
rect 2860 10218 2900 10303
rect 2763 9848 2805 9857
rect 2763 9808 2764 9848
rect 2804 9808 2805 9848
rect 2763 9799 2805 9808
rect 2763 9680 2805 9689
rect 2668 9640 2764 9680
rect 2804 9640 2805 9680
rect 2763 9631 2805 9640
rect 2668 9512 2708 9521
rect 2668 9101 2708 9472
rect 2764 9512 2804 9631
rect 2764 9463 2804 9472
rect 2763 9344 2805 9353
rect 2763 9304 2764 9344
rect 2804 9304 2805 9344
rect 2763 9295 2805 9304
rect 2667 9092 2709 9101
rect 2667 9052 2668 9092
rect 2708 9052 2709 9092
rect 2667 9043 2709 9052
rect 2668 8840 2708 8849
rect 2572 8800 2668 8840
rect 2668 8791 2708 8800
rect 2516 8632 2612 8672
rect 2476 8623 2516 8632
rect 2379 8588 2421 8597
rect 2379 8548 2380 8588
rect 2420 8548 2421 8588
rect 2379 8539 2421 8548
rect 2187 7748 2229 7757
rect 2187 7708 2188 7748
rect 2228 7708 2229 7748
rect 2187 7699 2229 7708
rect 2187 6992 2229 7001
rect 2187 6952 2188 6992
rect 2228 6952 2229 6992
rect 2187 6943 2229 6952
rect 1900 5692 2036 5732
rect 2092 5732 2132 5741
rect 1900 4565 1940 5692
rect 1995 5564 2037 5573
rect 1995 5524 1996 5564
rect 2036 5524 2037 5564
rect 1995 5515 2037 5524
rect 1899 4556 1941 4565
rect 1899 4516 1900 4556
rect 1940 4516 1941 4556
rect 1899 4507 1941 4516
rect 1804 4096 1940 4136
rect 1803 3968 1845 3977
rect 1803 3928 1804 3968
rect 1844 3928 1845 3968
rect 1803 3919 1845 3928
rect 1708 3331 1748 3340
rect 1228 1903 1268 1912
rect 1324 3088 1460 3128
rect 1324 1112 1364 3088
rect 1420 2624 1460 2633
rect 1420 1457 1460 2584
rect 1419 1448 1461 1457
rect 1419 1408 1420 1448
rect 1460 1408 1461 1448
rect 1419 1399 1461 1408
rect 1324 1063 1364 1072
rect 1035 944 1077 953
rect 1035 904 1036 944
rect 1076 904 1077 944
rect 1035 895 1077 904
rect 1804 80 1844 3919
rect 1900 3809 1940 4096
rect 1899 3800 1941 3809
rect 1899 3760 1900 3800
rect 1940 3760 1941 3800
rect 1899 3751 1941 3760
rect 1900 3380 1940 3389
rect 1900 197 1940 3340
rect 1899 188 1941 197
rect 1899 148 1900 188
rect 1940 148 1941 188
rect 1899 139 1941 148
rect 1996 80 2036 5515
rect 2092 5405 2132 5692
rect 2091 5396 2133 5405
rect 2091 5356 2092 5396
rect 2132 5356 2133 5396
rect 2091 5347 2133 5356
rect 2188 4724 2228 6943
rect 2283 6656 2325 6665
rect 2283 6616 2284 6656
rect 2324 6616 2325 6656
rect 2283 6607 2325 6616
rect 2284 5648 2324 6607
rect 2380 6488 2420 8539
rect 2475 8336 2517 8345
rect 2475 8296 2476 8336
rect 2516 8296 2517 8336
rect 2475 8287 2517 8296
rect 2476 8009 2516 8287
rect 2475 8000 2517 8009
rect 2475 7960 2476 8000
rect 2516 7960 2517 8000
rect 2475 7951 2517 7960
rect 2475 7748 2517 7757
rect 2475 7708 2476 7748
rect 2516 7708 2517 7748
rect 2475 7699 2517 7708
rect 2476 6908 2516 7699
rect 2572 7169 2612 8632
rect 2668 8168 2708 8177
rect 2764 8168 2804 9295
rect 2859 8672 2901 8681
rect 2859 8632 2860 8672
rect 2900 8632 2901 8672
rect 2859 8623 2901 8632
rect 2860 8538 2900 8623
rect 2956 8504 2996 10975
rect 3052 10940 3092 10949
rect 3052 10613 3092 10900
rect 3148 10940 3188 11908
rect 3244 11864 3284 11873
rect 3244 11705 3284 11824
rect 3243 11696 3285 11705
rect 3243 11656 3244 11696
rect 3284 11656 3285 11696
rect 3243 11647 3285 11656
rect 3188 10900 3284 10940
rect 3148 10891 3188 10900
rect 3051 10604 3093 10613
rect 3051 10564 3052 10604
rect 3092 10564 3093 10604
rect 3051 10555 3093 10564
rect 3051 10268 3093 10277
rect 3051 10228 3052 10268
rect 3092 10228 3093 10268
rect 3051 10219 3093 10228
rect 3052 10134 3092 10219
rect 3147 9596 3189 9605
rect 3147 9556 3148 9596
rect 3188 9556 3189 9596
rect 3147 9547 3189 9556
rect 3051 9512 3093 9521
rect 3051 9472 3052 9512
rect 3092 9472 3093 9512
rect 3051 9463 3093 9472
rect 3148 9512 3188 9547
rect 3052 8681 3092 9463
rect 3148 9461 3188 9472
rect 3244 9512 3284 10900
rect 3244 9463 3284 9472
rect 3243 8840 3285 8849
rect 3243 8800 3244 8840
rect 3284 8800 3285 8840
rect 3243 8791 3285 8800
rect 3051 8672 3093 8681
rect 3051 8632 3052 8672
rect 3092 8632 3093 8672
rect 3051 8623 3093 8632
rect 2956 8464 3102 8504
rect 2859 8420 2901 8429
rect 2859 8380 2860 8420
rect 2900 8380 2901 8420
rect 2859 8371 2901 8380
rect 2708 8128 2804 8168
rect 2860 8168 2900 8371
rect 3062 8336 3102 8464
rect 3147 8420 3189 8429
rect 3147 8380 3148 8420
rect 3188 8380 3189 8420
rect 3147 8371 3189 8380
rect 2668 8119 2708 8128
rect 2860 8119 2900 8128
rect 2956 8296 3102 8336
rect 2667 8000 2709 8009
rect 2667 7960 2668 8000
rect 2708 7960 2709 8000
rect 2667 7951 2709 7960
rect 2571 7160 2613 7169
rect 2571 7120 2572 7160
rect 2612 7120 2613 7160
rect 2571 7111 2613 7120
rect 2476 6868 2612 6908
rect 2476 6488 2516 6497
rect 2380 6448 2476 6488
rect 2476 6439 2516 6448
rect 2380 5648 2420 5657
rect 2284 5608 2380 5648
rect 2380 5599 2420 5608
rect 2475 5312 2517 5321
rect 2475 5272 2476 5312
rect 2516 5272 2517 5312
rect 2475 5263 2517 5272
rect 2476 4976 2516 5263
rect 2572 5060 2612 6868
rect 2668 6656 2708 7951
rect 2956 7580 2996 8296
rect 3052 7916 3092 7925
rect 3148 7916 3188 8371
rect 3244 8168 3284 8791
rect 3244 8119 3284 8128
rect 3092 7876 3188 7916
rect 3052 7867 3092 7876
rect 2860 7540 2996 7580
rect 2763 7160 2805 7169
rect 2763 7120 2764 7160
rect 2804 7120 2805 7160
rect 2763 7111 2805 7120
rect 2668 6607 2708 6616
rect 2667 6320 2709 6329
rect 2667 6280 2668 6320
rect 2708 6280 2709 6320
rect 2667 6271 2709 6280
rect 2668 5741 2708 6271
rect 2667 5732 2709 5741
rect 2667 5692 2668 5732
rect 2708 5692 2709 5732
rect 2667 5683 2709 5692
rect 2764 5321 2804 7111
rect 2763 5312 2805 5321
rect 2763 5272 2764 5312
rect 2804 5272 2805 5312
rect 2763 5263 2805 5272
rect 2860 5144 2900 7540
rect 3340 7505 3380 12235
rect 3436 11780 3476 11789
rect 3436 10361 3476 11740
rect 3532 11024 3572 13168
rect 3820 12293 3860 13173
rect 4012 13040 4052 13049
rect 4012 12881 4052 13000
rect 4011 12872 4053 12881
rect 4011 12832 4012 12872
rect 4052 12832 4053 12872
rect 4011 12823 4053 12832
rect 4012 12536 4052 12545
rect 4012 12293 4052 12496
rect 3819 12284 3861 12293
rect 3819 12244 3820 12284
rect 3860 12244 3861 12284
rect 3819 12235 3861 12244
rect 4011 12284 4053 12293
rect 4011 12244 4012 12284
rect 4052 12244 4053 12284
rect 4011 12235 4053 12244
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 4108 11948 4148 13588
rect 4204 13292 4244 13301
rect 4204 12965 4244 13252
rect 4203 12956 4245 12965
rect 4203 12916 4204 12956
rect 4244 12916 4245 12956
rect 4203 12907 4245 12916
rect 4204 12620 4244 12629
rect 4300 12620 4340 16192
rect 4396 16064 4436 16073
rect 4396 15149 4436 16024
rect 4492 15989 4532 18712
rect 4683 17072 4725 17081
rect 4683 17032 4684 17072
rect 4724 17032 4725 17072
rect 4683 17023 4725 17032
rect 4491 15980 4533 15989
rect 4491 15940 4492 15980
rect 4532 15940 4533 15980
rect 4491 15931 4533 15940
rect 4395 15140 4437 15149
rect 4395 15100 4396 15140
rect 4436 15100 4437 15140
rect 4395 15091 4437 15100
rect 4684 15065 4724 17023
rect 4780 15560 4820 20056
rect 4972 20047 5012 20056
rect 5356 20096 5396 20105
rect 5356 19937 5396 20056
rect 5355 19928 5397 19937
rect 5355 19888 5356 19928
rect 5396 19888 5397 19928
rect 5355 19879 5397 19888
rect 5163 19844 5205 19853
rect 5163 19804 5164 19844
rect 5204 19804 5205 19844
rect 5163 19795 5205 19804
rect 5164 19710 5204 19795
rect 5452 19769 5492 20392
rect 5451 19760 5493 19769
rect 5451 19720 5452 19760
rect 5492 19720 5493 19760
rect 5451 19711 5493 19720
rect 5355 19592 5397 19601
rect 5355 19552 5356 19592
rect 5396 19552 5397 19592
rect 5355 19543 5397 19552
rect 5356 19256 5396 19543
rect 5356 18929 5396 19216
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 5355 18920 5397 18929
rect 5355 18880 5356 18920
rect 5396 18880 5397 18920
rect 5355 18871 5397 18880
rect 5451 18836 5493 18845
rect 5451 18796 5452 18836
rect 5492 18796 5493 18836
rect 5451 18787 5493 18796
rect 5452 17753 5492 18787
rect 5548 18712 5780 18752
rect 5451 17744 5493 17753
rect 5451 17704 5452 17744
rect 5492 17704 5493 17744
rect 5451 17695 5493 17704
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 5548 17081 5588 18712
rect 5644 18584 5684 18593
rect 5644 17996 5684 18544
rect 5740 18584 5780 18712
rect 5740 18535 5780 18544
rect 5836 18164 5876 20728
rect 6028 18845 6068 21391
rect 6219 21356 6261 21365
rect 6219 21316 6220 21356
rect 6260 21316 6261 21356
rect 6219 21307 6261 21316
rect 6123 21188 6165 21197
rect 6123 21148 6124 21188
rect 6164 21148 6165 21188
rect 6123 21139 6165 21148
rect 6124 19769 6164 21139
rect 6220 20768 6260 21307
rect 6315 20936 6357 20945
rect 6315 20896 6316 20936
rect 6356 20896 6357 20936
rect 6315 20887 6357 20896
rect 6316 20852 6356 20887
rect 6316 20801 6356 20812
rect 6123 19760 6165 19769
rect 6123 19720 6124 19760
rect 6164 19720 6165 19760
rect 6123 19711 6165 19720
rect 6027 18836 6069 18845
rect 6027 18796 6028 18836
rect 6068 18796 6069 18836
rect 6027 18787 6069 18796
rect 6220 18668 6260 20728
rect 6315 20684 6357 20693
rect 6315 20644 6316 20684
rect 6356 20644 6357 20684
rect 6315 20635 6357 20644
rect 6316 19097 6356 20635
rect 6315 19088 6357 19097
rect 6315 19048 6316 19088
rect 6356 19048 6357 19088
rect 6315 19039 6357 19048
rect 6028 18628 6260 18668
rect 6028 18257 6068 18628
rect 6316 18584 6356 19039
rect 6220 18544 6356 18584
rect 6124 18500 6164 18511
rect 6124 18425 6164 18460
rect 6220 18500 6260 18544
rect 6220 18451 6260 18460
rect 6123 18416 6165 18425
rect 6123 18376 6124 18416
rect 6164 18376 6165 18416
rect 6123 18367 6165 18376
rect 6027 18248 6069 18257
rect 6027 18208 6028 18248
rect 6068 18208 6069 18248
rect 6027 18199 6069 18208
rect 5836 18124 5972 18164
rect 5836 17996 5876 18005
rect 5644 17956 5836 17996
rect 5836 17947 5876 17956
rect 5643 17744 5685 17753
rect 5643 17704 5644 17744
rect 5684 17704 5685 17744
rect 5643 17695 5685 17704
rect 5260 17072 5300 17081
rect 5260 16232 5300 17032
rect 5355 17072 5397 17081
rect 5355 17032 5356 17072
rect 5396 17032 5397 17072
rect 5355 17023 5397 17032
rect 5547 17072 5589 17081
rect 5547 17032 5548 17072
rect 5588 17032 5589 17072
rect 5547 17023 5589 17032
rect 5356 16938 5396 17023
rect 5644 16400 5684 17695
rect 5740 16988 5780 16997
rect 5740 16577 5780 16948
rect 5835 16988 5877 16997
rect 5835 16948 5836 16988
rect 5876 16948 5877 16988
rect 5835 16939 5877 16948
rect 5836 16854 5876 16939
rect 5932 16745 5972 18124
rect 6027 17744 6069 17753
rect 6027 17704 6028 17744
rect 6068 17704 6069 17744
rect 6027 17695 6069 17704
rect 5931 16736 5973 16745
rect 5931 16696 5932 16736
rect 5972 16696 5973 16736
rect 5931 16687 5973 16696
rect 5739 16568 5781 16577
rect 5739 16528 5740 16568
rect 5780 16528 5781 16568
rect 5739 16519 5781 16528
rect 5644 16360 5876 16400
rect 5644 16232 5684 16241
rect 5260 16192 5396 16232
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 5164 15728 5204 15737
rect 5356 15728 5396 16192
rect 5204 15688 5396 15728
rect 5164 15679 5204 15688
rect 4971 15560 5013 15569
rect 5356 15560 5396 15569
rect 4780 15520 4972 15560
rect 5012 15520 5013 15560
rect 4971 15511 5013 15520
rect 5355 15520 5356 15560
rect 5355 15511 5396 15520
rect 4972 15426 5012 15511
rect 5259 15476 5301 15485
rect 5355 15476 5395 15511
rect 5259 15436 5260 15476
rect 5300 15436 5395 15476
rect 5259 15427 5301 15436
rect 4779 15308 4821 15317
rect 4779 15268 4780 15308
rect 4820 15268 4821 15308
rect 4779 15259 4821 15268
rect 4683 15056 4725 15065
rect 4683 15016 4684 15056
rect 4724 15016 4725 15056
rect 4683 15007 4725 15016
rect 4684 14561 4724 15007
rect 4683 14552 4725 14561
rect 4683 14512 4684 14552
rect 4724 14512 4725 14552
rect 4683 14503 4725 14512
rect 4684 14132 4724 14141
rect 4492 14034 4532 14043
rect 4395 13712 4437 13721
rect 4395 13672 4396 13712
rect 4436 13672 4437 13712
rect 4395 13663 4437 13672
rect 4396 13460 4436 13663
rect 4396 13411 4436 13420
rect 4244 12580 4340 12620
rect 4204 12571 4244 12580
rect 4492 12452 4532 13994
rect 4684 12797 4724 14092
rect 4683 12788 4725 12797
rect 4683 12748 4684 12788
rect 4724 12748 4725 12788
rect 4683 12739 4725 12748
rect 4684 12536 4724 12545
rect 4492 12412 4628 12452
rect 4491 12284 4533 12293
rect 4491 12244 4492 12284
rect 4532 12244 4533 12284
rect 4491 12235 4533 12244
rect 4012 11908 4148 11948
rect 3820 11780 3860 11789
rect 3627 11528 3669 11537
rect 3627 11488 3628 11528
rect 3668 11488 3669 11528
rect 3627 11479 3669 11488
rect 3628 11394 3668 11479
rect 3820 11033 3860 11740
rect 4012 11201 4052 11908
rect 4203 11864 4245 11873
rect 4203 11824 4204 11864
rect 4244 11824 4245 11864
rect 4203 11815 4245 11824
rect 4107 11696 4149 11705
rect 4107 11656 4108 11696
rect 4148 11656 4149 11696
rect 4107 11647 4149 11656
rect 4108 11562 4148 11647
rect 4204 11360 4244 11815
rect 4204 11320 4436 11360
rect 4011 11192 4053 11201
rect 4011 11152 4012 11192
rect 4052 11152 4053 11192
rect 4011 11143 4053 11152
rect 4300 11108 4340 11117
rect 4300 11033 4340 11068
rect 3628 11024 3668 11033
rect 3532 10984 3628 11024
rect 3532 10445 3572 10984
rect 3628 10975 3668 10984
rect 3819 11024 3861 11033
rect 3819 10984 3820 11024
rect 3860 10984 3861 11024
rect 4300 11024 4352 11033
rect 3819 10975 3861 10984
rect 4108 11010 4148 11019
rect 4300 10984 4311 11024
rect 4351 10984 4352 11024
rect 4310 10975 4352 10984
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 3531 10436 3573 10445
rect 3531 10396 3532 10436
rect 3572 10396 3573 10436
rect 3531 10387 3573 10396
rect 3819 10436 3861 10445
rect 3819 10396 3820 10436
rect 3860 10396 3861 10436
rect 3819 10387 3861 10396
rect 3435 10352 3477 10361
rect 3435 10312 3436 10352
rect 3476 10312 3477 10352
rect 3435 10303 3477 10312
rect 3723 10184 3765 10193
rect 3532 10142 3572 10151
rect 3531 10102 3532 10109
rect 3723 10144 3724 10184
rect 3764 10144 3765 10184
rect 3723 10135 3765 10144
rect 3572 10102 3573 10109
rect 3531 10100 3573 10102
rect 3531 10060 3532 10100
rect 3572 10060 3573 10100
rect 3531 10051 3573 10060
rect 3435 10016 3477 10025
rect 3435 9976 3436 10016
rect 3476 9976 3477 10016
rect 3532 10007 3572 10051
rect 3435 9967 3477 9976
rect 3436 8093 3476 9967
rect 3724 9689 3764 10135
rect 3723 9680 3765 9689
rect 3723 9640 3724 9680
rect 3764 9640 3765 9680
rect 3723 9631 3765 9640
rect 3723 9512 3765 9521
rect 3820 9512 3860 10387
rect 3723 9472 3724 9512
rect 3764 9472 3860 9512
rect 3723 9463 3765 9472
rect 3724 9378 3764 9463
rect 3531 9092 3573 9101
rect 3531 9052 3532 9092
rect 3572 9052 3573 9092
rect 3531 9043 3573 9052
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3532 8177 3572 9043
rect 3627 8924 3669 8933
rect 3627 8884 3628 8924
rect 3668 8884 3669 8924
rect 3627 8875 3669 8884
rect 3628 8513 3668 8875
rect 4108 8849 4148 10970
rect 4203 10940 4245 10949
rect 4203 10900 4204 10940
rect 4244 10900 4245 10940
rect 4203 10891 4245 10900
rect 4204 9848 4244 10891
rect 4396 10856 4436 11320
rect 4492 10949 4532 12235
rect 4491 10940 4533 10949
rect 4491 10900 4492 10940
rect 4532 10900 4533 10940
rect 4491 10891 4533 10900
rect 4300 10816 4436 10856
rect 4300 10025 4340 10816
rect 4491 10772 4533 10781
rect 4491 10732 4492 10772
rect 4532 10732 4533 10772
rect 4491 10723 4533 10732
rect 4492 10638 4532 10723
rect 4395 10604 4437 10613
rect 4395 10564 4396 10604
rect 4436 10564 4437 10604
rect 4395 10555 4437 10564
rect 4299 10016 4341 10025
rect 4299 9976 4300 10016
rect 4340 9976 4341 10016
rect 4299 9967 4341 9976
rect 4204 9808 4340 9848
rect 4204 9521 4244 9602
rect 4203 9512 4245 9521
rect 4203 9467 4204 9512
rect 4244 9467 4245 9512
rect 4203 9463 4245 9467
rect 4204 9458 4244 9463
rect 4300 9344 4340 9808
rect 4396 9680 4436 10555
rect 4588 10529 4628 12412
rect 4684 12125 4724 12496
rect 4683 12116 4725 12125
rect 4683 12076 4684 12116
rect 4724 12076 4725 12116
rect 4683 12067 4725 12076
rect 4684 10940 4724 10949
rect 4684 10781 4724 10900
rect 4683 10772 4725 10781
rect 4683 10732 4684 10772
rect 4724 10732 4725 10772
rect 4683 10723 4725 10732
rect 4587 10520 4629 10529
rect 4587 10480 4588 10520
rect 4628 10480 4629 10520
rect 4587 10471 4629 10480
rect 4780 10352 4820 15259
rect 5355 15140 5397 15149
rect 5355 15100 5356 15140
rect 5396 15100 5397 15140
rect 5355 15091 5397 15100
rect 5547 15140 5589 15149
rect 5547 15100 5548 15140
rect 5588 15100 5589 15140
rect 5547 15091 5589 15100
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 5259 12620 5301 12629
rect 5259 12580 5260 12620
rect 5300 12580 5301 12620
rect 5259 12571 5301 12580
rect 5260 11696 5300 12571
rect 5356 11864 5396 15091
rect 5451 14720 5493 14729
rect 5451 14680 5452 14720
rect 5492 14680 5493 14720
rect 5451 14671 5493 14680
rect 5452 14586 5492 14671
rect 5452 13208 5492 13217
rect 5452 12368 5492 13168
rect 5548 13208 5588 15091
rect 5644 14972 5684 16192
rect 5740 16232 5780 16241
rect 5740 15989 5780 16192
rect 5739 15980 5781 15989
rect 5739 15940 5740 15980
rect 5780 15940 5781 15980
rect 5739 15931 5781 15940
rect 5644 14923 5684 14932
rect 5588 13168 5684 13208
rect 5548 13159 5588 13168
rect 5452 12328 5588 12368
rect 5548 11948 5588 12328
rect 5548 11899 5588 11908
rect 5356 11824 5492 11864
rect 5356 11696 5396 11705
rect 5260 11656 5356 11696
rect 5356 11647 5396 11656
rect 4928 11360 5296 11369
rect 5452 11360 5492 11824
rect 5644 11360 5684 13168
rect 5739 12872 5781 12881
rect 5739 12832 5740 12872
rect 5780 12832 5781 12872
rect 5739 12823 5781 12832
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 5356 11320 5492 11360
rect 5548 11320 5684 11360
rect 5259 11024 5301 11033
rect 5259 10984 5260 11024
rect 5300 10984 5301 11024
rect 5259 10975 5301 10984
rect 4875 10940 4917 10949
rect 4875 10900 4876 10940
rect 4916 10900 4917 10940
rect 4875 10891 4917 10900
rect 4876 10806 4916 10891
rect 5068 10772 5108 10781
rect 4971 10520 5013 10529
rect 4971 10480 4972 10520
rect 5012 10480 5013 10520
rect 4971 10471 5013 10480
rect 4972 10436 5012 10471
rect 4972 10385 5012 10396
rect 4396 9631 4436 9640
rect 4492 10312 4820 10352
rect 4395 9512 4437 9521
rect 4395 9472 4396 9512
rect 4436 9472 4437 9512
rect 4395 9463 4437 9472
rect 4204 9304 4340 9344
rect 4107 8840 4149 8849
rect 4107 8800 4108 8840
rect 4148 8800 4149 8840
rect 4107 8791 4149 8800
rect 3819 8756 3861 8765
rect 3819 8716 3820 8756
rect 3860 8716 3861 8756
rect 3819 8707 3861 8716
rect 3627 8504 3669 8513
rect 3627 8464 3628 8504
rect 3668 8464 3669 8504
rect 3627 8455 3669 8464
rect 3531 8168 3573 8177
rect 3531 8128 3532 8168
rect 3572 8128 3573 8168
rect 3531 8119 3573 8128
rect 3435 8084 3477 8093
rect 3435 8044 3436 8084
rect 3476 8044 3477 8084
rect 3435 8035 3477 8044
rect 3435 7916 3477 7925
rect 3435 7876 3436 7916
rect 3476 7876 3477 7916
rect 3435 7867 3477 7876
rect 3820 7916 3860 8707
rect 4108 8672 4148 8683
rect 4108 8597 4148 8632
rect 4107 8588 4149 8597
rect 4107 8548 4108 8588
rect 4148 8548 4149 8588
rect 4107 8539 4149 8548
rect 4204 8345 4244 9304
rect 4299 8840 4341 8849
rect 4299 8800 4300 8840
rect 4340 8800 4341 8840
rect 4299 8791 4341 8800
rect 4300 8706 4340 8791
rect 4203 8336 4245 8345
rect 4203 8296 4204 8336
rect 4244 8296 4245 8336
rect 4203 8287 4245 8296
rect 4203 8000 4245 8009
rect 4203 7960 4204 8000
rect 4244 7960 4245 8000
rect 4203 7951 4245 7960
rect 3820 7867 3860 7876
rect 3436 7782 3476 7867
rect 4012 7841 4052 7926
rect 4204 7866 4244 7951
rect 4011 7832 4053 7841
rect 4011 7792 4012 7832
rect 4052 7792 4053 7832
rect 4011 7783 4053 7792
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3339 7496 3381 7505
rect 3339 7456 3340 7496
rect 3380 7456 3381 7496
rect 3339 7447 3381 7456
rect 2955 7412 2997 7421
rect 2955 7372 2956 7412
rect 2996 7372 2997 7412
rect 2955 7363 2997 7372
rect 3819 7412 3861 7421
rect 4396 7412 4436 9463
rect 3819 7372 3820 7412
rect 3860 7372 3861 7412
rect 3819 7363 3861 7372
rect 4204 7372 4436 7412
rect 2956 7278 2996 7363
rect 3723 7328 3765 7337
rect 3723 7288 3724 7328
rect 3764 7288 3765 7328
rect 3723 7279 3765 7288
rect 3724 7244 3764 7279
rect 3244 7160 3284 7169
rect 3147 6824 3189 6833
rect 3147 6784 3148 6824
rect 3188 6784 3189 6824
rect 3147 6775 3189 6784
rect 3051 6488 3093 6497
rect 3051 6448 3052 6488
rect 3092 6448 3093 6488
rect 3051 6439 3093 6448
rect 3148 6488 3188 6775
rect 3148 6439 3188 6448
rect 3052 6354 3092 6439
rect 3051 5732 3093 5741
rect 3051 5692 3052 5732
rect 3092 5692 3093 5732
rect 3051 5683 3093 5692
rect 2764 5104 2900 5144
rect 2668 5060 2708 5069
rect 2572 5020 2668 5060
rect 2668 5011 2708 5020
rect 2188 4684 2420 4724
rect 2187 4556 2229 4565
rect 2187 4516 2188 4556
rect 2228 4516 2229 4556
rect 2187 4507 2229 4516
rect 2091 3632 2133 3641
rect 2091 3592 2092 3632
rect 2132 3592 2133 3632
rect 2091 3583 2133 3592
rect 2092 3498 2132 3583
rect 2188 80 2228 4507
rect 2283 3464 2325 3473
rect 2283 3424 2284 3464
rect 2324 3424 2325 3464
rect 2283 3415 2325 3424
rect 2284 3330 2324 3415
rect 2380 80 2420 4684
rect 2476 4136 2516 4936
rect 2668 4388 2708 4397
rect 2764 4388 2804 5104
rect 2860 4976 2900 4985
rect 2860 4649 2900 4936
rect 2955 4892 2997 4901
rect 2955 4852 2956 4892
rect 2996 4852 2997 4892
rect 2955 4843 2997 4852
rect 2859 4640 2901 4649
rect 2859 4600 2860 4640
rect 2900 4600 2901 4640
rect 2859 4591 2901 4600
rect 2708 4348 2804 4388
rect 2668 4339 2708 4348
rect 2859 4304 2901 4313
rect 2859 4264 2860 4304
rect 2900 4264 2901 4304
rect 2859 4255 2901 4264
rect 2860 4170 2900 4255
rect 2476 3641 2516 4096
rect 2571 3884 2613 3893
rect 2571 3844 2572 3884
rect 2612 3844 2613 3884
rect 2571 3835 2613 3844
rect 2475 3632 2517 3641
rect 2475 3592 2476 3632
rect 2516 3592 2517 3632
rect 2475 3583 2517 3592
rect 2572 3464 2612 3835
rect 2763 3548 2805 3557
rect 2763 3508 2764 3548
rect 2804 3508 2805 3548
rect 2763 3499 2805 3508
rect 2476 3424 2612 3464
rect 2476 1952 2516 3424
rect 2764 3053 2804 3499
rect 2763 3044 2805 3053
rect 2763 3004 2764 3044
rect 2804 3004 2805 3044
rect 2763 2995 2805 3004
rect 2668 2624 2708 2633
rect 2668 2549 2708 2584
rect 2667 2540 2709 2549
rect 2667 2500 2668 2540
rect 2708 2500 2709 2540
rect 2667 2491 2709 2500
rect 2668 2489 2708 2491
rect 2667 2120 2709 2129
rect 2667 2080 2668 2120
rect 2708 2080 2709 2120
rect 2667 2071 2709 2080
rect 2668 1986 2708 2071
rect 2476 1903 2516 1912
rect 2764 1448 2804 2995
rect 2859 2792 2901 2801
rect 2859 2752 2860 2792
rect 2900 2752 2901 2792
rect 2859 2743 2901 2752
rect 2860 2658 2900 2743
rect 2859 2204 2901 2213
rect 2859 2164 2860 2204
rect 2900 2164 2901 2204
rect 2859 2155 2901 2164
rect 2860 2120 2900 2155
rect 2860 2069 2900 2080
rect 2668 1408 2804 1448
rect 2572 1121 2612 1206
rect 2571 1112 2613 1121
rect 2571 1072 2572 1112
rect 2612 1072 2613 1112
rect 2571 1063 2613 1072
rect 2668 944 2708 1408
rect 2764 1280 2804 1289
rect 2956 1280 2996 4843
rect 3052 3296 3092 5683
rect 3244 4901 3284 7120
rect 3339 7160 3381 7169
rect 3339 7120 3340 7160
rect 3380 7120 3381 7160
rect 3339 7111 3381 7120
rect 3627 7160 3669 7169
rect 3627 7120 3628 7160
rect 3668 7120 3669 7160
rect 3627 7111 3669 7120
rect 3340 7026 3380 7111
rect 3628 6833 3668 7111
rect 3627 6824 3669 6833
rect 3627 6784 3628 6824
rect 3668 6784 3669 6824
rect 3627 6775 3669 6784
rect 3435 6740 3477 6749
rect 3435 6700 3436 6740
rect 3476 6700 3477 6740
rect 3435 6691 3477 6700
rect 3243 4892 3285 4901
rect 3243 4852 3244 4892
rect 3284 4852 3285 4892
rect 3243 4843 3285 4852
rect 3436 4388 3476 6691
rect 3724 6656 3764 7204
rect 3532 6616 3764 6656
rect 3820 7244 3860 7363
rect 3532 6488 3572 6616
rect 3532 6439 3572 6448
rect 3628 6488 3668 6497
rect 3820 6488 3860 7204
rect 4011 7160 4053 7169
rect 4011 7120 4012 7160
rect 4052 7120 4053 7160
rect 4011 7111 4053 7120
rect 3668 6448 3860 6488
rect 4012 6488 4052 7111
rect 4204 6992 4244 7372
rect 4300 7169 4340 7254
rect 4299 7160 4341 7169
rect 4492 7160 4532 10312
rect 4780 10184 4820 10193
rect 4683 10100 4725 10109
rect 4683 10060 4684 10100
rect 4724 10060 4725 10100
rect 4683 10051 4725 10060
rect 4588 9260 4628 9269
rect 4588 8933 4628 9220
rect 4587 8924 4629 8933
rect 4587 8884 4588 8924
rect 4628 8884 4629 8924
rect 4587 8875 4629 8884
rect 4587 8756 4629 8765
rect 4587 8716 4588 8756
rect 4628 8716 4629 8756
rect 4587 8707 4629 8716
rect 4684 8756 4724 10051
rect 4780 10025 4820 10144
rect 5068 10025 5108 10732
rect 5163 10688 5205 10697
rect 5163 10648 5164 10688
rect 5204 10648 5205 10688
rect 5163 10639 5205 10648
rect 5164 10436 5204 10639
rect 5164 10387 5204 10396
rect 5260 10100 5300 10975
rect 5356 10268 5396 11320
rect 5548 11033 5588 11320
rect 5643 11192 5685 11201
rect 5643 11152 5644 11192
rect 5684 11152 5685 11192
rect 5643 11143 5685 11152
rect 5356 10219 5396 10228
rect 5452 11024 5492 11033
rect 5260 10060 5396 10100
rect 4779 10016 4821 10025
rect 4779 9976 4780 10016
rect 4820 9976 4821 10016
rect 4779 9967 4821 9976
rect 5067 10016 5109 10025
rect 5067 9976 5068 10016
rect 5108 9976 5109 10016
rect 5067 9967 5109 9976
rect 4780 9532 4820 9967
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4780 9492 4916 9532
rect 4684 8707 4724 8716
rect 4780 9428 4820 9437
rect 4588 8597 4628 8707
rect 4587 8588 4629 8597
rect 4587 8548 4588 8588
rect 4628 8548 4629 8588
rect 4587 8539 4629 8548
rect 4588 7757 4628 8539
rect 4780 8168 4820 9388
rect 4876 8765 4916 9492
rect 5164 9428 5204 9437
rect 4971 9260 5013 9269
rect 4971 9220 4972 9260
rect 5012 9220 5013 9260
rect 4971 9211 5013 9220
rect 4972 9126 5012 9211
rect 5164 8933 5204 9388
rect 5163 8924 5205 8933
rect 5163 8884 5164 8924
rect 5204 8884 5205 8924
rect 5163 8875 5205 8884
rect 4875 8756 4917 8765
rect 4875 8716 4876 8756
rect 4916 8716 4917 8756
rect 4875 8707 4917 8716
rect 5164 8672 5204 8681
rect 4876 8513 4916 8598
rect 4875 8504 4917 8513
rect 4875 8464 4876 8504
rect 4916 8464 4917 8504
rect 5164 8504 5204 8632
rect 5260 8672 5300 8681
rect 5356 8672 5396 10060
rect 5452 8849 5492 10984
rect 5547 11024 5589 11033
rect 5547 10984 5548 11024
rect 5588 10984 5589 11024
rect 5547 10975 5589 10984
rect 5644 10856 5684 11143
rect 5548 10816 5684 10856
rect 5451 8840 5493 8849
rect 5451 8800 5452 8840
rect 5492 8800 5493 8840
rect 5451 8791 5493 8800
rect 5300 8632 5492 8672
rect 5260 8623 5300 8632
rect 5164 8464 5396 8504
rect 4875 8455 4917 8464
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 5259 8168 5301 8177
rect 4780 8128 4916 8168
rect 4587 7748 4629 7757
rect 4587 7708 4588 7748
rect 4628 7708 4629 7748
rect 4587 7699 4629 7708
rect 4299 7120 4300 7160
rect 4340 7120 4532 7160
rect 4780 7165 4820 7174
rect 4299 7111 4341 7120
rect 4204 6952 4340 6992
rect 4108 6488 4148 6497
rect 4012 6448 4108 6488
rect 3628 6439 3668 6448
rect 4108 6439 4148 6448
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3819 5900 3861 5909
rect 3819 5860 3820 5900
rect 3860 5860 3861 5900
rect 3819 5851 3861 5860
rect 3820 5766 3860 5851
rect 4204 5816 4244 5825
rect 4012 5732 4052 5741
rect 3628 5648 3668 5657
rect 3628 5321 3668 5608
rect 3627 5312 3669 5321
rect 3627 5272 3628 5312
rect 3668 5272 3669 5312
rect 3627 5263 3669 5272
rect 4012 4733 4052 5692
rect 4204 5657 4244 5776
rect 4203 5648 4245 5657
rect 4203 5608 4204 5648
rect 4244 5608 4245 5648
rect 4203 5599 4245 5608
rect 4203 5144 4245 5153
rect 4203 5104 4204 5144
rect 4244 5104 4245 5144
rect 4203 5095 4245 5104
rect 4108 4976 4148 4985
rect 4011 4724 4053 4733
rect 4011 4684 4012 4724
rect 4052 4684 4053 4724
rect 4011 4675 4053 4684
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 3436 4348 3764 4388
rect 3147 4220 3189 4229
rect 3147 4180 3148 4220
rect 3188 4180 3189 4220
rect 3147 4171 3189 4180
rect 3148 4136 3188 4171
rect 3148 3725 3188 4096
rect 3147 3716 3189 3725
rect 3147 3676 3148 3716
rect 3188 3676 3189 3716
rect 3147 3667 3189 3676
rect 3531 3632 3573 3641
rect 3531 3592 3532 3632
rect 3572 3592 3573 3632
rect 3531 3583 3573 3592
rect 3724 3632 3764 4348
rect 4108 3893 4148 4936
rect 4204 4892 4244 5095
rect 4300 5060 4340 6952
rect 4780 6833 4820 7125
rect 4876 7076 4916 8128
rect 5259 8128 5260 8168
rect 5300 8128 5301 8168
rect 5259 8119 5301 8128
rect 5163 7496 5205 7505
rect 5163 7456 5164 7496
rect 5204 7456 5205 7496
rect 5163 7447 5205 7456
rect 5164 7160 5204 7447
rect 5260 7253 5300 8119
rect 5259 7244 5301 7253
rect 5259 7204 5260 7244
rect 5300 7204 5301 7244
rect 5259 7195 5301 7204
rect 5164 7111 5204 7120
rect 4972 7076 5012 7085
rect 4876 7036 4972 7076
rect 4972 7027 5012 7036
rect 4779 6824 4821 6833
rect 4779 6784 4780 6824
rect 4820 6784 4821 6824
rect 4779 6775 4821 6784
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5259 6656 5301 6665
rect 5259 6616 5260 6656
rect 5300 6616 5301 6656
rect 5259 6607 5301 6616
rect 4780 6572 4820 6581
rect 4684 6532 4780 6572
rect 4588 6474 4628 6483
rect 4396 5993 4436 5995
rect 4395 5984 4437 5993
rect 4395 5944 4396 5984
rect 4436 5944 4437 5984
rect 4395 5935 4437 5944
rect 4396 5900 4436 5935
rect 4588 5900 4628 6434
rect 4396 5851 4436 5860
rect 4492 5860 4628 5900
rect 4395 5144 4437 5153
rect 4395 5104 4396 5144
rect 4436 5104 4437 5144
rect 4395 5095 4437 5104
rect 4300 5011 4340 5020
rect 4204 4852 4340 4892
rect 4203 4724 4245 4733
rect 4203 4684 4204 4724
rect 4244 4684 4245 4724
rect 4203 4675 4245 4684
rect 4204 3977 4244 4675
rect 4203 3968 4245 3977
rect 4203 3928 4204 3968
rect 4244 3928 4245 3968
rect 4300 3968 4340 4852
rect 4396 4136 4436 5095
rect 4492 4976 4532 5860
rect 4588 5732 4628 5741
rect 4684 5732 4724 6532
rect 4780 6523 4820 6532
rect 5163 6572 5205 6581
rect 5163 6532 5164 6572
rect 5204 6532 5205 6572
rect 5163 6523 5205 6532
rect 5164 6404 5204 6523
rect 5260 6404 5300 6607
rect 5356 6572 5396 8464
rect 5452 8177 5492 8632
rect 5451 8168 5493 8177
rect 5451 8128 5452 8168
rect 5492 8128 5493 8168
rect 5451 8119 5493 8128
rect 5452 8000 5492 8009
rect 5452 7757 5492 7960
rect 5451 7748 5493 7757
rect 5451 7708 5452 7748
rect 5492 7708 5493 7748
rect 5451 7699 5493 7708
rect 5548 6581 5588 10816
rect 5643 10520 5685 10529
rect 5643 10480 5644 10520
rect 5684 10480 5685 10520
rect 5643 10471 5685 10480
rect 5644 10184 5684 10471
rect 5644 10135 5684 10144
rect 5643 9512 5685 9521
rect 5643 9472 5644 9512
rect 5684 9472 5685 9512
rect 5643 9463 5685 9472
rect 5644 9378 5684 9463
rect 5643 8756 5685 8765
rect 5643 8716 5644 8756
rect 5684 8716 5685 8756
rect 5643 8707 5685 8716
rect 5740 8756 5780 12823
rect 5836 12620 5876 16360
rect 6028 16325 6068 17695
rect 6124 16997 6164 18367
rect 6219 18332 6261 18341
rect 6219 18292 6220 18332
rect 6260 18292 6261 18332
rect 6219 18283 6261 18292
rect 6123 16988 6165 16997
rect 6123 16948 6124 16988
rect 6164 16948 6165 16988
rect 6123 16939 6165 16948
rect 6027 16316 6069 16325
rect 6124 16316 6164 16325
rect 6027 16276 6028 16316
rect 6068 16276 6124 16316
rect 6027 16267 6069 16276
rect 6124 16267 6164 16276
rect 6220 16316 6260 18283
rect 6315 17072 6357 17081
rect 6412 17072 6452 24004
rect 6507 23876 6549 23885
rect 6507 23836 6508 23876
rect 6548 23836 6549 23876
rect 6507 23827 6549 23836
rect 6508 23792 6548 23827
rect 6508 23741 6548 23752
rect 6700 22289 6740 25087
rect 6892 25002 6932 25087
rect 7083 24800 7125 24809
rect 7083 24760 7084 24800
rect 7124 24760 7125 24800
rect 7083 24751 7125 24760
rect 6795 24212 6837 24221
rect 6795 24172 6796 24212
rect 6836 24172 6837 24212
rect 6795 24163 6837 24172
rect 6796 23129 6836 24163
rect 6795 23120 6837 23129
rect 6795 23080 6796 23120
rect 6836 23080 6837 23120
rect 6795 23071 6837 23080
rect 6699 22280 6741 22289
rect 6699 22240 6700 22280
rect 6740 22240 6741 22280
rect 6699 22231 6741 22240
rect 6507 22112 6549 22121
rect 6507 22072 6508 22112
rect 6548 22072 6549 22112
rect 6507 22063 6549 22072
rect 6508 21978 6548 22063
rect 7084 21365 7124 24751
rect 7083 21356 7125 21365
rect 7083 21316 7084 21356
rect 7124 21316 7125 21356
rect 7083 21307 7125 21316
rect 6795 20768 6837 20777
rect 6795 20728 6796 20768
rect 6836 20728 6837 20768
rect 6795 20719 6837 20728
rect 6796 20634 6836 20719
rect 7180 20693 7220 26356
rect 7371 26228 7413 26237
rect 7371 26188 7372 26228
rect 7412 26188 7413 26228
rect 7371 26179 7413 26188
rect 7275 26144 7317 26153
rect 7275 26104 7276 26144
rect 7316 26104 7317 26144
rect 7275 26095 7317 26104
rect 7372 26144 7412 26179
rect 7276 20945 7316 26095
rect 7372 26093 7412 26104
rect 7468 26069 7508 26767
rect 7563 26648 7605 26657
rect 7563 26608 7564 26648
rect 7604 26608 7605 26648
rect 7563 26599 7605 26608
rect 7564 26312 7604 26599
rect 7660 26573 7700 29128
rect 7756 29093 7796 32152
rect 7852 29681 7892 32824
rect 7948 32908 8180 32948
rect 7851 29672 7893 29681
rect 7851 29632 7852 29672
rect 7892 29632 7893 29672
rect 7851 29623 7893 29632
rect 7852 29513 7892 29623
rect 7851 29504 7893 29513
rect 7851 29464 7852 29504
rect 7892 29464 7893 29504
rect 7851 29455 7893 29464
rect 7851 29168 7893 29177
rect 7851 29128 7852 29168
rect 7892 29128 7893 29168
rect 7851 29119 7893 29128
rect 7755 29084 7797 29093
rect 7755 29044 7756 29084
rect 7796 29044 7797 29084
rect 7755 29035 7797 29044
rect 7852 28664 7892 29119
rect 7948 28748 7988 32908
rect 8139 32780 8181 32789
rect 8139 32740 8140 32780
rect 8180 32740 8181 32780
rect 8139 32731 8181 32740
rect 8043 31688 8085 31697
rect 8043 31648 8044 31688
rect 8084 31648 8085 31688
rect 8043 31639 8085 31648
rect 8044 31436 8084 31639
rect 8044 31387 8084 31396
rect 8140 31352 8180 32731
rect 8140 31268 8180 31312
rect 8044 31228 8180 31268
rect 8044 29849 8084 31228
rect 8236 31184 8276 33151
rect 8140 31144 8276 31184
rect 8043 29840 8085 29849
rect 8043 29800 8044 29840
rect 8084 29800 8085 29840
rect 8043 29791 8085 29800
rect 8140 29000 8180 31144
rect 8235 30680 8277 30689
rect 8235 30640 8236 30680
rect 8276 30640 8277 30680
rect 8235 30631 8277 30640
rect 8236 30546 8276 30631
rect 8140 28960 8276 29000
rect 7948 28708 8180 28748
rect 7852 28624 7988 28664
rect 7755 28412 7797 28421
rect 7755 28372 7756 28412
rect 7796 28372 7797 28412
rect 7755 28363 7797 28372
rect 7756 28328 7796 28363
rect 7756 28277 7796 28288
rect 7851 28328 7893 28337
rect 7851 28288 7852 28328
rect 7892 28288 7893 28328
rect 7851 28279 7893 28288
rect 7948 28328 7988 28624
rect 7948 28279 7988 28288
rect 7852 28194 7892 28279
rect 8044 28160 8084 28169
rect 7755 27908 7797 27917
rect 7755 27868 7756 27908
rect 7796 27868 7797 27908
rect 7755 27859 7797 27868
rect 7756 26816 7796 27859
rect 8044 27665 8084 28120
rect 8043 27656 8085 27665
rect 8043 27616 8044 27656
rect 8084 27616 8085 27656
rect 8043 27607 8085 27616
rect 7659 26564 7701 26573
rect 7659 26524 7660 26564
rect 7700 26524 7701 26564
rect 7659 26515 7701 26524
rect 7564 26263 7604 26272
rect 7659 26144 7701 26153
rect 7659 26104 7660 26144
rect 7700 26104 7701 26144
rect 7659 26095 7701 26104
rect 7467 26060 7509 26069
rect 7467 26020 7468 26060
rect 7508 26020 7509 26060
rect 7467 26011 7509 26020
rect 7660 26010 7700 26095
rect 7563 25724 7605 25733
rect 7563 25684 7564 25724
rect 7604 25684 7605 25724
rect 7563 25675 7605 25684
rect 7371 24968 7413 24977
rect 7371 24928 7372 24968
rect 7412 24928 7413 24968
rect 7371 24919 7413 24928
rect 7372 24632 7412 24919
rect 7564 24884 7604 25675
rect 7372 23801 7412 24592
rect 7468 24844 7604 24884
rect 7468 24548 7508 24844
rect 7756 24809 7796 26776
rect 8043 26564 8085 26573
rect 8043 26524 8044 26564
rect 8084 26524 8085 26564
rect 8043 26515 8085 26524
rect 7851 26396 7893 26405
rect 7851 26356 7852 26396
rect 7892 26356 7893 26396
rect 7851 26347 7893 26356
rect 7852 26144 7892 26347
rect 7947 26228 7989 26237
rect 7947 26188 7948 26228
rect 7988 26188 7989 26228
rect 7947 26179 7989 26188
rect 7852 26069 7892 26104
rect 7851 26060 7893 26069
rect 7851 26020 7852 26060
rect 7892 26020 7893 26060
rect 7851 26011 7893 26020
rect 7755 24800 7797 24809
rect 7755 24760 7756 24800
rect 7796 24760 7797 24800
rect 7755 24751 7797 24760
rect 7564 24716 7604 24725
rect 7604 24676 7700 24716
rect 7564 24667 7604 24676
rect 7660 24548 7700 24676
rect 7852 24632 7892 24641
rect 7852 24548 7892 24592
rect 7948 24632 7988 26179
rect 7948 24583 7988 24592
rect 7468 24508 7604 24548
rect 7660 24508 7892 24548
rect 7371 23792 7413 23801
rect 7371 23752 7372 23792
rect 7412 23752 7413 23792
rect 7371 23743 7413 23752
rect 7372 23120 7412 23743
rect 7564 23549 7604 24508
rect 8044 23885 8084 26515
rect 7851 23876 7893 23885
rect 7851 23836 7852 23876
rect 7892 23836 7893 23876
rect 7851 23827 7893 23836
rect 8043 23876 8085 23885
rect 8043 23836 8044 23876
rect 8084 23836 8085 23876
rect 8043 23827 8085 23836
rect 7755 23792 7797 23801
rect 7755 23752 7756 23792
rect 7796 23752 7797 23792
rect 7755 23743 7797 23752
rect 7756 23658 7796 23743
rect 7563 23540 7605 23549
rect 7563 23500 7564 23540
rect 7604 23500 7605 23540
rect 7563 23491 7605 23500
rect 7564 23120 7604 23129
rect 7372 23080 7564 23120
rect 7372 22541 7412 23080
rect 7564 23071 7604 23080
rect 7756 22868 7796 22877
rect 7371 22532 7413 22541
rect 7371 22492 7372 22532
rect 7412 22492 7413 22532
rect 7371 22483 7413 22492
rect 7756 22280 7796 22828
rect 7852 22709 7892 23827
rect 7947 23708 7989 23717
rect 7947 23668 7948 23708
rect 7988 23668 7989 23708
rect 7947 23659 7989 23668
rect 7948 23574 7988 23659
rect 8043 23372 8085 23381
rect 8043 23332 8044 23372
rect 8084 23332 8085 23372
rect 8043 23323 8085 23332
rect 8044 23129 8084 23323
rect 8043 23120 8085 23129
rect 8043 23080 8044 23120
rect 8084 23080 8085 23120
rect 8043 23071 8085 23080
rect 7851 22700 7893 22709
rect 7851 22660 7852 22700
rect 7892 22660 7893 22700
rect 7851 22651 7893 22660
rect 7756 22231 7796 22240
rect 7852 22280 7892 22289
rect 7852 21953 7892 22240
rect 7659 21944 7701 21953
rect 7659 21904 7660 21944
rect 7700 21904 7701 21944
rect 7659 21895 7701 21904
rect 7851 21944 7893 21953
rect 7851 21904 7852 21944
rect 7892 21904 7893 21944
rect 7851 21895 7893 21904
rect 7275 20936 7317 20945
rect 7275 20896 7276 20936
rect 7316 20896 7317 20936
rect 7275 20887 7317 20896
rect 7276 20773 7316 20782
rect 7179 20684 7221 20693
rect 7179 20644 7180 20684
rect 7220 20644 7221 20684
rect 7179 20635 7221 20644
rect 7276 20516 7316 20733
rect 6796 20476 7316 20516
rect 7468 20600 7508 20609
rect 6796 20264 6836 20476
rect 6796 20215 6836 20224
rect 6604 20096 6644 20105
rect 6604 19769 6644 20056
rect 6987 20096 7029 20105
rect 6987 20056 6988 20096
rect 7028 20056 7029 20096
rect 6987 20047 7029 20056
rect 6988 19962 7028 20047
rect 6603 19760 6645 19769
rect 6603 19720 6604 19760
rect 6644 19720 6645 19760
rect 6603 19711 6645 19720
rect 6987 19340 7029 19349
rect 6987 19300 6988 19340
rect 7028 19300 7029 19340
rect 6987 19291 7029 19300
rect 6604 19256 6644 19265
rect 6604 18845 6644 19216
rect 6988 19256 7028 19291
rect 6988 19205 7028 19216
rect 6699 19172 6741 19181
rect 6699 19132 6700 19172
rect 6740 19132 6741 19172
rect 6699 19123 6741 19132
rect 6603 18836 6645 18845
rect 6603 18796 6604 18836
rect 6644 18796 6645 18836
rect 6603 18787 6645 18796
rect 6700 18752 6740 19123
rect 6796 19088 6836 19097
rect 6836 19048 7220 19088
rect 6796 19039 6836 19048
rect 7083 18920 7125 18929
rect 7083 18880 7084 18920
rect 7124 18880 7125 18920
rect 7083 18871 7125 18880
rect 6700 18712 6836 18752
rect 6700 18584 6740 18595
rect 6700 18509 6740 18544
rect 6699 18500 6741 18509
rect 6699 18460 6700 18500
rect 6740 18460 6741 18500
rect 6699 18451 6741 18460
rect 6700 17417 6740 18451
rect 6699 17408 6741 17417
rect 6699 17368 6700 17408
rect 6740 17368 6741 17408
rect 6699 17359 6741 17368
rect 6796 17156 6836 18712
rect 7084 17744 7124 18871
rect 7180 18579 7220 19048
rect 7372 18668 7412 18677
rect 7180 18530 7220 18539
rect 7276 18628 7372 18668
rect 7084 17695 7124 17704
rect 6988 17156 7028 17165
rect 6315 17032 6316 17072
rect 6356 17032 6452 17072
rect 6700 17116 6836 17156
rect 6892 17116 6988 17156
rect 6315 17023 6357 17032
rect 6316 16938 6356 17023
rect 6507 16820 6549 16829
rect 6507 16780 6508 16820
rect 6548 16780 6549 16820
rect 6507 16771 6549 16780
rect 6411 16400 6453 16409
rect 6411 16360 6412 16400
rect 6452 16360 6453 16400
rect 6411 16351 6453 16360
rect 6028 16182 6068 16267
rect 6220 15905 6260 16276
rect 6219 15896 6261 15905
rect 6219 15856 6220 15896
rect 6260 15856 6261 15896
rect 6219 15847 6261 15856
rect 6412 15317 6452 16351
rect 6411 15308 6453 15317
rect 6411 15268 6412 15308
rect 6452 15268 6453 15308
rect 6411 15259 6453 15268
rect 6027 14972 6069 14981
rect 6027 14932 6028 14972
rect 6068 14932 6069 14972
rect 6027 14923 6069 14932
rect 6028 14720 6068 14923
rect 6028 14671 6068 14680
rect 6315 14300 6357 14309
rect 6315 14260 6316 14300
rect 6356 14260 6357 14300
rect 6315 14251 6357 14260
rect 6220 14048 6260 14057
rect 5931 13376 5973 13385
rect 5931 13336 5932 13376
rect 5972 13336 5973 13376
rect 5931 13327 5973 13336
rect 5932 13292 5972 13327
rect 5932 13040 5972 13252
rect 6028 13208 6068 13217
rect 6068 13168 6164 13208
rect 6028 13159 6068 13168
rect 5932 13000 6068 13040
rect 5931 12620 5973 12629
rect 5836 12580 5932 12620
rect 5972 12580 5973 12620
rect 5931 12571 5973 12580
rect 5932 12536 5972 12571
rect 5932 12485 5972 12496
rect 5740 8707 5780 8716
rect 5836 11696 5876 11705
rect 5644 8622 5684 8707
rect 5644 8168 5684 8177
rect 5836 8168 5876 11656
rect 5931 11696 5973 11705
rect 5931 11656 5932 11696
rect 5972 11656 5973 11696
rect 5931 11647 5973 11656
rect 5932 11562 5972 11647
rect 5931 11276 5973 11285
rect 5931 11236 5932 11276
rect 5972 11236 5973 11276
rect 5931 11227 5973 11236
rect 5932 11024 5972 11227
rect 5932 9605 5972 10984
rect 6028 11024 6068 13000
rect 6124 12881 6164 13168
rect 6123 12872 6165 12881
rect 6123 12832 6124 12872
rect 6164 12832 6165 12872
rect 6123 12823 6165 12832
rect 6124 12620 6164 12629
rect 6220 12620 6260 14008
rect 6164 12580 6260 12620
rect 6316 14048 6356 14251
rect 6124 12571 6164 12580
rect 6316 11864 6356 14008
rect 6411 14048 6453 14057
rect 6411 14008 6412 14048
rect 6452 14008 6453 14048
rect 6411 13999 6453 14008
rect 6124 11824 6356 11864
rect 6124 11705 6164 11824
rect 6412 11780 6452 13999
rect 6508 13889 6548 16771
rect 6700 16661 6740 17116
rect 6796 17058 6836 17067
rect 6699 16652 6741 16661
rect 6699 16612 6700 16652
rect 6740 16612 6741 16652
rect 6699 16603 6741 16612
rect 6699 16400 6741 16409
rect 6699 16360 6700 16400
rect 6740 16360 6741 16400
rect 6699 16351 6741 16360
rect 6700 16232 6740 16351
rect 6700 16183 6740 16192
rect 6796 15728 6836 17018
rect 6796 15679 6836 15688
rect 6892 15644 6932 17116
rect 6988 17107 7028 17116
rect 7179 16820 7221 16829
rect 7179 16780 7180 16820
rect 7220 16780 7221 16820
rect 7179 16771 7221 16780
rect 7180 16686 7220 16771
rect 7276 16568 7316 18628
rect 7372 18619 7412 18628
rect 7371 17240 7413 17249
rect 7371 17200 7372 17240
rect 7412 17200 7413 17240
rect 7371 17191 7413 17200
rect 7372 17072 7412 17191
rect 7372 17023 7412 17032
rect 6879 15604 6932 15644
rect 7084 16528 7316 16568
rect 6603 15560 6645 15569
rect 6879 15560 6919 15604
rect 6603 15520 6604 15560
rect 6644 15520 6645 15560
rect 6603 15511 6645 15520
rect 6796 15520 6919 15560
rect 6604 15426 6644 15511
rect 6796 14384 6836 15520
rect 6988 15518 7028 15527
rect 6988 14897 7028 15478
rect 6987 14888 7029 14897
rect 6987 14848 6988 14888
rect 7028 14848 7029 14888
rect 6987 14839 7029 14848
rect 7084 14813 7124 16528
rect 7228 16241 7268 16250
rect 7268 16201 7316 16232
rect 7228 16192 7316 16201
rect 7179 15308 7221 15317
rect 7179 15268 7180 15308
rect 7220 15268 7221 15308
rect 7276 15308 7316 16192
rect 7371 16064 7413 16073
rect 7371 16024 7372 16064
rect 7412 16024 7413 16064
rect 7371 16015 7413 16024
rect 7372 15930 7412 16015
rect 7468 15485 7508 20560
rect 7563 20348 7605 20357
rect 7563 20308 7564 20348
rect 7604 20308 7605 20348
rect 7563 20299 7605 20308
rect 7564 20189 7604 20299
rect 7563 20180 7605 20189
rect 7563 20140 7564 20180
rect 7604 20140 7605 20180
rect 7563 20131 7605 20140
rect 7563 18248 7605 18257
rect 7563 18208 7564 18248
rect 7604 18208 7605 18248
rect 7563 18199 7605 18208
rect 7467 15476 7509 15485
rect 7467 15436 7468 15476
rect 7508 15436 7509 15476
rect 7467 15427 7509 15436
rect 7276 15268 7508 15308
rect 7179 15259 7221 15268
rect 7083 14804 7125 14813
rect 7083 14764 7084 14804
rect 7124 14764 7125 14804
rect 7083 14755 7125 14764
rect 6604 14344 6836 14384
rect 6987 14384 7029 14393
rect 6987 14344 6988 14384
rect 7028 14344 7029 14384
rect 6507 13880 6549 13889
rect 6507 13840 6508 13880
rect 6548 13840 6549 13880
rect 6507 13831 6549 13840
rect 6507 13712 6549 13721
rect 6507 13672 6508 13712
rect 6548 13672 6549 13712
rect 6507 13663 6549 13672
rect 6508 13208 6548 13663
rect 6508 13159 6548 13168
rect 6412 11731 6452 11740
rect 6123 11696 6165 11705
rect 6123 11656 6124 11696
rect 6164 11656 6165 11696
rect 6123 11647 6165 11656
rect 6315 11696 6357 11705
rect 6315 11656 6316 11696
rect 6356 11656 6357 11696
rect 6315 11647 6357 11656
rect 6028 10975 6068 10984
rect 6124 10109 6164 11647
rect 6316 11562 6356 11647
rect 6508 11024 6548 11033
rect 6508 10697 6548 10984
rect 6507 10688 6549 10697
rect 6507 10648 6508 10688
rect 6548 10648 6549 10688
rect 6507 10639 6549 10648
rect 6219 10520 6261 10529
rect 6219 10480 6220 10520
rect 6260 10480 6261 10520
rect 6219 10471 6261 10480
rect 6220 10193 6260 10471
rect 6508 10445 6548 10639
rect 6507 10436 6549 10445
rect 6507 10396 6508 10436
rect 6548 10396 6549 10436
rect 6507 10387 6549 10396
rect 6315 10352 6357 10361
rect 6315 10312 6316 10352
rect 6356 10312 6357 10352
rect 6315 10303 6357 10312
rect 6219 10184 6261 10193
rect 6219 10144 6220 10184
rect 6260 10144 6261 10184
rect 6219 10135 6261 10144
rect 6123 10100 6165 10109
rect 6123 10060 6124 10100
rect 6164 10060 6165 10100
rect 6123 10051 6165 10060
rect 6219 10016 6261 10025
rect 6219 9976 6220 10016
rect 6260 9976 6261 10016
rect 6219 9967 6261 9976
rect 5931 9596 5973 9605
rect 5931 9556 5932 9596
rect 5972 9556 5973 9596
rect 5931 9547 5973 9556
rect 5932 8765 5972 9547
rect 6123 9512 6165 9521
rect 6123 9472 6124 9512
rect 6164 9472 6165 9512
rect 6123 9463 6165 9472
rect 5931 8756 5973 8765
rect 5931 8716 5932 8756
rect 5972 8716 5973 8756
rect 5931 8707 5973 8716
rect 5931 8588 5973 8597
rect 5931 8548 5932 8588
rect 5972 8548 5973 8588
rect 5931 8539 5973 8548
rect 5684 8128 5876 8168
rect 5644 8119 5684 8128
rect 5739 8000 5781 8009
rect 5836 8000 5876 8009
rect 5739 7960 5740 8000
rect 5780 7960 5836 8000
rect 5739 7951 5781 7960
rect 5836 7951 5876 7960
rect 5740 6749 5780 7951
rect 5835 7412 5877 7421
rect 5835 7372 5836 7412
rect 5876 7372 5877 7412
rect 5835 7363 5877 7372
rect 5739 6740 5781 6749
rect 5739 6700 5740 6740
rect 5780 6700 5781 6740
rect 5739 6691 5781 6700
rect 5547 6572 5589 6581
rect 5356 6532 5492 6572
rect 5356 6404 5396 6413
rect 5260 6364 5356 6404
rect 5164 6355 5204 6364
rect 5356 6355 5396 6364
rect 4971 6320 5013 6329
rect 4971 6280 4972 6320
rect 5012 6280 5013 6320
rect 4971 6271 5013 6280
rect 4972 6186 5012 6271
rect 4628 5692 4724 5732
rect 4875 5732 4917 5741
rect 4875 5692 4876 5732
rect 4916 5692 4917 5732
rect 4588 5683 4628 5692
rect 4875 5683 4917 5692
rect 4876 5598 4916 5683
rect 5067 5648 5109 5657
rect 5067 5608 5068 5648
rect 5108 5608 5109 5648
rect 5067 5599 5109 5608
rect 5068 5514 5108 5599
rect 4779 5312 4821 5321
rect 4779 5272 4780 5312
rect 4820 5272 4821 5312
rect 4779 5263 4821 5272
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 4780 5144 4820 5263
rect 5452 5144 5492 6532
rect 5547 6532 5548 6572
rect 5588 6532 5589 6572
rect 5547 6523 5589 6532
rect 5739 6572 5781 6581
rect 5739 6532 5740 6572
rect 5780 6532 5781 6572
rect 5739 6523 5781 6532
rect 5548 6320 5588 6329
rect 5740 6320 5780 6523
rect 5588 6280 5780 6320
rect 5548 6271 5588 6280
rect 5547 6152 5589 6161
rect 5547 6112 5548 6152
rect 5588 6112 5589 6152
rect 5547 6103 5589 6112
rect 4780 5095 4820 5104
rect 5356 5104 5492 5144
rect 4492 4936 4724 4976
rect 4587 4808 4629 4817
rect 4587 4768 4588 4808
rect 4628 4768 4629 4808
rect 4587 4759 4629 4768
rect 4588 4674 4628 4759
rect 4587 4388 4629 4397
rect 4587 4348 4588 4388
rect 4628 4348 4629 4388
rect 4587 4339 4629 4348
rect 4588 4254 4628 4339
rect 4396 4087 4436 4096
rect 4491 3968 4533 3977
rect 4300 3928 4436 3968
rect 4203 3919 4245 3928
rect 4107 3884 4149 3893
rect 4107 3844 4108 3884
rect 4148 3844 4149 3884
rect 4107 3835 4149 3844
rect 3724 3583 3764 3592
rect 3532 3464 3572 3583
rect 4204 3557 4244 3559
rect 4203 3548 4245 3557
rect 4203 3508 4204 3548
rect 4244 3508 4245 3548
rect 4203 3499 4245 3508
rect 3532 3415 3572 3424
rect 4108 3464 4148 3473
rect 3052 3256 3188 3296
rect 3051 3128 3093 3137
rect 3051 3088 3052 3128
rect 3092 3088 3093 3128
rect 3051 3079 3093 3088
rect 3052 1868 3092 3079
rect 3148 2540 3188 3256
rect 3531 3044 3573 3053
rect 3531 3004 3532 3044
rect 3572 3004 3573 3044
rect 3531 2995 3573 3004
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 3435 2876 3477 2885
rect 3435 2836 3436 2876
rect 3476 2836 3477 2876
rect 3435 2827 3477 2836
rect 3436 2742 3476 2827
rect 3244 2708 3284 2717
rect 3284 2668 3380 2708
rect 3244 2659 3284 2668
rect 3243 2540 3285 2549
rect 3148 2500 3244 2540
rect 3284 2500 3285 2540
rect 3243 2491 3285 2500
rect 3243 2288 3285 2297
rect 3243 2248 3244 2288
rect 3284 2248 3285 2288
rect 3243 2239 3285 2248
rect 3052 1819 3092 1828
rect 3147 1868 3189 1877
rect 3147 1828 3148 1868
rect 3188 1828 3189 1868
rect 3147 1819 3189 1828
rect 2804 1240 2996 1280
rect 2764 1231 2804 1240
rect 3148 1196 3188 1819
rect 3148 1147 3188 1156
rect 2763 1112 2805 1121
rect 2763 1072 2764 1112
rect 2804 1072 2805 1112
rect 2763 1063 2805 1072
rect 2572 904 2708 944
rect 2572 80 2612 904
rect 2764 80 2804 1063
rect 3147 1028 3189 1037
rect 3147 988 3148 1028
rect 3188 988 3189 1028
rect 3147 979 3189 988
rect 2955 944 2997 953
rect 2955 904 2956 944
rect 2996 904 2997 944
rect 2955 895 2997 904
rect 2956 810 2996 895
rect 2955 608 2997 617
rect 2955 568 2956 608
rect 2996 568 2997 608
rect 2955 559 2997 568
rect 2956 80 2996 559
rect 3148 80 3188 979
rect 3244 944 3284 2239
rect 3340 2129 3380 2668
rect 3532 2624 3572 2995
rect 4108 2960 4148 3424
rect 4204 3464 4244 3499
rect 4204 3415 4244 3424
rect 4396 3221 4436 3928
rect 4491 3928 4492 3968
rect 4532 3928 4533 3968
rect 4491 3919 4533 3928
rect 4395 3212 4437 3221
rect 4395 3172 4396 3212
rect 4436 3172 4437 3212
rect 4395 3163 4437 3172
rect 4203 2960 4245 2969
rect 4108 2920 4204 2960
rect 4244 2920 4245 2960
rect 4203 2911 4245 2920
rect 3627 2792 3669 2801
rect 3627 2752 3628 2792
rect 3668 2752 3669 2792
rect 3627 2743 3669 2752
rect 4011 2792 4053 2801
rect 4011 2752 4012 2792
rect 4052 2752 4053 2792
rect 4011 2743 4053 2752
rect 3436 2584 3572 2624
rect 3628 2666 3668 2743
rect 3628 2617 3668 2626
rect 3339 2120 3381 2129
rect 3339 2080 3340 2120
rect 3380 2080 3381 2120
rect 3339 2071 3381 2080
rect 3339 1952 3381 1961
rect 3339 1912 3340 1952
rect 3380 1912 3381 1952
rect 3339 1903 3381 1912
rect 3436 1952 3476 2584
rect 3531 2204 3573 2213
rect 3531 2164 3532 2204
rect 3572 2164 3573 2204
rect 3531 2155 3573 2164
rect 3436 1903 3476 1912
rect 3340 1818 3380 1903
rect 3532 1112 3572 2155
rect 3916 1952 3956 1961
rect 4012 1952 4052 2743
rect 4395 2372 4437 2381
rect 4395 2332 4396 2372
rect 4436 2332 4437 2372
rect 4395 2323 4437 2332
rect 3956 1912 4052 1952
rect 4396 1952 4436 2323
rect 3916 1903 3956 1912
rect 4396 1903 4436 1912
rect 3820 1868 3860 1877
rect 3820 1700 3860 1828
rect 4299 1784 4341 1793
rect 4299 1744 4300 1784
rect 4340 1744 4341 1784
rect 4299 1735 4341 1744
rect 3820 1660 4148 1700
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 3723 1280 3765 1289
rect 3723 1240 3724 1280
rect 3764 1240 3765 1280
rect 3723 1231 3765 1240
rect 3532 1063 3572 1072
rect 3244 904 3572 944
rect 3339 524 3381 533
rect 3339 484 3340 524
rect 3380 484 3381 524
rect 3339 475 3381 484
rect 3340 80 3380 475
rect 3532 80 3572 904
rect 3724 80 3764 1231
rect 3915 692 3957 701
rect 3915 652 3916 692
rect 3956 652 3957 692
rect 3915 643 3957 652
rect 3916 80 3956 643
rect 4108 80 4148 1660
rect 4300 80 4340 1735
rect 4492 1037 4532 3919
rect 4684 3548 4724 4936
rect 4924 4934 4964 4943
rect 4924 4892 4964 4894
rect 4780 4852 4964 4892
rect 4780 3632 4820 4852
rect 4971 4556 5013 4565
rect 4971 4516 4972 4556
rect 5012 4516 5013 4556
rect 4971 4507 5013 4516
rect 4972 4220 5012 4507
rect 5356 4397 5396 5104
rect 5451 4976 5493 4985
rect 5451 4936 5452 4976
rect 5492 4936 5493 4976
rect 5451 4927 5493 4936
rect 5452 4842 5492 4927
rect 5355 4388 5397 4397
rect 5355 4348 5356 4388
rect 5396 4348 5397 4388
rect 5355 4339 5397 4348
rect 4972 4171 5012 4180
rect 5356 4136 5396 4145
rect 5548 4136 5588 6103
rect 5643 5648 5685 5657
rect 5643 5608 5644 5648
rect 5684 5608 5685 5648
rect 5643 5599 5685 5608
rect 5396 4096 5588 4136
rect 5356 4087 5396 4096
rect 5164 3977 5204 4062
rect 5163 3968 5205 3977
rect 5163 3928 5164 3968
rect 5204 3928 5205 3968
rect 5163 3919 5205 3928
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 5451 3632 5493 3641
rect 4780 3592 5108 3632
rect 4684 3508 4820 3548
rect 4588 3380 4628 3389
rect 4588 2960 4628 3340
rect 4684 3380 4724 3389
rect 4684 3221 4724 3340
rect 4683 3212 4725 3221
rect 4683 3172 4684 3212
rect 4724 3172 4725 3212
rect 4683 3163 4725 3172
rect 4588 2920 4724 2960
rect 4684 1793 4724 2920
rect 4780 2120 4820 3508
rect 5068 2876 5108 3592
rect 5451 3592 5452 3632
rect 5492 3592 5493 3632
rect 5451 3583 5493 3592
rect 5164 3464 5204 3473
rect 5164 3305 5204 3424
rect 5259 3464 5301 3473
rect 5259 3424 5260 3464
rect 5300 3424 5301 3464
rect 5259 3415 5301 3424
rect 5163 3296 5205 3305
rect 5163 3256 5164 3296
rect 5204 3256 5205 3296
rect 5163 3247 5205 3256
rect 5068 2827 5108 2836
rect 4875 2624 4917 2633
rect 4875 2584 4876 2624
rect 4916 2584 4917 2624
rect 4875 2575 4917 2584
rect 5260 2624 5300 3415
rect 5355 3296 5397 3305
rect 5355 3256 5356 3296
rect 5396 3256 5397 3296
rect 5355 3247 5397 3256
rect 5260 2575 5300 2584
rect 4876 2490 4916 2575
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5068 2120 5108 2129
rect 5356 2120 5396 3247
rect 4780 2080 5012 2120
rect 4876 1938 4916 1947
rect 4683 1784 4725 1793
rect 4683 1744 4684 1784
rect 4724 1744 4725 1784
rect 4683 1735 4725 1744
rect 4876 1625 4916 1898
rect 4875 1616 4917 1625
rect 4875 1576 4876 1616
rect 4916 1576 4917 1616
rect 4875 1567 4917 1576
rect 4683 1532 4725 1541
rect 4683 1492 4684 1532
rect 4724 1492 4725 1532
rect 4683 1483 4725 1492
rect 4684 1373 4724 1483
rect 4683 1364 4725 1373
rect 4683 1324 4684 1364
rect 4724 1324 4725 1364
rect 4683 1315 4725 1324
rect 4875 1364 4917 1373
rect 4875 1324 4876 1364
rect 4916 1324 4917 1364
rect 4875 1315 4917 1324
rect 4684 1112 4724 1315
rect 4780 1112 4820 1121
rect 4684 1072 4780 1112
rect 4780 1063 4820 1072
rect 4491 1028 4533 1037
rect 4491 988 4492 1028
rect 4532 988 4533 1028
rect 4491 979 4533 988
rect 4683 944 4725 953
rect 4876 944 4916 1315
rect 4972 1280 5012 2080
rect 5108 2080 5396 2120
rect 5068 2071 5108 2080
rect 5259 1952 5301 1961
rect 5259 1912 5260 1952
rect 5300 1912 5301 1952
rect 5259 1903 5301 1912
rect 5260 1818 5300 1903
rect 4972 1231 5012 1240
rect 5259 1280 5301 1289
rect 5259 1240 5260 1280
rect 5300 1240 5301 1280
rect 5259 1231 5301 1240
rect 5260 1112 5300 1231
rect 5260 1063 5300 1072
rect 4683 904 4684 944
rect 4724 904 4725 944
rect 4683 895 4725 904
rect 4780 904 4916 944
rect 4491 860 4533 869
rect 4491 820 4492 860
rect 4532 820 4533 860
rect 4491 811 4533 820
rect 4492 80 4532 811
rect 4684 80 4724 895
rect 4780 608 4820 904
rect 5355 860 5397 869
rect 5355 820 5356 860
rect 5396 820 5397 860
rect 5355 811 5397 820
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 5067 608 5109 617
rect 4780 568 4916 608
rect 4876 80 4916 568
rect 5067 568 5068 608
rect 5108 568 5109 608
rect 5067 559 5109 568
rect 5068 80 5108 559
rect 5356 440 5396 811
rect 5260 400 5396 440
rect 5260 80 5300 400
rect 5452 80 5492 3583
rect 5644 3548 5684 5599
rect 5739 5564 5781 5573
rect 5739 5524 5740 5564
rect 5780 5524 5781 5564
rect 5739 5515 5781 5524
rect 5548 3508 5684 3548
rect 5548 3389 5588 3508
rect 5644 3450 5684 3459
rect 5547 3380 5589 3389
rect 5547 3340 5548 3380
rect 5588 3340 5589 3380
rect 5547 3331 5589 3340
rect 5644 2960 5684 3410
rect 5548 2920 5684 2960
rect 5548 953 5588 2920
rect 5740 2540 5780 5515
rect 5836 3632 5876 7363
rect 5932 5573 5972 8539
rect 6124 8093 6164 9463
rect 6220 9101 6260 9967
rect 6219 9092 6261 9101
rect 6219 9052 6220 9092
rect 6260 9052 6261 9092
rect 6219 9043 6261 9052
rect 6219 8840 6261 8849
rect 6219 8800 6220 8840
rect 6260 8800 6261 8840
rect 6219 8791 6261 8800
rect 6220 8672 6260 8791
rect 6123 8084 6165 8093
rect 6123 8044 6124 8084
rect 6164 8044 6165 8084
rect 6123 8035 6165 8044
rect 6027 7580 6069 7589
rect 6027 7540 6028 7580
rect 6068 7540 6069 7580
rect 6027 7531 6069 7540
rect 6028 6488 6068 7531
rect 6220 7421 6260 8632
rect 6219 7412 6261 7421
rect 6219 7372 6220 7412
rect 6260 7372 6261 7412
rect 6219 7363 6261 7372
rect 6316 7001 6356 10303
rect 6411 10016 6453 10025
rect 6411 9976 6412 10016
rect 6452 9976 6453 10016
rect 6411 9967 6453 9976
rect 6412 8177 6452 9967
rect 6411 8168 6453 8177
rect 6411 8128 6412 8168
rect 6452 8128 6453 8168
rect 6411 8119 6453 8128
rect 6604 7757 6644 14344
rect 6987 14335 7029 14344
rect 6699 14216 6741 14225
rect 6699 14176 6700 14216
rect 6740 14176 6741 14216
rect 6699 14167 6741 14176
rect 6700 14048 6740 14167
rect 6700 13385 6740 14008
rect 6795 14048 6837 14057
rect 6988 14048 7028 14335
rect 6795 14008 6796 14048
rect 6836 14008 7028 14048
rect 7180 14048 7220 15259
rect 7468 14972 7508 15268
rect 7468 14923 7508 14932
rect 7371 14804 7413 14813
rect 7371 14764 7372 14804
rect 7412 14764 7413 14804
rect 7371 14755 7413 14764
rect 7275 14720 7317 14729
rect 7275 14680 7276 14720
rect 7316 14680 7317 14720
rect 7275 14671 7317 14680
rect 7276 14586 7316 14671
rect 7276 14048 7316 14057
rect 7180 14008 7276 14048
rect 6795 13999 6837 14008
rect 7276 13999 7316 14008
rect 6796 13914 6836 13999
rect 7372 13889 7412 14755
rect 7371 13880 7413 13889
rect 7371 13840 7372 13880
rect 7412 13840 7413 13880
rect 7371 13831 7413 13840
rect 6795 13796 6837 13805
rect 6795 13756 6796 13796
rect 6836 13756 6837 13796
rect 6795 13747 6837 13756
rect 6699 13376 6741 13385
rect 6699 13336 6700 13376
rect 6740 13336 6741 13376
rect 6699 13327 6741 13336
rect 6796 12536 6836 13747
rect 7036 13217 7076 13226
rect 7467 13208 7509 13217
rect 7076 13177 7124 13208
rect 7036 13168 7124 13177
rect 6796 9185 6836 12496
rect 6891 11864 6933 11873
rect 6891 11824 6892 11864
rect 6932 11824 6933 11864
rect 6891 11815 6933 11824
rect 6892 11696 6932 11815
rect 6892 11647 6932 11656
rect 6891 11444 6933 11453
rect 6891 11404 6892 11444
rect 6932 11404 6933 11444
rect 6891 11395 6933 11404
rect 6892 10184 6932 11395
rect 6892 10135 6932 10144
rect 6988 11010 7028 11019
rect 6892 9521 6932 9606
rect 6891 9512 6933 9521
rect 6891 9472 6892 9512
rect 6932 9472 6933 9512
rect 6891 9463 6933 9472
rect 6891 9344 6933 9353
rect 6891 9304 6892 9344
rect 6932 9304 6933 9344
rect 6891 9295 6933 9304
rect 6795 9176 6837 9185
rect 6795 9136 6796 9176
rect 6836 9136 6837 9176
rect 6795 9127 6837 9136
rect 6892 9008 6932 9295
rect 6796 8968 6932 9008
rect 6700 8677 6740 8686
rect 6603 7748 6645 7757
rect 6603 7708 6604 7748
rect 6644 7708 6645 7748
rect 6603 7699 6645 7708
rect 6700 7580 6740 8637
rect 6796 7589 6836 8968
rect 6892 8504 6932 8513
rect 6892 7925 6932 8464
rect 6988 8177 7028 10970
rect 7084 10436 7124 13168
rect 7467 13168 7468 13208
rect 7508 13168 7509 13208
rect 7467 13159 7509 13168
rect 7179 13124 7221 13133
rect 7179 13084 7180 13124
rect 7220 13084 7221 13124
rect 7179 13075 7221 13084
rect 7180 12990 7220 13075
rect 7468 13074 7508 13159
rect 7275 12956 7317 12965
rect 7275 12916 7276 12956
rect 7316 12916 7317 12956
rect 7564 12956 7604 18199
rect 7660 16241 7700 21895
rect 7851 21608 7893 21617
rect 7756 21568 7852 21608
rect 7892 21568 7893 21608
rect 7756 18257 7796 21568
rect 7851 21559 7893 21568
rect 7852 21474 7892 21559
rect 7851 20096 7893 20105
rect 7851 20056 7852 20096
rect 7892 20056 7893 20096
rect 7851 20047 7893 20056
rect 7755 18248 7797 18257
rect 7755 18208 7756 18248
rect 7796 18208 7797 18248
rect 7755 18199 7797 18208
rect 7755 18080 7797 18089
rect 7755 18040 7756 18080
rect 7796 18040 7797 18080
rect 7755 18031 7797 18040
rect 7659 16232 7701 16241
rect 7659 16192 7660 16232
rect 7700 16192 7701 16232
rect 7659 16183 7701 16192
rect 7756 14132 7796 18031
rect 7852 16913 7892 20047
rect 7851 16904 7893 16913
rect 7851 16864 7852 16904
rect 7892 16864 7893 16904
rect 7851 16855 7893 16864
rect 7947 15224 7989 15233
rect 7947 15184 7948 15224
rect 7988 15184 7989 15224
rect 7947 15175 7989 15184
rect 7948 14216 7988 15175
rect 8044 14225 8084 23071
rect 8140 20180 8180 28708
rect 8236 25733 8276 28960
rect 8332 26237 8372 33664
rect 8428 33653 8468 33664
rect 8524 33704 8564 33713
rect 8716 33704 8756 33739
rect 8564 33664 8660 33704
rect 8524 33655 8564 33664
rect 8524 33536 8564 33545
rect 8427 33200 8469 33209
rect 8427 33160 8428 33200
rect 8468 33160 8469 33200
rect 8427 33151 8469 33160
rect 8428 32369 8468 33151
rect 8427 32360 8469 32369
rect 8427 32320 8428 32360
rect 8468 32320 8469 32360
rect 8427 32311 8469 32320
rect 8524 32201 8564 33496
rect 8620 33209 8660 33664
rect 8619 33200 8661 33209
rect 8619 33160 8620 33200
rect 8660 33160 8661 33200
rect 8619 33151 8661 33160
rect 8619 33032 8661 33041
rect 8619 32992 8620 33032
rect 8660 32992 8661 33032
rect 8619 32983 8661 32992
rect 8523 32192 8565 32201
rect 8523 32152 8524 32192
rect 8564 32152 8565 32192
rect 8523 32143 8565 32152
rect 8620 31520 8660 32983
rect 8716 32789 8756 33664
rect 8812 33704 8852 33713
rect 8812 33545 8852 33664
rect 8811 33536 8853 33545
rect 8811 33496 8812 33536
rect 8852 33496 8853 33536
rect 8811 33487 8853 33496
rect 8811 33368 8853 33377
rect 8811 33328 8812 33368
rect 8852 33328 8853 33368
rect 8811 33319 8853 33328
rect 8715 32780 8757 32789
rect 8715 32740 8716 32780
rect 8756 32740 8757 32780
rect 8715 32731 8757 32740
rect 8428 31480 8660 31520
rect 8331 26228 8373 26237
rect 8331 26188 8332 26228
rect 8372 26188 8373 26228
rect 8331 26179 8373 26188
rect 8235 25724 8277 25733
rect 8235 25684 8236 25724
rect 8276 25684 8277 25724
rect 8235 25675 8277 25684
rect 8428 25472 8468 31480
rect 8619 31352 8661 31361
rect 8619 31312 8620 31352
rect 8660 31312 8661 31352
rect 8619 31303 8661 31312
rect 8620 31218 8660 31303
rect 8523 30680 8565 30689
rect 8523 30640 8524 30680
rect 8564 30640 8565 30680
rect 8523 30631 8565 30640
rect 8524 27581 8564 30631
rect 8812 30437 8852 33319
rect 9004 32864 9044 32873
rect 9004 32621 9044 32824
rect 9003 32612 9045 32621
rect 9003 32572 9004 32612
rect 9044 32572 9045 32612
rect 9003 32563 9045 32572
rect 8908 32192 8948 32201
rect 9004 32192 9044 32563
rect 9100 32537 9140 33832
rect 9196 33704 9236 35671
rect 9292 34460 9332 35923
rect 9388 34544 9428 36688
rect 9675 36560 9717 36569
rect 9675 36520 9676 36560
rect 9716 36520 9717 36560
rect 9675 36511 9717 36520
rect 9483 36308 9525 36317
rect 9483 36268 9484 36308
rect 9524 36268 9525 36308
rect 9483 36259 9525 36268
rect 9484 35888 9524 36259
rect 9579 35972 9621 35981
rect 9579 35932 9580 35972
rect 9620 35932 9621 35972
rect 9579 35923 9621 35932
rect 9484 35839 9524 35848
rect 9580 35888 9620 35923
rect 9580 35837 9620 35848
rect 9676 35720 9716 36511
rect 9580 35680 9716 35720
rect 9388 34504 9524 34544
rect 9292 34420 9428 34460
rect 9388 34376 9428 34420
rect 9292 34356 9332 34365
rect 9292 34049 9332 34316
rect 9291 34040 9333 34049
rect 9291 34000 9292 34040
rect 9332 34000 9333 34040
rect 9291 33991 9333 34000
rect 9236 33664 9332 33704
rect 9196 33655 9236 33664
rect 9196 33041 9236 33126
rect 9292 33116 9332 33664
rect 9388 33377 9428 34336
rect 9387 33368 9429 33377
rect 9387 33328 9388 33368
rect 9428 33328 9429 33368
rect 9387 33319 9429 33328
rect 9387 33200 9429 33209
rect 9387 33160 9388 33200
rect 9428 33160 9429 33200
rect 9387 33151 9429 33160
rect 9292 33076 9337 33116
rect 9195 33032 9237 33041
rect 9297 33032 9337 33076
rect 9195 32992 9196 33032
rect 9236 32992 9237 33032
rect 9195 32983 9237 32992
rect 9292 32992 9337 33032
rect 9292 32864 9332 32992
rect 9388 32873 9428 33151
rect 9196 32824 9332 32864
rect 9099 32528 9141 32537
rect 9099 32488 9100 32528
rect 9140 32488 9141 32528
rect 9099 32479 9141 32488
rect 9099 32360 9141 32369
rect 9099 32320 9100 32360
rect 9140 32320 9141 32360
rect 9099 32311 9141 32320
rect 9100 32226 9140 32311
rect 8948 32152 9044 32192
rect 8908 31949 8948 32152
rect 8907 31940 8949 31949
rect 8907 31900 8908 31940
rect 8948 31900 8949 31940
rect 8907 31891 8949 31900
rect 9100 31357 9140 31366
rect 8907 30680 8949 30689
rect 8907 30640 8908 30680
rect 8948 30640 8949 30680
rect 8907 30631 8949 30640
rect 8811 30428 8853 30437
rect 8811 30388 8812 30428
rect 8852 30388 8853 30428
rect 8811 30379 8853 30388
rect 8811 30260 8853 30269
rect 8811 30220 8812 30260
rect 8852 30220 8853 30260
rect 8811 30211 8853 30220
rect 8812 29840 8852 30211
rect 8812 29336 8852 29800
rect 8716 29296 8852 29336
rect 8716 27665 8756 29296
rect 8812 29168 8852 29177
rect 8908 29168 8948 30631
rect 9004 30092 9044 30101
rect 9100 30092 9140 31317
rect 9196 30269 9236 32824
rect 9292 32705 9332 32824
rect 9387 32864 9429 32873
rect 9387 32824 9388 32864
rect 9428 32824 9429 32864
rect 9387 32815 9429 32824
rect 9388 32730 9428 32815
rect 9291 32696 9333 32705
rect 9291 32656 9292 32696
rect 9332 32656 9333 32696
rect 9291 32647 9333 32656
rect 9387 32528 9429 32537
rect 9387 32488 9388 32528
rect 9428 32488 9429 32528
rect 9387 32479 9429 32488
rect 9292 32201 9332 32286
rect 9291 32192 9333 32201
rect 9291 32152 9292 32192
rect 9332 32152 9333 32192
rect 9291 32143 9333 32152
rect 9388 32192 9428 32479
rect 9484 32360 9524 34504
rect 9580 33041 9620 35680
rect 9675 35300 9717 35309
rect 9675 35260 9676 35300
rect 9716 35260 9717 35300
rect 9675 35251 9717 35260
rect 9676 35216 9716 35251
rect 9676 35165 9716 35176
rect 9772 34544 9812 36688
rect 9868 36723 9908 37192
rect 10060 36896 10100 39376
rect 10251 39248 10293 39257
rect 10251 39208 10252 39248
rect 10292 39208 10293 39248
rect 10251 39199 10293 39208
rect 10060 36847 10100 36856
rect 9868 36674 9908 36683
rect 9867 36140 9909 36149
rect 9867 36100 9868 36140
rect 9908 36100 9909 36140
rect 9867 36091 9909 36100
rect 9868 35981 9908 36091
rect 9867 35972 9909 35981
rect 9867 35932 9868 35972
rect 9908 35932 9909 35972
rect 9867 35923 9909 35932
rect 9676 34504 9812 34544
rect 9964 35888 10004 35897
rect 9579 33032 9621 33041
rect 9579 32992 9580 33032
rect 9620 32992 9621 33032
rect 9579 32983 9621 32992
rect 9676 32621 9716 34504
rect 9964 34385 10004 35848
rect 10060 35888 10100 35897
rect 9771 34376 9813 34385
rect 9771 34336 9772 34376
rect 9812 34336 9813 34376
rect 9771 34327 9813 34336
rect 9868 34376 9908 34385
rect 9772 34242 9812 34327
rect 9771 33368 9813 33377
rect 9771 33328 9772 33368
rect 9812 33328 9813 33368
rect 9771 33319 9813 33328
rect 9772 32948 9812 33319
rect 9868 33125 9908 34336
rect 9963 34376 10005 34385
rect 9963 34336 9964 34376
rect 10004 34336 10005 34376
rect 9963 34327 10005 34336
rect 9867 33116 9909 33125
rect 9867 33076 9868 33116
rect 9908 33076 9909 33116
rect 9867 33067 9909 33076
rect 9772 32908 9908 32948
rect 9771 32780 9813 32789
rect 9771 32740 9772 32780
rect 9812 32740 9813 32780
rect 9771 32731 9813 32740
rect 9675 32612 9717 32621
rect 9675 32572 9676 32612
rect 9716 32572 9717 32612
rect 9675 32563 9717 32572
rect 9484 32311 9524 32320
rect 9579 32360 9621 32369
rect 9579 32320 9580 32360
rect 9620 32320 9621 32360
rect 9579 32311 9621 32320
rect 9388 32143 9428 32152
rect 9580 32192 9620 32311
rect 9772 32201 9812 32731
rect 9580 32143 9620 32152
rect 9675 32192 9717 32201
rect 9675 32152 9676 32192
rect 9716 32152 9717 32192
rect 9772 32192 9817 32201
rect 9772 32152 9777 32192
rect 9675 32143 9717 32152
rect 9777 32143 9817 32152
rect 9676 32058 9716 32143
rect 9292 31940 9332 31949
rect 9868 31940 9908 32908
rect 9292 31361 9332 31900
rect 9676 31900 9908 31940
rect 9676 31520 9716 31900
rect 9388 31480 9716 31520
rect 9291 31352 9333 31361
rect 9291 31312 9292 31352
rect 9332 31312 9333 31352
rect 9291 31303 9333 31312
rect 9291 31184 9333 31193
rect 9291 31144 9292 31184
rect 9332 31144 9333 31184
rect 9291 31135 9333 31144
rect 9292 31050 9332 31135
rect 9195 30260 9237 30269
rect 9195 30220 9196 30260
rect 9236 30220 9237 30260
rect 9195 30211 9237 30220
rect 9044 30052 9140 30092
rect 9004 30043 9044 30052
rect 9003 29336 9045 29345
rect 9003 29296 9004 29336
rect 9044 29296 9045 29336
rect 9003 29287 9045 29296
rect 9291 29336 9333 29345
rect 9291 29296 9292 29336
rect 9332 29296 9333 29336
rect 9291 29287 9333 29296
rect 9004 29202 9044 29287
rect 8852 29128 8948 29168
rect 9292 29168 9332 29287
rect 9388 29177 9428 31480
rect 9580 31352 9620 31361
rect 9580 30848 9620 31312
rect 9676 31352 9716 31480
rect 9676 31303 9716 31312
rect 9964 31436 10004 34327
rect 10060 32789 10100 35848
rect 10155 33116 10197 33125
rect 10155 33076 10156 33116
rect 10196 33076 10197 33116
rect 10155 33067 10197 33076
rect 10059 32780 10101 32789
rect 10059 32740 10060 32780
rect 10100 32740 10101 32780
rect 10059 32731 10101 32740
rect 10156 32360 10196 33067
rect 10060 32320 10196 32360
rect 10060 32192 10100 32320
rect 10060 31781 10100 32152
rect 10155 32192 10197 32201
rect 10155 32152 10156 32192
rect 10196 32152 10197 32192
rect 10155 32143 10197 32152
rect 10156 32058 10196 32143
rect 10059 31772 10101 31781
rect 10059 31732 10060 31772
rect 10100 31732 10101 31772
rect 10059 31723 10101 31732
rect 10155 31688 10197 31697
rect 10155 31648 10156 31688
rect 10196 31648 10197 31688
rect 10155 31639 10197 31648
rect 10060 31436 10100 31445
rect 9964 31396 10060 31436
rect 9676 30848 9716 30857
rect 9580 30808 9676 30848
rect 9676 30799 9716 30808
rect 9484 30689 9524 30774
rect 9867 30764 9909 30773
rect 9867 30724 9868 30764
rect 9908 30724 9909 30764
rect 9867 30715 9909 30724
rect 9483 30680 9525 30689
rect 9483 30640 9484 30680
rect 9524 30640 9525 30680
rect 9483 30631 9525 30640
rect 9868 30680 9908 30715
rect 9868 30629 9908 30640
rect 9483 30428 9525 30437
rect 9483 30388 9484 30428
rect 9524 30388 9620 30428
rect 9483 30379 9525 30388
rect 9483 30260 9525 30269
rect 9483 30220 9484 30260
rect 9524 30220 9525 30260
rect 9483 30211 9525 30220
rect 8812 29119 8852 29128
rect 9292 29119 9332 29128
rect 9387 29168 9429 29177
rect 9387 29128 9388 29168
rect 9428 29128 9429 29168
rect 9387 29119 9429 29128
rect 9388 29034 9428 29119
rect 9291 29000 9333 29009
rect 9291 28960 9292 29000
rect 9332 28960 9333 29000
rect 9291 28951 9333 28960
rect 8811 28244 8853 28253
rect 8811 28204 8812 28244
rect 8852 28204 8853 28244
rect 8811 28195 8853 28204
rect 8715 27656 8757 27665
rect 8715 27616 8716 27656
rect 8756 27616 8757 27656
rect 8715 27607 8757 27616
rect 8523 27572 8565 27581
rect 8523 27532 8524 27572
rect 8564 27532 8565 27572
rect 8523 27523 8565 27532
rect 8524 26993 8564 27523
rect 8716 27522 8756 27607
rect 8523 26984 8565 26993
rect 8523 26944 8524 26984
rect 8564 26944 8565 26984
rect 8812 26984 8852 28195
rect 8908 27740 8948 27749
rect 8948 27700 9236 27740
rect 8908 27691 8948 27700
rect 9196 27656 9236 27700
rect 9196 27607 9236 27616
rect 9292 27656 9332 28951
rect 8812 26944 8948 26984
rect 8523 26935 8565 26944
rect 8524 26816 8564 26825
rect 8524 26573 8564 26776
rect 8716 26816 8756 26825
rect 8619 26648 8661 26657
rect 8619 26608 8620 26648
rect 8660 26608 8661 26648
rect 8619 26599 8661 26608
rect 8523 26564 8565 26573
rect 8523 26524 8524 26564
rect 8564 26524 8565 26564
rect 8523 26515 8565 26524
rect 8620 26514 8660 26599
rect 8619 26228 8661 26237
rect 8619 26188 8620 26228
rect 8660 26188 8661 26228
rect 8619 26179 8661 26188
rect 8523 26144 8565 26153
rect 8523 26104 8524 26144
rect 8564 26104 8565 26144
rect 8523 26095 8565 26104
rect 8524 25556 8564 26095
rect 8524 25507 8564 25516
rect 8236 25432 8468 25472
rect 8236 23960 8276 25432
rect 8331 25304 8373 25313
rect 8331 25264 8332 25304
rect 8372 25264 8373 25304
rect 8331 25255 8373 25264
rect 8332 25170 8372 25255
rect 8427 25220 8469 25229
rect 8427 25180 8428 25220
rect 8468 25180 8469 25220
rect 8427 25171 8469 25180
rect 8428 25052 8468 25171
rect 8332 25012 8468 25052
rect 8523 25052 8565 25061
rect 8523 25012 8524 25052
rect 8564 25012 8565 25052
rect 8332 24632 8372 25012
rect 8523 25003 8565 25012
rect 8332 24583 8372 24592
rect 8427 24632 8469 24641
rect 8427 24592 8428 24632
rect 8468 24592 8469 24632
rect 8427 24583 8469 24592
rect 8428 24498 8468 24583
rect 8427 23960 8469 23969
rect 8236 23920 8428 23960
rect 8468 23920 8469 23960
rect 8427 23911 8469 23920
rect 8332 23792 8372 23803
rect 8332 23717 8372 23752
rect 8428 23792 8468 23911
rect 8428 23743 8468 23752
rect 8331 23708 8373 23717
rect 8331 23668 8332 23708
rect 8372 23668 8373 23708
rect 8331 23659 8373 23668
rect 8235 23540 8277 23549
rect 8235 23500 8236 23540
rect 8276 23500 8277 23540
rect 8235 23491 8277 23500
rect 8236 22280 8276 23491
rect 8428 23120 8468 23129
rect 8524 23120 8564 25003
rect 8468 23080 8564 23120
rect 8331 22448 8373 22457
rect 8331 22408 8332 22448
rect 8372 22408 8373 22448
rect 8331 22399 8373 22408
rect 8332 22364 8372 22399
rect 8332 22313 8372 22324
rect 8236 21281 8276 22240
rect 8428 22112 8468 23080
rect 8332 22072 8468 22112
rect 8235 21272 8277 21281
rect 8235 21232 8236 21272
rect 8276 21232 8277 21272
rect 8235 21223 8277 21232
rect 8140 20140 8276 20180
rect 8236 20096 8276 20140
rect 8236 19256 8276 20056
rect 8332 19937 8372 22072
rect 8524 20768 8564 20777
rect 8428 20264 8468 20273
rect 8524 20264 8564 20728
rect 8468 20224 8564 20264
rect 8620 20768 8660 26179
rect 8716 25817 8756 26776
rect 8812 26816 8852 26825
rect 8812 26153 8852 26776
rect 8811 26144 8853 26153
rect 8811 26104 8812 26144
rect 8852 26104 8853 26144
rect 8811 26095 8853 26104
rect 8715 25808 8757 25817
rect 8715 25768 8716 25808
rect 8756 25768 8757 25808
rect 8715 25759 8757 25768
rect 8908 25472 8948 26944
rect 9003 26900 9045 26909
rect 9003 26860 9004 26900
rect 9044 26860 9045 26900
rect 9003 26851 9045 26860
rect 9004 26816 9044 26851
rect 9004 25976 9044 26776
rect 9292 26489 9332 27616
rect 9388 28328 9428 28337
rect 9484 28328 9524 30211
rect 9428 28288 9524 28328
rect 9291 26480 9333 26489
rect 9291 26440 9292 26480
rect 9332 26440 9333 26480
rect 9291 26431 9333 26440
rect 9291 26228 9333 26237
rect 9291 26188 9292 26228
rect 9332 26188 9333 26228
rect 9291 26179 9333 26188
rect 9100 26144 9140 26153
rect 9100 26060 9140 26104
rect 9292 26094 9332 26179
rect 9195 26060 9237 26069
rect 9100 26020 9196 26060
rect 9236 26020 9237 26060
rect 9195 26011 9237 26020
rect 9004 25936 9140 25976
rect 9003 25808 9045 25817
rect 9003 25768 9004 25808
rect 9044 25768 9045 25808
rect 9003 25759 9045 25768
rect 8812 25432 8948 25472
rect 8715 25220 8757 25229
rect 8715 25180 8716 25220
rect 8756 25180 8757 25220
rect 8715 25171 8757 25180
rect 8716 25086 8756 25171
rect 8812 24464 8852 25432
rect 8908 25304 8948 25313
rect 8908 24977 8948 25264
rect 8907 24968 8949 24977
rect 8907 24928 8908 24968
rect 8948 24928 8949 24968
rect 8907 24919 8949 24928
rect 8908 24632 8948 24641
rect 9004 24632 9044 25759
rect 9100 24884 9140 25936
rect 9196 25313 9236 26011
rect 9388 25388 9428 28288
rect 9483 27656 9525 27665
rect 9483 27616 9484 27656
rect 9524 27616 9525 27656
rect 9483 27607 9525 27616
rect 9484 26825 9524 27607
rect 9483 26816 9525 26825
rect 9483 26776 9484 26816
rect 9524 26776 9525 26816
rect 9483 26767 9525 26776
rect 9292 25348 9428 25388
rect 9195 25304 9237 25313
rect 9195 25264 9196 25304
rect 9236 25264 9237 25304
rect 9195 25255 9237 25264
rect 9292 25061 9332 25348
rect 9387 25220 9429 25229
rect 9387 25180 9388 25220
rect 9428 25180 9429 25220
rect 9387 25171 9429 25180
rect 9291 25052 9333 25061
rect 9291 25012 9292 25052
rect 9332 25012 9333 25052
rect 9291 25003 9333 25012
rect 9100 24844 9332 24884
rect 8948 24592 9236 24632
rect 8908 24583 8948 24592
rect 8812 24424 8948 24464
rect 8811 23792 8853 23801
rect 8811 23752 8812 23792
rect 8852 23752 8853 23792
rect 8811 23743 8853 23752
rect 8908 23792 8948 24424
rect 8812 23658 8852 23743
rect 8908 23717 8948 23752
rect 8907 23708 8949 23717
rect 8907 23668 8908 23708
rect 8948 23668 8949 23708
rect 8907 23659 8949 23668
rect 8811 23456 8853 23465
rect 8811 23416 8812 23456
rect 8852 23416 8853 23456
rect 8811 23407 8853 23416
rect 8428 20215 8468 20224
rect 8331 19928 8373 19937
rect 8331 19888 8332 19928
rect 8372 19888 8373 19928
rect 8331 19879 8373 19888
rect 8332 19517 8372 19879
rect 8331 19508 8373 19517
rect 8331 19468 8332 19508
rect 8372 19468 8373 19508
rect 8331 19459 8373 19468
rect 8620 19424 8660 20728
rect 8812 22280 8852 23407
rect 9099 22532 9141 22541
rect 9099 22492 9100 22532
rect 9140 22492 9141 22532
rect 9099 22483 9141 22492
rect 8812 20180 8852 22240
rect 9100 21617 9140 22483
rect 9099 21608 9141 21617
rect 9099 21568 9100 21608
rect 9140 21568 9141 21608
rect 9099 21559 9141 21568
rect 9100 21474 9140 21559
rect 9099 20852 9141 20861
rect 9099 20812 9100 20852
rect 9140 20812 9141 20852
rect 9099 20803 9141 20812
rect 9004 20768 9044 20777
rect 9004 20180 9044 20728
rect 9100 20718 9140 20803
rect 8812 20140 8948 20180
rect 9004 20140 9140 20180
rect 8715 20096 8757 20105
rect 8715 20056 8716 20096
rect 8756 20056 8757 20096
rect 8715 20047 8757 20056
rect 8716 19962 8756 20047
rect 8620 19384 8852 19424
rect 8236 19013 8276 19216
rect 8716 19256 8756 19265
rect 8428 19172 8468 19181
rect 8716 19172 8756 19216
rect 8812 19256 8852 19384
rect 8908 19340 8948 20140
rect 8908 19300 9044 19340
rect 8852 19216 8948 19256
rect 8812 19207 8852 19216
rect 8468 19132 8756 19172
rect 8428 19123 8468 19132
rect 8235 19004 8277 19013
rect 8235 18964 8236 19004
rect 8276 18964 8277 19004
rect 8235 18955 8277 18964
rect 8332 17744 8372 17753
rect 8332 17249 8372 17704
rect 8812 17744 8852 17753
rect 8524 17660 8564 17669
rect 8812 17660 8852 17704
rect 8564 17620 8852 17660
rect 8908 17744 8948 19216
rect 9004 18257 9044 19300
rect 9100 19256 9140 20140
rect 9196 19433 9236 24592
rect 9292 23213 9332 24844
rect 9388 24627 9428 25171
rect 9484 24977 9524 26767
rect 9580 26312 9620 30388
rect 9868 29177 9908 29262
rect 9867 29168 9909 29177
rect 9867 29128 9868 29168
rect 9908 29128 9909 29168
rect 9867 29119 9909 29128
rect 9772 29084 9812 29093
rect 9772 29000 9812 29044
rect 9964 29000 10004 31396
rect 10060 31387 10100 31396
rect 10156 31436 10196 31639
rect 10156 31387 10196 31396
rect 10059 29504 10101 29513
rect 10059 29464 10060 29504
rect 10100 29464 10101 29504
rect 10059 29455 10101 29464
rect 9772 28960 10004 29000
rect 9771 27656 9813 27665
rect 9771 27616 9772 27656
rect 9812 27616 9813 27656
rect 9771 27607 9813 27616
rect 9675 27572 9717 27581
rect 9675 27532 9676 27572
rect 9716 27532 9717 27572
rect 9675 27523 9717 27532
rect 9676 27245 9716 27523
rect 9772 27522 9812 27607
rect 9868 27497 9908 28960
rect 10060 27908 10100 29455
rect 9964 27868 10100 27908
rect 9867 27488 9909 27497
rect 9867 27448 9868 27488
rect 9908 27448 9909 27488
rect 9867 27439 9909 27448
rect 9964 27320 10004 27868
rect 10252 27824 10292 39199
rect 10348 38249 10388 39460
rect 10732 38921 10772 39712
rect 10731 38912 10773 38921
rect 10731 38872 10732 38912
rect 10772 38872 10773 38912
rect 10731 38863 10773 38872
rect 10539 38576 10581 38585
rect 10539 38536 10540 38576
rect 10580 38536 10581 38576
rect 10539 38527 10581 38536
rect 10347 38240 10389 38249
rect 10347 38200 10348 38240
rect 10388 38200 10389 38240
rect 10347 38191 10389 38200
rect 10540 38240 10580 38527
rect 10732 38408 10772 38863
rect 10827 38492 10869 38501
rect 10827 38452 10828 38492
rect 10868 38452 10869 38492
rect 10827 38443 10869 38452
rect 10732 38359 10772 38368
rect 10580 38200 10676 38240
rect 10540 38191 10580 38200
rect 10636 38081 10676 38200
rect 10635 38072 10677 38081
rect 10635 38032 10636 38072
rect 10676 38032 10677 38072
rect 10635 38023 10677 38032
rect 10539 37988 10581 37997
rect 10539 37948 10540 37988
rect 10580 37948 10581 37988
rect 10539 37939 10581 37948
rect 10540 37400 10580 37939
rect 10580 37360 10676 37400
rect 10540 37351 10580 37360
rect 10347 36308 10389 36317
rect 10347 36268 10348 36308
rect 10388 36268 10389 36308
rect 10347 36259 10389 36268
rect 10348 35813 10388 36259
rect 10540 35888 10580 35897
rect 10347 35804 10389 35813
rect 10347 35764 10348 35804
rect 10388 35764 10389 35804
rect 10347 35755 10389 35764
rect 10443 35216 10485 35225
rect 10443 35176 10444 35216
rect 10484 35176 10485 35216
rect 10443 35167 10485 35176
rect 10347 35048 10389 35057
rect 10347 35008 10348 35048
rect 10388 35008 10389 35048
rect 10347 34999 10389 35008
rect 10348 34376 10388 34999
rect 10348 32948 10388 34336
rect 10444 33704 10484 35167
rect 10444 33655 10484 33664
rect 10348 32908 10484 32948
rect 10347 32780 10389 32789
rect 10347 32740 10348 32780
rect 10388 32740 10389 32780
rect 10347 32731 10389 32740
rect 10348 31697 10388 32731
rect 10347 31688 10389 31697
rect 10347 31648 10348 31688
rect 10388 31648 10389 31688
rect 10347 31639 10389 31648
rect 10348 29168 10388 29177
rect 10444 29168 10484 32908
rect 10540 31604 10580 35848
rect 10636 34217 10676 37360
rect 10828 36728 10868 38443
rect 10828 36149 10868 36688
rect 10827 36140 10869 36149
rect 10827 36100 10828 36140
rect 10868 36100 10869 36140
rect 10827 36091 10869 36100
rect 10924 35384 10964 40627
rect 11308 39920 11348 41635
rect 11404 40508 11444 46087
rect 11788 46061 11828 48355
rect 11884 48161 11924 48532
rect 11980 48532 12076 48572
rect 11883 48152 11925 48161
rect 11883 48112 11884 48152
rect 11924 48112 11925 48152
rect 11883 48103 11925 48112
rect 11980 47312 12020 48532
rect 12076 48523 12116 48532
rect 12171 48236 12213 48245
rect 12171 48196 12172 48236
rect 12212 48196 12213 48236
rect 12171 48187 12213 48196
rect 12075 47480 12117 47489
rect 12075 47440 12076 47480
rect 12116 47440 12117 47480
rect 12075 47431 12117 47440
rect 12076 47346 12116 47431
rect 11932 47302 12020 47312
rect 11972 47272 12020 47302
rect 11932 47253 11972 47262
rect 12172 46640 12212 48187
rect 12268 47984 12308 49456
rect 12460 49447 12500 49456
rect 12652 49456 12940 49496
rect 12652 49412 12692 49456
rect 12940 49447 12980 49456
rect 13036 49496 13076 49867
rect 13420 49496 13460 50119
rect 12652 49363 12692 49372
rect 13036 49328 13076 49456
rect 12844 49288 13076 49328
rect 13228 49456 13420 49496
rect 12268 47935 12308 47944
rect 12748 47984 12788 47993
rect 12460 47900 12500 47909
rect 12748 47900 12788 47944
rect 12500 47860 12788 47900
rect 12844 47984 12884 49288
rect 13131 48824 13173 48833
rect 13131 48784 13132 48824
rect 13172 48784 13173 48824
rect 13131 48775 13173 48784
rect 13132 48690 13172 48775
rect 13228 47984 13268 49456
rect 13420 49447 13460 49456
rect 13516 49496 13556 50203
rect 13612 49505 13652 50296
rect 13516 48572 13556 49456
rect 13611 49496 13653 49505
rect 13611 49456 13612 49496
rect 13652 49456 13653 49496
rect 13611 49447 13653 49456
rect 13611 49244 13653 49253
rect 13611 49204 13612 49244
rect 13652 49204 13653 49244
rect 13611 49195 13653 49204
rect 13420 48532 13556 48572
rect 12460 47851 12500 47860
rect 12267 47312 12309 47321
rect 12267 47272 12268 47312
rect 12308 47272 12309 47312
rect 12267 47263 12309 47272
rect 12076 46600 12212 46640
rect 11787 46052 11829 46061
rect 11787 46012 11788 46052
rect 11828 46012 11829 46052
rect 11787 46003 11829 46012
rect 11596 45800 11636 45809
rect 11636 45760 11732 45800
rect 11596 45751 11636 45760
rect 11595 45380 11637 45389
rect 11595 45340 11596 45380
rect 11636 45340 11637 45380
rect 11595 45331 11637 45340
rect 11499 45296 11541 45305
rect 11499 45256 11500 45296
rect 11540 45256 11541 45296
rect 11499 45247 11541 45256
rect 11500 44288 11540 45247
rect 11500 44239 11540 44248
rect 11596 43532 11636 45331
rect 11692 45305 11732 45760
rect 11788 45548 11828 45557
rect 11691 45296 11733 45305
rect 11691 45256 11692 45296
rect 11732 45256 11733 45296
rect 11691 45247 11733 45256
rect 11788 45044 11828 45508
rect 11740 45004 11828 45044
rect 11740 45002 11780 45004
rect 11740 44953 11780 44962
rect 11884 44792 11924 44801
rect 11884 44549 11924 44752
rect 11883 44540 11925 44549
rect 11883 44500 11884 44540
rect 11924 44500 11925 44540
rect 11883 44491 11925 44500
rect 12076 44456 12116 46600
rect 12172 46472 12212 46500
rect 12268 46472 12308 47263
rect 12844 46640 12884 47944
rect 13132 47944 13228 47984
rect 12940 47312 12980 47321
rect 12940 47069 12980 47272
rect 12939 47060 12981 47069
rect 12939 47020 12940 47060
rect 12980 47020 12981 47060
rect 12939 47011 12981 47020
rect 12939 46892 12981 46901
rect 12939 46852 12940 46892
rect 12980 46852 12981 46892
rect 12939 46843 12981 46852
rect 12748 46600 12884 46640
rect 12212 46432 12308 46472
rect 12172 46423 12212 46432
rect 12171 46052 12213 46061
rect 12171 46012 12172 46052
rect 12212 46012 12213 46052
rect 12171 46003 12213 46012
rect 12172 44960 12212 46003
rect 12172 44911 12212 44920
rect 12076 44416 12212 44456
rect 11692 44372 11732 44381
rect 11732 44332 12020 44372
rect 11692 44323 11732 44332
rect 11980 44288 12020 44332
rect 11980 44239 12020 44248
rect 12075 44288 12117 44297
rect 12075 44248 12076 44288
rect 12116 44248 12117 44288
rect 12075 44239 12117 44248
rect 12076 44154 12116 44239
rect 11884 43532 11924 43541
rect 11596 43492 11884 43532
rect 11884 43483 11924 43492
rect 11692 43280 11732 43289
rect 11692 42869 11732 43240
rect 11691 42860 11733 42869
rect 11691 42820 11692 42860
rect 11732 42820 11733 42860
rect 11691 42811 11733 42820
rect 11500 42776 11540 42785
rect 11500 42617 11540 42736
rect 12075 42776 12117 42785
rect 12075 42736 12076 42776
rect 12116 42736 12117 42776
rect 12075 42727 12117 42736
rect 11499 42608 11541 42617
rect 11499 42568 11500 42608
rect 11540 42568 11541 42608
rect 11499 42559 11541 42568
rect 11500 42029 11540 42559
rect 11691 42356 11733 42365
rect 11691 42316 11692 42356
rect 11732 42316 11733 42356
rect 11691 42307 11733 42316
rect 11499 42020 11541 42029
rect 11499 41980 11500 42020
rect 11540 41980 11541 42020
rect 11499 41971 11541 41980
rect 11500 40517 11540 40561
rect 11499 40508 11541 40517
rect 11404 40468 11500 40508
rect 11540 40468 11541 40508
rect 11499 40466 11541 40468
rect 11499 40459 11500 40466
rect 11540 40459 11541 40466
rect 11500 40417 11540 40426
rect 11212 39880 11348 39920
rect 11212 39080 11252 39880
rect 11308 39752 11348 39761
rect 11308 39341 11348 39712
rect 11307 39332 11349 39341
rect 11307 39292 11308 39332
rect 11348 39292 11349 39332
rect 11307 39283 11349 39292
rect 11020 39040 11252 39080
rect 11020 37820 11060 39040
rect 11212 38912 11252 38921
rect 11212 38669 11252 38872
rect 11404 38744 11444 38755
rect 11596 38744 11636 38753
rect 11404 38669 11444 38704
rect 11500 38704 11596 38744
rect 11211 38660 11253 38669
rect 11211 38620 11212 38660
rect 11252 38620 11253 38660
rect 11211 38611 11253 38620
rect 11403 38660 11445 38669
rect 11403 38620 11404 38660
rect 11444 38620 11445 38660
rect 11403 38611 11445 38620
rect 11115 38576 11157 38585
rect 11115 38536 11116 38576
rect 11156 38536 11157 38576
rect 11115 38527 11157 38536
rect 11116 38240 11156 38527
rect 11500 38492 11540 38704
rect 11596 38695 11636 38704
rect 11308 38452 11540 38492
rect 11116 38191 11156 38200
rect 11211 38240 11253 38249
rect 11211 38200 11212 38240
rect 11252 38200 11253 38240
rect 11211 38191 11253 38200
rect 11308 38240 11348 38452
rect 11692 38249 11732 42307
rect 11883 38996 11925 39005
rect 11883 38956 11884 38996
rect 11924 38956 11925 38996
rect 11883 38947 11925 38956
rect 11788 38912 11828 38921
rect 11788 38669 11828 38872
rect 11884 38912 11924 38947
rect 11787 38660 11829 38669
rect 11787 38620 11788 38660
rect 11828 38620 11829 38660
rect 11787 38611 11829 38620
rect 11308 38191 11348 38200
rect 11404 38240 11444 38249
rect 11212 38106 11252 38191
rect 11307 38072 11349 38081
rect 11307 38032 11308 38072
rect 11348 38032 11349 38072
rect 11307 38023 11349 38032
rect 11020 37780 11252 37820
rect 11068 35897 11108 35906
rect 11108 35857 11156 35888
rect 11068 35848 11156 35857
rect 11116 35384 11156 35848
rect 11212 35804 11252 37780
rect 11212 35755 11252 35764
rect 11211 35636 11253 35645
rect 11211 35596 11212 35636
rect 11252 35596 11253 35636
rect 11211 35587 11253 35596
rect 10924 35344 11060 35384
rect 10923 35216 10965 35225
rect 10923 35176 10924 35216
rect 10964 35176 10965 35216
rect 10923 35167 10965 35176
rect 10924 35082 10964 35167
rect 11020 34889 11060 35344
rect 11116 35335 11156 35344
rect 11019 34880 11061 34889
rect 11019 34840 11020 34880
rect 11060 34840 11061 34880
rect 11019 34831 11061 34840
rect 11019 34628 11061 34637
rect 11019 34588 11020 34628
rect 11060 34588 11061 34628
rect 11019 34579 11061 34588
rect 10828 34381 10868 34390
rect 10732 34341 10828 34381
rect 10635 34208 10677 34217
rect 10635 34168 10636 34208
rect 10676 34168 10677 34208
rect 10635 34159 10677 34168
rect 10636 33872 10676 33881
rect 10732 33872 10772 34341
rect 10828 34332 10868 34341
rect 11020 34292 11060 34579
rect 11020 34243 11060 34252
rect 10676 33832 10772 33872
rect 10636 33823 10676 33832
rect 11020 33797 11060 33828
rect 11019 33788 11061 33797
rect 11019 33748 11020 33788
rect 11060 33748 11061 33788
rect 11019 33739 11061 33748
rect 10924 33704 10964 33713
rect 10828 33032 10868 33041
rect 10924 33032 10964 33664
rect 11020 33704 11060 33739
rect 11020 33293 11060 33664
rect 11019 33284 11061 33293
rect 11019 33244 11020 33284
rect 11060 33244 11061 33284
rect 11019 33235 11061 33244
rect 10868 32992 10964 33032
rect 10828 32983 10868 32992
rect 10635 32948 10677 32957
rect 11020 32948 11060 33235
rect 10635 32908 10636 32948
rect 10676 32908 10677 32948
rect 10635 32899 10677 32908
rect 10924 32908 11060 32948
rect 10636 32864 10676 32899
rect 10636 32813 10676 32824
rect 10731 32696 10773 32705
rect 10731 32656 10732 32696
rect 10772 32656 10773 32696
rect 10731 32647 10773 32656
rect 10732 32192 10772 32647
rect 10635 31604 10677 31613
rect 10540 31564 10636 31604
rect 10676 31564 10677 31604
rect 10635 31555 10677 31564
rect 10636 31352 10676 31555
rect 10636 31303 10676 31312
rect 10539 30680 10581 30689
rect 10539 30640 10540 30680
rect 10580 30640 10581 30680
rect 10539 30631 10581 30640
rect 10388 29128 10484 29168
rect 10348 28337 10388 29128
rect 10347 28328 10389 28337
rect 10347 28288 10348 28328
rect 10388 28288 10389 28328
rect 10540 28328 10580 30631
rect 10732 30521 10772 32152
rect 10731 30512 10773 30521
rect 10731 30472 10732 30512
rect 10772 30472 10773 30512
rect 10731 30463 10773 30472
rect 10635 29924 10677 29933
rect 10635 29884 10636 29924
rect 10676 29884 10677 29924
rect 10635 29875 10677 29884
rect 10636 29000 10676 29875
rect 10924 29513 10964 32908
rect 11020 32822 11060 32831
rect 11020 32705 11060 32782
rect 11019 32696 11061 32705
rect 11019 32656 11020 32696
rect 11060 32656 11061 32696
rect 11019 32647 11061 32656
rect 11212 31520 11252 35587
rect 11020 31480 11252 31520
rect 11020 29933 11060 31480
rect 11164 31361 11204 31370
rect 11308 31361 11348 38023
rect 11404 36317 11444 38200
rect 11691 38240 11733 38249
rect 11691 38200 11692 38240
rect 11732 38200 11733 38240
rect 11691 38191 11733 38200
rect 11595 37568 11637 37577
rect 11595 37528 11596 37568
rect 11636 37528 11637 37568
rect 11595 37519 11637 37528
rect 11403 36308 11445 36317
rect 11403 36268 11404 36308
rect 11444 36268 11445 36308
rect 11403 36259 11445 36268
rect 11403 36140 11445 36149
rect 11403 36100 11404 36140
rect 11444 36100 11445 36140
rect 11403 36091 11445 36100
rect 11404 35888 11444 36091
rect 11404 35839 11444 35848
rect 11403 34796 11445 34805
rect 11403 34756 11404 34796
rect 11444 34756 11445 34796
rect 11403 34747 11445 34756
rect 11404 33881 11444 34747
rect 11499 33956 11541 33965
rect 11499 33916 11500 33956
rect 11540 33916 11541 33956
rect 11499 33907 11541 33916
rect 11403 33872 11445 33881
rect 11403 33832 11404 33872
rect 11444 33832 11445 33872
rect 11403 33823 11445 33832
rect 11404 33704 11444 33823
rect 11404 33655 11444 33664
rect 11500 33629 11540 33907
rect 11499 33620 11541 33629
rect 11499 33580 11500 33620
rect 11540 33580 11541 33620
rect 11499 33571 11541 33580
rect 11500 33486 11540 33571
rect 11596 32957 11636 37519
rect 11692 37400 11732 38191
rect 11884 38165 11924 38872
rect 11979 38912 12021 38921
rect 11979 38872 11980 38912
rect 12020 38872 12021 38912
rect 11979 38863 12021 38872
rect 11980 38778 12020 38863
rect 11883 38156 11925 38165
rect 11883 38116 11884 38156
rect 11924 38116 11925 38156
rect 11883 38107 11925 38116
rect 12076 37577 12116 42727
rect 12075 37568 12117 37577
rect 12075 37528 12076 37568
rect 12116 37528 12117 37568
rect 12075 37519 12117 37528
rect 11788 37400 11828 37409
rect 11692 37360 11788 37400
rect 11828 37360 12116 37400
rect 11788 37351 11828 37360
rect 11980 37232 12020 37241
rect 11787 36812 11829 36821
rect 11787 36772 11788 36812
rect 11828 36772 11829 36812
rect 11787 36763 11829 36772
rect 11691 36476 11733 36485
rect 11691 36436 11692 36476
rect 11732 36436 11733 36476
rect 11691 36427 11733 36436
rect 11595 32948 11637 32957
rect 11595 32908 11596 32948
rect 11636 32908 11637 32948
rect 11595 32899 11637 32908
rect 11307 31352 11349 31361
rect 11204 31321 11252 31352
rect 11164 31312 11252 31321
rect 11212 30848 11252 31312
rect 11307 31312 11308 31352
rect 11348 31312 11349 31352
rect 11307 31303 11349 31312
rect 11308 31184 11348 31193
rect 11348 31144 11540 31184
rect 11308 31135 11348 31144
rect 11500 30941 11540 31144
rect 11499 30932 11541 30941
rect 11499 30892 11500 30932
rect 11540 30892 11541 30932
rect 11499 30883 11541 30892
rect 11308 30848 11348 30857
rect 11212 30808 11308 30848
rect 11308 30799 11348 30808
rect 11115 30680 11157 30689
rect 11115 30640 11116 30680
rect 11156 30640 11157 30680
rect 11115 30631 11157 30640
rect 11403 30680 11445 30689
rect 11403 30640 11404 30680
rect 11444 30640 11445 30680
rect 11403 30631 11445 30640
rect 11500 30680 11540 30691
rect 11116 30546 11156 30631
rect 11211 30512 11253 30521
rect 11211 30472 11212 30512
rect 11252 30472 11253 30512
rect 11211 30463 11253 30472
rect 11115 30260 11157 30269
rect 11115 30220 11116 30260
rect 11156 30220 11157 30260
rect 11115 30211 11157 30220
rect 11019 29924 11061 29933
rect 11019 29884 11020 29924
rect 11060 29884 11061 29924
rect 11019 29875 11061 29884
rect 10923 29504 10965 29513
rect 10923 29464 10924 29504
rect 10964 29464 10965 29504
rect 10923 29455 10965 29464
rect 10828 29154 10868 29163
rect 10636 28960 10772 29000
rect 10732 28412 10772 28960
rect 10828 28580 10868 29114
rect 10924 29093 10964 29455
rect 11020 29252 11060 29261
rect 10923 29084 10965 29093
rect 10923 29044 10924 29084
rect 10964 29044 10965 29084
rect 10923 29035 10965 29044
rect 10828 28531 10868 28540
rect 11020 28505 11060 29212
rect 11116 28757 11156 30211
rect 11115 28748 11157 28757
rect 11115 28708 11116 28748
rect 11156 28708 11157 28748
rect 11115 28699 11157 28708
rect 11019 28496 11061 28505
rect 11019 28456 11020 28496
rect 11060 28456 11061 28496
rect 11019 28447 11061 28456
rect 10732 28372 10868 28412
rect 10636 28328 10676 28337
rect 10540 28288 10636 28328
rect 10347 28279 10389 28288
rect 10636 28279 10676 28288
rect 9868 27280 10004 27320
rect 10060 27784 10292 27824
rect 9675 27236 9717 27245
rect 9675 27196 9676 27236
rect 9716 27196 9717 27236
rect 9675 27187 9717 27196
rect 9580 26272 9716 26312
rect 9579 26144 9621 26153
rect 9579 26104 9580 26144
rect 9620 26104 9621 26144
rect 9579 26095 9621 26104
rect 9676 26144 9716 26272
rect 9771 26228 9813 26237
rect 9771 26188 9772 26228
rect 9812 26188 9813 26228
rect 9771 26179 9813 26188
rect 9580 26010 9620 26095
rect 9483 24968 9525 24977
rect 9483 24928 9484 24968
rect 9524 24928 9525 24968
rect 9483 24919 9525 24928
rect 9579 24716 9621 24725
rect 9579 24676 9580 24716
rect 9620 24676 9621 24716
rect 9579 24667 9621 24676
rect 9388 24578 9428 24587
rect 9580 24582 9620 24667
rect 9483 24464 9525 24473
rect 9483 24424 9484 24464
rect 9524 24424 9525 24464
rect 9483 24415 9525 24424
rect 9388 23792 9428 23801
rect 9291 23204 9333 23213
rect 9291 23164 9292 23204
rect 9332 23164 9333 23204
rect 9291 23155 9333 23164
rect 9292 22285 9332 22294
rect 9292 21776 9332 22245
rect 9292 21727 9332 21736
rect 9291 20852 9333 20861
rect 9291 20812 9292 20852
rect 9332 20812 9333 20852
rect 9291 20803 9333 20812
rect 9195 19424 9237 19433
rect 9195 19384 9196 19424
rect 9236 19384 9237 19424
rect 9195 19375 9237 19384
rect 9196 19256 9236 19265
rect 9100 19216 9196 19256
rect 9100 18584 9140 18593
rect 9100 18509 9140 18544
rect 9099 18500 9141 18509
rect 9099 18460 9100 18500
rect 9140 18460 9141 18500
rect 9099 18451 9141 18460
rect 9003 18248 9045 18257
rect 9003 18208 9004 18248
rect 9044 18208 9045 18248
rect 9003 18199 9045 18208
rect 9100 17837 9140 18451
rect 9099 17828 9141 17837
rect 9099 17788 9100 17828
rect 9140 17788 9141 17828
rect 9099 17779 9141 17788
rect 9196 17744 9236 19216
rect 9292 19256 9332 20803
rect 9388 20105 9428 23752
rect 9484 23129 9524 24415
rect 9676 23465 9716 26104
rect 9772 26144 9812 26179
rect 9772 26093 9812 26104
rect 9868 25733 9908 27280
rect 9964 26312 10004 26321
rect 9964 26153 10004 26272
rect 9963 26144 10005 26153
rect 9963 26104 9964 26144
rect 10004 26104 10005 26144
rect 9963 26095 10005 26104
rect 9867 25724 9909 25733
rect 9867 25684 9868 25724
rect 9908 25684 9909 25724
rect 9867 25675 9909 25684
rect 9771 25304 9813 25313
rect 9771 25264 9772 25304
rect 9812 25264 9813 25304
rect 9771 25255 9813 25264
rect 9675 23456 9717 23465
rect 9675 23416 9676 23456
rect 9716 23416 9717 23456
rect 9675 23407 9717 23416
rect 9483 23120 9525 23129
rect 9676 23120 9716 23129
rect 9483 23080 9484 23120
rect 9524 23080 9525 23120
rect 9483 23071 9525 23080
rect 9580 23080 9676 23120
rect 9580 22541 9620 23080
rect 9676 23071 9716 23080
rect 9772 22952 9812 25255
rect 9964 24632 10004 24641
rect 9964 23969 10004 24592
rect 10060 24212 10100 27784
rect 10252 27656 10292 27665
rect 10252 27413 10292 27616
rect 10251 27404 10293 27413
rect 10251 27364 10252 27404
rect 10292 27364 10293 27404
rect 10251 27355 10293 27364
rect 10252 26825 10292 26910
rect 10251 26816 10293 26825
rect 10251 26776 10252 26816
rect 10292 26776 10293 26816
rect 10251 26767 10293 26776
rect 10251 26648 10293 26657
rect 10251 26608 10252 26648
rect 10292 26608 10293 26648
rect 10251 26599 10293 26608
rect 10155 26228 10197 26237
rect 10155 26188 10156 26228
rect 10196 26188 10197 26228
rect 10155 26179 10197 26188
rect 10156 26144 10196 26179
rect 10156 26093 10196 26104
rect 10252 26144 10292 26599
rect 10348 26489 10388 28279
rect 10732 27642 10772 27651
rect 10732 27152 10772 27602
rect 10444 27112 10772 27152
rect 10444 27068 10484 27112
rect 10828 27068 10868 28372
rect 10923 27740 10965 27749
rect 10923 27700 10924 27740
rect 10964 27700 10965 27740
rect 10923 27691 10965 27700
rect 10924 27606 10964 27691
rect 10444 27019 10484 27028
rect 10732 27028 10868 27068
rect 10636 26816 10676 26825
rect 10636 26489 10676 26776
rect 10347 26480 10389 26489
rect 10347 26440 10348 26480
rect 10388 26440 10389 26480
rect 10347 26431 10389 26440
rect 10635 26480 10677 26489
rect 10635 26440 10636 26480
rect 10676 26440 10677 26480
rect 10635 26431 10677 26440
rect 10443 26228 10485 26237
rect 10443 26188 10444 26228
rect 10484 26188 10485 26228
rect 10443 26179 10485 26188
rect 10252 26095 10292 26104
rect 10347 26144 10389 26153
rect 10347 26104 10348 26144
rect 10388 26104 10389 26144
rect 10347 26095 10389 26104
rect 10348 26010 10388 26095
rect 10444 26094 10484 26179
rect 10635 26144 10677 26153
rect 10635 26104 10636 26144
rect 10676 26104 10677 26144
rect 10635 26095 10677 26104
rect 10636 26010 10676 26095
rect 10155 25724 10197 25733
rect 10155 25684 10156 25724
rect 10196 25684 10197 25724
rect 10155 25675 10197 25684
rect 10156 25313 10196 25675
rect 10155 25304 10197 25313
rect 10155 25264 10156 25304
rect 10196 25264 10197 25304
rect 10155 25255 10197 25264
rect 10156 25170 10196 25255
rect 10732 24800 10772 27028
rect 11116 26648 11156 28699
rect 10924 26608 11156 26648
rect 10636 24760 10772 24800
rect 10828 25304 10868 25313
rect 10252 24641 10292 24726
rect 10251 24632 10293 24641
rect 10251 24592 10252 24632
rect 10292 24592 10293 24632
rect 10251 24583 10293 24592
rect 10444 24632 10484 24641
rect 10636 24632 10676 24760
rect 10484 24592 10676 24632
rect 10731 24632 10773 24641
rect 10731 24592 10732 24632
rect 10772 24592 10773 24632
rect 10444 24583 10484 24592
rect 10252 24380 10292 24389
rect 10292 24340 10388 24380
rect 10252 24331 10292 24340
rect 10060 24172 10292 24212
rect 9963 23960 10005 23969
rect 9963 23920 9964 23960
rect 10004 23920 10005 23960
rect 9963 23911 10005 23920
rect 9868 23797 9908 23806
rect 9868 23288 9908 23757
rect 9868 23239 9908 23248
rect 9867 23120 9909 23129
rect 9867 23080 9868 23120
rect 9908 23080 9909 23120
rect 9867 23071 9909 23080
rect 9676 22912 9812 22952
rect 9579 22532 9621 22541
rect 9579 22492 9580 22532
rect 9620 22492 9621 22532
rect 9579 22483 9621 22492
rect 9483 22112 9525 22121
rect 9483 22072 9484 22112
rect 9524 22072 9525 22112
rect 9483 22063 9525 22072
rect 9484 21978 9524 22063
rect 9484 21608 9524 21617
rect 9484 21029 9524 21568
rect 9483 21020 9525 21029
rect 9483 20980 9484 21020
rect 9524 20980 9525 21020
rect 9483 20971 9525 20980
rect 9387 20096 9429 20105
rect 9387 20056 9388 20096
rect 9428 20056 9429 20096
rect 9387 20047 9429 20056
rect 9332 19216 9428 19256
rect 9292 19207 9332 19216
rect 9292 17744 9332 17753
rect 9196 17704 9292 17744
rect 8524 17611 8564 17620
rect 8908 17576 8948 17704
rect 8716 17536 8948 17576
rect 8716 17324 8756 17536
rect 9292 17324 9332 17704
rect 8524 17284 8756 17324
rect 9100 17284 9332 17324
rect 9388 17744 9428 19216
rect 8331 17240 8373 17249
rect 8331 17200 8332 17240
rect 8372 17200 8373 17240
rect 8331 17191 8373 17200
rect 8139 16904 8181 16913
rect 8139 16864 8140 16904
rect 8180 16864 8181 16904
rect 8139 16855 8181 16864
rect 7948 14167 7988 14176
rect 8043 14216 8085 14225
rect 8043 14176 8044 14216
rect 8084 14176 8085 14216
rect 8043 14167 8085 14176
rect 7660 14092 7796 14132
rect 7660 13040 7700 14092
rect 7756 14034 7796 14043
rect 7756 13217 7796 13994
rect 7755 13208 7797 13217
rect 7755 13168 7756 13208
rect 7796 13168 7797 13208
rect 7755 13159 7797 13168
rect 7660 13000 7892 13040
rect 7564 12916 7796 12956
rect 7275 12907 7317 12916
rect 7179 11108 7221 11117
rect 7179 11068 7180 11108
rect 7220 11068 7221 11108
rect 7179 11059 7221 11068
rect 7180 10974 7220 11059
rect 7084 10387 7124 10396
rect 7276 10184 7316 12907
rect 7563 11780 7605 11789
rect 7563 11740 7564 11780
rect 7604 11740 7605 11780
rect 7563 11731 7605 11740
rect 7180 10144 7316 10184
rect 7372 11701 7412 11710
rect 7084 9689 7124 9774
rect 7083 9680 7125 9689
rect 7083 9640 7084 9680
rect 7124 9640 7125 9680
rect 7083 9631 7125 9640
rect 7083 9512 7125 9521
rect 7083 9472 7084 9512
rect 7124 9472 7125 9512
rect 7083 9463 7125 9472
rect 7084 8849 7124 9463
rect 7083 8840 7125 8849
rect 7083 8800 7084 8840
rect 7124 8800 7125 8840
rect 7083 8791 7125 8800
rect 6987 8168 7029 8177
rect 6987 8128 6988 8168
rect 7028 8128 7029 8168
rect 6987 8119 7029 8128
rect 7084 8000 7124 8791
rect 7084 7925 7124 7960
rect 6891 7916 6933 7925
rect 6891 7876 6892 7916
rect 6932 7876 6933 7916
rect 6891 7867 6933 7876
rect 7083 7916 7125 7925
rect 7083 7876 7084 7916
rect 7124 7876 7125 7916
rect 7083 7867 7125 7876
rect 7083 7748 7125 7757
rect 7083 7708 7084 7748
rect 7124 7708 7125 7748
rect 7083 7699 7125 7708
rect 6508 7540 6740 7580
rect 6795 7580 6837 7589
rect 6795 7540 6796 7580
rect 6836 7540 6837 7580
rect 6411 7160 6453 7169
rect 6411 7120 6412 7160
rect 6452 7120 6453 7160
rect 6411 7111 6453 7120
rect 6412 7026 6452 7111
rect 6315 6992 6357 7001
rect 6315 6952 6316 6992
rect 6356 6952 6357 6992
rect 6315 6943 6357 6952
rect 6123 6824 6165 6833
rect 6123 6784 6124 6824
rect 6164 6784 6165 6824
rect 6123 6775 6165 6784
rect 5931 5564 5973 5573
rect 5931 5524 5932 5564
rect 5972 5524 5973 5564
rect 5931 5515 5973 5524
rect 6028 5237 6068 6448
rect 6027 5228 6069 5237
rect 6027 5188 6028 5228
rect 6068 5188 6069 5228
rect 6027 5179 6069 5188
rect 5932 4901 5972 4986
rect 5931 4892 5973 4901
rect 5931 4852 5932 4892
rect 5972 4852 5973 4892
rect 5931 4843 5973 4852
rect 6028 4892 6068 4901
rect 5931 4640 5973 4649
rect 5931 4600 5932 4640
rect 5972 4600 5973 4640
rect 5931 4591 5973 4600
rect 5836 3583 5876 3592
rect 5932 3464 5972 4591
rect 5644 2500 5780 2540
rect 5836 3424 5972 3464
rect 5547 944 5589 953
rect 5547 904 5548 944
rect 5588 904 5589 944
rect 5547 895 5589 904
rect 5644 80 5684 2500
rect 5836 80 5876 3424
rect 6028 3380 6068 4852
rect 5932 3340 6068 3380
rect 5932 617 5972 3340
rect 6027 3212 6069 3221
rect 6027 3172 6028 3212
rect 6068 3172 6069 3212
rect 6027 3163 6069 3172
rect 6028 3078 6068 3163
rect 6124 2540 6164 6775
rect 6411 6236 6453 6245
rect 6411 6196 6412 6236
rect 6452 6196 6453 6236
rect 6411 6187 6453 6196
rect 6219 5984 6261 5993
rect 6219 5944 6220 5984
rect 6260 5944 6261 5984
rect 6219 5935 6261 5944
rect 6220 4649 6260 5935
rect 6316 5648 6356 5657
rect 6412 5648 6452 6187
rect 6508 5900 6548 7540
rect 6795 7531 6837 7540
rect 6988 7165 7028 7174
rect 6604 6992 6644 7001
rect 6604 6749 6644 6952
rect 6795 6992 6837 7001
rect 6795 6952 6796 6992
rect 6836 6952 6837 6992
rect 6795 6943 6837 6952
rect 6796 6858 6836 6943
rect 6988 6749 7028 7125
rect 6603 6740 6645 6749
rect 6603 6700 6604 6740
rect 6644 6700 6645 6740
rect 6603 6691 6645 6700
rect 6987 6740 7029 6749
rect 6987 6700 6988 6740
rect 7028 6700 7029 6740
rect 6987 6691 7029 6700
rect 6508 5851 6548 5860
rect 6796 5648 6836 5657
rect 6356 5608 6452 5648
rect 6700 5608 6796 5648
rect 6316 5321 6356 5608
rect 6315 5312 6357 5321
rect 6315 5272 6316 5312
rect 6356 5272 6357 5312
rect 6315 5263 6357 5272
rect 6508 4976 6548 4985
rect 6412 4957 6452 4966
rect 6412 4817 6452 4917
rect 6411 4808 6453 4817
rect 6411 4768 6412 4808
rect 6452 4768 6453 4808
rect 6411 4759 6453 4768
rect 6219 4640 6261 4649
rect 6219 4600 6220 4640
rect 6260 4600 6261 4640
rect 6219 4591 6261 4600
rect 6315 4220 6357 4229
rect 6508 4220 6548 4936
rect 6315 4180 6316 4220
rect 6356 4180 6357 4220
rect 6315 4171 6357 4180
rect 6412 4180 6548 4220
rect 6220 3464 6260 3473
rect 6220 2633 6260 3424
rect 6219 2624 6261 2633
rect 6219 2584 6220 2624
rect 6260 2584 6261 2624
rect 6219 2575 6261 2584
rect 6028 2500 6164 2540
rect 5931 608 5973 617
rect 5931 568 5932 608
rect 5972 568 5973 608
rect 5931 559 5973 568
rect 6028 80 6068 2500
rect 6123 2120 6165 2129
rect 6123 2080 6124 2120
rect 6164 2080 6165 2120
rect 6123 2071 6165 2080
rect 6124 281 6164 2071
rect 6220 2036 6260 2575
rect 6316 2213 6356 4171
rect 6412 3221 6452 4180
rect 6604 4136 6644 4145
rect 6508 4096 6604 4136
rect 6411 3212 6453 3221
rect 6411 3172 6412 3212
rect 6452 3172 6453 3212
rect 6411 3163 6453 3172
rect 6508 2624 6548 4096
rect 6604 4087 6644 4096
rect 6700 2876 6740 5608
rect 6796 5599 6836 5608
rect 6891 5648 6933 5657
rect 6891 5608 6892 5648
rect 6932 5608 6933 5648
rect 6891 5599 6933 5608
rect 6892 5514 6932 5599
rect 7084 5060 7124 7699
rect 7180 5480 7220 10144
rect 7275 10016 7317 10025
rect 7275 9976 7276 10016
rect 7316 9976 7317 10016
rect 7275 9967 7317 9976
rect 7276 9882 7316 9967
rect 7372 9689 7412 11661
rect 7564 11612 7604 11731
rect 7756 11621 7796 12916
rect 7852 11705 7892 13000
rect 7947 12788 7989 12797
rect 7947 12748 7948 12788
rect 7988 12748 7989 12788
rect 7947 12739 7989 12748
rect 7851 11696 7893 11705
rect 7851 11656 7852 11696
rect 7892 11656 7893 11696
rect 7851 11647 7893 11656
rect 7564 11563 7604 11572
rect 7755 11612 7797 11621
rect 7755 11572 7756 11612
rect 7796 11572 7797 11612
rect 7755 11563 7797 11572
rect 7467 10940 7509 10949
rect 7467 10900 7468 10940
rect 7508 10900 7509 10940
rect 7467 10891 7509 10900
rect 7468 10268 7508 10891
rect 7468 10219 7508 10228
rect 7467 10100 7509 10109
rect 7467 10060 7468 10100
rect 7508 10060 7509 10100
rect 7467 10051 7509 10060
rect 7371 9680 7413 9689
rect 7371 9640 7372 9680
rect 7412 9640 7413 9680
rect 7371 9631 7413 9640
rect 7276 9512 7316 9521
rect 7276 9353 7316 9472
rect 7275 9344 7317 9353
rect 7275 9304 7276 9344
rect 7316 9304 7317 9344
rect 7275 9295 7317 9304
rect 7372 8672 7412 8681
rect 7275 8168 7317 8177
rect 7275 8128 7276 8168
rect 7316 8128 7317 8168
rect 7275 8119 7317 8128
rect 7276 8034 7316 8119
rect 7275 7160 7317 7169
rect 7275 7120 7276 7160
rect 7316 7120 7317 7160
rect 7275 7111 7317 7120
rect 7276 6665 7316 7111
rect 7275 6656 7317 6665
rect 7275 6616 7276 6656
rect 7316 6616 7317 6656
rect 7372 6656 7412 8632
rect 7468 8672 7508 10051
rect 7756 9353 7796 11563
rect 7755 9344 7797 9353
rect 7755 9304 7756 9344
rect 7796 9304 7797 9344
rect 7755 9295 7797 9304
rect 7852 8756 7892 11647
rect 7468 8623 7508 8632
rect 7563 8672 7605 8681
rect 7563 8632 7564 8672
rect 7604 8632 7605 8672
rect 7563 8623 7605 8632
rect 7467 7748 7509 7757
rect 7467 7708 7468 7748
rect 7508 7708 7509 7748
rect 7467 7699 7509 7708
rect 7468 7614 7508 7699
rect 7467 7160 7509 7169
rect 7467 7120 7468 7160
rect 7508 7120 7509 7160
rect 7467 7111 7509 7120
rect 7468 7026 7508 7111
rect 7468 6656 7508 6665
rect 7372 6616 7468 6656
rect 7275 6607 7317 6616
rect 7468 6607 7508 6616
rect 7276 6488 7316 6607
rect 7276 6439 7316 6448
rect 7371 5900 7413 5909
rect 7371 5860 7372 5900
rect 7412 5860 7413 5900
rect 7371 5851 7413 5860
rect 7275 5732 7317 5741
rect 7275 5692 7276 5732
rect 7316 5692 7317 5732
rect 7275 5683 7317 5692
rect 7372 5732 7412 5851
rect 7372 5683 7412 5692
rect 7276 5598 7316 5683
rect 7180 5440 7316 5480
rect 7180 5153 7220 5238
rect 7179 5144 7221 5153
rect 7179 5104 7180 5144
rect 7220 5104 7221 5144
rect 7179 5095 7221 5104
rect 6892 5020 7124 5060
rect 6795 4808 6837 4817
rect 6795 4768 6796 4808
rect 6836 4768 6837 4808
rect 6795 4759 6837 4768
rect 6796 4674 6836 4759
rect 6795 4388 6837 4397
rect 6795 4348 6796 4388
rect 6836 4348 6837 4388
rect 6795 4339 6837 4348
rect 6796 4254 6836 4339
rect 6700 2827 6740 2836
rect 6795 2792 6837 2801
rect 6795 2752 6796 2792
rect 6836 2752 6837 2792
rect 6795 2743 6837 2752
rect 6411 2540 6453 2549
rect 6411 2500 6412 2540
rect 6452 2500 6453 2540
rect 6411 2491 6453 2500
rect 6315 2204 6357 2213
rect 6315 2164 6316 2204
rect 6356 2164 6357 2204
rect 6315 2155 6357 2164
rect 6220 1996 6356 2036
rect 6316 1364 6356 1996
rect 6412 1709 6452 2491
rect 6508 1952 6548 2584
rect 6699 2120 6741 2129
rect 6699 2080 6700 2120
rect 6740 2080 6741 2120
rect 6699 2071 6741 2080
rect 6700 1986 6740 2071
rect 6411 1700 6453 1709
rect 6411 1660 6412 1700
rect 6452 1660 6453 1700
rect 6411 1651 6453 1660
rect 6508 1541 6548 1912
rect 6507 1532 6549 1541
rect 6507 1492 6508 1532
rect 6548 1492 6549 1532
rect 6507 1483 6549 1492
rect 6316 1324 6548 1364
rect 6411 1196 6453 1205
rect 6411 1156 6412 1196
rect 6452 1156 6453 1196
rect 6411 1147 6453 1156
rect 6123 272 6165 281
rect 6123 232 6124 272
rect 6164 232 6165 272
rect 6123 223 6165 232
rect 6219 188 6261 197
rect 6219 148 6220 188
rect 6260 148 6261 188
rect 6219 139 6261 148
rect 6220 80 6260 139
rect 6412 80 6452 1147
rect 6508 1112 6548 1324
rect 6700 1280 6740 1289
rect 6796 1280 6836 2743
rect 6892 2549 6932 5020
rect 7179 4976 7221 4985
rect 7179 4936 7180 4976
rect 7220 4936 7221 4976
rect 7179 4927 7221 4936
rect 6988 4892 7028 4901
rect 7028 4852 7124 4892
rect 6988 4843 7028 4852
rect 6987 4724 7029 4733
rect 6987 4684 6988 4724
rect 7028 4684 7029 4724
rect 6987 4675 7029 4684
rect 6988 4136 7028 4675
rect 6988 4087 7028 4096
rect 7084 3137 7124 4852
rect 7083 3128 7125 3137
rect 7083 3088 7084 3128
rect 7124 3088 7125 3128
rect 7083 3079 7125 3088
rect 6987 2708 7029 2717
rect 6987 2668 6988 2708
rect 7028 2668 7029 2708
rect 6987 2659 7029 2668
rect 6988 2624 7028 2659
rect 7084 2633 7124 2718
rect 6988 2573 7028 2584
rect 7083 2624 7125 2633
rect 7083 2584 7084 2624
rect 7124 2584 7125 2624
rect 7083 2575 7125 2584
rect 6891 2540 6933 2549
rect 6891 2500 6892 2540
rect 6932 2500 6933 2540
rect 6891 2491 6933 2500
rect 7180 2456 7220 4927
rect 7276 4724 7316 5440
rect 7467 5312 7509 5321
rect 7467 5272 7468 5312
rect 7508 5272 7509 5312
rect 7467 5263 7509 5272
rect 7468 5069 7508 5263
rect 7467 5060 7509 5069
rect 7467 5020 7468 5060
rect 7508 5020 7509 5060
rect 7467 5011 7509 5020
rect 7372 4901 7412 4986
rect 7564 4976 7604 8623
rect 7660 7916 7700 7925
rect 7852 7916 7892 8716
rect 7948 8756 7988 12739
rect 8044 12629 8084 12660
rect 8043 12620 8085 12629
rect 8043 12580 8044 12620
rect 8084 12580 8085 12620
rect 8043 12571 8085 12580
rect 8044 12536 8084 12571
rect 8044 11453 8084 12496
rect 8140 11873 8180 16855
rect 8236 16232 8276 16241
rect 8236 15728 8276 16192
rect 8332 16232 8372 16241
rect 8524 16232 8564 17284
rect 8619 17072 8661 17081
rect 8619 17032 8620 17072
rect 8660 17032 8661 17072
rect 8619 17023 8661 17032
rect 8620 16938 8660 17023
rect 9100 16241 9140 17284
rect 9195 17156 9237 17165
rect 9195 17116 9196 17156
rect 9236 17116 9237 17156
rect 9195 17107 9237 17116
rect 9196 17072 9236 17107
rect 9196 17021 9236 17032
rect 9388 16904 9428 17704
rect 9484 17165 9524 20971
rect 9579 20768 9621 20777
rect 9579 20728 9580 20768
rect 9620 20728 9621 20768
rect 9579 20719 9621 20728
rect 9580 20634 9620 20719
rect 9579 18668 9621 18677
rect 9579 18628 9580 18668
rect 9620 18628 9621 18668
rect 9579 18619 9621 18628
rect 9483 17156 9525 17165
rect 9483 17116 9484 17156
rect 9524 17116 9525 17156
rect 9483 17107 9525 17116
rect 9196 16864 9428 16904
rect 8372 16192 8564 16232
rect 8332 16183 8372 16192
rect 8428 15728 8468 15737
rect 8236 15688 8428 15728
rect 8428 15679 8468 15688
rect 8236 15560 8276 15571
rect 8236 15485 8276 15520
rect 8235 15476 8277 15485
rect 8235 15436 8236 15476
rect 8276 15436 8277 15476
rect 8235 15427 8277 15436
rect 8427 14972 8469 14981
rect 8427 14932 8428 14972
rect 8468 14932 8469 14972
rect 8427 14923 8469 14932
rect 8428 14729 8468 14923
rect 8427 14720 8469 14729
rect 8427 14680 8428 14720
rect 8468 14680 8469 14720
rect 8427 14671 8469 14680
rect 8427 14216 8469 14225
rect 8427 14176 8428 14216
rect 8468 14176 8469 14216
rect 8427 14167 8469 14176
rect 8331 14048 8373 14057
rect 8331 14008 8332 14048
rect 8372 14008 8373 14048
rect 8331 13999 8373 14008
rect 8235 13208 8277 13217
rect 8235 13168 8236 13208
rect 8276 13168 8277 13208
rect 8235 13159 8277 13168
rect 8236 12620 8276 13159
rect 8236 12571 8276 12580
rect 8139 11864 8181 11873
rect 8139 11824 8140 11864
rect 8180 11824 8181 11864
rect 8139 11815 8181 11824
rect 8139 11696 8181 11705
rect 8139 11656 8140 11696
rect 8180 11656 8181 11696
rect 8139 11647 8181 11656
rect 8043 11444 8085 11453
rect 8043 11404 8044 11444
rect 8084 11404 8085 11444
rect 8043 11395 8085 11404
rect 8043 11024 8085 11033
rect 8043 10984 8044 11024
rect 8084 10984 8085 11024
rect 8043 10975 8085 10984
rect 7948 8707 7988 8716
rect 8044 8177 8084 10975
rect 8043 8168 8085 8177
rect 8043 8128 8044 8168
rect 8084 8128 8085 8168
rect 8043 8119 8085 8128
rect 8044 7916 8084 7925
rect 7700 7876 7796 7916
rect 7852 7876 7988 7916
rect 7660 7867 7700 7876
rect 7659 7160 7701 7169
rect 7659 7120 7660 7160
rect 7700 7120 7701 7160
rect 7659 7111 7701 7120
rect 7660 6749 7700 7111
rect 7659 6740 7701 6749
rect 7659 6700 7660 6740
rect 7700 6700 7701 6740
rect 7659 6691 7701 6700
rect 7660 6488 7700 6497
rect 7660 6329 7700 6448
rect 7659 6320 7701 6329
rect 7659 6280 7660 6320
rect 7700 6280 7701 6320
rect 7659 6271 7701 6280
rect 7659 6068 7701 6077
rect 7659 6028 7660 6068
rect 7700 6028 7701 6068
rect 7659 6019 7701 6028
rect 7371 4892 7413 4901
rect 7371 4852 7372 4892
rect 7412 4852 7413 4892
rect 7371 4843 7413 4852
rect 7564 4817 7604 4936
rect 7563 4808 7605 4817
rect 7563 4768 7564 4808
rect 7604 4768 7605 4808
rect 7563 4759 7605 4768
rect 7276 4684 7412 4724
rect 7275 4556 7317 4565
rect 7275 4516 7276 4556
rect 7316 4516 7317 4556
rect 7275 4507 7317 4516
rect 6988 2416 7220 2456
rect 6988 2372 7028 2416
rect 6740 1240 6836 1280
rect 6892 2332 7028 2372
rect 6700 1231 6740 1240
rect 6508 785 6548 1072
rect 6795 1112 6837 1121
rect 6795 1072 6796 1112
rect 6836 1072 6837 1112
rect 6795 1063 6837 1072
rect 6507 776 6549 785
rect 6507 736 6508 776
rect 6548 736 6549 776
rect 6507 727 6549 736
rect 6603 692 6645 701
rect 6603 652 6604 692
rect 6644 652 6645 692
rect 6603 643 6645 652
rect 6604 80 6644 643
rect 6796 80 6836 1063
rect 6892 617 6932 2332
rect 7083 2288 7125 2297
rect 7083 2248 7084 2288
rect 7124 2248 7125 2288
rect 7083 2239 7125 2248
rect 6987 2204 7029 2213
rect 6987 2164 6988 2204
rect 7028 2164 7029 2204
rect 6987 2155 7029 2164
rect 6988 2120 7028 2155
rect 6988 1280 7028 2080
rect 6988 1231 7028 1240
rect 7084 944 7124 2239
rect 7180 1952 7220 1961
rect 7180 1793 7220 1912
rect 7179 1784 7221 1793
rect 7179 1744 7180 1784
rect 7220 1744 7221 1784
rect 7179 1735 7221 1744
rect 7180 1112 7220 1121
rect 7276 1112 7316 4507
rect 7220 1072 7316 1112
rect 7180 1063 7220 1072
rect 7084 904 7220 944
rect 6891 608 6933 617
rect 6891 568 6892 608
rect 6932 568 6933 608
rect 6891 559 6933 568
rect 6987 356 7029 365
rect 6987 316 6988 356
rect 7028 316 7029 356
rect 6987 307 7029 316
rect 6988 80 7028 307
rect 7180 80 7220 904
rect 7372 80 7412 4684
rect 7563 4136 7605 4145
rect 7563 4096 7564 4136
rect 7604 4096 7605 4136
rect 7563 4087 7605 4096
rect 7467 3716 7509 3725
rect 7467 3676 7468 3716
rect 7508 3676 7509 3716
rect 7467 3667 7509 3676
rect 7468 3473 7508 3667
rect 7467 3464 7509 3473
rect 7467 3424 7468 3464
rect 7508 3424 7509 3464
rect 7467 3415 7509 3424
rect 7468 3330 7508 3415
rect 7564 3296 7604 4087
rect 7660 3473 7700 6019
rect 7756 3977 7796 7876
rect 7852 7748 7892 7757
rect 7852 7085 7892 7708
rect 7948 7337 7988 7876
rect 8044 7757 8084 7876
rect 8043 7748 8085 7757
rect 8043 7708 8044 7748
rect 8084 7708 8085 7748
rect 8043 7699 8085 7708
rect 7947 7328 7989 7337
rect 7947 7288 7948 7328
rect 7988 7288 7989 7328
rect 7947 7279 7989 7288
rect 7947 7160 7989 7169
rect 7947 7120 7948 7160
rect 7988 7120 7989 7160
rect 7947 7111 7989 7120
rect 8044 7160 8084 7171
rect 7851 7076 7893 7085
rect 7851 7036 7852 7076
rect 7892 7036 7893 7076
rect 7851 7027 7893 7036
rect 7948 7026 7988 7111
rect 8044 7085 8084 7120
rect 8043 7076 8085 7085
rect 8043 7036 8044 7076
rect 8084 7036 8085 7076
rect 8043 7027 8085 7036
rect 7851 6740 7893 6749
rect 7851 6700 7852 6740
rect 7892 6700 7893 6740
rect 7851 6691 7893 6700
rect 7852 5648 7892 6691
rect 7947 6320 7989 6329
rect 7947 6280 7948 6320
rect 7988 6280 7989 6320
rect 7947 6271 7989 6280
rect 7755 3968 7797 3977
rect 7755 3928 7756 3968
rect 7796 3928 7797 3968
rect 7755 3919 7797 3928
rect 7659 3464 7701 3473
rect 7659 3424 7660 3464
rect 7700 3424 7701 3464
rect 7659 3415 7701 3424
rect 7755 3380 7797 3389
rect 7755 3340 7756 3380
rect 7796 3340 7797 3380
rect 7755 3331 7797 3340
rect 7564 3256 7700 3296
rect 7563 2708 7605 2717
rect 7563 2668 7564 2708
rect 7604 2668 7605 2708
rect 7563 2659 7605 2668
rect 7468 2624 7508 2633
rect 7468 1373 7508 2584
rect 7564 2574 7604 2659
rect 7467 1364 7509 1373
rect 7467 1324 7468 1364
rect 7508 1324 7509 1364
rect 7467 1315 7509 1324
rect 7660 1205 7700 3256
rect 7756 3246 7796 3331
rect 7852 3221 7892 5608
rect 7948 4649 7988 6271
rect 8044 5741 8084 7027
rect 8140 6833 8180 11647
rect 8332 8345 8372 13999
rect 8428 11024 8468 14167
rect 8524 14057 8564 16192
rect 8715 16232 8757 16241
rect 8715 16192 8716 16232
rect 8756 16192 8757 16232
rect 8715 16183 8757 16192
rect 8812 16232 8852 16241
rect 8619 15392 8661 15401
rect 8619 15352 8620 15392
rect 8660 15352 8661 15392
rect 8619 15343 8661 15352
rect 8620 14897 8660 15343
rect 8619 14888 8661 14897
rect 8619 14848 8620 14888
rect 8660 14848 8661 14888
rect 8619 14839 8661 14848
rect 8716 14216 8756 16183
rect 8812 16148 8852 16192
rect 9099 16232 9141 16241
rect 9099 16192 9100 16232
rect 9140 16192 9141 16232
rect 9099 16183 9141 16192
rect 8812 16108 9044 16148
rect 9004 16064 9044 16108
rect 9196 16064 9236 16864
rect 9387 16736 9429 16745
rect 9387 16696 9388 16736
rect 9428 16696 9429 16736
rect 9387 16687 9429 16696
rect 9291 16652 9333 16661
rect 9291 16612 9292 16652
rect 9332 16612 9333 16652
rect 9291 16603 9333 16612
rect 9004 16024 9236 16064
rect 8907 15980 8949 15989
rect 8907 15940 8908 15980
rect 8948 15940 8949 15980
rect 8907 15931 8949 15940
rect 8812 15560 8852 15569
rect 8812 15401 8852 15520
rect 8811 15392 8853 15401
rect 8811 15352 8812 15392
rect 8852 15352 8853 15392
rect 8811 15343 8853 15352
rect 8716 14176 8852 14216
rect 8523 14048 8565 14057
rect 8523 14008 8524 14048
rect 8564 14008 8565 14048
rect 8523 13999 8565 14008
rect 8620 14048 8660 14057
rect 8620 13637 8660 14008
rect 8715 14048 8757 14057
rect 8715 14008 8716 14048
rect 8756 14008 8757 14048
rect 8715 13999 8757 14008
rect 8716 13914 8756 13999
rect 8812 13796 8852 14176
rect 8716 13756 8852 13796
rect 8619 13628 8661 13637
rect 8619 13588 8620 13628
rect 8660 13588 8661 13628
rect 8619 13579 8661 13588
rect 8716 13460 8756 13756
rect 8908 13721 8948 15931
rect 9099 14132 9141 14141
rect 9099 14092 9100 14132
rect 9140 14092 9141 14132
rect 9099 14083 9141 14092
rect 9100 14048 9140 14083
rect 9100 13997 9140 14008
rect 9196 14048 9236 16024
rect 9196 13999 9236 14008
rect 9292 16232 9332 16603
rect 9292 13880 9332 16192
rect 9004 13840 9332 13880
rect 8907 13712 8949 13721
rect 8907 13672 8908 13712
rect 8948 13672 8949 13712
rect 8907 13663 8949 13672
rect 8811 13628 8853 13637
rect 8811 13588 8812 13628
rect 8852 13588 8853 13628
rect 8811 13579 8853 13588
rect 8524 13420 8756 13460
rect 8812 13460 8852 13579
rect 8908 13460 8948 13469
rect 8812 13420 8908 13460
rect 8524 12032 8564 13420
rect 8908 13411 8948 13420
rect 8716 13208 8756 13217
rect 8716 12629 8756 13168
rect 8715 12620 8757 12629
rect 8715 12580 8716 12620
rect 8756 12580 8757 12620
rect 8715 12571 8757 12580
rect 8716 12293 8756 12571
rect 8812 12536 8852 12545
rect 8715 12284 8757 12293
rect 8715 12244 8716 12284
rect 8756 12244 8757 12284
rect 8715 12235 8757 12244
rect 8524 11992 8660 12032
rect 8620 11705 8660 11992
rect 8715 11864 8757 11873
rect 8715 11824 8716 11864
rect 8756 11824 8757 11864
rect 8715 11815 8757 11824
rect 8524 11696 8564 11705
rect 8524 11360 8564 11656
rect 8619 11696 8661 11705
rect 8619 11656 8620 11696
rect 8660 11656 8661 11696
rect 8619 11647 8661 11656
rect 8620 11562 8660 11647
rect 8524 11320 8660 11360
rect 8523 11024 8565 11033
rect 8428 10984 8524 11024
rect 8564 10984 8565 11024
rect 8523 10975 8565 10984
rect 8427 10688 8469 10697
rect 8427 10648 8428 10688
rect 8468 10648 8469 10688
rect 8427 10639 8469 10648
rect 8428 8672 8468 10639
rect 8524 10613 8564 10975
rect 8523 10604 8565 10613
rect 8523 10564 8524 10604
rect 8564 10564 8565 10604
rect 8523 10555 8565 10564
rect 8620 9680 8660 11320
rect 8716 10184 8756 11815
rect 8716 9848 8756 10144
rect 8812 10025 8852 12496
rect 8907 12368 8949 12377
rect 8907 12328 8908 12368
rect 8948 12328 8949 12368
rect 8907 12319 8949 12328
rect 8811 10016 8853 10025
rect 8811 9976 8812 10016
rect 8852 9976 8853 10016
rect 8811 9967 8853 9976
rect 8908 9941 8948 12319
rect 9004 11780 9044 13840
rect 9099 13376 9141 13385
rect 9099 13336 9100 13376
rect 9140 13336 9141 13376
rect 9099 13327 9141 13336
rect 9100 12881 9140 13327
rect 9388 13208 9428 16687
rect 9484 16325 9524 17107
rect 9483 16316 9525 16325
rect 9483 16276 9484 16316
rect 9524 16276 9525 16316
rect 9483 16267 9525 16276
rect 9580 15224 9620 18619
rect 9676 16232 9716 22912
rect 9771 20768 9813 20777
rect 9771 20728 9772 20768
rect 9812 20728 9813 20768
rect 9771 20719 9813 20728
rect 9772 19256 9812 20719
rect 9772 17744 9812 19216
rect 9868 18509 9908 23071
rect 9964 20861 10004 23911
rect 10059 23708 10101 23717
rect 10059 23668 10060 23708
rect 10100 23668 10101 23708
rect 10059 23659 10101 23668
rect 10060 23574 10100 23659
rect 10155 23624 10197 23633
rect 10155 23584 10156 23624
rect 10196 23584 10197 23624
rect 10155 23575 10197 23584
rect 10059 23120 10101 23129
rect 10059 23080 10060 23120
rect 10100 23080 10101 23120
rect 10059 23071 10101 23080
rect 10060 22986 10100 23071
rect 10156 22289 10196 23575
rect 10252 22541 10292 24172
rect 10348 23792 10388 24340
rect 10540 24221 10580 24592
rect 10731 24583 10773 24592
rect 10539 24212 10581 24221
rect 10539 24172 10540 24212
rect 10580 24172 10581 24212
rect 10539 24163 10581 24172
rect 10732 23969 10772 24583
rect 10828 24389 10868 25264
rect 10827 24380 10869 24389
rect 10827 24340 10828 24380
rect 10868 24340 10869 24380
rect 10827 24331 10869 24340
rect 10731 23960 10773 23969
rect 10924 23960 10964 26608
rect 11019 26480 11061 26489
rect 11019 26440 11020 26480
rect 11060 26440 11061 26480
rect 11019 26431 11061 26440
rect 11020 25481 11060 26431
rect 11019 25472 11061 25481
rect 11019 25432 11020 25472
rect 11060 25432 11061 25472
rect 11019 25423 11061 25432
rect 10731 23920 10732 23960
rect 10772 23920 10773 23960
rect 10731 23911 10773 23920
rect 10828 23920 10964 23960
rect 10444 23792 10484 23801
rect 10348 23752 10444 23792
rect 10444 23743 10484 23752
rect 10635 23792 10677 23801
rect 10635 23752 10636 23792
rect 10676 23752 10677 23792
rect 10635 23743 10677 23752
rect 10732 23792 10772 23911
rect 10732 23743 10772 23752
rect 10540 23624 10580 23633
rect 10540 23129 10580 23584
rect 10539 23120 10581 23129
rect 10539 23080 10540 23120
rect 10580 23080 10581 23120
rect 10539 23071 10581 23080
rect 10636 22793 10676 23743
rect 10635 22784 10677 22793
rect 10635 22744 10636 22784
rect 10676 22744 10677 22784
rect 10635 22735 10677 22744
rect 10251 22532 10293 22541
rect 10251 22492 10252 22532
rect 10292 22492 10293 22532
rect 10251 22483 10293 22492
rect 10155 22280 10197 22289
rect 10540 22280 10580 22289
rect 10828 22280 10868 23920
rect 10923 23792 10965 23801
rect 10923 23752 10924 23792
rect 10964 23752 10965 23792
rect 10923 23743 10965 23752
rect 10924 23658 10964 23743
rect 10155 22240 10156 22280
rect 10196 22240 10197 22280
rect 10155 22231 10197 22240
rect 10348 22240 10540 22280
rect 10580 22240 10868 22280
rect 9963 20852 10005 20861
rect 9963 20812 9964 20852
rect 10004 20812 10005 20852
rect 9963 20803 10005 20812
rect 10108 20777 10148 20786
rect 10148 20737 10196 20768
rect 10108 20728 10196 20737
rect 10156 20264 10196 20728
rect 10252 20693 10292 20778
rect 10251 20684 10293 20693
rect 10251 20644 10252 20684
rect 10292 20644 10293 20684
rect 10251 20635 10293 20644
rect 10251 20516 10293 20525
rect 10251 20476 10252 20516
rect 10292 20476 10293 20516
rect 10251 20467 10293 20476
rect 10156 20215 10196 20224
rect 9964 20096 10004 20105
rect 10252 20096 10292 20467
rect 9964 19013 10004 20056
rect 10156 20056 10292 20096
rect 10059 19424 10101 19433
rect 10059 19384 10060 19424
rect 10100 19384 10101 19424
rect 10059 19375 10101 19384
rect 9963 19004 10005 19013
rect 9963 18964 9964 19004
rect 10004 18964 10005 19004
rect 9963 18955 10005 18964
rect 9867 18500 9909 18509
rect 9867 18460 9868 18500
rect 9908 18460 9909 18500
rect 9867 18451 9909 18460
rect 9868 17744 9908 17753
rect 9772 17704 9868 17744
rect 9868 16661 9908 17704
rect 9963 16988 10005 16997
rect 9963 16948 9964 16988
rect 10004 16948 10005 16988
rect 9963 16939 10005 16948
rect 9867 16652 9909 16661
rect 9867 16612 9868 16652
rect 9908 16612 9909 16652
rect 9867 16603 9909 16612
rect 9964 16325 10004 16939
rect 9963 16316 10005 16325
rect 9963 16276 9964 16316
rect 10004 16276 10005 16316
rect 9963 16267 10005 16276
rect 9820 16241 9860 16250
rect 9676 16192 9727 16232
rect 9860 16201 9908 16232
rect 9820 16192 9908 16201
rect 9687 16148 9727 16192
rect 9687 16108 9812 16148
rect 9675 15980 9717 15989
rect 9675 15940 9676 15980
rect 9716 15940 9717 15980
rect 9675 15931 9717 15940
rect 9676 15485 9716 15931
rect 9675 15476 9717 15485
rect 9675 15436 9676 15476
rect 9716 15436 9717 15476
rect 9675 15427 9717 15436
rect 9484 15184 9620 15224
rect 9484 13385 9524 15184
rect 9676 14720 9716 15427
rect 9772 15401 9812 16108
rect 9771 15392 9813 15401
rect 9771 15352 9772 15392
rect 9812 15352 9813 15392
rect 9771 15343 9813 15352
rect 9771 15056 9813 15065
rect 9771 15016 9772 15056
rect 9812 15016 9813 15056
rect 9771 15007 9813 15016
rect 9676 14671 9716 14680
rect 9772 14552 9812 15007
rect 9868 14972 9908 16192
rect 9964 16148 10004 16267
rect 9964 16099 10004 16108
rect 10060 15896 10100 19375
rect 10156 17333 10196 20056
rect 10252 19265 10292 19270
rect 10251 19261 10293 19265
rect 10251 19216 10252 19261
rect 10292 19216 10293 19261
rect 10251 19207 10293 19216
rect 10252 19126 10292 19207
rect 10251 19004 10293 19013
rect 10251 18964 10252 19004
rect 10292 18964 10293 19004
rect 10251 18955 10293 18964
rect 10252 18845 10292 18955
rect 10251 18836 10293 18845
rect 10251 18796 10252 18836
rect 10292 18796 10293 18836
rect 10251 18787 10293 18796
rect 10252 18584 10292 18787
rect 10348 18761 10388 22240
rect 10540 22231 10580 22240
rect 10731 21608 10773 21617
rect 10731 21568 10732 21608
rect 10772 21568 10773 21608
rect 10731 21559 10773 21568
rect 10732 21474 10772 21559
rect 10924 21356 10964 21365
rect 10540 21316 10924 21356
rect 10540 20768 10580 21316
rect 10924 21307 10964 21316
rect 10731 21188 10773 21197
rect 11020 21188 11060 25423
rect 11115 24212 11157 24221
rect 11115 24172 11116 24212
rect 11156 24172 11157 24212
rect 11115 24163 11157 24172
rect 11116 24053 11156 24163
rect 11115 24044 11157 24053
rect 11115 24004 11116 24044
rect 11156 24004 11157 24044
rect 11115 23995 11157 24004
rect 10731 21148 10732 21188
rect 10772 21148 10773 21188
rect 10731 21139 10773 21148
rect 10924 21148 11060 21188
rect 10540 20719 10580 20728
rect 10636 20768 10676 20777
rect 10636 20525 10676 20728
rect 10635 20516 10677 20525
rect 10635 20476 10636 20516
rect 10676 20476 10677 20516
rect 10635 20467 10677 20476
rect 10732 19844 10772 21139
rect 10828 20096 10868 20105
rect 10828 20021 10868 20056
rect 10827 20012 10869 20021
rect 10827 19972 10828 20012
rect 10868 19972 10869 20012
rect 10827 19963 10869 19972
rect 10636 19804 10772 19844
rect 10539 19256 10581 19265
rect 10539 19216 10540 19256
rect 10580 19216 10581 19256
rect 10539 19207 10581 19216
rect 10444 19046 10484 19055
rect 10443 19006 10444 19013
rect 10484 19006 10485 19013
rect 10443 19004 10485 19006
rect 10443 18964 10444 19004
rect 10484 18964 10485 19004
rect 10443 18955 10485 18964
rect 10444 18911 10484 18955
rect 10347 18752 10389 18761
rect 10347 18712 10348 18752
rect 10388 18712 10389 18752
rect 10347 18703 10389 18712
rect 10540 18752 10580 19207
rect 10636 18752 10676 19804
rect 10828 19760 10868 19963
rect 10732 19720 10868 19760
rect 10732 18929 10772 19720
rect 10827 19592 10869 19601
rect 10827 19552 10828 19592
rect 10868 19552 10869 19592
rect 10827 19543 10869 19552
rect 10828 19256 10868 19543
rect 10828 19207 10868 19216
rect 10731 18920 10773 18929
rect 10731 18880 10732 18920
rect 10772 18880 10773 18920
rect 10731 18871 10773 18880
rect 10924 18836 10964 21148
rect 11116 21104 11156 23995
rect 11212 21281 11252 30463
rect 11404 29840 11444 30631
rect 11500 30605 11540 30640
rect 11499 30596 11541 30605
rect 11499 30556 11500 30596
rect 11540 30556 11541 30596
rect 11499 30547 11541 30556
rect 11596 30437 11636 32899
rect 11595 30428 11637 30437
rect 11595 30388 11596 30428
rect 11636 30388 11637 30428
rect 11595 30379 11637 30388
rect 11404 29791 11444 29800
rect 11596 29840 11636 29849
rect 11692 29840 11732 36427
rect 11636 29800 11732 29840
rect 11596 29791 11636 29800
rect 11308 29672 11348 29681
rect 11308 29345 11348 29632
rect 11307 29336 11349 29345
rect 11307 29296 11308 29336
rect 11348 29296 11349 29336
rect 11307 29287 11349 29296
rect 11320 29177 11360 29196
rect 11308 29168 11360 29177
rect 11403 29168 11445 29177
rect 11348 29128 11404 29168
rect 11444 29128 11445 29168
rect 11308 29119 11348 29128
rect 11403 29119 11445 29128
rect 11499 28076 11541 28085
rect 11499 28036 11500 28076
rect 11540 28036 11541 28076
rect 11499 28027 11541 28036
rect 11403 27908 11445 27917
rect 11403 27868 11404 27908
rect 11444 27868 11445 27908
rect 11403 27859 11445 27868
rect 11307 23540 11349 23549
rect 11307 23500 11308 23540
rect 11348 23500 11349 23540
rect 11307 23491 11349 23500
rect 11308 23120 11348 23491
rect 11308 23071 11348 23080
rect 11307 22784 11349 22793
rect 11307 22744 11308 22784
rect 11348 22744 11349 22784
rect 11307 22735 11349 22744
rect 11211 21272 11253 21281
rect 11211 21232 11212 21272
rect 11252 21232 11253 21272
rect 11211 21223 11253 21232
rect 11116 21064 11252 21104
rect 11115 20852 11157 20861
rect 11115 20812 11116 20852
rect 11156 20812 11157 20852
rect 11115 20803 11157 20812
rect 11019 20768 11061 20777
rect 11019 20728 11020 20768
rect 11060 20728 11061 20768
rect 11019 20719 11061 20728
rect 11020 20273 11060 20719
rect 11019 20264 11061 20273
rect 11019 20224 11020 20264
rect 11060 20224 11061 20264
rect 11019 20215 11061 20224
rect 10924 18796 11060 18836
rect 10827 18752 10869 18761
rect 10636 18712 10772 18752
rect 10540 18703 10580 18712
rect 10348 18584 10388 18593
rect 10252 18544 10348 18584
rect 10155 17324 10197 17333
rect 10155 17284 10156 17324
rect 10196 17284 10197 17324
rect 10155 17275 10197 17284
rect 10155 17072 10197 17081
rect 10155 17032 10156 17072
rect 10196 17032 10197 17072
rect 10155 17023 10197 17032
rect 10156 15989 10196 17023
rect 10252 16409 10292 18544
rect 10348 18535 10388 18544
rect 10396 17753 10436 17762
rect 10436 17713 10676 17744
rect 10396 17704 10676 17713
rect 10540 17576 10580 17585
rect 10443 17240 10485 17249
rect 10443 17200 10444 17240
rect 10484 17200 10485 17240
rect 10443 17191 10485 17200
rect 10444 17072 10484 17191
rect 10444 17023 10484 17032
rect 10251 16400 10293 16409
rect 10251 16360 10252 16400
rect 10292 16360 10293 16400
rect 10251 16351 10293 16360
rect 10252 16232 10292 16241
rect 10155 15980 10197 15989
rect 10155 15940 10156 15980
rect 10196 15940 10197 15980
rect 10155 15931 10197 15940
rect 9964 15856 10100 15896
rect 9964 14981 10004 15856
rect 10252 15728 10292 16192
rect 10252 15679 10292 15688
rect 10348 16232 10388 16241
rect 10348 15569 10388 16192
rect 10540 16157 10580 17536
rect 10636 17240 10676 17704
rect 10636 17191 10676 17200
rect 10732 17081 10772 18712
rect 10827 18712 10828 18752
rect 10868 18712 10869 18752
rect 10827 18703 10869 18712
rect 10731 17072 10773 17081
rect 10731 17032 10732 17072
rect 10772 17032 10773 17072
rect 10731 17023 10773 17032
rect 10828 16484 10868 18703
rect 10636 16444 10868 16484
rect 11020 18584 11060 18796
rect 10539 16148 10581 16157
rect 10539 16108 10540 16148
rect 10580 16108 10581 16148
rect 10539 16099 10581 16108
rect 10540 15905 10580 16099
rect 10539 15896 10581 15905
rect 10539 15856 10540 15896
rect 10580 15856 10581 15896
rect 10539 15847 10581 15856
rect 10059 15560 10101 15569
rect 10059 15520 10060 15560
rect 10100 15520 10101 15560
rect 10059 15511 10101 15520
rect 10347 15560 10389 15569
rect 10347 15520 10348 15560
rect 10388 15520 10389 15560
rect 10347 15511 10389 15520
rect 10060 15401 10100 15511
rect 10059 15392 10101 15401
rect 10059 15352 10060 15392
rect 10100 15352 10101 15392
rect 10059 15343 10101 15352
rect 9868 14923 9908 14932
rect 9963 14972 10005 14981
rect 9963 14932 9964 14972
rect 10004 14932 10005 14972
rect 9963 14923 10005 14932
rect 10636 14813 10676 16444
rect 10827 16316 10869 16325
rect 10827 16276 10828 16316
rect 10868 16276 10869 16316
rect 10827 16267 10869 16276
rect 10731 16232 10773 16241
rect 10731 16192 10732 16232
rect 10772 16192 10773 16232
rect 10731 16183 10773 16192
rect 10732 16098 10772 16183
rect 10828 16182 10868 16267
rect 11020 16064 11060 18544
rect 11116 17585 11156 20803
rect 11115 17576 11157 17585
rect 11115 17536 11116 17576
rect 11156 17536 11157 17576
rect 11115 17527 11157 17536
rect 11115 17408 11157 17417
rect 11115 17368 11116 17408
rect 11156 17368 11157 17408
rect 11115 17359 11157 17368
rect 10828 16024 11060 16064
rect 10731 15896 10773 15905
rect 10731 15856 10732 15896
rect 10772 15856 10773 15896
rect 10731 15847 10773 15856
rect 10635 14804 10677 14813
rect 10635 14764 10636 14804
rect 10676 14764 10677 14804
rect 10635 14755 10677 14764
rect 10539 14720 10581 14729
rect 10539 14680 10540 14720
rect 10580 14680 10581 14720
rect 10539 14671 10581 14680
rect 10540 14586 10580 14671
rect 9676 14512 9812 14552
rect 9676 14048 9716 14512
rect 10348 14132 10388 14141
rect 9676 13999 9716 14008
rect 10156 14034 10196 14043
rect 9483 13376 9525 13385
rect 9483 13336 9484 13376
rect 9524 13336 9525 13376
rect 9483 13327 9525 13336
rect 9484 13208 9524 13217
rect 9388 13168 9484 13208
rect 9099 12872 9141 12881
rect 9099 12832 9100 12872
rect 9140 12832 9141 12872
rect 9099 12823 9141 12832
rect 9004 11731 9044 11740
rect 9100 11780 9140 12823
rect 9484 11957 9524 13168
rect 9579 12788 9621 12797
rect 9579 12748 9580 12788
rect 9620 12748 9621 12788
rect 9579 12739 9621 12748
rect 9483 11948 9525 11957
rect 9483 11908 9484 11948
rect 9524 11908 9525 11948
rect 9483 11899 9525 11908
rect 9100 11731 9140 11740
rect 9195 11696 9237 11705
rect 9195 11656 9196 11696
rect 9236 11656 9237 11696
rect 9195 11647 9237 11656
rect 9580 11696 9620 12739
rect 10156 12704 10196 13994
rect 10348 13301 10388 14092
rect 10732 13880 10772 15847
rect 10636 13840 10772 13880
rect 10347 13292 10389 13301
rect 10347 13252 10348 13292
rect 10388 13252 10389 13292
rect 10347 13243 10389 13252
rect 10636 12965 10676 13840
rect 10731 13208 10773 13217
rect 10731 13168 10732 13208
rect 10772 13168 10773 13208
rect 10731 13159 10773 13168
rect 10635 12956 10677 12965
rect 10635 12916 10636 12956
rect 10676 12916 10677 12956
rect 10635 12907 10677 12916
rect 10252 12704 10292 12713
rect 10156 12664 10252 12704
rect 10252 12655 10292 12664
rect 10443 12704 10485 12713
rect 10443 12664 10444 12704
rect 10484 12664 10485 12704
rect 10443 12655 10485 12664
rect 10059 12620 10101 12629
rect 10059 12580 10060 12620
rect 10100 12580 10101 12620
rect 10059 12571 10101 12580
rect 10060 12536 10100 12571
rect 10444 12570 10484 12655
rect 10732 12629 10772 13159
rect 10731 12620 10773 12629
rect 10731 12580 10732 12620
rect 10772 12580 10773 12620
rect 10731 12571 10773 12580
rect 10060 12485 10100 12496
rect 10636 12452 10676 12461
rect 10348 12412 10636 12452
rect 9580 11647 9620 11656
rect 10060 11701 10100 11710
rect 9196 11360 9236 11647
rect 9867 11444 9909 11453
rect 9867 11404 9868 11444
rect 9908 11404 9909 11444
rect 9867 11395 9909 11404
rect 9196 11320 9428 11360
rect 9099 10016 9141 10025
rect 9099 9976 9100 10016
rect 9140 9976 9141 10016
rect 9099 9967 9141 9976
rect 8907 9932 8949 9941
rect 8907 9892 8908 9932
rect 8948 9892 8949 9932
rect 8907 9883 8949 9892
rect 8716 9808 8852 9848
rect 8716 9680 8756 9689
rect 8620 9640 8716 9680
rect 8716 9631 8756 9640
rect 8524 9512 8564 9521
rect 8812 9512 8852 9808
rect 8564 9472 8660 9512
rect 8524 9463 8564 9472
rect 8523 9260 8565 9269
rect 8523 9220 8524 9260
rect 8564 9220 8565 9260
rect 8523 9211 8565 9220
rect 8428 8623 8468 8632
rect 8524 8504 8564 9211
rect 8620 8849 8660 9472
rect 8716 9472 8852 9512
rect 8619 8840 8661 8849
rect 8619 8800 8620 8840
rect 8660 8800 8661 8840
rect 8619 8791 8661 8800
rect 8428 8464 8564 8504
rect 8331 8336 8373 8345
rect 8331 8296 8332 8336
rect 8372 8296 8373 8336
rect 8331 8287 8373 8296
rect 8235 8252 8277 8261
rect 8235 8212 8236 8252
rect 8276 8212 8277 8252
rect 8235 8203 8277 8212
rect 8236 8000 8276 8203
rect 8236 7951 8276 7960
rect 8331 7160 8373 7169
rect 8331 7120 8332 7160
rect 8372 7120 8373 7160
rect 8331 7111 8373 7120
rect 8428 7160 8468 8464
rect 8716 7505 8756 9472
rect 9100 9185 9140 9967
rect 9099 9176 9141 9185
rect 9099 9136 9100 9176
rect 9140 9136 9141 9176
rect 9099 9127 9141 9136
rect 8811 9092 8853 9101
rect 8811 9052 8812 9092
rect 8852 9052 8853 9092
rect 8811 9043 8853 9052
rect 8715 7496 8757 7505
rect 8715 7456 8716 7496
rect 8756 7456 8757 7496
rect 8715 7447 8757 7456
rect 8812 7412 8852 9043
rect 8956 8681 8996 8690
rect 9100 8681 9140 9127
rect 9099 8672 9141 8681
rect 8996 8641 9044 8672
rect 8956 8632 9044 8641
rect 9004 7496 9044 8632
rect 9099 8632 9100 8672
rect 9140 8632 9141 8672
rect 9099 8623 9141 8632
rect 9100 8504 9140 8513
rect 9140 8464 9332 8504
rect 9100 8455 9140 8464
rect 9004 7456 9140 7496
rect 8812 7372 8948 7412
rect 8811 7244 8853 7253
rect 8811 7204 8812 7244
rect 8852 7204 8853 7244
rect 8811 7195 8853 7204
rect 8139 6824 8181 6833
rect 8139 6784 8140 6824
rect 8180 6784 8181 6824
rect 8139 6775 8181 6784
rect 8235 6320 8277 6329
rect 8235 6280 8236 6320
rect 8276 6280 8277 6320
rect 8235 6271 8277 6280
rect 8043 5732 8085 5741
rect 8043 5692 8044 5732
rect 8084 5692 8085 5732
rect 8043 5683 8085 5692
rect 8043 4892 8085 4901
rect 8043 4852 8044 4892
rect 8084 4852 8085 4892
rect 8043 4843 8085 4852
rect 7947 4640 7989 4649
rect 7947 4600 7948 4640
rect 7988 4600 7989 4640
rect 7947 4591 7989 4600
rect 7851 3212 7893 3221
rect 7851 3172 7852 3212
rect 7892 3172 7893 3212
rect 7851 3163 7893 3172
rect 7948 3212 7988 3221
rect 8044 3212 8084 4843
rect 8236 4304 8276 6271
rect 8332 5909 8372 7111
rect 8331 5900 8373 5909
rect 8331 5860 8332 5900
rect 8372 5860 8373 5900
rect 8331 5851 8373 5860
rect 8140 4264 8276 4304
rect 8332 5653 8372 5662
rect 8428 5657 8468 7120
rect 8524 7160 8564 7169
rect 8564 7120 8660 7160
rect 8524 7111 8564 7120
rect 8523 6992 8565 7001
rect 8523 6952 8524 6992
rect 8564 6952 8565 6992
rect 8523 6943 8565 6952
rect 8140 4145 8180 4264
rect 8139 4136 8181 4145
rect 8139 4096 8140 4136
rect 8180 4096 8181 4136
rect 8139 4087 8181 4096
rect 8236 4136 8276 4145
rect 8236 3893 8276 4096
rect 8235 3884 8277 3893
rect 8235 3844 8236 3884
rect 8276 3844 8277 3884
rect 8235 3835 8277 3844
rect 8139 3800 8181 3809
rect 8139 3760 8140 3800
rect 8180 3760 8181 3800
rect 8139 3751 8181 3760
rect 8140 3380 8180 3751
rect 8332 3380 8372 5613
rect 8427 5648 8469 5657
rect 8427 5608 8428 5648
rect 8468 5608 8469 5648
rect 8427 5599 8469 5608
rect 8524 5564 8564 6943
rect 8524 5515 8564 5524
rect 8620 4397 8660 7120
rect 8812 7110 8852 7195
rect 8908 6824 8948 7372
rect 8812 6784 8948 6824
rect 9004 6992 9044 7001
rect 8812 6740 8852 6784
rect 8716 6700 8852 6740
rect 8716 6245 8756 6700
rect 8907 6656 8949 6665
rect 8907 6616 8908 6656
rect 8948 6616 8949 6656
rect 8907 6607 8949 6616
rect 8811 6572 8853 6581
rect 8811 6532 8812 6572
rect 8852 6532 8853 6572
rect 8811 6523 8853 6532
rect 8715 6236 8757 6245
rect 8715 6196 8716 6236
rect 8756 6196 8757 6236
rect 8715 6187 8757 6196
rect 8812 5144 8852 6523
rect 8908 6488 8948 6607
rect 8908 6439 8948 6448
rect 9004 6077 9044 6952
rect 9100 6656 9140 7456
rect 9100 6607 9140 6616
rect 9196 6992 9236 7001
rect 9099 6236 9141 6245
rect 9099 6196 9100 6236
rect 9140 6196 9141 6236
rect 9099 6187 9141 6196
rect 9003 6068 9045 6077
rect 9003 6028 9004 6068
rect 9044 6028 9045 6068
rect 9003 6019 9045 6028
rect 8907 5732 8949 5741
rect 8907 5692 8908 5732
rect 8948 5692 8949 5732
rect 8907 5683 8949 5692
rect 8908 5598 8948 5683
rect 9100 5648 9140 6187
rect 9196 5825 9236 6952
rect 9292 6656 9332 8464
rect 9388 7832 9428 11320
rect 9772 11024 9812 11033
rect 9580 10984 9772 11024
rect 9580 8681 9620 10984
rect 9772 10975 9812 10984
rect 9868 10184 9908 11395
rect 9964 11192 10004 11201
rect 10060 11192 10100 11661
rect 10252 11612 10292 11621
rect 10348 11612 10388 12412
rect 10636 12403 10676 12412
rect 10539 12284 10581 12293
rect 10539 12244 10540 12284
rect 10580 12244 10581 12284
rect 10539 12235 10581 12244
rect 10443 11948 10485 11957
rect 10443 11908 10444 11948
rect 10484 11908 10485 11948
rect 10443 11899 10485 11908
rect 10292 11572 10388 11612
rect 10252 11563 10292 11572
rect 10004 11152 10100 11192
rect 9964 11143 10004 11152
rect 10252 11024 10292 11033
rect 10156 10436 10196 10445
rect 10252 10436 10292 10984
rect 10196 10396 10292 10436
rect 10348 11024 10388 11033
rect 10156 10387 10196 10396
rect 9964 10184 10004 10193
rect 9868 10144 9964 10184
rect 9964 10135 10004 10144
rect 10155 9680 10197 9689
rect 10155 9640 10156 9680
rect 10196 9640 10197 9680
rect 10155 9631 10197 9640
rect 9964 9512 10004 9521
rect 9676 9472 9964 9512
rect 9579 8672 9621 8681
rect 9484 8632 9580 8672
rect 9620 8632 9621 8672
rect 9484 8000 9524 8632
rect 9579 8623 9621 8632
rect 9579 8504 9621 8513
rect 9579 8464 9580 8504
rect 9620 8464 9621 8504
rect 9579 8455 9621 8464
rect 9484 7951 9524 7960
rect 9388 7792 9524 7832
rect 9388 7244 9428 7253
rect 9388 7001 9428 7204
rect 9387 6992 9429 7001
rect 9387 6952 9388 6992
rect 9428 6952 9429 6992
rect 9387 6943 9429 6952
rect 9292 6616 9428 6656
rect 9292 6488 9332 6497
rect 9292 6161 9332 6448
rect 9291 6152 9333 6161
rect 9291 6112 9292 6152
rect 9332 6112 9333 6152
rect 9291 6103 9333 6112
rect 9291 5900 9333 5909
rect 9291 5860 9292 5900
rect 9332 5860 9333 5900
rect 9291 5851 9333 5860
rect 9195 5816 9237 5825
rect 9195 5776 9196 5816
rect 9236 5776 9237 5816
rect 9195 5767 9237 5776
rect 9292 5816 9332 5851
rect 9292 5765 9332 5776
rect 9100 5608 9332 5648
rect 9100 5480 9140 5489
rect 9003 5144 9045 5153
rect 8812 5104 8948 5144
rect 8811 4976 8853 4985
rect 8811 4936 8812 4976
rect 8852 4936 8853 4976
rect 8811 4927 8853 4936
rect 8812 4842 8852 4927
rect 8619 4388 8661 4397
rect 8619 4348 8620 4388
rect 8660 4348 8661 4388
rect 8619 4339 8661 4348
rect 8764 4145 8804 4154
rect 8524 4105 8764 4136
rect 8524 4096 8804 4105
rect 8428 4052 8468 4061
rect 8524 4052 8564 4096
rect 8908 4052 8948 5104
rect 9003 5104 9004 5144
rect 9044 5104 9045 5144
rect 9003 5095 9045 5104
rect 9004 5010 9044 5095
rect 8468 4012 8564 4052
rect 8812 4012 8948 4052
rect 8428 4003 8468 4012
rect 8619 3968 8661 3977
rect 8619 3928 8620 3968
rect 8660 3928 8661 3968
rect 8619 3919 8661 3928
rect 8620 3834 8660 3919
rect 8715 3548 8757 3557
rect 8715 3508 8716 3548
rect 8756 3508 8757 3548
rect 8715 3499 8757 3508
rect 8620 3464 8660 3473
rect 8620 3380 8660 3424
rect 8716 3464 8756 3499
rect 8716 3413 8756 3424
rect 8140 3331 8180 3340
rect 8236 3340 8372 3380
rect 8428 3340 8660 3380
rect 8044 3172 8180 3212
rect 7755 3128 7797 3137
rect 7755 3088 7756 3128
rect 7796 3088 7797 3128
rect 7755 3079 7797 3088
rect 7659 1196 7701 1205
rect 7659 1156 7660 1196
rect 7700 1156 7701 1196
rect 7659 1147 7701 1156
rect 7563 1028 7605 1037
rect 7563 988 7564 1028
rect 7604 988 7605 1028
rect 7563 979 7605 988
rect 7564 80 7604 979
rect 7756 80 7796 3079
rect 7948 1289 7988 3172
rect 8044 2624 8084 2633
rect 8044 2549 8084 2584
rect 8043 2540 8085 2549
rect 8043 2500 8044 2540
rect 8084 2500 8085 2540
rect 8043 2491 8085 2500
rect 8044 2213 8084 2491
rect 8043 2204 8085 2213
rect 8043 2164 8044 2204
rect 8084 2164 8085 2204
rect 8043 2155 8085 2164
rect 7947 1280 7989 1289
rect 7947 1240 7948 1280
rect 7988 1240 7989 1280
rect 7947 1231 7989 1240
rect 7947 104 7989 113
rect 7947 80 7948 104
rect 1784 0 1864 80
rect 1976 0 2056 80
rect 2168 0 2248 80
rect 2360 0 2440 80
rect 2552 0 2632 80
rect 2744 0 2824 80
rect 2936 0 3016 80
rect 3128 0 3208 80
rect 3320 0 3400 80
rect 3512 0 3592 80
rect 3704 0 3784 80
rect 3896 0 3976 80
rect 4088 0 4168 80
rect 4280 0 4360 80
rect 4472 0 4552 80
rect 4664 0 4744 80
rect 4856 0 4936 80
rect 5048 0 5128 80
rect 5240 0 5320 80
rect 5432 0 5512 80
rect 5624 0 5704 80
rect 5816 0 5896 80
rect 6008 0 6088 80
rect 6200 0 6280 80
rect 6392 0 6472 80
rect 6584 0 6664 80
rect 6776 0 6856 80
rect 6968 0 7048 80
rect 7160 0 7240 80
rect 7352 0 7432 80
rect 7544 0 7624 80
rect 7736 0 7816 80
rect 7928 64 7948 80
rect 7988 80 7989 104
rect 8140 80 8180 3172
rect 8236 2549 8276 3340
rect 8331 3212 8373 3221
rect 8331 3172 8332 3212
rect 8372 3172 8373 3212
rect 8331 3163 8373 3172
rect 8332 3078 8372 3163
rect 8235 2540 8277 2549
rect 8235 2500 8236 2540
rect 8276 2500 8277 2540
rect 8235 2491 8277 2500
rect 8235 2372 8277 2381
rect 8235 2332 8236 2372
rect 8276 2332 8277 2372
rect 8235 2323 8277 2332
rect 8236 1280 8276 2323
rect 8428 2129 8468 3340
rect 8715 3128 8757 3137
rect 8715 3088 8716 3128
rect 8756 3088 8757 3128
rect 8715 3079 8757 3088
rect 8523 2792 8565 2801
rect 8523 2752 8524 2792
rect 8564 2752 8565 2792
rect 8523 2743 8565 2752
rect 8524 2638 8564 2743
rect 8524 2589 8564 2598
rect 8619 2540 8661 2549
rect 8619 2500 8620 2540
rect 8660 2500 8661 2540
rect 8619 2491 8661 2500
rect 8716 2540 8756 3079
rect 8716 2491 8756 2500
rect 8523 2204 8565 2213
rect 8523 2164 8524 2204
rect 8564 2164 8565 2204
rect 8523 2155 8565 2164
rect 8427 2120 8469 2129
rect 8427 2080 8428 2120
rect 8468 2080 8469 2120
rect 8427 2071 8469 2080
rect 8428 1952 8468 1961
rect 8524 1952 8564 2155
rect 8620 2120 8660 2491
rect 8812 2204 8852 4012
rect 9100 3968 9140 5440
rect 9292 5312 9332 5608
rect 9388 5489 9428 6616
rect 9484 6161 9524 7792
rect 9580 7580 9620 8455
rect 9676 8168 9716 9472
rect 9964 9463 10004 9472
rect 10060 9512 10100 9521
rect 9867 9344 9909 9353
rect 9867 9304 9868 9344
rect 9908 9304 9909 9344
rect 9867 9295 9909 9304
rect 9676 8119 9716 8128
rect 9868 8168 9908 9295
rect 10060 9269 10100 9472
rect 10059 9260 10101 9269
rect 10059 9220 10060 9260
rect 10100 9220 10101 9260
rect 10059 9211 10101 9220
rect 9868 8119 9908 8128
rect 10060 8009 10100 8090
rect 10059 8000 10101 8009
rect 10059 7955 10060 8000
rect 10100 7955 10101 8000
rect 10059 7951 10101 7955
rect 10060 7946 10100 7951
rect 10059 7664 10101 7673
rect 10059 7624 10060 7664
rect 10100 7624 10101 7664
rect 10059 7615 10101 7624
rect 9580 7540 9716 7580
rect 9579 7412 9621 7421
rect 9579 7372 9580 7412
rect 9620 7372 9621 7412
rect 9579 7363 9621 7372
rect 9580 7278 9620 7363
rect 9483 6152 9525 6161
rect 9483 6112 9484 6152
rect 9524 6112 9525 6152
rect 9483 6103 9525 6112
rect 9676 5816 9716 7540
rect 9772 7244 9812 7253
rect 9772 6068 9812 7204
rect 9772 6028 10004 6068
rect 9771 5900 9813 5909
rect 9771 5860 9772 5900
rect 9812 5860 9813 5900
rect 9771 5851 9813 5860
rect 9484 5776 9716 5816
rect 9387 5480 9429 5489
rect 9387 5440 9388 5480
rect 9428 5440 9429 5480
rect 9387 5431 9429 5440
rect 9292 5272 9428 5312
rect 9291 5060 9333 5069
rect 9291 5020 9292 5060
rect 9332 5020 9333 5060
rect 9291 5011 9333 5020
rect 9196 4976 9236 4985
rect 9196 4397 9236 4936
rect 9195 4388 9237 4397
rect 9195 4348 9196 4388
rect 9236 4348 9237 4388
rect 9195 4339 9237 4348
rect 9195 4220 9237 4229
rect 9195 4180 9196 4220
rect 9236 4180 9237 4220
rect 9195 4171 9237 4180
rect 9004 3928 9140 3968
rect 8907 2708 8949 2717
rect 8907 2668 8908 2708
rect 8948 2668 8949 2708
rect 8907 2659 8949 2668
rect 8908 2574 8948 2659
rect 8812 2164 8948 2204
rect 8620 2071 8660 2080
rect 8811 2036 8853 2045
rect 8811 1996 8812 2036
rect 8852 1996 8853 2036
rect 8811 1987 8853 1996
rect 8468 1912 8564 1952
rect 8428 1541 8468 1912
rect 8812 1902 8852 1987
rect 8908 1541 8948 2164
rect 9004 1700 9044 3928
rect 9196 3884 9236 4171
rect 9100 3844 9236 3884
rect 9292 4136 9332 5011
rect 9100 3464 9140 3844
rect 9292 3809 9332 4096
rect 9291 3800 9333 3809
rect 9291 3760 9292 3800
rect 9332 3760 9333 3800
rect 9291 3751 9333 3760
rect 9100 3415 9140 3424
rect 9291 3464 9333 3473
rect 9291 3424 9292 3464
rect 9332 3424 9333 3464
rect 9291 3415 9333 3424
rect 9195 3380 9237 3389
rect 9195 3340 9196 3380
rect 9236 3340 9237 3380
rect 9195 3331 9237 3340
rect 9196 3246 9236 3331
rect 9100 2792 9140 2801
rect 9100 2633 9140 2752
rect 9292 2708 9332 3415
rect 9292 2659 9332 2668
rect 9099 2624 9141 2633
rect 9099 2584 9100 2624
rect 9140 2584 9141 2624
rect 9099 2575 9141 2584
rect 9100 1877 9140 1962
rect 9099 1868 9141 1877
rect 9099 1828 9100 1868
rect 9140 1828 9141 1868
rect 9099 1819 9141 1828
rect 9291 1700 9333 1709
rect 9004 1660 9140 1700
rect 8427 1532 8469 1541
rect 8427 1492 8428 1532
rect 8468 1492 8469 1532
rect 8427 1483 8469 1492
rect 8907 1532 8949 1541
rect 8907 1492 8908 1532
rect 8948 1492 8949 1532
rect 8907 1483 8949 1492
rect 8620 1280 8660 1291
rect 8236 1240 8372 1280
rect 8332 80 8372 1240
rect 8620 1205 8660 1240
rect 8907 1280 8949 1289
rect 8907 1240 8908 1280
rect 8948 1240 8949 1280
rect 8907 1231 8949 1240
rect 8619 1196 8661 1205
rect 8619 1156 8620 1196
rect 8660 1156 8661 1196
rect 8619 1147 8661 1156
rect 8427 1112 8469 1121
rect 8427 1072 8428 1112
rect 8468 1072 8469 1112
rect 8427 1063 8469 1072
rect 8715 1112 8757 1121
rect 8715 1072 8716 1112
rect 8756 1072 8757 1112
rect 8715 1063 8757 1072
rect 8812 1112 8852 1121
rect 8428 533 8468 1063
rect 8427 524 8469 533
rect 8427 484 8428 524
rect 8468 484 8469 524
rect 8427 475 8469 484
rect 8523 272 8565 281
rect 8523 232 8524 272
rect 8564 232 8565 272
rect 8523 223 8565 232
rect 8524 80 8564 223
rect 8716 80 8756 1063
rect 8812 869 8852 1072
rect 8811 860 8853 869
rect 8811 820 8812 860
rect 8852 820 8853 860
rect 8811 811 8853 820
rect 8908 80 8948 1231
rect 9100 80 9140 1660
rect 9291 1660 9292 1700
rect 9332 1660 9333 1700
rect 9291 1651 9333 1660
rect 9292 1566 9332 1651
rect 9388 1037 9428 5272
rect 9484 3212 9524 5776
rect 9676 5648 9716 5657
rect 9676 5153 9716 5608
rect 9772 5648 9812 5851
rect 9772 5321 9812 5608
rect 9771 5312 9813 5321
rect 9771 5272 9772 5312
rect 9812 5272 9813 5312
rect 9771 5263 9813 5272
rect 9675 5144 9717 5153
rect 9675 5104 9676 5144
rect 9716 5104 9717 5144
rect 9675 5095 9717 5104
rect 9772 4220 9812 4229
rect 9580 4180 9772 4220
rect 9580 3389 9620 4180
rect 9772 4171 9812 4180
rect 9867 4220 9909 4229
rect 9867 4180 9868 4220
rect 9908 4180 9909 4220
rect 9867 4171 9909 4180
rect 9868 4086 9908 4171
rect 9964 3968 10004 6028
rect 9772 3928 10004 3968
rect 9675 3800 9717 3809
rect 9675 3760 9676 3800
rect 9716 3760 9717 3800
rect 9675 3751 9717 3760
rect 9676 3464 9716 3751
rect 9676 3415 9716 3424
rect 9579 3380 9621 3389
rect 9579 3340 9580 3380
rect 9620 3340 9621 3380
rect 9579 3331 9621 3340
rect 9484 3172 9620 3212
rect 9483 2876 9525 2885
rect 9483 2836 9484 2876
rect 9524 2836 9525 2876
rect 9483 2827 9525 2836
rect 9484 2742 9524 2827
rect 9484 1877 9524 1962
rect 9483 1868 9525 1877
rect 9483 1828 9484 1868
rect 9524 1828 9525 1868
rect 9483 1819 9525 1828
rect 9580 1700 9620 3172
rect 9675 2708 9717 2717
rect 9675 2668 9676 2708
rect 9716 2668 9717 2708
rect 9675 2659 9717 2668
rect 9676 2574 9716 2659
rect 9772 2381 9812 3928
rect 10060 3884 10100 7615
rect 10156 5993 10196 9631
rect 10348 9269 10388 10984
rect 10444 9428 10484 11899
rect 10540 11705 10580 12235
rect 10539 11696 10581 11705
rect 10539 11656 10540 11696
rect 10580 11656 10581 11696
rect 10539 11647 10581 11656
rect 10540 11562 10580 11647
rect 10828 11360 10868 16024
rect 11116 15905 11156 17359
rect 11115 15896 11157 15905
rect 11115 15856 11116 15896
rect 11156 15856 11157 15896
rect 11115 15847 11157 15856
rect 11020 15560 11060 15569
rect 11020 15317 11060 15520
rect 11115 15560 11157 15569
rect 11115 15520 11116 15560
rect 11156 15520 11157 15560
rect 11115 15511 11157 15520
rect 11019 15308 11061 15317
rect 11019 15268 11020 15308
rect 11060 15268 11061 15308
rect 11019 15259 11061 15268
rect 11116 15140 11156 15511
rect 11020 15100 11156 15140
rect 10923 14048 10965 14057
rect 10923 14008 10924 14048
rect 10964 14008 10965 14048
rect 10923 13999 10965 14008
rect 10924 13460 10964 13999
rect 10924 13411 10964 13420
rect 11020 13292 11060 15100
rect 11212 14468 11252 21064
rect 11308 20777 11348 22735
rect 11307 20768 11349 20777
rect 11307 20728 11308 20768
rect 11348 20728 11349 20768
rect 11307 20719 11349 20728
rect 11404 20180 11444 27859
rect 11500 27656 11540 28027
rect 11596 27665 11636 27750
rect 11500 27607 11540 27616
rect 11595 27656 11637 27665
rect 11595 27616 11596 27656
rect 11636 27616 11637 27656
rect 11595 27607 11637 27616
rect 11499 27488 11541 27497
rect 11692 27488 11732 29800
rect 11788 29093 11828 36763
rect 11980 36737 12020 37192
rect 11979 36728 12021 36737
rect 11979 36688 11980 36728
rect 12020 36688 12021 36728
rect 11979 36679 12021 36688
rect 12076 36728 12116 37360
rect 12076 35141 12116 36688
rect 12075 35132 12117 35141
rect 12075 35092 12076 35132
rect 12116 35092 12117 35132
rect 12075 35083 12117 35092
rect 11980 33704 12020 33713
rect 11884 33664 11980 33704
rect 11787 29084 11829 29093
rect 11787 29044 11788 29084
rect 11828 29044 11829 29084
rect 11787 29035 11829 29044
rect 11884 29000 11924 33664
rect 11980 33655 12020 33664
rect 12172 33368 12212 44416
rect 12268 39425 12308 46432
rect 12652 46472 12692 46481
rect 12364 46388 12404 46397
rect 12652 46388 12692 46432
rect 12404 46348 12692 46388
rect 12748 46472 12788 46600
rect 12364 46339 12404 46348
rect 12555 46220 12597 46229
rect 12555 46180 12556 46220
rect 12596 46180 12597 46220
rect 12555 46171 12597 46180
rect 12556 44288 12596 46171
rect 12651 44792 12693 44801
rect 12651 44752 12652 44792
rect 12692 44752 12693 44792
rect 12651 44743 12693 44752
rect 12556 44239 12596 44248
rect 12652 44213 12692 44743
rect 12748 44297 12788 46432
rect 12747 44288 12789 44297
rect 12747 44248 12748 44288
rect 12788 44248 12789 44288
rect 12747 44239 12789 44248
rect 12459 44204 12501 44213
rect 12459 44164 12460 44204
rect 12500 44164 12501 44204
rect 12459 44155 12501 44164
rect 12651 44204 12693 44213
rect 12651 44164 12652 44204
rect 12692 44164 12693 44204
rect 12651 44155 12693 44164
rect 12460 44070 12500 44155
rect 12459 42440 12501 42449
rect 12459 42400 12460 42440
rect 12500 42400 12501 42440
rect 12459 42391 12501 42400
rect 12267 39416 12309 39425
rect 12267 39376 12268 39416
rect 12308 39376 12309 39416
rect 12267 39367 12309 39376
rect 12267 39080 12309 39089
rect 12267 39040 12268 39080
rect 12308 39040 12309 39080
rect 12267 39031 12309 39040
rect 12268 38946 12308 39031
rect 12460 38996 12500 42391
rect 12556 41936 12596 41945
rect 12556 40853 12596 41896
rect 12555 40844 12597 40853
rect 12555 40804 12556 40844
rect 12596 40804 12597 40844
rect 12555 40795 12597 40804
rect 12556 40424 12596 40795
rect 12652 40601 12692 44155
rect 12747 42776 12789 42785
rect 12747 42736 12748 42776
rect 12788 42736 12789 42776
rect 12747 42727 12789 42736
rect 12748 42642 12788 42727
rect 12940 42692 12980 46843
rect 13132 46481 13172 47944
rect 13228 47935 13268 47944
rect 13324 47984 13364 47993
rect 13420 47984 13460 48532
rect 13612 48488 13652 49195
rect 13364 47944 13460 47984
rect 13516 48448 13652 48488
rect 13131 46472 13173 46481
rect 13131 46432 13132 46472
rect 13172 46432 13173 46472
rect 13131 46423 13173 46432
rect 13228 46472 13268 46481
rect 13324 46472 13364 47944
rect 13516 47405 13556 48448
rect 13611 47984 13653 47993
rect 13611 47944 13612 47984
rect 13652 47944 13653 47984
rect 13611 47935 13653 47944
rect 13515 47396 13557 47405
rect 13515 47356 13516 47396
rect 13556 47356 13557 47396
rect 13515 47347 13557 47356
rect 13612 46640 13652 47935
rect 13708 47816 13748 51127
rect 13804 50177 13844 51220
rect 13996 51176 14036 56587
rect 14092 56561 14132 56764
rect 14091 56552 14133 56561
rect 14091 56512 14092 56552
rect 14132 56512 14133 56552
rect 14091 56503 14133 56512
rect 14092 56225 14132 56503
rect 14091 56216 14133 56225
rect 14091 56176 14092 56216
rect 14132 56176 14133 56216
rect 14091 56167 14133 56176
rect 14091 54788 14133 54797
rect 14091 54748 14092 54788
rect 14132 54748 14133 54788
rect 14091 54739 14133 54748
rect 14092 53360 14132 54739
rect 14188 54209 14228 65071
rect 14284 60836 14324 65248
rect 14379 65248 14380 65288
rect 14420 65248 14421 65288
rect 14379 65239 14421 65248
rect 14476 64616 14516 64627
rect 14476 64541 14516 64576
rect 14475 64532 14517 64541
rect 14475 64492 14476 64532
rect 14516 64492 14517 64532
rect 14475 64483 14517 64492
rect 14572 63944 14612 65827
rect 14668 63953 14708 68692
rect 14955 68396 14997 68405
rect 14955 68356 14956 68396
rect 14996 68356 14997 68396
rect 14955 68347 14997 68356
rect 14763 67892 14805 67901
rect 14763 67852 14764 67892
rect 14804 67852 14805 67892
rect 14763 67843 14805 67852
rect 14764 66968 14804 67843
rect 14859 67724 14901 67733
rect 14859 67684 14860 67724
rect 14900 67684 14901 67724
rect 14859 67675 14901 67684
rect 14860 67640 14900 67675
rect 14860 67589 14900 67600
rect 14860 66968 14900 66977
rect 14764 66928 14860 66968
rect 14764 65456 14804 66928
rect 14860 66919 14900 66928
rect 14956 66968 14996 68347
rect 14859 66800 14901 66809
rect 14859 66760 14860 66800
rect 14900 66760 14901 66800
rect 14859 66751 14901 66760
rect 14860 65885 14900 66751
rect 14859 65876 14901 65885
rect 14859 65836 14860 65876
rect 14900 65836 14901 65876
rect 14859 65827 14901 65836
rect 14764 65381 14804 65416
rect 14860 65456 14900 65465
rect 14956 65456 14996 66928
rect 14900 65416 14996 65456
rect 14860 65407 14900 65416
rect 14763 65372 14805 65381
rect 14763 65332 14764 65372
rect 14804 65332 14805 65372
rect 14763 65323 14805 65332
rect 14764 65292 14804 65323
rect 14763 65204 14805 65213
rect 14763 65164 14764 65204
rect 14804 65164 14805 65204
rect 14763 65155 14805 65164
rect 14572 63895 14612 63904
rect 14667 63944 14709 63953
rect 14667 63904 14668 63944
rect 14708 63904 14709 63944
rect 14667 63895 14709 63904
rect 14476 63860 14516 63871
rect 14476 63785 14516 63820
rect 14475 63776 14517 63785
rect 14475 63736 14476 63776
rect 14516 63736 14517 63776
rect 14475 63727 14517 63736
rect 14380 62560 14708 62600
rect 14380 62432 14420 62560
rect 14380 62383 14420 62392
rect 14476 62432 14516 62441
rect 14476 61853 14516 62392
rect 14475 61844 14517 61853
rect 14475 61804 14476 61844
rect 14516 61804 14517 61844
rect 14475 61795 14517 61804
rect 14668 61844 14708 62560
rect 14668 61795 14708 61804
rect 14764 62432 14804 65155
rect 14956 65129 14996 65416
rect 14955 65120 14997 65129
rect 14955 65080 14956 65120
rect 14996 65080 14997 65120
rect 14955 65071 14997 65080
rect 15052 63944 15092 68860
rect 15052 63895 15092 63904
rect 14859 63356 14901 63365
rect 14859 63316 14860 63356
rect 14900 63316 14901 63356
rect 14859 63307 14901 63316
rect 14860 63104 14900 63307
rect 14860 63055 14900 63064
rect 14860 62432 14900 62441
rect 14764 62392 14860 62432
rect 14476 61592 14516 61603
rect 14476 61517 14516 61552
rect 14475 61508 14517 61517
rect 14475 61468 14476 61508
rect 14516 61468 14517 61508
rect 14475 61459 14517 61468
rect 14764 61088 14804 62392
rect 14860 62383 14900 62392
rect 14956 62348 14996 62357
rect 14859 61676 14901 61685
rect 14859 61636 14860 61676
rect 14900 61636 14901 61676
rect 14859 61627 14901 61636
rect 14860 61542 14900 61627
rect 14956 61340 14996 62308
rect 15148 61517 15188 70120
rect 15435 70111 15477 70120
rect 15532 70076 15572 70531
rect 15532 70036 15668 70076
rect 15339 69992 15381 70001
rect 15339 69952 15340 69992
rect 15380 69952 15381 69992
rect 15339 69943 15381 69952
rect 15340 66968 15380 69943
rect 15436 69908 15476 69917
rect 15436 69833 15476 69868
rect 15531 69908 15573 69917
rect 15531 69868 15532 69908
rect 15572 69868 15573 69908
rect 15531 69859 15573 69868
rect 15435 69824 15477 69833
rect 15435 69784 15436 69824
rect 15476 69784 15477 69824
rect 15435 69775 15477 69784
rect 15436 69152 15476 69775
rect 15532 69236 15572 69859
rect 15532 69187 15572 69196
rect 15436 68657 15476 69112
rect 15435 68648 15477 68657
rect 15435 68608 15436 68648
rect 15476 68608 15477 68648
rect 15435 68599 15477 68608
rect 15436 68480 15476 68489
rect 15476 68440 15572 68480
rect 15436 68431 15476 68440
rect 15436 66968 15476 66977
rect 15340 66928 15436 66968
rect 15243 65540 15285 65549
rect 15243 65500 15244 65540
rect 15284 65500 15285 65540
rect 15243 65491 15285 65500
rect 15147 61508 15189 61517
rect 15147 61468 15148 61508
rect 15188 61468 15189 61508
rect 15147 61459 15189 61468
rect 14860 61300 14996 61340
rect 15052 61424 15092 61433
rect 14860 61181 14900 61300
rect 14859 61172 14901 61181
rect 14859 61132 14860 61172
rect 14900 61132 14901 61172
rect 14859 61123 14901 61132
rect 14956 61097 14996 61182
rect 15052 61181 15092 61384
rect 15051 61172 15093 61181
rect 15051 61132 15052 61172
rect 15092 61132 15093 61172
rect 15051 61123 15093 61132
rect 14668 61048 14804 61088
rect 14955 61088 14997 61097
rect 15244 61088 15284 65491
rect 15340 65465 15380 66928
rect 15436 66919 15476 66928
rect 15435 66800 15477 66809
rect 15435 66760 15436 66800
rect 15476 66760 15477 66800
rect 15435 66751 15477 66760
rect 15339 65456 15381 65465
rect 15339 65416 15340 65456
rect 15380 65416 15381 65456
rect 15339 65407 15381 65416
rect 15340 65322 15380 65407
rect 15436 64280 15476 66751
rect 15532 65717 15572 68440
rect 15531 65708 15573 65717
rect 15531 65668 15532 65708
rect 15572 65668 15573 65708
rect 15531 65659 15573 65668
rect 15531 64448 15573 64457
rect 15531 64408 15532 64448
rect 15572 64408 15573 64448
rect 15531 64399 15573 64408
rect 15340 64240 15476 64280
rect 15340 62273 15380 64240
rect 15532 63939 15572 64399
rect 15532 63890 15572 63899
rect 15531 63272 15573 63281
rect 15531 63232 15532 63272
rect 15572 63232 15573 63272
rect 15531 63223 15573 63232
rect 15532 62525 15572 63223
rect 15531 62516 15573 62525
rect 15531 62476 15532 62516
rect 15572 62476 15573 62516
rect 15531 62467 15573 62476
rect 15436 62432 15476 62441
rect 15339 62264 15381 62273
rect 15339 62224 15340 62264
rect 15380 62224 15381 62264
rect 15339 62215 15381 62224
rect 15339 61256 15381 61265
rect 15339 61216 15340 61256
rect 15380 61216 15381 61256
rect 15339 61207 15381 61216
rect 14955 61048 14956 61088
rect 14996 61048 14997 61088
rect 14476 60920 14516 60931
rect 14476 60845 14516 60880
rect 14571 60920 14613 60929
rect 14571 60880 14572 60920
rect 14612 60880 14613 60920
rect 14571 60871 14613 60880
rect 14475 60836 14517 60845
rect 14284 60796 14420 60836
rect 14284 60668 14324 60677
rect 14380 60668 14420 60796
rect 14475 60796 14476 60836
rect 14516 60796 14517 60836
rect 14475 60787 14517 60796
rect 14572 60786 14612 60871
rect 14380 60628 14612 60668
rect 14284 60080 14324 60628
rect 14475 60416 14517 60425
rect 14475 60376 14476 60416
rect 14516 60376 14517 60416
rect 14475 60367 14517 60376
rect 14380 60080 14420 60089
rect 14284 60040 14380 60080
rect 14380 60031 14420 60040
rect 14476 60080 14516 60367
rect 14379 59912 14421 59921
rect 14379 59872 14380 59912
rect 14420 59872 14421 59912
rect 14379 59863 14421 59872
rect 14283 59744 14325 59753
rect 14283 59704 14284 59744
rect 14324 59704 14325 59744
rect 14283 59695 14325 59704
rect 14284 56393 14324 59695
rect 14283 56384 14325 56393
rect 14283 56344 14284 56384
rect 14324 56344 14325 56384
rect 14283 56335 14325 56344
rect 14283 56132 14325 56141
rect 14283 56092 14284 56132
rect 14324 56092 14325 56132
rect 14283 56083 14325 56092
rect 14187 54200 14229 54209
rect 14187 54160 14188 54200
rect 14228 54160 14229 54200
rect 14187 54151 14229 54160
rect 14284 53444 14324 56083
rect 14380 55049 14420 59863
rect 14476 59753 14516 60040
rect 14475 59744 14517 59753
rect 14475 59704 14476 59744
rect 14516 59704 14517 59744
rect 14475 59695 14517 59704
rect 14475 59492 14517 59501
rect 14475 59452 14476 59492
rect 14516 59452 14517 59492
rect 14475 59443 14517 59452
rect 14476 59408 14516 59443
rect 14476 59333 14516 59368
rect 14475 59324 14517 59333
rect 14475 59284 14476 59324
rect 14516 59284 14517 59324
rect 14475 59275 14517 59284
rect 14476 55553 14516 59275
rect 14572 59249 14612 60628
rect 14668 59585 14708 61048
rect 14955 61039 14997 61048
rect 15148 61048 15284 61088
rect 14764 60920 14804 60929
rect 14764 60509 14804 60880
rect 14860 60920 14900 60929
rect 14763 60500 14805 60509
rect 14763 60460 14764 60500
rect 14804 60460 14805 60500
rect 14763 60451 14805 60460
rect 14860 60248 14900 60880
rect 15017 60905 15057 60914
rect 15017 60593 15057 60865
rect 15016 60584 15058 60593
rect 15016 60544 15017 60584
rect 15057 60544 15058 60584
rect 15016 60535 15058 60544
rect 14955 60416 14997 60425
rect 14955 60376 14956 60416
rect 14996 60376 14997 60416
rect 14955 60367 14997 60376
rect 14764 60208 14900 60248
rect 14667 59576 14709 59585
rect 14667 59536 14668 59576
rect 14708 59536 14709 59576
rect 14667 59527 14709 59536
rect 14764 59576 14804 60208
rect 14859 60080 14901 60089
rect 14859 60040 14860 60080
rect 14900 60040 14901 60080
rect 14859 60031 14901 60040
rect 14956 60080 14996 60367
rect 14996 60040 15092 60080
rect 14956 60031 14996 60040
rect 14860 59946 14900 60031
rect 14955 59828 14997 59837
rect 14955 59788 14956 59828
rect 14996 59788 14997 59828
rect 14955 59779 14997 59788
rect 14764 59527 14804 59536
rect 14667 59408 14709 59417
rect 14667 59368 14668 59408
rect 14708 59368 14709 59408
rect 14667 59359 14709 59368
rect 14956 59408 14996 59779
rect 14956 59359 14996 59368
rect 14571 59240 14613 59249
rect 14571 59200 14572 59240
rect 14612 59200 14613 59240
rect 14571 59191 14613 59200
rect 14571 57056 14613 57065
rect 14571 57016 14572 57056
rect 14612 57016 14613 57056
rect 14571 57007 14613 57016
rect 14572 56922 14612 57007
rect 14475 55544 14517 55553
rect 14475 55504 14476 55544
rect 14516 55504 14517 55544
rect 14475 55495 14517 55504
rect 14668 55460 14708 59359
rect 15052 58820 15092 60040
rect 14764 58780 15092 58820
rect 14764 55973 14804 58780
rect 15148 58736 15188 61048
rect 15244 60920 15284 60929
rect 15244 60593 15284 60880
rect 15340 60920 15380 61207
rect 15436 61097 15476 62392
rect 15435 61088 15477 61097
rect 15435 61048 15436 61088
rect 15476 61048 15477 61088
rect 15435 61039 15477 61048
rect 15532 61088 15572 61097
rect 15340 60871 15380 60880
rect 15243 60584 15285 60593
rect 15243 60544 15244 60584
rect 15284 60544 15285 60584
rect 15243 60535 15285 60544
rect 15436 60080 15476 61039
rect 15532 60929 15572 61048
rect 15531 60920 15573 60929
rect 15531 60880 15532 60920
rect 15572 60880 15573 60920
rect 15531 60871 15573 60880
rect 15436 60031 15476 60040
rect 15243 59576 15285 59585
rect 15243 59536 15244 59576
rect 15284 59536 15285 59576
rect 15243 59527 15285 59536
rect 14860 58696 15188 58736
rect 14860 56477 14900 58696
rect 14956 58568 14996 58577
rect 14956 56729 14996 58528
rect 15148 58400 15188 58409
rect 15148 57233 15188 58360
rect 15147 57224 15189 57233
rect 15147 57184 15148 57224
rect 15188 57184 15189 57224
rect 15147 57175 15189 57184
rect 15052 57065 15092 57074
rect 15051 57016 15052 57065
rect 15092 57016 15093 57065
rect 15244 57056 15284 59527
rect 15339 58988 15381 58997
rect 15339 58948 15340 58988
rect 15380 58948 15381 58988
rect 15339 58939 15381 58948
rect 15340 58661 15380 58939
rect 15339 58652 15381 58661
rect 15339 58612 15340 58652
rect 15380 58612 15381 58652
rect 15339 58603 15381 58612
rect 15340 58568 15380 58603
rect 15340 58518 15380 58528
rect 15340 57896 15380 57905
rect 15340 57728 15380 57856
rect 15435 57728 15477 57737
rect 15340 57688 15436 57728
rect 15476 57688 15477 57728
rect 15435 57679 15477 57688
rect 15244 57016 15380 57056
rect 15051 57007 15093 57016
rect 15052 56932 15092 57007
rect 15147 56972 15189 56981
rect 15147 56932 15148 56972
rect 15188 56932 15189 56972
rect 15147 56923 15189 56932
rect 14955 56720 14997 56729
rect 14955 56680 14956 56720
rect 14996 56680 14997 56720
rect 14955 56671 14997 56680
rect 15051 56552 15093 56561
rect 15051 56512 15052 56552
rect 15092 56512 15093 56552
rect 15051 56503 15093 56512
rect 14859 56468 14901 56477
rect 14859 56428 14860 56468
rect 14900 56428 14901 56468
rect 14859 56419 14901 56428
rect 14763 55964 14805 55973
rect 14763 55924 14764 55964
rect 14804 55924 14805 55964
rect 14763 55915 14805 55924
rect 14668 55420 14804 55460
rect 14475 55376 14517 55385
rect 14475 55336 14476 55376
rect 14516 55336 14517 55376
rect 14475 55327 14517 55336
rect 14379 55040 14421 55049
rect 14379 55000 14380 55040
rect 14420 55000 14421 55040
rect 14379 54991 14421 55000
rect 14476 54881 14516 55327
rect 14571 55124 14613 55133
rect 14571 55084 14572 55124
rect 14612 55084 14613 55124
rect 14571 55075 14613 55084
rect 14380 54872 14420 54881
rect 14380 54293 14420 54832
rect 14475 54872 14517 54881
rect 14475 54832 14476 54872
rect 14516 54832 14517 54872
rect 14475 54823 14517 54832
rect 14476 54738 14516 54823
rect 14379 54284 14421 54293
rect 14379 54244 14380 54284
rect 14420 54244 14421 54284
rect 14379 54235 14421 54244
rect 14475 54032 14517 54041
rect 14475 53992 14476 54032
rect 14516 53992 14517 54032
rect 14475 53983 14517 53992
rect 14476 53453 14516 53983
rect 14475 53444 14517 53453
rect 14284 53404 14420 53444
rect 14188 53360 14228 53369
rect 14092 53320 14188 53360
rect 14188 53311 14228 53320
rect 14283 53276 14325 53285
rect 14283 53236 14284 53276
rect 14324 53236 14325 53276
rect 14283 53227 14325 53236
rect 14187 53192 14229 53201
rect 14187 53152 14188 53192
rect 14228 53152 14229 53192
rect 14187 53143 14229 53152
rect 14188 52688 14228 53143
rect 14284 53142 14324 53227
rect 14380 52856 14420 53404
rect 14475 53404 14476 53444
rect 14516 53404 14517 53444
rect 14475 53395 14517 53404
rect 14380 52816 14516 52856
rect 14379 52688 14421 52697
rect 14188 52648 14324 52688
rect 14188 52520 14228 52531
rect 14188 52445 14228 52480
rect 14187 52436 14229 52445
rect 14187 52396 14188 52436
rect 14228 52396 14229 52436
rect 14187 52387 14229 52396
rect 14092 51857 14132 51942
rect 14091 51848 14133 51857
rect 14091 51808 14092 51848
rect 14132 51808 14133 51848
rect 14091 51799 14133 51808
rect 14188 51764 14228 51773
rect 14091 51512 14133 51521
rect 14091 51472 14092 51512
rect 14132 51472 14133 51512
rect 14091 51463 14133 51472
rect 13900 51136 14036 51176
rect 13803 50168 13845 50177
rect 13803 50128 13804 50168
rect 13844 50128 13845 50168
rect 13803 50119 13845 50128
rect 13803 49496 13845 49505
rect 13803 49456 13804 49496
rect 13844 49456 13845 49496
rect 13803 49447 13845 49456
rect 13804 47993 13844 49447
rect 13803 47984 13845 47993
rect 13803 47944 13804 47984
rect 13844 47944 13845 47984
rect 13803 47935 13845 47944
rect 13708 47776 13844 47816
rect 13612 46600 13748 46640
rect 13268 46432 13364 46472
rect 13708 46472 13748 46600
rect 13132 46338 13172 46423
rect 13228 46229 13268 46432
rect 13708 46423 13748 46432
rect 13227 46220 13269 46229
rect 13227 46180 13228 46220
rect 13268 46180 13269 46220
rect 13227 46171 13269 46180
rect 13804 46052 13844 47776
rect 13516 46012 13844 46052
rect 13419 45296 13461 45305
rect 13419 45256 13420 45296
rect 13460 45256 13461 45296
rect 13419 45247 13461 45256
rect 13420 44960 13460 45247
rect 13420 44911 13460 44920
rect 13516 44372 13556 46012
rect 13707 45800 13749 45809
rect 13707 45760 13708 45800
rect 13748 45760 13749 45800
rect 13707 45758 13749 45760
rect 13707 45751 13708 45758
rect 13748 45751 13749 45758
rect 13708 45296 13748 45718
rect 13708 45256 13844 45296
rect 13420 44332 13556 44372
rect 13612 44792 13652 44801
rect 13036 44288 13076 44299
rect 13036 44213 13076 44248
rect 13227 44288 13269 44297
rect 13227 44248 13228 44288
rect 13268 44248 13269 44288
rect 13227 44239 13269 44248
rect 13035 44204 13077 44213
rect 13035 44164 13036 44204
rect 13076 44164 13077 44204
rect 13035 44155 13077 44164
rect 13131 43616 13173 43625
rect 13131 43576 13132 43616
rect 13172 43576 13173 43616
rect 13131 43567 13173 43576
rect 13132 43482 13172 43567
rect 13132 42776 13172 42787
rect 13132 42701 13172 42736
rect 12844 42652 12980 42692
rect 13131 42692 13173 42701
rect 13131 42652 13132 42692
rect 13172 42652 13173 42692
rect 12748 41768 12788 41777
rect 12748 41609 12788 41728
rect 12747 41600 12789 41609
rect 12747 41560 12748 41600
rect 12788 41560 12789 41600
rect 12747 41551 12789 41560
rect 12651 40592 12693 40601
rect 12651 40552 12652 40592
rect 12692 40552 12693 40592
rect 12651 40543 12693 40552
rect 12748 40424 12788 40433
rect 12556 40384 12748 40424
rect 12556 39752 12596 40384
rect 12748 40375 12788 40384
rect 12748 39836 12788 39847
rect 12748 39761 12788 39796
rect 12747 39752 12789 39761
rect 12556 39703 12596 39712
rect 12652 39712 12748 39752
rect 12788 39712 12789 39752
rect 12555 39584 12597 39593
rect 12555 39544 12556 39584
rect 12596 39544 12597 39584
rect 12555 39535 12597 39544
rect 12556 39164 12596 39535
rect 12556 39115 12596 39124
rect 12460 38956 12596 38996
rect 12363 38912 12405 38921
rect 12363 38872 12364 38912
rect 12404 38872 12405 38912
rect 12363 38863 12405 38872
rect 12364 38778 12404 38863
rect 12459 38408 12501 38417
rect 12459 38368 12460 38408
rect 12500 38368 12501 38408
rect 12459 38359 12501 38368
rect 12268 37400 12308 37409
rect 12268 36896 12308 37360
rect 12268 36847 12308 36856
rect 12364 37400 12404 37409
rect 12364 35981 12404 37360
rect 12460 36485 12500 38359
rect 12459 36476 12501 36485
rect 12459 36436 12460 36476
rect 12500 36436 12501 36476
rect 12459 36427 12501 36436
rect 12363 35972 12405 35981
rect 12363 35932 12364 35972
rect 12404 35932 12405 35972
rect 12363 35923 12405 35932
rect 12267 35720 12309 35729
rect 12267 35680 12268 35720
rect 12308 35680 12309 35720
rect 12267 35671 12309 35680
rect 12268 35216 12308 35671
rect 12268 35167 12308 35176
rect 12364 35216 12404 35923
rect 12364 35167 12404 35176
rect 12556 34889 12596 38956
rect 12652 38912 12692 39712
rect 12747 39703 12789 39712
rect 12844 39080 12884 42652
rect 13131 42643 13173 42652
rect 12940 42524 12980 42533
rect 12980 42484 13076 42524
rect 12940 42475 12980 42484
rect 13036 41936 13076 42484
rect 13132 42281 13172 42643
rect 13131 42272 13173 42281
rect 13131 42232 13132 42272
rect 13172 42232 13173 42272
rect 13131 42223 13173 42232
rect 13132 41945 13172 42030
rect 13036 41887 13076 41896
rect 13131 41936 13173 41945
rect 13131 41896 13132 41936
rect 13172 41896 13173 41936
rect 13131 41887 13173 41896
rect 13228 41768 13268 44239
rect 13420 43709 13460 44332
rect 13612 44288 13652 44752
rect 13564 44278 13652 44288
rect 13604 44248 13652 44278
rect 13708 44372 13748 44381
rect 13564 44229 13604 44238
rect 13419 43700 13461 43709
rect 13419 43660 13420 43700
rect 13460 43660 13461 43700
rect 13419 43651 13461 43660
rect 13324 43532 13364 43541
rect 13708 43532 13748 44332
rect 13364 43492 13748 43532
rect 13324 43483 13364 43492
rect 13804 43448 13844 45256
rect 13804 43399 13844 43408
rect 13516 41936 13556 41947
rect 13516 41861 13556 41896
rect 13612 41936 13652 41945
rect 13652 41896 13748 41936
rect 13612 41887 13652 41896
rect 13515 41852 13557 41861
rect 13515 41812 13516 41852
rect 13556 41812 13557 41852
rect 13515 41803 13557 41812
rect 13036 41728 13268 41768
rect 12940 40256 12980 40265
rect 12940 39752 12980 40216
rect 13036 40013 13076 41728
rect 13611 41600 13653 41609
rect 13611 41560 13612 41600
rect 13652 41560 13653 41600
rect 13611 41551 13653 41560
rect 13228 41264 13268 41273
rect 13420 41264 13460 41273
rect 13132 41224 13228 41264
rect 13035 40004 13077 40013
rect 13035 39964 13036 40004
rect 13076 39964 13077 40004
rect 13035 39955 13077 39964
rect 13132 39929 13172 41224
rect 13228 41215 13268 41224
rect 13324 41224 13420 41264
rect 13324 40928 13364 41224
rect 13420 41215 13460 41224
rect 13612 41264 13652 41551
rect 13708 41441 13748 41896
rect 13900 41768 13940 51136
rect 13995 51008 14037 51017
rect 13995 50968 13996 51008
rect 14036 50968 14037 51008
rect 13995 50959 14037 50968
rect 13996 50597 14036 50959
rect 13995 50588 14037 50597
rect 13995 50548 13996 50588
rect 14036 50548 14037 50588
rect 13995 50539 14037 50548
rect 14092 50420 14132 51463
rect 14188 51017 14228 51724
rect 14187 51008 14229 51017
rect 14187 50968 14188 51008
rect 14228 50968 14229 51008
rect 14187 50959 14229 50968
rect 13996 50380 14132 50420
rect 14188 50840 14228 50849
rect 13996 50168 14036 50380
rect 14188 50336 14228 50800
rect 14284 50588 14324 52648
rect 14379 52648 14380 52688
rect 14420 52648 14421 52688
rect 14379 52639 14421 52648
rect 14380 51848 14420 52639
rect 14380 51008 14420 51808
rect 14476 51521 14516 52816
rect 14572 51941 14612 55075
rect 14667 54284 14709 54293
rect 14667 54244 14668 54284
rect 14708 54244 14709 54284
rect 14667 54235 14709 54244
rect 14668 54150 14708 54235
rect 14764 54200 14804 55420
rect 14955 55040 14997 55049
rect 14955 55000 14956 55040
rect 14996 55000 14997 55040
rect 14955 54991 14997 55000
rect 14956 54872 14996 54991
rect 14956 54823 14996 54832
rect 14859 54788 14901 54797
rect 14859 54748 14860 54788
rect 14900 54748 14901 54788
rect 14859 54739 14901 54748
rect 14860 54654 14900 54739
rect 14764 54160 14996 54200
rect 14860 54032 14900 54041
rect 14763 53864 14805 53873
rect 14763 53824 14764 53864
rect 14804 53824 14805 53864
rect 14763 53815 14805 53824
rect 14667 53360 14709 53369
rect 14667 53320 14668 53360
rect 14708 53320 14709 53360
rect 14667 53311 14709 53320
rect 14764 53360 14804 53815
rect 14860 53789 14900 53992
rect 14859 53780 14901 53789
rect 14859 53740 14860 53780
rect 14900 53740 14901 53780
rect 14859 53731 14901 53740
rect 14764 53311 14804 53320
rect 14571 51932 14613 51941
rect 14571 51892 14572 51932
rect 14612 51892 14613 51932
rect 14571 51883 14613 51892
rect 14572 51848 14612 51883
rect 14572 51797 14612 51808
rect 14571 51680 14613 51689
rect 14571 51640 14572 51680
rect 14612 51640 14613 51680
rect 14571 51631 14613 51640
rect 14475 51512 14517 51521
rect 14475 51472 14476 51512
rect 14516 51472 14517 51512
rect 14475 51463 14517 51472
rect 14476 51008 14516 51017
rect 14380 50968 14476 51008
rect 14476 50959 14516 50968
rect 14572 51008 14612 51631
rect 14572 50959 14612 50968
rect 14668 51008 14708 53311
rect 14860 53201 14900 53731
rect 14859 53192 14901 53201
rect 14859 53152 14860 53192
rect 14900 53152 14901 53192
rect 14859 53143 14901 53152
rect 14859 52688 14901 52697
rect 14859 52648 14860 52688
rect 14900 52648 14901 52688
rect 14859 52639 14901 52648
rect 14860 52520 14900 52639
rect 14860 52471 14900 52480
rect 14859 51848 14901 51857
rect 14859 51808 14860 51848
rect 14900 51808 14901 51848
rect 14859 51799 14901 51808
rect 14860 51689 14900 51799
rect 14859 51680 14901 51689
rect 14859 51640 14860 51680
rect 14900 51640 14901 51680
rect 14859 51631 14901 51640
rect 14956 51428 14996 54160
rect 15052 52865 15092 56503
rect 15051 52856 15093 52865
rect 15051 52816 15052 52856
rect 15092 52816 15093 52856
rect 15051 52807 15093 52816
rect 15148 52688 15188 56923
rect 15243 56888 15285 56897
rect 15243 56848 15244 56888
rect 15284 56848 15285 56888
rect 15243 56839 15285 56848
rect 15244 56754 15284 56839
rect 15340 56645 15380 57016
rect 15436 56981 15476 57679
rect 15532 57653 15572 57738
rect 15531 57644 15573 57653
rect 15531 57604 15532 57644
rect 15572 57604 15573 57644
rect 15531 57595 15573 57604
rect 15628 57476 15668 70036
rect 15820 68480 15860 70867
rect 15916 69161 15956 72883
rect 16011 71252 16053 71261
rect 16011 71212 16012 71252
rect 16052 71212 16053 71252
rect 16011 71203 16053 71212
rect 16012 71118 16052 71203
rect 16011 71000 16053 71009
rect 16011 70960 16012 71000
rect 16052 70960 16053 71000
rect 16011 70951 16053 70960
rect 16012 69992 16052 70951
rect 16108 70496 16148 73723
rect 16204 73100 16244 74311
rect 16300 73184 16340 77512
rect 16395 77512 16396 77552
rect 16436 77512 16437 77552
rect 16395 77503 16437 77512
rect 16396 73613 16436 77503
rect 16492 75032 16532 79183
rect 16588 78485 16628 80704
rect 16876 80576 16916 80587
rect 16876 80501 16916 80536
rect 16875 80492 16917 80501
rect 16875 80452 16876 80492
rect 16916 80452 16917 80492
rect 16875 80443 16917 80452
rect 16684 80324 16724 80333
rect 16724 80284 16820 80324
rect 16684 80275 16724 80284
rect 16683 79988 16725 79997
rect 16683 79948 16684 79988
rect 16724 79948 16725 79988
rect 16683 79939 16725 79948
rect 16684 79661 16724 79939
rect 16683 79652 16725 79661
rect 16683 79612 16684 79652
rect 16724 79612 16725 79652
rect 16683 79603 16725 79612
rect 16683 79484 16725 79493
rect 16683 79444 16684 79484
rect 16724 79444 16725 79484
rect 16683 79435 16725 79444
rect 16587 78476 16629 78485
rect 16587 78436 16588 78476
rect 16628 78436 16629 78476
rect 16587 78427 16629 78436
rect 16684 77384 16724 79435
rect 16780 79316 16820 80284
rect 16876 79997 16916 80443
rect 16875 79988 16917 79997
rect 16875 79948 16876 79988
rect 16916 79948 16917 79988
rect 16875 79939 16917 79948
rect 16876 79736 16916 79745
rect 16876 79493 16916 79696
rect 16875 79484 16917 79493
rect 16875 79444 16876 79484
rect 16916 79444 16917 79484
rect 16875 79435 16917 79444
rect 16780 79276 16916 79316
rect 16876 78238 16916 79276
rect 16876 78189 16916 78198
rect 16972 78149 17012 80704
rect 17068 79829 17108 82720
rect 17067 79820 17109 79829
rect 17067 79780 17068 79820
rect 17108 79780 17109 79820
rect 17067 79771 17109 79780
rect 17067 79652 17109 79661
rect 17067 79612 17068 79652
rect 17108 79612 17109 79652
rect 17067 79603 17109 79612
rect 17068 79064 17108 79603
rect 17164 79232 17204 85936
rect 17260 84272 17300 84281
rect 17260 84029 17300 84232
rect 17259 84020 17301 84029
rect 17259 83980 17260 84020
rect 17300 83980 17301 84020
rect 17259 83971 17301 83980
rect 17260 83273 17300 83971
rect 17259 83264 17301 83273
rect 17259 83224 17260 83264
rect 17300 83224 17301 83264
rect 17259 83215 17301 83224
rect 17356 83189 17396 85936
rect 17355 83180 17397 83189
rect 17355 83140 17356 83180
rect 17396 83140 17397 83180
rect 17355 83131 17397 83140
rect 17451 82760 17493 82769
rect 17451 82720 17452 82760
rect 17492 82720 17493 82760
rect 17451 82711 17493 82720
rect 17452 82626 17492 82711
rect 17260 82592 17300 82601
rect 17260 81920 17300 82552
rect 17548 81920 17588 85936
rect 17740 84533 17780 85936
rect 17739 84524 17781 84533
rect 17739 84484 17740 84524
rect 17780 84484 17781 84524
rect 17739 84475 17781 84484
rect 17932 84449 17972 85936
rect 18124 84785 18164 85936
rect 18219 85028 18261 85037
rect 18219 84988 18220 85028
rect 18260 84988 18261 85028
rect 18219 84979 18261 84988
rect 18123 84776 18165 84785
rect 18123 84736 18124 84776
rect 18164 84736 18165 84776
rect 18123 84727 18165 84736
rect 17931 84440 17973 84449
rect 17931 84400 17932 84440
rect 17972 84400 17973 84440
rect 17931 84391 17973 84400
rect 18027 84272 18069 84281
rect 18027 84232 18028 84272
rect 18068 84232 18069 84272
rect 18027 84223 18069 84232
rect 17739 83684 17781 83693
rect 17739 83644 17740 83684
rect 17780 83644 17781 83684
rect 17739 83635 17781 83644
rect 17740 83600 17780 83635
rect 17740 82769 17780 83560
rect 17932 83348 17972 83357
rect 17836 83308 17932 83348
rect 17739 82760 17781 82769
rect 17739 82720 17740 82760
rect 17780 82720 17781 82760
rect 17739 82711 17781 82720
rect 17836 82592 17876 83308
rect 17932 83299 17972 83308
rect 17260 81880 17396 81920
rect 17259 80660 17301 80669
rect 17259 80620 17260 80660
rect 17300 80620 17301 80660
rect 17259 80611 17301 80620
rect 17260 79652 17300 80611
rect 17356 79750 17396 81880
rect 17356 79701 17396 79710
rect 17452 81880 17588 81920
rect 17644 82552 17876 82592
rect 17260 79612 17396 79652
rect 17164 79192 17300 79232
rect 17164 79064 17204 79073
rect 17068 79024 17164 79064
rect 17068 78737 17108 79024
rect 17164 79015 17204 79024
rect 17163 78812 17205 78821
rect 17163 78772 17164 78812
rect 17204 78772 17205 78812
rect 17163 78763 17205 78772
rect 17067 78728 17109 78737
rect 17067 78688 17068 78728
rect 17108 78688 17109 78728
rect 17067 78679 17109 78688
rect 17067 78560 17109 78569
rect 17067 78520 17068 78560
rect 17108 78520 17109 78560
rect 17067 78511 17109 78520
rect 16971 78140 17013 78149
rect 16971 78100 16972 78140
rect 17012 78100 17013 78140
rect 16971 78091 17013 78100
rect 17068 78056 17108 78511
rect 17068 77804 17108 78016
rect 16876 77764 17108 77804
rect 16779 77552 16821 77561
rect 16779 77512 16780 77552
rect 16820 77512 16821 77552
rect 16779 77503 16821 77512
rect 16780 77418 16820 77503
rect 16588 77344 16724 77384
rect 16588 75209 16628 77344
rect 16683 75872 16725 75881
rect 16683 75832 16684 75872
rect 16724 75832 16725 75872
rect 16683 75823 16725 75832
rect 16587 75200 16629 75209
rect 16587 75160 16588 75200
rect 16628 75160 16629 75200
rect 16587 75151 16629 75160
rect 16684 75200 16724 75823
rect 16876 75704 16916 77764
rect 17164 77636 17204 78763
rect 17260 78233 17300 79192
rect 17356 79054 17396 79612
rect 17452 79325 17492 81880
rect 17644 79829 17684 82552
rect 18028 82172 18068 84223
rect 18124 83357 18164 83442
rect 18123 83348 18165 83357
rect 18123 83308 18124 83348
rect 18164 83308 18165 83348
rect 18220 83348 18260 84979
rect 18316 84113 18356 85936
rect 18411 84692 18453 84701
rect 18411 84652 18412 84692
rect 18452 84652 18453 84692
rect 18411 84643 18453 84652
rect 18315 84104 18357 84113
rect 18315 84064 18316 84104
rect 18356 84064 18357 84104
rect 18315 84055 18357 84064
rect 18315 83936 18357 83945
rect 18315 83896 18316 83936
rect 18356 83896 18357 83936
rect 18315 83887 18357 83896
rect 18316 83516 18356 83887
rect 18316 83467 18356 83476
rect 18220 83308 18356 83348
rect 18123 83299 18165 83308
rect 18219 83180 18261 83189
rect 18219 83140 18220 83180
rect 18260 83140 18261 83180
rect 18219 83131 18261 83140
rect 18123 83096 18165 83105
rect 18123 83056 18124 83096
rect 18164 83056 18165 83096
rect 18123 83047 18165 83056
rect 17836 82132 18068 82172
rect 17739 80408 17781 80417
rect 17739 80368 17740 80408
rect 17780 80368 17781 80408
rect 17739 80359 17781 80368
rect 17740 79997 17780 80359
rect 17739 79988 17781 79997
rect 17739 79948 17740 79988
rect 17780 79948 17781 79988
rect 17739 79939 17781 79948
rect 17643 79820 17685 79829
rect 17643 79780 17644 79820
rect 17684 79780 17685 79820
rect 17643 79771 17685 79780
rect 17547 79568 17589 79577
rect 17547 79528 17548 79568
rect 17588 79528 17589 79568
rect 17547 79519 17589 79528
rect 17548 79434 17588 79519
rect 17548 79325 17588 79327
rect 17440 79316 17492 79325
rect 17440 79276 17441 79316
rect 17481 79276 17492 79316
rect 17547 79316 17589 79325
rect 17547 79276 17548 79316
rect 17588 79276 17589 79316
rect 17440 79267 17482 79276
rect 17547 79267 17589 79276
rect 17548 79232 17588 79267
rect 17548 79183 17588 79192
rect 17644 79064 17684 79771
rect 17739 79652 17781 79661
rect 17739 79612 17740 79652
rect 17780 79612 17781 79652
rect 17739 79603 17781 79612
rect 17740 79518 17780 79603
rect 17836 79400 17876 82132
rect 18028 82088 18068 82132
rect 18028 82039 18068 82048
rect 17931 81920 17973 81929
rect 17931 81880 17932 81920
rect 17972 81880 17973 81920
rect 17931 81871 17973 81880
rect 17932 80417 17972 81871
rect 18028 81248 18068 81257
rect 18028 80669 18068 81208
rect 18124 80744 18164 83047
rect 18220 82013 18260 83131
rect 18219 82004 18261 82013
rect 18219 81964 18220 82004
rect 18260 81964 18261 82004
rect 18219 81955 18261 81964
rect 18316 81920 18356 83308
rect 18412 83189 18452 84643
rect 18508 84524 18548 85936
rect 18700 84701 18740 85936
rect 18892 84860 18932 85936
rect 19084 85037 19124 85936
rect 19276 85121 19316 85936
rect 19275 85112 19317 85121
rect 19275 85072 19276 85112
rect 19316 85072 19317 85112
rect 19275 85063 19317 85072
rect 19083 85028 19125 85037
rect 19083 84988 19084 85028
rect 19124 84988 19125 85028
rect 19083 84979 19125 84988
rect 19468 84953 19508 85936
rect 19467 84944 19509 84953
rect 19467 84904 19468 84944
rect 19508 84904 19509 84944
rect 19467 84895 19509 84904
rect 19563 84860 19605 84869
rect 18892 84820 19412 84860
rect 18699 84692 18741 84701
rect 18699 84652 18700 84692
rect 18740 84652 18741 84692
rect 18699 84643 18741 84652
rect 18808 84692 19176 84701
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 18808 84643 19176 84652
rect 18891 84524 18933 84533
rect 18508 84484 18740 84524
rect 18700 84281 18740 84484
rect 18891 84484 18892 84524
rect 18932 84484 18933 84524
rect 18891 84475 18933 84484
rect 18892 84390 18932 84475
rect 19275 84440 19317 84449
rect 19275 84400 19276 84440
rect 19316 84400 19317 84440
rect 19275 84391 19317 84400
rect 19084 84356 19124 84365
rect 18507 84272 18549 84281
rect 18507 84232 18508 84272
rect 18548 84232 18549 84272
rect 18507 84223 18549 84232
rect 18699 84272 18741 84281
rect 18699 84232 18700 84272
rect 18740 84232 18741 84272
rect 18699 84223 18741 84232
rect 18508 84138 18548 84223
rect 19084 84197 19124 84316
rect 19276 84306 19316 84391
rect 19083 84188 19125 84197
rect 19083 84148 19084 84188
rect 19124 84148 19125 84188
rect 19372 84188 19412 84820
rect 19563 84820 19564 84860
rect 19604 84820 19605 84860
rect 19563 84811 19605 84820
rect 19468 84365 19508 84450
rect 19467 84356 19509 84365
rect 19467 84316 19468 84356
rect 19508 84316 19509 84356
rect 19467 84307 19509 84316
rect 19372 84148 19508 84188
rect 19083 84139 19125 84148
rect 18700 84104 18740 84113
rect 18604 84064 18700 84104
rect 18507 83768 18549 83777
rect 18507 83728 18508 83768
rect 18548 83728 18549 83768
rect 18507 83719 18549 83728
rect 18508 83634 18548 83719
rect 18411 83180 18453 83189
rect 18411 83140 18412 83180
rect 18452 83140 18453 83180
rect 18411 83131 18453 83140
rect 18507 83012 18549 83021
rect 18507 82972 18508 83012
rect 18548 82972 18549 83012
rect 18604 83012 18644 84064
rect 18700 84055 18740 84064
rect 18892 83644 19124 83684
rect 18700 83525 18740 83610
rect 18699 83516 18741 83525
rect 18699 83476 18700 83516
rect 18740 83476 18741 83516
rect 18699 83467 18741 83476
rect 18892 83348 18932 83644
rect 19084 83642 19124 83644
rect 19084 83593 19124 83602
rect 19276 83600 19316 83609
rect 19084 83441 19124 83526
rect 19083 83432 19125 83441
rect 19083 83392 19084 83432
rect 19124 83392 19125 83432
rect 19083 83383 19125 83392
rect 18700 83308 18932 83348
rect 18700 83189 18740 83308
rect 18699 83180 18741 83189
rect 18699 83140 18700 83180
rect 18740 83140 18741 83180
rect 18699 83131 18741 83140
rect 18808 83180 19176 83189
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 18808 83131 19176 83140
rect 19083 83012 19125 83021
rect 18604 82972 18836 83012
rect 18507 82963 18549 82972
rect 18508 82088 18548 82963
rect 18699 82760 18741 82769
rect 18699 82720 18700 82760
rect 18740 82720 18741 82760
rect 18699 82711 18741 82720
rect 18700 82626 18740 82711
rect 18604 82088 18644 82097
rect 18508 82048 18604 82088
rect 18604 82039 18644 82048
rect 18316 81880 18452 81920
rect 18220 81836 18260 81845
rect 18260 81796 18356 81836
rect 18220 81787 18260 81796
rect 18219 81080 18261 81089
rect 18219 81040 18220 81080
rect 18260 81040 18261 81080
rect 18219 81031 18261 81040
rect 18220 80946 18260 81031
rect 18124 80704 18260 80744
rect 18027 80660 18069 80669
rect 18027 80620 18028 80660
rect 18068 80620 18069 80660
rect 18027 80611 18069 80620
rect 18123 80576 18165 80585
rect 18123 80536 18124 80576
rect 18164 80536 18165 80576
rect 18123 80527 18165 80536
rect 18124 80442 18164 80527
rect 17931 80408 17973 80417
rect 17931 80368 17932 80408
rect 17972 80368 17973 80408
rect 17931 80359 17973 80368
rect 18123 79988 18165 79997
rect 18123 79948 18124 79988
rect 18164 79948 18165 79988
rect 18123 79939 18165 79948
rect 17931 79904 17973 79913
rect 17931 79864 17932 79904
rect 17972 79864 17973 79904
rect 17931 79855 17973 79864
rect 17932 79750 17972 79855
rect 17932 79701 17972 79710
rect 18124 79661 18164 79939
rect 18123 79652 18165 79661
rect 18123 79612 18124 79652
rect 18164 79612 18165 79652
rect 18123 79603 18165 79612
rect 17356 79014 17492 79054
rect 17644 79015 17684 79024
rect 17740 79360 17876 79400
rect 17356 78821 17396 78906
rect 17355 78812 17397 78821
rect 17355 78772 17356 78812
rect 17396 78772 17397 78812
rect 17355 78763 17397 78772
rect 17452 78308 17492 79014
rect 17740 78812 17780 79360
rect 17931 79232 17973 79241
rect 17931 79192 17932 79232
rect 17972 79192 17973 79232
rect 17931 79183 17973 79192
rect 18124 79232 18164 79241
rect 18220 79232 18260 80704
rect 18164 79192 18260 79232
rect 18124 79183 18164 79192
rect 17835 79064 17877 79073
rect 17835 79024 17836 79064
rect 17876 79024 17877 79064
rect 17835 79015 17877 79024
rect 17932 79064 17972 79183
rect 17932 79015 17972 79024
rect 18027 79064 18069 79073
rect 18027 79024 18028 79064
rect 18068 79024 18069 79064
rect 18027 79015 18069 79024
rect 18316 79045 18356 81796
rect 18412 79988 18452 81880
rect 18796 81845 18836 82972
rect 19083 82972 19084 83012
rect 19124 82972 19125 83012
rect 19083 82963 19125 82972
rect 19084 82878 19124 82963
rect 18891 82676 18933 82685
rect 18891 82636 18892 82676
rect 18932 82636 18933 82676
rect 18891 82627 18933 82636
rect 18892 82542 18932 82627
rect 19276 81929 19316 83560
rect 19372 83600 19412 83609
rect 19372 83021 19412 83560
rect 19468 83180 19508 84148
rect 19564 83768 19604 84811
rect 19755 84776 19797 84785
rect 19755 84736 19756 84776
rect 19796 84736 19797 84776
rect 19755 84727 19797 84736
rect 19659 84104 19701 84113
rect 19659 84064 19660 84104
rect 19700 84064 19701 84104
rect 19659 84055 19701 84064
rect 19660 83970 19700 84055
rect 19564 83719 19604 83728
rect 19756 83684 19796 84727
rect 20043 84608 20085 84617
rect 20043 84568 20044 84608
rect 20084 84568 20085 84608
rect 20043 84559 20085 84568
rect 20044 84440 20084 84559
rect 20044 84391 20084 84400
rect 19851 84356 19893 84365
rect 19851 84316 19852 84356
rect 19892 84316 19893 84356
rect 19851 84307 19893 84316
rect 20236 84356 20276 84365
rect 20276 84316 20660 84356
rect 20236 84307 20276 84316
rect 19852 84222 19892 84307
rect 19947 84272 19989 84281
rect 19947 84232 19948 84272
rect 19988 84232 19989 84272
rect 19947 84223 19989 84232
rect 19948 83768 19988 84223
rect 20048 83936 20416 83945
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20048 83887 20416 83896
rect 19948 83719 19988 83728
rect 19756 83644 19892 83684
rect 19755 83516 19797 83525
rect 19755 83476 19756 83516
rect 19796 83476 19797 83516
rect 19755 83467 19797 83476
rect 19756 83382 19796 83467
rect 19852 83180 19892 83644
rect 20121 83513 20161 83522
rect 20121 83273 20161 83473
rect 20120 83264 20162 83273
rect 20120 83224 20121 83264
rect 20161 83224 20162 83264
rect 20120 83215 20162 83224
rect 19468 83140 19604 83180
rect 19852 83140 20084 83180
rect 19371 83012 19413 83021
rect 19371 82972 19372 83012
rect 19412 82972 19413 83012
rect 19371 82963 19413 82972
rect 19468 82760 19508 82769
rect 19372 82676 19412 82687
rect 19372 82601 19412 82636
rect 19371 82592 19413 82601
rect 19371 82552 19372 82592
rect 19412 82552 19413 82592
rect 19371 82543 19413 82552
rect 19468 82517 19508 82720
rect 19467 82508 19509 82517
rect 19467 82468 19468 82508
rect 19508 82468 19509 82508
rect 19467 82459 19509 82468
rect 19275 81920 19317 81929
rect 19275 81880 19276 81920
rect 19316 81880 19317 81920
rect 19275 81871 19317 81880
rect 18795 81836 18837 81845
rect 18795 81796 18796 81836
rect 18836 81796 18837 81836
rect 18795 81787 18837 81796
rect 19275 81752 19317 81761
rect 19275 81712 19276 81752
rect 19316 81712 19317 81752
rect 19275 81703 19317 81712
rect 18808 81668 19176 81677
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 18808 81619 19176 81628
rect 18603 81416 18645 81425
rect 18603 81376 18604 81416
rect 18644 81376 18645 81416
rect 18603 81367 18645 81376
rect 18604 81282 18644 81367
rect 18795 81248 18837 81257
rect 18795 81208 18796 81248
rect 18836 81208 18837 81248
rect 18795 81199 18837 81208
rect 18796 81114 18836 81199
rect 18508 81080 18548 81091
rect 18508 81005 18548 81040
rect 18603 81080 18645 81089
rect 18603 81040 18604 81080
rect 18644 81040 18645 81080
rect 18603 81031 18645 81040
rect 18507 80996 18549 81005
rect 18507 80956 18508 80996
rect 18548 80956 18549 80996
rect 18507 80947 18549 80956
rect 18507 80408 18549 80417
rect 18507 80368 18508 80408
rect 18548 80368 18549 80408
rect 18507 80359 18549 80368
rect 18508 80274 18548 80359
rect 18412 79948 18548 79988
rect 18412 79736 18452 79747
rect 18412 79661 18452 79696
rect 18411 79652 18453 79661
rect 18411 79612 18412 79652
rect 18452 79612 18453 79652
rect 18411 79603 18453 79612
rect 18508 79157 18548 79948
rect 18507 79148 18549 79157
rect 18507 79108 18508 79148
rect 18548 79108 18549 79148
rect 18507 79099 18549 79108
rect 18412 79045 18452 79054
rect 17836 78930 17876 79015
rect 18028 78930 18068 79015
rect 18316 79005 18412 79045
rect 18412 78996 18452 79005
rect 18508 79045 18548 79054
rect 18508 78989 18548 79005
rect 18219 78980 18261 78989
rect 18219 78940 18220 78980
rect 18260 78940 18261 78980
rect 18219 78931 18261 78940
rect 18507 78980 18549 78989
rect 18507 78940 18508 78980
rect 18548 78940 18549 78980
rect 18507 78931 18549 78940
rect 17740 78772 17876 78812
rect 17643 78476 17685 78485
rect 17643 78436 17644 78476
rect 17684 78436 17685 78476
rect 17643 78427 17685 78436
rect 17644 78342 17684 78427
rect 17836 78308 17876 78772
rect 18123 78644 18165 78653
rect 18123 78604 18124 78644
rect 18164 78604 18165 78644
rect 18123 78595 18165 78604
rect 17259 78224 17301 78233
rect 17259 78184 17260 78224
rect 17300 78184 17301 78224
rect 17259 78175 17301 78184
rect 17259 78056 17301 78065
rect 17259 78016 17260 78056
rect 17300 78016 17301 78056
rect 17259 78007 17301 78016
rect 17260 77922 17300 78007
rect 17355 77720 17397 77729
rect 17355 77680 17356 77720
rect 17396 77680 17397 77720
rect 17355 77671 17397 77680
rect 17164 77596 17300 77636
rect 17163 77468 17205 77477
rect 17163 77428 17164 77468
rect 17204 77428 17205 77468
rect 17163 77419 17205 77428
rect 17164 77334 17204 77419
rect 16972 77300 17012 77309
rect 16972 75881 17012 77260
rect 16971 75872 17013 75881
rect 16971 75832 16972 75872
rect 17012 75832 17013 75872
rect 16971 75823 17013 75832
rect 16876 75664 17012 75704
rect 16875 75452 16917 75461
rect 16875 75412 16876 75452
rect 16916 75412 16917 75452
rect 16875 75403 16917 75412
rect 16684 75151 16724 75160
rect 16780 75200 16820 75209
rect 16780 75032 16820 75160
rect 16492 74992 16820 75032
rect 16491 74528 16533 74537
rect 16491 74488 16492 74528
rect 16532 74488 16533 74528
rect 16491 74479 16533 74488
rect 16492 74394 16532 74479
rect 16395 73604 16437 73613
rect 16395 73564 16396 73604
rect 16436 73564 16437 73604
rect 16395 73555 16437 73564
rect 16300 73144 16436 73184
rect 16204 73060 16340 73100
rect 16204 72932 16244 72941
rect 16204 72176 16244 72892
rect 16300 72932 16340 73060
rect 16396 72941 16436 73144
rect 16300 72260 16340 72892
rect 16395 72932 16437 72941
rect 16395 72892 16396 72932
rect 16436 72892 16437 72932
rect 16395 72883 16437 72892
rect 16300 72211 16340 72220
rect 16204 71672 16244 72136
rect 16395 72008 16437 72017
rect 16395 71968 16396 72008
rect 16436 71968 16437 72008
rect 16395 71959 16437 71968
rect 16204 71632 16340 71672
rect 16204 71504 16244 71513
rect 16204 71429 16244 71464
rect 16203 71420 16245 71429
rect 16203 71380 16204 71420
rect 16244 71380 16245 71420
rect 16203 71371 16245 71380
rect 16204 70664 16244 71371
rect 16204 70615 16244 70624
rect 16108 70456 16244 70496
rect 15915 69152 15957 69161
rect 15915 69112 15916 69152
rect 15956 69112 15957 69152
rect 15915 69103 15957 69112
rect 16012 69152 16052 69952
rect 15916 68480 15956 68489
rect 15820 68440 15916 68480
rect 15916 67640 15956 68440
rect 15916 67556 15956 67600
rect 15820 67516 15956 67556
rect 15820 66632 15860 67516
rect 15915 67220 15957 67229
rect 15915 67180 15916 67220
rect 15956 67180 15957 67220
rect 15915 67171 15957 67180
rect 15916 66963 15956 67171
rect 15916 66914 15956 66923
rect 16012 66809 16052 69112
rect 16107 68984 16149 68993
rect 16107 68944 16108 68984
rect 16148 68944 16149 68984
rect 16107 68935 16149 68944
rect 16108 67229 16148 68935
rect 16107 67220 16149 67229
rect 16107 67180 16108 67220
rect 16148 67180 16149 67220
rect 16107 67171 16149 67180
rect 16107 67052 16149 67061
rect 16107 67012 16108 67052
rect 16148 67012 16149 67052
rect 16107 67003 16149 67012
rect 16108 66918 16148 67003
rect 16011 66800 16053 66809
rect 16011 66760 16012 66800
rect 16052 66760 16053 66800
rect 16011 66751 16053 66760
rect 15820 66592 16148 66632
rect 15723 66128 15765 66137
rect 15723 66088 15724 66128
rect 15764 66088 15765 66128
rect 15723 66079 15765 66088
rect 15724 65994 15764 66079
rect 15916 65960 15956 65969
rect 15916 65456 15956 65920
rect 16011 65540 16053 65549
rect 16011 65500 16012 65540
rect 16052 65500 16053 65540
rect 16011 65491 16053 65500
rect 15868 65446 15956 65456
rect 15908 65416 15956 65446
rect 16012 65406 16052 65491
rect 15868 65397 15908 65406
rect 15723 64616 15765 64625
rect 15723 64576 15724 64616
rect 15764 64576 15765 64616
rect 15723 64567 15765 64576
rect 15724 64482 15764 64567
rect 15915 64448 15957 64457
rect 15915 64408 15916 64448
rect 15956 64408 15957 64448
rect 15915 64399 15957 64408
rect 15916 64314 15956 64399
rect 16108 64373 16148 66592
rect 16107 64364 16149 64373
rect 16107 64324 16108 64364
rect 16148 64324 16149 64364
rect 16107 64315 16149 64324
rect 15819 64280 15861 64289
rect 15819 64240 15820 64280
rect 15860 64240 15861 64280
rect 15819 64231 15861 64240
rect 15724 64028 15764 64037
rect 15724 63281 15764 63988
rect 15723 63272 15765 63281
rect 15723 63232 15724 63272
rect 15764 63232 15765 63272
rect 15723 63223 15765 63232
rect 15723 63104 15765 63113
rect 15723 63064 15724 63104
rect 15764 63064 15765 63104
rect 15723 63055 15765 63064
rect 15724 58064 15764 63055
rect 15820 58400 15860 64231
rect 16204 63113 16244 70456
rect 16300 69917 16340 71632
rect 16299 69908 16341 69917
rect 16299 69868 16300 69908
rect 16340 69868 16341 69908
rect 16299 69859 16341 69868
rect 16396 69824 16436 71959
rect 16491 71252 16533 71261
rect 16491 71212 16492 71252
rect 16532 71212 16533 71252
rect 16491 71203 16533 71212
rect 16492 69987 16532 71203
rect 16684 70337 16724 74992
rect 16780 74528 16820 74537
rect 16876 74528 16916 75403
rect 16972 75189 17012 75664
rect 17164 75293 17204 75378
rect 17260 75377 17300 77596
rect 17356 77586 17396 77671
rect 17452 76712 17492 78268
rect 17835 78268 17836 78308
rect 17835 78259 17876 78268
rect 18027 78308 18069 78317
rect 18027 78268 18028 78308
rect 18068 78268 18069 78308
rect 18027 78259 18069 78268
rect 17547 78224 17589 78233
rect 17547 78184 17548 78224
rect 17588 78184 17589 78224
rect 17547 78175 17589 78184
rect 17548 77720 17588 78175
rect 17835 78140 17875 78259
rect 18028 78174 18068 78259
rect 18124 78149 18164 78595
rect 17931 78140 17973 78149
rect 17835 78100 17876 78140
rect 17548 77671 17588 77680
rect 17739 77552 17781 77561
rect 17739 77512 17740 77552
rect 17780 77512 17781 77552
rect 17739 77503 17781 77512
rect 17740 77468 17780 77503
rect 17740 77417 17780 77428
rect 17492 76672 17588 76712
rect 17452 76663 17492 76672
rect 17451 76040 17493 76049
rect 17451 76000 17452 76040
rect 17492 76000 17493 76040
rect 17451 75991 17493 76000
rect 17452 75906 17492 75991
rect 17355 75620 17397 75629
rect 17355 75580 17356 75620
rect 17396 75580 17397 75620
rect 17355 75571 17397 75580
rect 17259 75368 17301 75377
rect 17259 75328 17260 75368
rect 17300 75328 17301 75368
rect 17259 75319 17301 75328
rect 17163 75284 17205 75293
rect 17163 75244 17164 75284
rect 17204 75244 17205 75284
rect 17163 75235 17205 75244
rect 17260 75200 17300 75209
rect 16972 75160 17260 75189
rect 16972 75149 17300 75160
rect 16820 74488 16916 74528
rect 16780 74479 16820 74488
rect 16876 73688 16916 74488
rect 16971 74528 17013 74537
rect 16971 74488 16972 74528
rect 17012 74488 17013 74528
rect 16971 74479 17013 74488
rect 16876 73639 16916 73648
rect 16780 73016 16820 73025
rect 16780 72176 16820 72976
rect 16875 72932 16917 72941
rect 16875 72892 16876 72932
rect 16916 72892 16917 72932
rect 16875 72883 16917 72892
rect 16780 71933 16820 72136
rect 16779 71924 16821 71933
rect 16779 71884 16780 71924
rect 16820 71884 16821 71924
rect 16779 71875 16821 71884
rect 16683 70328 16725 70337
rect 16683 70288 16684 70328
rect 16724 70288 16725 70328
rect 16683 70279 16725 70288
rect 16684 70076 16724 70085
rect 16492 69938 16532 69947
rect 16588 70036 16684 70076
rect 16396 69784 16532 69824
rect 16395 69656 16437 69665
rect 16395 69616 16396 69656
rect 16436 69616 16437 69656
rect 16395 69607 16437 69616
rect 16299 69152 16341 69161
rect 16299 69112 16300 69152
rect 16340 69112 16341 69152
rect 16299 69103 16341 69112
rect 16300 64121 16340 69103
rect 16299 64112 16341 64121
rect 16299 64072 16300 64112
rect 16340 64072 16341 64112
rect 16299 64063 16341 64072
rect 16300 63944 16340 63955
rect 16300 63869 16340 63904
rect 16299 63860 16341 63869
rect 16299 63820 16300 63860
rect 16340 63820 16341 63860
rect 16299 63811 16341 63820
rect 16108 63104 16148 63113
rect 15915 63020 15957 63029
rect 16108 63020 16148 63064
rect 16203 63104 16245 63113
rect 16203 63064 16204 63104
rect 16244 63064 16245 63104
rect 16203 63055 16245 63064
rect 15915 62980 15916 63020
rect 15956 62980 16148 63020
rect 15915 62971 15957 62980
rect 16300 62936 16340 62945
rect 16012 62896 16300 62936
rect 16012 62432 16052 62896
rect 16300 62887 16340 62896
rect 16107 62600 16149 62609
rect 16107 62560 16108 62600
rect 16148 62560 16149 62600
rect 16107 62551 16149 62560
rect 16108 62466 16148 62551
rect 15964 62422 16052 62432
rect 16004 62392 16052 62422
rect 15964 62373 16004 62382
rect 16203 61844 16245 61853
rect 16203 61804 16204 61844
rect 16244 61804 16245 61844
rect 16203 61795 16245 61804
rect 16107 61760 16149 61769
rect 16107 61720 16108 61760
rect 16148 61720 16149 61760
rect 16107 61711 16149 61720
rect 15916 61676 15956 61685
rect 15916 61433 15956 61636
rect 16108 61626 16148 61711
rect 15915 61424 15957 61433
rect 15915 61384 15916 61424
rect 15956 61384 15957 61424
rect 15915 61375 15957 61384
rect 16204 60836 16244 61795
rect 16300 61685 16340 61716
rect 16299 61676 16341 61685
rect 16299 61636 16300 61676
rect 16340 61636 16341 61676
rect 16299 61627 16341 61636
rect 16300 61592 16340 61627
rect 16300 61349 16340 61552
rect 16299 61340 16341 61349
rect 16299 61300 16300 61340
rect 16340 61300 16341 61340
rect 16299 61291 16341 61300
rect 16300 60962 16340 61291
rect 16300 60913 16340 60922
rect 16204 60796 16340 60836
rect 16203 60668 16245 60677
rect 16203 60628 16204 60668
rect 16244 60628 16245 60668
rect 16203 60619 16245 60628
rect 15916 60085 15956 60094
rect 15916 59585 15956 60045
rect 16107 59912 16149 59921
rect 16107 59872 16108 59912
rect 16148 59872 16149 59912
rect 16107 59863 16149 59872
rect 16108 59778 16148 59863
rect 15915 59576 15957 59585
rect 15915 59536 15916 59576
rect 15956 59536 15957 59576
rect 15915 59527 15957 59536
rect 16204 59408 16244 60619
rect 16204 59359 16244 59368
rect 15820 58360 16148 58400
rect 15724 58024 15860 58064
rect 15723 57896 15765 57905
rect 15723 57856 15724 57896
rect 15764 57856 15765 57896
rect 15723 57847 15765 57856
rect 15724 57762 15764 57847
rect 15723 57644 15765 57653
rect 15723 57604 15724 57644
rect 15764 57604 15765 57644
rect 15723 57595 15765 57604
rect 15532 57436 15668 57476
rect 15435 56972 15477 56981
rect 15435 56932 15436 56972
rect 15476 56932 15477 56972
rect 15435 56923 15477 56932
rect 15339 56636 15381 56645
rect 15339 56596 15340 56636
rect 15380 56596 15381 56636
rect 15339 56587 15381 56596
rect 15244 56384 15284 56393
rect 15244 56225 15284 56344
rect 15339 56384 15381 56393
rect 15339 56344 15340 56384
rect 15380 56344 15381 56384
rect 15339 56335 15381 56344
rect 15243 56216 15285 56225
rect 15243 56176 15244 56216
rect 15284 56176 15285 56216
rect 15243 56167 15285 56176
rect 15340 55124 15380 56335
rect 15532 55553 15572 57436
rect 15724 57392 15764 57595
rect 15628 57352 15764 57392
rect 15628 57056 15668 57352
rect 15628 56225 15668 57016
rect 15723 57056 15765 57065
rect 15723 57016 15724 57056
rect 15764 57016 15765 57056
rect 15723 57007 15765 57016
rect 15724 56922 15764 57007
rect 15820 56888 15860 58024
rect 15915 57476 15957 57485
rect 15915 57436 15916 57476
rect 15956 57436 15957 57476
rect 15915 57427 15957 57436
rect 15916 57056 15956 57427
rect 16011 57140 16053 57149
rect 16011 57100 16012 57140
rect 16052 57100 16053 57140
rect 16011 57091 16053 57100
rect 15916 57007 15956 57016
rect 16012 57006 16052 57091
rect 15820 56848 15956 56888
rect 15723 56636 15765 56645
rect 15723 56596 15724 56636
rect 15764 56596 15765 56636
rect 15723 56587 15765 56596
rect 15724 56384 15764 56587
rect 15627 56216 15669 56225
rect 15627 56176 15628 56216
rect 15668 56176 15669 56216
rect 15627 56167 15669 56176
rect 15531 55544 15573 55553
rect 15531 55504 15532 55544
rect 15572 55504 15573 55544
rect 15531 55495 15573 55504
rect 15340 55084 15572 55124
rect 15339 54956 15381 54965
rect 15339 54916 15340 54956
rect 15380 54916 15381 54956
rect 15339 54907 15381 54916
rect 15244 53346 15284 53355
rect 15244 52697 15284 53306
rect 15052 52648 15188 52688
rect 15243 52688 15285 52697
rect 15243 52648 15244 52688
rect 15284 52648 15285 52688
rect 15052 52445 15092 52648
rect 15243 52639 15285 52648
rect 15148 52520 15188 52529
rect 15051 52436 15093 52445
rect 15051 52396 15052 52436
rect 15092 52396 15093 52436
rect 15051 52387 15093 52396
rect 15052 51773 15092 52387
rect 15148 52361 15188 52480
rect 15243 52520 15285 52529
rect 15243 52480 15244 52520
rect 15284 52480 15285 52520
rect 15243 52471 15285 52480
rect 15244 52386 15284 52471
rect 15147 52352 15189 52361
rect 15147 52312 15148 52352
rect 15188 52312 15189 52352
rect 15147 52303 15189 52312
rect 15051 51764 15093 51773
rect 15051 51724 15052 51764
rect 15092 51724 15093 51764
rect 15051 51715 15093 51724
rect 15147 51680 15189 51689
rect 15147 51640 15148 51680
rect 15188 51640 15189 51680
rect 15147 51631 15189 51640
rect 14860 51388 14996 51428
rect 14763 51176 14805 51185
rect 14763 51136 14764 51176
rect 14804 51136 14805 51176
rect 14763 51127 14805 51136
rect 14668 50959 14708 50968
rect 14764 51008 14804 51127
rect 14764 50959 14804 50968
rect 14284 50548 14612 50588
rect 14140 50326 14228 50336
rect 14180 50296 14228 50326
rect 14284 50420 14324 50429
rect 14140 50277 14180 50286
rect 14187 50168 14229 50177
rect 13996 50128 14132 50168
rect 13995 49496 14037 49505
rect 13995 49456 13996 49496
rect 14036 49456 14037 49496
rect 13995 49447 14037 49456
rect 13996 49362 14036 49447
rect 13995 49160 14037 49169
rect 13995 49120 13996 49160
rect 14036 49120 14037 49160
rect 13995 49111 14037 49120
rect 13996 48077 14036 49111
rect 13995 48068 14037 48077
rect 13995 48028 13996 48068
rect 14036 48028 14037 48068
rect 13995 48019 14037 48028
rect 14092 42785 14132 50128
rect 14187 50128 14188 50168
rect 14228 50128 14229 50168
rect 14187 50119 14229 50128
rect 14188 47321 14228 50119
rect 14284 50093 14324 50380
rect 14379 50336 14421 50345
rect 14476 50336 14516 50345
rect 14379 50296 14380 50336
rect 14420 50296 14476 50336
rect 14379 50287 14421 50296
rect 14476 50287 14516 50296
rect 14283 50084 14325 50093
rect 14283 50044 14284 50084
rect 14324 50044 14325 50084
rect 14283 50035 14325 50044
rect 14284 49505 14324 50035
rect 14283 49496 14325 49505
rect 14283 49456 14284 49496
rect 14324 49456 14325 49496
rect 14283 49447 14325 49456
rect 14380 49412 14420 50287
rect 14572 50093 14612 50548
rect 14571 50084 14613 50093
rect 14571 50044 14572 50084
rect 14612 50044 14613 50084
rect 14571 50035 14613 50044
rect 14572 49841 14612 50035
rect 14571 49832 14613 49841
rect 14571 49792 14572 49832
rect 14612 49792 14613 49832
rect 14571 49783 14613 49792
rect 14860 49580 14900 51388
rect 15051 51176 15093 51185
rect 15051 51136 15052 51176
rect 15092 51136 15093 51176
rect 15051 51127 15093 51136
rect 14956 51017 14996 51102
rect 14955 51008 14997 51017
rect 14955 50968 14956 51008
rect 14996 50968 14997 51008
rect 14955 50959 14997 50968
rect 15052 51008 15092 51127
rect 15052 50959 15092 50968
rect 15148 51008 15188 51631
rect 15340 51353 15380 54907
rect 15436 54872 15476 54883
rect 15436 54797 15476 54832
rect 15435 54788 15477 54797
rect 15435 54748 15436 54788
rect 15476 54748 15477 54788
rect 15435 54739 15477 54748
rect 15435 53444 15477 53453
rect 15435 53404 15436 53444
rect 15476 53404 15477 53444
rect 15435 53395 15477 53404
rect 15436 53310 15476 53395
rect 15532 52865 15572 55084
rect 15627 53360 15669 53369
rect 15627 53320 15628 53360
rect 15668 53320 15669 53360
rect 15627 53311 15669 53320
rect 15628 53226 15668 53311
rect 15724 53285 15764 56344
rect 15819 56300 15861 56309
rect 15819 56260 15820 56300
rect 15860 56260 15861 56300
rect 15819 56251 15861 56260
rect 15820 56166 15860 56251
rect 15819 55796 15861 55805
rect 15819 55756 15820 55796
rect 15860 55756 15861 55796
rect 15819 55747 15861 55756
rect 15820 55544 15860 55747
rect 15820 55495 15860 55504
rect 15819 55376 15861 55385
rect 15819 55336 15820 55376
rect 15860 55336 15861 55376
rect 15819 55327 15861 55336
rect 15723 53276 15765 53285
rect 15723 53236 15724 53276
rect 15764 53236 15765 53276
rect 15723 53227 15765 53236
rect 15724 53108 15764 53117
rect 15628 53068 15724 53108
rect 15531 52856 15573 52865
rect 15531 52816 15532 52856
rect 15572 52816 15573 52856
rect 15531 52807 15573 52816
rect 15532 52688 15572 52697
rect 15339 51344 15381 51353
rect 15339 51304 15340 51344
rect 15380 51304 15381 51344
rect 15339 51295 15381 51304
rect 15436 51269 15476 51354
rect 15435 51260 15477 51269
rect 15435 51220 15436 51260
rect 15476 51220 15477 51260
rect 15435 51211 15477 51220
rect 15532 51017 15572 52648
rect 15148 50959 15188 50968
rect 15244 51008 15284 51017
rect 15436 51008 15476 51017
rect 15284 50968 15436 51008
rect 15244 50959 15284 50968
rect 15436 50959 15476 50968
rect 15531 51008 15573 51017
rect 15531 50968 15532 51008
rect 15572 50968 15573 51008
rect 15531 50959 15573 50968
rect 15628 51008 15668 53068
rect 15724 53059 15764 53068
rect 15723 52520 15765 52529
rect 15723 52480 15724 52520
rect 15764 52480 15765 52520
rect 15723 52471 15765 52480
rect 15724 51941 15764 52471
rect 15820 52016 15860 55327
rect 15916 55049 15956 56848
rect 16011 56300 16053 56309
rect 16011 56260 16012 56300
rect 16052 56260 16053 56300
rect 16011 56251 16053 56260
rect 16012 55469 16052 56251
rect 16011 55460 16053 55469
rect 16011 55420 16012 55460
rect 16052 55420 16053 55460
rect 16011 55411 16053 55420
rect 16108 55133 16148 58360
rect 16203 57224 16245 57233
rect 16203 57184 16204 57224
rect 16244 57184 16245 57224
rect 16203 57175 16245 57184
rect 16204 57056 16244 57175
rect 16204 56729 16244 57016
rect 16203 56720 16245 56729
rect 16203 56680 16204 56720
rect 16244 56680 16245 56720
rect 16203 56671 16245 56680
rect 16300 56552 16340 60796
rect 16396 59753 16436 69607
rect 16492 69166 16532 69784
rect 16492 69117 16532 69126
rect 16492 65372 16532 65381
rect 16492 64625 16532 65332
rect 16491 64616 16533 64625
rect 16491 64576 16492 64616
rect 16532 64576 16533 64616
rect 16491 64567 16533 64576
rect 16491 63020 16533 63029
rect 16491 62980 16492 63020
rect 16532 62980 16533 63020
rect 16491 62971 16533 62980
rect 16395 59744 16437 59753
rect 16395 59704 16396 59744
rect 16436 59704 16437 59744
rect 16395 59695 16437 59704
rect 16395 59576 16437 59585
rect 16395 59536 16396 59576
rect 16436 59536 16437 59576
rect 16395 59527 16437 59536
rect 16396 59442 16436 59527
rect 16492 57989 16532 62971
rect 16588 60332 16628 70036
rect 16684 70027 16724 70036
rect 16876 69665 16916 72883
rect 16875 69656 16917 69665
rect 16875 69616 16876 69656
rect 16916 69616 16917 69656
rect 16875 69607 16917 69616
rect 16875 69488 16917 69497
rect 16875 69448 16876 69488
rect 16916 69448 16917 69488
rect 16875 69439 16917 69448
rect 16684 68984 16724 68993
rect 16724 68944 16820 68984
rect 16684 68935 16724 68944
rect 16683 66968 16725 66977
rect 16683 66928 16684 66968
rect 16724 66928 16725 66968
rect 16683 66919 16725 66928
rect 16684 66834 16724 66919
rect 16684 66128 16724 66137
rect 16684 65969 16724 66088
rect 16683 65960 16725 65969
rect 16683 65920 16684 65960
rect 16724 65920 16725 65960
rect 16683 65911 16725 65920
rect 16683 65288 16725 65297
rect 16683 65248 16684 65288
rect 16724 65248 16725 65288
rect 16683 65239 16725 65248
rect 16684 65154 16724 65239
rect 16684 62348 16724 62357
rect 16684 61601 16724 62308
rect 16780 62021 16820 68944
rect 16876 63281 16916 69439
rect 16972 66800 17012 74479
rect 17068 66893 17108 75149
rect 17259 73016 17301 73025
rect 17259 72971 17260 73016
rect 17300 72971 17301 73016
rect 17259 72967 17301 72971
rect 17260 72881 17300 72967
rect 17356 72764 17396 75571
rect 17548 73193 17588 76672
rect 17644 76544 17684 76553
rect 17684 76504 17780 76544
rect 17644 76495 17684 76504
rect 17644 75788 17684 75797
rect 17644 75629 17684 75748
rect 17643 75620 17685 75629
rect 17643 75580 17644 75620
rect 17684 75580 17685 75620
rect 17643 75571 17685 75580
rect 17740 75452 17780 76504
rect 17836 76049 17876 78100
rect 17931 78100 17932 78140
rect 17972 78100 17973 78140
rect 17931 78091 17973 78100
rect 18123 78140 18165 78149
rect 18123 78100 18124 78140
rect 18164 78100 18165 78140
rect 18123 78091 18165 78100
rect 17932 77720 17972 78091
rect 18220 77897 18260 78931
rect 18508 78910 18548 78931
rect 18604 78569 18644 81031
rect 18891 80660 18933 80669
rect 18891 80620 18892 80660
rect 18932 80620 18933 80660
rect 18891 80611 18933 80620
rect 18892 80576 18932 80611
rect 18892 80525 18932 80536
rect 18700 80324 18740 80333
rect 18603 78560 18645 78569
rect 18603 78520 18604 78560
rect 18644 78520 18645 78560
rect 18603 78511 18645 78520
rect 18507 78476 18549 78485
rect 18507 78436 18508 78476
rect 18548 78436 18549 78476
rect 18507 78427 18549 78436
rect 18508 78342 18548 78427
rect 18603 78392 18645 78401
rect 18603 78352 18604 78392
rect 18644 78352 18645 78392
rect 18700 78392 18740 80284
rect 18808 80156 19176 80165
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 18808 80107 19176 80116
rect 19179 79988 19221 79997
rect 19179 79948 19180 79988
rect 19220 79948 19221 79988
rect 19179 79939 19221 79948
rect 18892 79736 18932 79745
rect 18796 79696 18892 79736
rect 18796 79409 18836 79696
rect 18892 79687 18932 79696
rect 18987 79736 19029 79745
rect 18987 79696 18988 79736
rect 19028 79696 19029 79736
rect 18987 79687 19029 79696
rect 18988 79602 19028 79687
rect 18795 79400 18837 79409
rect 18795 79360 18796 79400
rect 18836 79360 18837 79400
rect 18795 79351 18837 79360
rect 19180 79325 19220 79939
rect 19276 79568 19316 81703
rect 19564 81509 19604 83140
rect 20044 83012 20084 83140
rect 20044 82963 20084 82972
rect 20236 82844 20276 82853
rect 19756 82760 19796 82771
rect 19756 82685 19796 82720
rect 19755 82676 19797 82685
rect 19755 82636 19756 82676
rect 19796 82636 19797 82676
rect 19755 82627 19797 82636
rect 19659 81836 19701 81845
rect 19659 81796 19660 81836
rect 19700 81796 19701 81836
rect 19659 81787 19701 81796
rect 19563 81500 19605 81509
rect 19563 81460 19564 81500
rect 19604 81460 19605 81500
rect 19563 81451 19605 81460
rect 19468 79829 19508 79850
rect 19467 79820 19509 79829
rect 19467 79780 19468 79820
rect 19508 79780 19509 79820
rect 19467 79771 19509 79780
rect 19468 79755 19508 79771
rect 19372 79736 19412 79745
rect 19468 79706 19508 79715
rect 19372 79652 19412 79696
rect 19372 79612 19508 79652
rect 19276 79528 19412 79568
rect 19179 79316 19221 79325
rect 19179 79276 19180 79316
rect 19220 79276 19221 79316
rect 19179 79267 19221 79276
rect 19372 79073 19412 79528
rect 19468 79493 19508 79612
rect 19467 79484 19509 79493
rect 19467 79444 19468 79484
rect 19508 79444 19509 79484
rect 19467 79435 19509 79444
rect 19563 79400 19605 79409
rect 19563 79360 19564 79400
rect 19604 79360 19605 79400
rect 19563 79351 19605 79360
rect 19371 79064 19413 79073
rect 19371 79024 19372 79064
rect 19412 79024 19413 79064
rect 19371 79015 19413 79024
rect 19468 79064 19508 79073
rect 19564 79064 19604 79351
rect 19508 79024 19604 79064
rect 18891 78980 18933 78989
rect 18891 78940 18892 78980
rect 18932 78940 18933 78980
rect 18891 78931 18933 78940
rect 18988 78980 19028 78991
rect 18892 78846 18932 78931
rect 18988 78905 19028 78940
rect 18987 78896 19029 78905
rect 18987 78856 18988 78896
rect 19028 78856 19029 78896
rect 18987 78847 19029 78856
rect 19275 78896 19317 78905
rect 19275 78856 19276 78896
rect 19316 78856 19317 78896
rect 19275 78847 19317 78856
rect 18808 78644 19176 78653
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 18808 78595 19176 78604
rect 18700 78352 18836 78392
rect 18603 78343 18645 78352
rect 18316 78308 18356 78317
rect 18219 77888 18261 77897
rect 18219 77848 18220 77888
rect 18260 77848 18261 77888
rect 18219 77839 18261 77848
rect 17932 77671 17972 77680
rect 18219 77720 18261 77729
rect 18219 77680 18220 77720
rect 18260 77680 18261 77720
rect 18219 77671 18261 77680
rect 18124 77468 18164 77477
rect 18028 77428 18124 77468
rect 17931 76880 17973 76889
rect 17931 76840 17932 76880
rect 17972 76840 17973 76880
rect 17931 76831 17973 76840
rect 17932 76746 17972 76831
rect 18028 76721 18068 77428
rect 18124 77419 18164 77428
rect 18123 76796 18165 76805
rect 18123 76756 18124 76796
rect 18164 76756 18165 76796
rect 18123 76747 18165 76756
rect 18027 76712 18069 76721
rect 18027 76672 18028 76712
rect 18068 76672 18069 76712
rect 18027 76663 18069 76672
rect 18124 76662 18164 76747
rect 17835 76040 17877 76049
rect 17835 76000 17836 76040
rect 17876 76000 17877 76040
rect 17835 75991 17877 76000
rect 18027 76040 18069 76049
rect 18027 76000 18028 76040
rect 18068 76000 18069 76040
rect 18027 75991 18069 76000
rect 17644 75412 17780 75452
rect 17836 75788 17876 75797
rect 17547 73184 17589 73193
rect 17547 73144 17548 73184
rect 17588 73144 17589 73184
rect 17547 73135 17589 73144
rect 17644 73109 17684 75412
rect 17740 75209 17780 75294
rect 17739 75200 17781 75209
rect 17739 75160 17740 75200
rect 17780 75160 17781 75200
rect 17739 75151 17781 75160
rect 17739 75032 17781 75041
rect 17739 74992 17740 75032
rect 17780 74992 17781 75032
rect 17739 74983 17781 74992
rect 17452 73100 17492 73109
rect 17452 72941 17492 73060
rect 17643 73100 17685 73109
rect 17643 73060 17644 73100
rect 17684 73060 17685 73100
rect 17643 73051 17685 73060
rect 17451 72932 17493 72941
rect 17451 72892 17452 72932
rect 17492 72892 17493 72932
rect 17451 72883 17493 72892
rect 17547 72848 17589 72857
rect 17547 72808 17548 72848
rect 17588 72808 17589 72848
rect 17547 72799 17589 72808
rect 17260 72724 17396 72764
rect 17260 72190 17300 72724
rect 17260 72141 17300 72150
rect 17451 72008 17493 72017
rect 17451 71968 17452 72008
rect 17492 71968 17493 72008
rect 17451 71959 17493 71968
rect 17452 71874 17492 71959
rect 17163 71504 17205 71513
rect 17163 71464 17164 71504
rect 17204 71464 17205 71504
rect 17163 71455 17205 71464
rect 17451 71504 17493 71513
rect 17451 71464 17452 71504
rect 17492 71464 17493 71504
rect 17451 71455 17493 71464
rect 17164 68489 17204 71455
rect 17452 71370 17492 71455
rect 17548 71009 17588 72799
rect 17644 71252 17684 71261
rect 17259 71000 17301 71009
rect 17259 70960 17260 71000
rect 17300 70960 17301 71000
rect 17259 70951 17301 70960
rect 17547 71000 17589 71009
rect 17547 70960 17548 71000
rect 17588 70960 17589 71000
rect 17547 70951 17589 70960
rect 17260 70664 17300 70951
rect 17644 70748 17684 71212
rect 17548 70708 17684 70748
rect 17452 70664 17492 70673
rect 17260 70624 17452 70664
rect 17163 68480 17205 68489
rect 17163 68440 17164 68480
rect 17204 68440 17205 68480
rect 17163 68431 17205 68440
rect 17260 68312 17300 70624
rect 17452 70615 17492 70624
rect 17451 70328 17493 70337
rect 17451 70288 17452 70328
rect 17492 70288 17493 70328
rect 17548 70328 17588 70708
rect 17643 70580 17685 70589
rect 17643 70540 17644 70580
rect 17684 70540 17685 70580
rect 17643 70531 17685 70540
rect 17644 70446 17684 70531
rect 17740 70496 17780 74983
rect 17836 73529 17876 75748
rect 18028 74537 18068 75991
rect 18220 75713 18260 77671
rect 18316 77393 18356 78268
rect 18411 78308 18453 78317
rect 18411 78268 18412 78308
rect 18452 78268 18453 78308
rect 18411 78259 18453 78268
rect 18315 77384 18357 77393
rect 18315 77344 18316 77384
rect 18356 77344 18357 77384
rect 18315 77335 18357 77344
rect 18316 77250 18356 77335
rect 18315 77132 18357 77141
rect 18315 77092 18316 77132
rect 18356 77092 18357 77132
rect 18315 77083 18357 77092
rect 18219 75704 18261 75713
rect 18219 75664 18220 75704
rect 18260 75664 18261 75704
rect 18219 75655 18261 75664
rect 18219 75368 18261 75377
rect 18219 75328 18220 75368
rect 18260 75328 18261 75368
rect 18219 75319 18261 75328
rect 18220 75214 18260 75319
rect 18220 75165 18260 75174
rect 18027 74528 18069 74537
rect 18027 74488 18028 74528
rect 18068 74488 18069 74528
rect 18027 74479 18069 74488
rect 17931 74444 17973 74453
rect 17931 74404 17932 74444
rect 17972 74404 17973 74444
rect 17931 74395 17973 74404
rect 17835 73520 17877 73529
rect 17835 73480 17836 73520
rect 17876 73480 17877 73520
rect 17835 73471 17877 73480
rect 17932 70673 17972 74395
rect 18028 74394 18068 74479
rect 18220 74276 18260 74285
rect 18028 74236 18220 74276
rect 17931 70664 17973 70673
rect 17931 70624 17932 70664
rect 17972 70624 17973 70664
rect 17931 70615 17973 70624
rect 17740 70456 17972 70496
rect 17835 70328 17877 70337
rect 17548 70288 17780 70328
rect 17451 70279 17493 70288
rect 17164 68272 17300 68312
rect 17164 67640 17204 68272
rect 17356 68228 17396 68237
rect 17067 66884 17109 66893
rect 17067 66844 17068 66884
rect 17108 66844 17109 66884
rect 17067 66835 17109 66844
rect 16972 64280 17012 66760
rect 17164 66137 17204 67600
rect 17260 68188 17356 68228
rect 17163 66128 17205 66137
rect 17163 66088 17164 66128
rect 17204 66088 17205 66128
rect 17163 66079 17205 66088
rect 17164 64280 17204 66079
rect 17260 64616 17300 68188
rect 17356 68179 17396 68188
rect 17452 67649 17492 70279
rect 17740 68984 17780 70288
rect 17835 70288 17836 70328
rect 17876 70288 17877 70328
rect 17835 70279 17877 70288
rect 17836 69068 17876 70279
rect 17932 69245 17972 70456
rect 18028 69665 18068 74236
rect 18220 74227 18260 74236
rect 18123 73688 18165 73697
rect 18123 73648 18124 73688
rect 18164 73648 18165 73688
rect 18316 73688 18356 77083
rect 18412 76712 18452 78259
rect 18604 78224 18644 78343
rect 18700 78224 18740 78233
rect 18604 78184 18700 78224
rect 18700 78175 18740 78184
rect 18507 78140 18549 78149
rect 18507 78100 18508 78140
rect 18548 78100 18644 78140
rect 18507 78091 18549 78100
rect 18507 77888 18549 77897
rect 18507 77848 18508 77888
rect 18548 77848 18549 77888
rect 18507 77839 18549 77848
rect 18508 76889 18548 77839
rect 18604 77552 18644 78100
rect 18604 77477 18644 77512
rect 18603 77468 18645 77477
rect 18603 77428 18604 77468
rect 18644 77428 18645 77468
rect 18603 77419 18645 77428
rect 18604 77388 18644 77419
rect 18796 77300 18836 78352
rect 18604 77260 18836 77300
rect 18507 76880 18549 76889
rect 18507 76840 18508 76880
rect 18548 76840 18549 76880
rect 18507 76831 18549 76840
rect 18412 76663 18452 76672
rect 18508 76712 18548 76831
rect 18508 76663 18548 76672
rect 18604 76544 18644 77260
rect 18808 77132 19176 77141
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 18808 77083 19176 77092
rect 19276 76964 19316 78847
rect 18988 76924 19316 76964
rect 18699 76880 18741 76889
rect 18699 76840 18700 76880
rect 18740 76840 18741 76880
rect 18699 76831 18741 76840
rect 18891 76880 18933 76889
rect 18891 76840 18892 76880
rect 18932 76840 18933 76880
rect 18891 76831 18933 76840
rect 18508 76504 18644 76544
rect 18411 75032 18453 75041
rect 18411 74992 18412 75032
rect 18452 74992 18453 75032
rect 18411 74983 18453 74992
rect 18412 74898 18452 74983
rect 18508 74528 18548 76504
rect 18700 76292 18740 76831
rect 18892 76796 18932 76831
rect 18892 76745 18932 76756
rect 18988 76796 19028 76924
rect 18988 76747 19028 76756
rect 19371 76796 19413 76805
rect 19371 76756 19372 76796
rect 19412 76756 19413 76796
rect 19371 76747 19413 76756
rect 18508 74479 18548 74488
rect 18604 76252 18740 76292
rect 18604 74528 18644 76252
rect 19276 76040 19316 76049
rect 19276 75797 19316 76000
rect 19275 75788 19317 75797
rect 19275 75748 19276 75788
rect 19316 75748 19317 75788
rect 19275 75739 19317 75748
rect 18808 75620 19176 75629
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 18808 75571 19176 75580
rect 19372 75452 19412 76747
rect 19468 76712 19508 79024
rect 19660 78812 19700 81787
rect 19756 79913 19796 82627
rect 20236 82592 20276 82804
rect 20236 82552 20564 82592
rect 20048 82424 20416 82433
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20048 82375 20416 82384
rect 19852 82088 19892 82097
rect 19852 81920 19892 82048
rect 19852 81880 19988 81920
rect 19948 81248 19988 81880
rect 20043 81836 20085 81845
rect 20043 81796 20044 81836
rect 20084 81796 20085 81836
rect 20043 81787 20085 81796
rect 20044 81702 20084 81787
rect 20524 81425 20564 82552
rect 20523 81416 20565 81425
rect 20523 81376 20524 81416
rect 20564 81376 20565 81416
rect 20523 81367 20565 81376
rect 20044 81248 20084 81257
rect 19948 81208 20044 81248
rect 19948 80669 19988 81208
rect 20044 81199 20084 81208
rect 20236 81080 20276 81089
rect 20276 81040 20564 81080
rect 20236 81031 20276 81040
rect 20048 80912 20416 80921
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20048 80863 20416 80872
rect 19947 80660 19989 80669
rect 19947 80620 19948 80660
rect 19988 80620 19989 80660
rect 19947 80611 19989 80620
rect 20140 80534 20180 80543
rect 20140 80417 20180 80494
rect 20139 80408 20181 80417
rect 20139 80368 20140 80408
rect 20180 80368 20181 80408
rect 20139 80359 20181 80368
rect 19851 80324 19893 80333
rect 19851 80284 19852 80324
rect 19892 80284 19893 80324
rect 19851 80275 19893 80284
rect 19755 79904 19797 79913
rect 19755 79864 19756 79904
rect 19796 79864 19797 79904
rect 19755 79855 19797 79864
rect 19756 79736 19796 79855
rect 19756 79687 19796 79696
rect 19852 79736 19892 80275
rect 19947 79820 19989 79829
rect 19947 79780 19948 79820
rect 19988 79780 19989 79820
rect 19947 79771 19989 79780
rect 19852 79687 19892 79696
rect 19948 79736 19988 79771
rect 19948 79685 19988 79696
rect 20044 79568 20084 79577
rect 19948 79528 20044 79568
rect 19948 79241 19988 79528
rect 20044 79519 20084 79528
rect 20048 79400 20416 79409
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20048 79351 20416 79360
rect 19947 79232 19989 79241
rect 19947 79192 19948 79232
rect 19988 79192 19989 79232
rect 20524 79232 20564 81040
rect 20620 80501 20660 84316
rect 20619 80492 20661 80501
rect 20619 80452 20620 80492
rect 20660 80452 20661 80492
rect 20619 80443 20661 80452
rect 20524 79192 20756 79232
rect 19947 79183 19989 79192
rect 20140 79148 20180 79157
rect 20180 79108 20660 79148
rect 20140 79099 20180 79108
rect 19947 79064 19989 79073
rect 19947 79019 19948 79064
rect 19988 79019 19989 79064
rect 19947 79015 19989 79019
rect 19948 78929 19988 79015
rect 19660 78772 20084 78812
rect 19948 78224 19988 78233
rect 19852 78184 19948 78224
rect 19755 77888 19797 77897
rect 19755 77848 19756 77888
rect 19796 77848 19797 77888
rect 19755 77839 19797 77848
rect 19563 77300 19605 77309
rect 19563 77260 19564 77300
rect 19604 77260 19605 77300
rect 19563 77251 19605 77260
rect 19468 76663 19508 76672
rect 18508 73688 18548 73697
rect 18316 73648 18508 73688
rect 18123 73639 18165 73648
rect 18124 73193 18164 73639
rect 18316 73520 18356 73529
rect 18123 73184 18165 73193
rect 18123 73144 18124 73184
rect 18164 73144 18165 73184
rect 18123 73135 18165 73144
rect 18124 72857 18164 73135
rect 18316 73100 18356 73480
rect 18412 73445 18452 73648
rect 18508 73639 18548 73648
rect 18507 73520 18549 73529
rect 18507 73480 18508 73520
rect 18548 73480 18549 73520
rect 18507 73471 18549 73480
rect 18411 73436 18453 73445
rect 18411 73396 18412 73436
rect 18452 73396 18453 73436
rect 18411 73387 18453 73396
rect 18220 73060 18356 73100
rect 18123 72848 18165 72857
rect 18123 72808 18124 72848
rect 18164 72808 18165 72848
rect 18123 72799 18165 72808
rect 18123 70496 18165 70505
rect 18123 70456 18124 70496
rect 18164 70456 18165 70496
rect 18123 70447 18165 70456
rect 18027 69656 18069 69665
rect 18027 69616 18028 69656
rect 18068 69616 18069 69656
rect 18027 69607 18069 69616
rect 17931 69236 17973 69245
rect 17931 69196 17932 69236
rect 17972 69196 17973 69236
rect 17931 69187 17973 69196
rect 17836 69028 17972 69068
rect 17740 68944 17876 68984
rect 17643 68480 17685 68489
rect 17643 68440 17644 68480
rect 17684 68440 17685 68480
rect 17643 68431 17685 68440
rect 17451 67640 17493 67649
rect 17451 67600 17452 67640
rect 17492 67600 17493 67640
rect 17451 67591 17493 67600
rect 17356 67472 17396 67481
rect 17356 65456 17396 67432
rect 17644 66305 17684 68431
rect 17836 66968 17876 68944
rect 17932 67640 17972 69028
rect 18124 68480 18164 70447
rect 18220 69992 18260 73060
rect 18412 73016 18452 73025
rect 18316 72976 18412 73016
rect 18316 71504 18356 72976
rect 18412 72967 18452 72976
rect 18508 72176 18548 73471
rect 18508 72127 18548 72136
rect 18604 72176 18644 74488
rect 18988 75412 19412 75452
rect 18988 74528 19028 75412
rect 18988 74479 19028 74488
rect 19084 74444 19124 74453
rect 19084 74285 19124 74404
rect 19083 74276 19125 74285
rect 19083 74236 19084 74276
rect 19124 74236 19125 74276
rect 19083 74227 19125 74236
rect 19275 74276 19317 74285
rect 19275 74236 19276 74276
rect 19316 74236 19317 74276
rect 19275 74227 19317 74236
rect 18808 74108 19176 74117
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 18808 74059 19176 74068
rect 18699 73436 18741 73445
rect 18699 73396 18700 73436
rect 18740 73396 18741 73436
rect 18699 73387 18741 73396
rect 18604 72127 18644 72136
rect 18316 71261 18356 71464
rect 18603 71336 18645 71345
rect 18603 71296 18604 71336
rect 18644 71296 18645 71336
rect 18603 71287 18645 71296
rect 18315 71252 18357 71261
rect 18315 71212 18316 71252
rect 18356 71212 18357 71252
rect 18315 71203 18357 71212
rect 18508 70664 18548 70675
rect 18508 70505 18548 70624
rect 18507 70496 18549 70505
rect 18507 70456 18508 70496
rect 18548 70456 18549 70496
rect 18507 70447 18549 70456
rect 18604 70328 18644 71287
rect 18700 70337 18740 73387
rect 18808 72596 19176 72605
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 18808 72547 19176 72556
rect 19084 72260 19124 72269
rect 19276 72260 19316 74227
rect 19124 72220 19316 72260
rect 19084 72211 19124 72220
rect 18988 72176 19028 72187
rect 18988 72101 19028 72136
rect 19372 72101 19412 75412
rect 19564 75200 19604 77251
rect 19659 76292 19701 76301
rect 19659 76252 19660 76292
rect 19700 76252 19701 76292
rect 19659 76243 19701 76252
rect 19660 76208 19700 76243
rect 19660 76157 19700 76168
rect 19659 75704 19701 75713
rect 19659 75664 19660 75704
rect 19700 75664 19701 75704
rect 19659 75655 19701 75664
rect 19468 75160 19604 75200
rect 18987 72092 19029 72101
rect 18987 72052 18988 72092
rect 19028 72052 19029 72092
rect 18987 72043 19029 72052
rect 19371 72092 19413 72101
rect 19371 72052 19372 72092
rect 19412 72052 19413 72092
rect 19371 72043 19413 72052
rect 18808 71084 19176 71093
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 18808 71035 19176 71044
rect 19371 70496 19413 70505
rect 19371 70456 19372 70496
rect 19412 70456 19413 70496
rect 19371 70447 19413 70456
rect 18508 70288 18644 70328
rect 18699 70328 18741 70337
rect 18699 70288 18700 70328
rect 18740 70288 18741 70328
rect 18220 69943 18260 69952
rect 18316 69992 18356 70001
rect 18508 69992 18548 70288
rect 18699 70279 18741 70288
rect 18700 69992 18740 70001
rect 18356 69952 18452 69992
rect 18316 69943 18356 69952
rect 18315 69656 18357 69665
rect 18315 69616 18316 69656
rect 18356 69616 18357 69656
rect 18315 69607 18357 69616
rect 18316 69152 18356 69607
rect 18316 69103 18356 69112
rect 18412 69152 18452 69952
rect 18508 69952 18700 69992
rect 18508 69320 18548 69952
rect 18700 69943 18740 69952
rect 18795 69992 18837 70001
rect 18795 69952 18796 69992
rect 18836 69952 18837 69992
rect 18795 69943 18837 69952
rect 19276 69992 19316 70001
rect 18796 69740 18836 69943
rect 18700 69700 18836 69740
rect 18700 69404 18740 69700
rect 18808 69572 19176 69581
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 18808 69523 19176 69532
rect 19276 69404 19316 69952
rect 18700 69364 18932 69404
rect 18508 69280 18836 69320
rect 18796 69152 18836 69280
rect 18892 69236 18932 69364
rect 18892 69187 18932 69196
rect 19180 69364 19316 69404
rect 19180 69161 19220 69364
rect 19372 69320 19412 70447
rect 19468 69833 19508 75160
rect 19564 74528 19604 74537
rect 19660 74528 19700 75655
rect 19604 74488 19700 74528
rect 19564 72176 19604 74488
rect 19659 74360 19701 74369
rect 19659 74320 19660 74360
rect 19700 74320 19701 74360
rect 19659 74311 19701 74320
rect 19564 72127 19604 72136
rect 19660 73016 19700 74311
rect 19756 73856 19796 77839
rect 19852 77552 19892 78184
rect 19948 78175 19988 78184
rect 20044 78056 20084 78772
rect 20140 78065 20180 78150
rect 19852 76049 19892 77512
rect 19948 78016 20084 78056
rect 20139 78056 20181 78065
rect 20139 78016 20140 78056
rect 20180 78016 20181 78056
rect 19948 76726 19988 78016
rect 20139 78007 20181 78016
rect 20048 77888 20416 77897
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20048 77839 20416 77848
rect 20044 77309 20084 77394
rect 20043 77300 20085 77309
rect 20043 77260 20044 77300
rect 20084 77260 20085 77300
rect 20043 77251 20085 77260
rect 20043 77132 20085 77141
rect 20043 77092 20044 77132
rect 20084 77092 20085 77132
rect 20043 77083 20085 77092
rect 19948 76677 19988 76686
rect 20044 76628 20084 77083
rect 19948 76588 20084 76628
rect 19851 76040 19893 76049
rect 19851 76000 19852 76040
rect 19892 76000 19893 76040
rect 19851 75991 19893 76000
rect 19948 74696 19988 76588
rect 20140 76553 20180 76638
rect 20139 76544 20181 76553
rect 20139 76504 20140 76544
rect 20180 76504 20181 76544
rect 20139 76495 20181 76504
rect 20048 76376 20416 76385
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20048 76327 20416 76336
rect 20043 76208 20085 76217
rect 20043 76168 20044 76208
rect 20084 76168 20085 76208
rect 20043 76159 20085 76168
rect 20044 76074 20084 76159
rect 20236 75956 20276 75965
rect 20140 75368 20180 75377
rect 20236 75368 20276 75916
rect 20180 75328 20276 75368
rect 20140 75300 20180 75328
rect 20044 75041 20084 75126
rect 20043 75032 20085 75041
rect 20043 74992 20044 75032
rect 20084 74992 20085 75032
rect 20043 74983 20085 74992
rect 20048 74864 20416 74873
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20048 74815 20416 74824
rect 19948 74656 20084 74696
rect 20044 74523 20084 74656
rect 20235 74612 20277 74621
rect 20235 74572 20236 74612
rect 20276 74572 20277 74612
rect 20235 74563 20277 74572
rect 20044 74474 20084 74483
rect 20236 74478 20276 74563
rect 19756 73816 19892 73856
rect 19755 73688 19797 73697
rect 19755 73648 19756 73688
rect 19796 73648 19797 73688
rect 19755 73639 19797 73648
rect 19756 73554 19796 73639
rect 19852 73193 19892 73816
rect 19948 73520 19988 73529
rect 19851 73184 19893 73193
rect 19851 73144 19852 73184
rect 19892 73144 19893 73184
rect 19851 73135 19893 73144
rect 19660 71513 19700 72976
rect 19851 72764 19893 72773
rect 19851 72724 19852 72764
rect 19892 72724 19893 72764
rect 19851 72715 19893 72724
rect 19852 72630 19892 72715
rect 19564 71504 19604 71513
rect 19564 71009 19604 71464
rect 19659 71504 19701 71513
rect 19948 71504 19988 73480
rect 20048 73352 20416 73361
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20048 73303 20416 73312
rect 20043 73184 20085 73193
rect 20043 73144 20044 73184
rect 20084 73144 20085 73184
rect 20043 73135 20085 73144
rect 20044 72190 20084 73135
rect 20620 72512 20660 79108
rect 20716 77141 20756 79192
rect 20715 77132 20757 77141
rect 20715 77092 20716 77132
rect 20756 77092 20757 77132
rect 20715 77083 20757 77092
rect 21291 74612 21333 74621
rect 21291 74572 21292 74612
rect 21332 74572 21333 74612
rect 21291 74563 21333 74572
rect 21099 72512 21141 72521
rect 20620 72472 20756 72512
rect 20044 72141 20084 72150
rect 20236 72008 20276 72017
rect 20276 71968 20564 72008
rect 20236 71959 20276 71968
rect 20048 71840 20416 71849
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20048 71791 20416 71800
rect 19659 71464 19660 71504
rect 19700 71464 19701 71504
rect 19659 71455 19701 71464
rect 19852 71464 19988 71504
rect 19563 71000 19605 71009
rect 19563 70960 19564 71000
rect 19604 70960 19605 71000
rect 19563 70951 19605 70960
rect 19660 70916 19700 71455
rect 19756 71252 19796 71261
rect 19756 71093 19796 71212
rect 19755 71084 19797 71093
rect 19755 71044 19756 71084
rect 19796 71044 19797 71084
rect 19755 71035 19797 71044
rect 19660 70876 19796 70916
rect 19659 70748 19701 70757
rect 19659 70708 19660 70748
rect 19700 70708 19701 70748
rect 19659 70699 19701 70708
rect 19467 69824 19509 69833
rect 19467 69784 19468 69824
rect 19508 69784 19509 69824
rect 19467 69775 19509 69784
rect 19276 69280 19412 69320
rect 18452 69112 18548 69152
rect 18412 69103 18452 69112
rect 18412 68480 18452 68489
rect 18124 68440 18412 68480
rect 17932 67591 17972 67600
rect 18027 67640 18069 67649
rect 18027 67600 18028 67640
rect 18068 67600 18069 67640
rect 18027 67591 18069 67600
rect 17932 66968 17972 66977
rect 17836 66928 17932 66968
rect 17932 66919 17972 66928
rect 18028 66968 18068 67591
rect 18123 67136 18165 67145
rect 18123 67096 18124 67136
rect 18164 67096 18165 67136
rect 18123 67087 18165 67096
rect 18028 66919 18068 66928
rect 18124 66800 18164 67087
rect 18028 66760 18164 66800
rect 18316 66800 18356 68440
rect 18412 68431 18452 68440
rect 18411 68228 18453 68237
rect 18508 68228 18548 69112
rect 18796 68816 18836 69112
rect 19179 69152 19221 69161
rect 19179 69112 19180 69152
rect 19220 69112 19221 69152
rect 19179 69103 19221 69112
rect 18411 68188 18412 68228
rect 18452 68188 18548 68228
rect 18700 68776 18836 68816
rect 18411 68179 18453 68188
rect 18412 67724 18452 68179
rect 18412 66968 18452 67684
rect 18412 66919 18452 66928
rect 18508 67640 18548 67649
rect 18700 67640 18740 68776
rect 18808 68060 19176 68069
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 18808 68011 19176 68020
rect 18548 67600 18740 67640
rect 18988 67640 19028 67649
rect 18508 66968 18548 67600
rect 18603 67304 18645 67313
rect 18603 67264 18604 67304
rect 18644 67264 18645 67304
rect 18603 67255 18645 67264
rect 18508 66919 18548 66928
rect 18316 66760 18452 66800
rect 17643 66296 17685 66305
rect 17643 66256 17644 66296
rect 17684 66256 17685 66296
rect 17643 66247 17685 66256
rect 17931 66296 17973 66305
rect 17931 66256 17932 66296
rect 17972 66256 17973 66296
rect 17931 66247 17973 66256
rect 17932 66128 17972 66247
rect 17932 65540 17972 66088
rect 17836 65500 17972 65540
rect 17452 65456 17492 65465
rect 17356 65416 17452 65456
rect 17452 65407 17492 65416
rect 17548 65456 17588 65467
rect 17548 65381 17588 65416
rect 17547 65372 17589 65381
rect 17547 65332 17548 65372
rect 17588 65332 17684 65372
rect 17547 65323 17589 65332
rect 17548 64616 17588 64625
rect 17260 64576 17548 64616
rect 17548 64567 17588 64576
rect 17644 64616 17684 65332
rect 17644 64567 17684 64576
rect 17836 64532 17876 65500
rect 18028 65456 18068 66760
rect 18219 66212 18261 66221
rect 18219 66172 18220 66212
rect 18260 66172 18261 66212
rect 18219 66163 18261 66172
rect 18124 65960 18164 65969
rect 18124 65549 18164 65920
rect 18123 65540 18165 65549
rect 18123 65500 18124 65540
rect 18164 65500 18165 65540
rect 18123 65491 18165 65500
rect 17932 65372 17972 65381
rect 18028 65372 18068 65416
rect 18028 65332 18164 65372
rect 17932 65129 17972 65332
rect 17931 65120 17973 65129
rect 17931 65080 17932 65120
rect 17972 65080 17973 65120
rect 17931 65071 17973 65080
rect 17932 64700 17972 65071
rect 18028 64700 18068 64709
rect 17932 64660 18028 64700
rect 18028 64651 18068 64660
rect 18124 64700 18164 65332
rect 18124 64651 18164 64660
rect 17836 64492 18164 64532
rect 16972 64240 17108 64280
rect 17164 64240 17588 64280
rect 16875 63272 16917 63281
rect 16875 63232 16876 63272
rect 16916 63232 16917 63272
rect 16875 63223 16917 63232
rect 16875 62600 16917 62609
rect 16875 62560 16876 62600
rect 16916 62560 16917 62600
rect 16875 62551 16917 62560
rect 16876 62466 16916 62551
rect 16779 62012 16821 62021
rect 16779 61972 16780 62012
rect 16820 61972 16821 62012
rect 16779 61963 16821 61972
rect 16683 61592 16725 61601
rect 16683 61552 16684 61592
rect 16724 61552 16725 61592
rect 16683 61543 16725 61552
rect 16971 61004 17013 61013
rect 16971 60964 16972 61004
rect 17012 60964 17013 61004
rect 16971 60955 17013 60964
rect 16875 60500 16917 60509
rect 16875 60460 16876 60500
rect 16916 60460 16917 60500
rect 16875 60451 16917 60460
rect 16588 60292 16724 60332
rect 16588 60164 16628 60173
rect 16588 59501 16628 60124
rect 16587 59492 16629 59501
rect 16587 59452 16588 59492
rect 16628 59452 16629 59492
rect 16587 59443 16629 59452
rect 16684 59249 16724 60292
rect 16779 60080 16821 60089
rect 16779 60040 16780 60080
rect 16820 60040 16821 60080
rect 16779 60031 16821 60040
rect 16780 59912 16820 60031
rect 16780 59863 16820 59872
rect 16779 59744 16821 59753
rect 16779 59704 16780 59744
rect 16820 59704 16821 59744
rect 16779 59695 16821 59704
rect 16683 59240 16725 59249
rect 16683 59200 16684 59240
rect 16724 59200 16725 59240
rect 16683 59191 16725 59200
rect 16588 58568 16628 58577
rect 16780 58568 16820 59695
rect 16876 59324 16916 60451
rect 16972 60164 17012 60955
rect 16972 60115 17012 60124
rect 16972 59324 17012 59333
rect 16876 59284 16972 59324
rect 16972 59275 17012 59284
rect 16491 57980 16533 57989
rect 16491 57940 16492 57980
rect 16532 57940 16533 57980
rect 16491 57931 16533 57940
rect 16588 57737 16628 58528
rect 16684 58528 16820 58568
rect 16684 58157 16724 58528
rect 16780 58400 16820 58409
rect 16683 58148 16725 58157
rect 16683 58108 16684 58148
rect 16724 58108 16725 58148
rect 16683 58099 16725 58108
rect 16587 57728 16629 57737
rect 16587 57688 16588 57728
rect 16628 57688 16629 57728
rect 16587 57679 16629 57688
rect 16780 57233 16820 58360
rect 17068 57905 17108 64240
rect 17356 60929 17396 64240
rect 17548 63944 17588 64240
rect 17548 63895 17588 63904
rect 18124 63944 18164 64492
rect 17740 63692 17780 63701
rect 17932 63692 17972 63701
rect 17780 63652 17876 63692
rect 17740 63643 17780 63652
rect 17739 63440 17781 63449
rect 17739 63400 17740 63440
rect 17780 63400 17781 63440
rect 17739 63391 17781 63400
rect 17740 62432 17780 63391
rect 17836 63272 17876 63652
rect 17932 63449 17972 63652
rect 17931 63440 17973 63449
rect 17931 63400 17932 63440
rect 17972 63400 17973 63440
rect 17931 63391 17973 63400
rect 17836 63232 17972 63272
rect 17932 63104 17972 63232
rect 18027 63188 18069 63197
rect 18027 63148 18028 63188
rect 18068 63148 18069 63188
rect 18027 63139 18069 63148
rect 17932 63055 17972 63064
rect 18028 63104 18068 63139
rect 17932 62432 17972 62441
rect 17740 62392 17932 62432
rect 17932 62383 17972 62392
rect 18028 62432 18068 63064
rect 17547 61592 17589 61601
rect 17547 61552 17548 61592
rect 17588 61552 17589 61592
rect 17547 61543 17589 61552
rect 17548 61458 17588 61543
rect 17451 61424 17493 61433
rect 17740 61424 17780 61433
rect 17451 61384 17452 61424
rect 17492 61384 17493 61424
rect 17451 61375 17493 61384
rect 17644 61384 17740 61424
rect 17355 60920 17397 60929
rect 17355 60880 17356 60920
rect 17396 60880 17397 60920
rect 17355 60871 17397 60880
rect 17163 60752 17205 60761
rect 17163 60712 17164 60752
rect 17204 60712 17205 60752
rect 17163 60703 17205 60712
rect 17164 60332 17204 60703
rect 17164 60283 17204 60292
rect 17355 60164 17397 60173
rect 17355 60124 17356 60164
rect 17396 60124 17397 60164
rect 17355 60115 17397 60124
rect 17356 60030 17396 60115
rect 17356 59324 17396 59333
rect 17163 59240 17205 59249
rect 17163 59200 17164 59240
rect 17204 59200 17205 59240
rect 17163 59191 17205 59200
rect 17164 59106 17204 59191
rect 17259 58652 17301 58661
rect 17259 58612 17260 58652
rect 17300 58612 17301 58652
rect 17259 58603 17301 58612
rect 17260 58518 17300 58603
rect 17356 58073 17396 59284
rect 17452 58904 17492 61375
rect 17547 60920 17589 60929
rect 17547 60880 17548 60920
rect 17588 60880 17589 60920
rect 17547 60871 17589 60880
rect 17548 60786 17588 60871
rect 17547 60416 17589 60425
rect 17547 60376 17548 60416
rect 17588 60376 17589 60416
rect 17547 60367 17589 60376
rect 17548 60332 17588 60367
rect 17548 60281 17588 60292
rect 17644 59408 17684 61384
rect 17740 61375 17780 61384
rect 17740 60668 17780 60677
rect 17740 60080 17780 60628
rect 17836 60080 17876 60089
rect 17740 60040 17836 60080
rect 17836 60031 17876 60040
rect 17932 60080 17972 60089
rect 18028 60080 18068 62392
rect 18124 61760 18164 63904
rect 18220 63197 18260 66163
rect 18316 66128 18356 66137
rect 18316 65969 18356 66088
rect 18315 65960 18357 65969
rect 18315 65920 18316 65960
rect 18356 65920 18357 65960
rect 18315 65911 18357 65920
rect 18412 65792 18452 66760
rect 18316 65752 18452 65792
rect 18316 64541 18356 65752
rect 18508 65456 18548 65465
rect 18412 65416 18508 65456
rect 18412 65045 18452 65416
rect 18508 65407 18548 65416
rect 18604 65288 18644 67255
rect 18988 66968 19028 67600
rect 18988 66893 19028 66928
rect 18987 66884 19029 66893
rect 18987 66844 18988 66884
rect 19028 66844 19029 66884
rect 18987 66835 19029 66844
rect 18808 66548 19176 66557
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 18808 66499 19176 66508
rect 18987 66212 19029 66221
rect 18987 66172 18988 66212
rect 19028 66172 19029 66212
rect 18987 66163 19029 66172
rect 18988 65451 19028 66163
rect 18988 65402 19028 65411
rect 19180 65540 19220 65549
rect 18508 65248 18644 65288
rect 18411 65036 18453 65045
rect 18411 64996 18412 65036
rect 18452 64996 18453 65036
rect 18411 64987 18453 64996
rect 18315 64532 18357 64541
rect 18315 64492 18316 64532
rect 18356 64492 18357 64532
rect 18315 64483 18357 64492
rect 18316 63533 18356 64483
rect 18315 63524 18357 63533
rect 18315 63484 18316 63524
rect 18356 63484 18357 63524
rect 18315 63475 18357 63484
rect 18411 63272 18453 63281
rect 18411 63232 18412 63272
rect 18452 63232 18453 63272
rect 18411 63223 18453 63232
rect 18219 63188 18261 63197
rect 18219 63148 18220 63188
rect 18260 63148 18261 63188
rect 18219 63139 18261 63148
rect 18412 63188 18452 63223
rect 18412 62432 18452 63148
rect 18316 62392 18412 62432
rect 18124 61720 18260 61760
rect 17972 60040 18068 60080
rect 18124 61592 18164 61601
rect 18124 60920 18164 61552
rect 18220 61517 18260 61720
rect 18219 61508 18261 61517
rect 18219 61468 18220 61508
rect 18260 61468 18261 61508
rect 18219 61459 18261 61468
rect 17836 59408 17876 59417
rect 17644 59368 17836 59408
rect 17836 59359 17876 59368
rect 17932 59408 17972 60040
rect 17932 59359 17972 59368
rect 17547 59156 17589 59165
rect 17547 59116 17548 59156
rect 17588 59116 17589 59156
rect 17547 59107 17589 59116
rect 17548 59022 17588 59107
rect 17452 58864 17588 58904
rect 17451 58400 17493 58409
rect 17451 58360 17452 58400
rect 17492 58360 17493 58400
rect 17451 58351 17493 58360
rect 17452 58266 17492 58351
rect 17548 58148 17588 58864
rect 17644 58652 17684 58663
rect 17644 58577 17684 58612
rect 18124 58577 18164 60880
rect 18316 60164 18356 62392
rect 18412 62383 18452 62392
rect 18508 63188 18548 65248
rect 19180 65213 19220 65500
rect 19179 65204 19221 65213
rect 19179 65164 19180 65204
rect 19220 65164 19221 65204
rect 19179 65155 19221 65164
rect 18603 65036 18645 65045
rect 18603 64996 18604 65036
rect 18644 64996 18645 65036
rect 18603 64987 18645 64996
rect 18808 65036 19176 65045
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 18808 64987 19176 64996
rect 18604 64616 18644 64987
rect 19132 64625 19172 64634
rect 19276 64616 19316 69280
rect 19371 69152 19413 69161
rect 19371 69112 19372 69152
rect 19412 69112 19413 69152
rect 19371 69103 19413 69112
rect 19372 69018 19412 69103
rect 19467 69068 19509 69077
rect 19467 69028 19468 69068
rect 19508 69028 19509 69068
rect 19467 69019 19509 69028
rect 19371 68648 19413 68657
rect 19371 68608 19372 68648
rect 19412 68608 19413 68648
rect 19371 68599 19413 68608
rect 19372 67556 19412 68599
rect 19468 67654 19508 69019
rect 19660 68657 19700 70699
rect 19756 70664 19796 70876
rect 19756 70615 19796 70624
rect 19852 69992 19892 71464
rect 19947 70496 19989 70505
rect 19947 70456 19948 70496
rect 19988 70456 19989 70496
rect 19947 70447 19989 70456
rect 19948 70362 19988 70447
rect 20048 70328 20416 70337
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20048 70279 20416 70288
rect 20524 70253 20564 71968
rect 20523 70244 20565 70253
rect 20523 70204 20524 70244
rect 20564 70204 20565 70244
rect 20523 70195 20565 70204
rect 19947 70076 19989 70085
rect 19947 70036 19948 70076
rect 19988 70036 19989 70076
rect 19947 70027 19989 70036
rect 19804 69982 19892 69992
rect 19844 69952 19892 69982
rect 19948 69942 19988 70027
rect 19804 69933 19844 69942
rect 19851 69824 19893 69833
rect 19851 69784 19852 69824
rect 19892 69784 19893 69824
rect 19851 69775 19893 69784
rect 19852 69166 19892 69775
rect 19852 69117 19892 69126
rect 20523 69152 20565 69161
rect 20523 69112 20524 69152
rect 20564 69112 20565 69152
rect 20523 69103 20565 69112
rect 20044 68993 20084 69078
rect 20043 68984 20085 68993
rect 20043 68944 20044 68984
rect 20084 68944 20085 68984
rect 20043 68935 20085 68944
rect 20048 68816 20416 68825
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20048 68767 20416 68776
rect 19659 68648 19701 68657
rect 19659 68608 19660 68648
rect 19700 68608 19701 68648
rect 19659 68599 19701 68608
rect 19468 67605 19508 67614
rect 19660 68480 19700 68489
rect 19660 67556 19700 68440
rect 19852 68228 19892 68237
rect 19372 67516 19508 67556
rect 19468 66963 19508 67516
rect 19468 66914 19508 66923
rect 19564 67516 19700 67556
rect 19756 68188 19852 68228
rect 19467 66128 19509 66137
rect 19564 66128 19604 67516
rect 19660 67430 19700 67439
rect 19660 67229 19700 67390
rect 19659 67220 19701 67229
rect 19659 67180 19660 67220
rect 19700 67180 19701 67220
rect 19659 67171 19701 67180
rect 19659 67052 19701 67061
rect 19659 67012 19660 67052
rect 19700 67012 19701 67052
rect 19659 67003 19701 67012
rect 19660 66918 19700 67003
rect 19756 66221 19796 68188
rect 19852 68179 19892 68188
rect 20048 67304 20416 67313
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20048 67255 20416 67264
rect 19851 67220 19893 67229
rect 19851 67180 19852 67220
rect 19892 67180 19893 67220
rect 19851 67171 19893 67180
rect 19755 66212 19797 66221
rect 19755 66172 19756 66212
rect 19796 66172 19797 66212
rect 19755 66163 19797 66172
rect 19467 66088 19468 66128
rect 19508 66088 19564 66128
rect 19467 66079 19509 66088
rect 19564 66079 19604 66088
rect 19756 65960 19796 65969
rect 19564 65920 19756 65960
rect 19371 65540 19413 65549
rect 19371 65500 19372 65540
rect 19412 65500 19413 65540
rect 19371 65491 19413 65500
rect 19172 64585 19316 64616
rect 19132 64576 19316 64585
rect 18604 64567 18644 64576
rect 19275 64448 19317 64457
rect 19275 64408 19276 64448
rect 19316 64408 19317 64448
rect 19275 64399 19317 64408
rect 19276 64314 19316 64399
rect 19372 64112 19412 65491
rect 19276 64072 19412 64112
rect 18603 63608 18645 63617
rect 18603 63568 18604 63608
rect 18644 63568 18645 63608
rect 18603 63559 18645 63568
rect 18508 62432 18548 63148
rect 18508 62383 18548 62392
rect 18507 60836 18549 60845
rect 18507 60796 18508 60836
rect 18548 60796 18549 60836
rect 18507 60787 18549 60796
rect 18411 60248 18453 60257
rect 18411 60208 18412 60248
rect 18452 60208 18453 60248
rect 18411 60199 18453 60208
rect 18219 59408 18261 59417
rect 18219 59368 18220 59408
rect 18260 59368 18261 59408
rect 18219 59359 18261 59368
rect 18316 59408 18356 60124
rect 18316 59359 18356 59368
rect 18412 60164 18452 60199
rect 18412 59408 18452 60124
rect 18412 59359 18452 59368
rect 17643 58568 17685 58577
rect 17643 58528 17644 58568
rect 17684 58528 17685 58568
rect 17643 58519 17685 58528
rect 18028 58568 18068 58577
rect 17452 58108 17588 58148
rect 17836 58400 17876 58409
rect 17355 58064 17397 58073
rect 17355 58024 17356 58064
rect 17396 58024 17397 58064
rect 17355 58015 17397 58024
rect 16972 57896 17012 57905
rect 16972 57737 17012 57856
rect 17067 57896 17109 57905
rect 17067 57856 17068 57896
rect 17108 57856 17109 57896
rect 17067 57847 17109 57856
rect 16971 57728 17013 57737
rect 16971 57688 16972 57728
rect 17012 57688 17013 57728
rect 16971 57679 17013 57688
rect 17164 57644 17204 57653
rect 17068 57604 17164 57644
rect 16779 57224 16821 57233
rect 16779 57184 16780 57224
rect 16820 57184 16821 57224
rect 16779 57175 16821 57184
rect 17068 57224 17108 57604
rect 17164 57595 17204 57604
rect 17355 57644 17397 57653
rect 17355 57604 17356 57644
rect 17396 57604 17397 57644
rect 17355 57595 17397 57604
rect 17356 57510 17396 57595
rect 17452 57224 17492 58108
rect 17547 57980 17589 57989
rect 17547 57940 17548 57980
rect 17588 57940 17589 57980
rect 17547 57931 17589 57940
rect 17548 57896 17588 57931
rect 17548 57845 17588 57856
rect 17836 57821 17876 58360
rect 18028 58148 18068 58528
rect 18123 58568 18165 58577
rect 18123 58528 18124 58568
rect 18164 58528 18165 58568
rect 18123 58519 18165 58528
rect 18028 58108 18164 58148
rect 17835 57812 17877 57821
rect 17835 57772 17836 57812
rect 17876 57772 17877 57812
rect 17835 57763 17877 57772
rect 17835 57644 17877 57653
rect 17835 57604 17836 57644
rect 17876 57604 17877 57644
rect 17835 57595 17877 57604
rect 17068 57184 17396 57224
rect 17452 57184 17780 57224
rect 16875 57140 16917 57149
rect 16875 57100 16876 57140
rect 16916 57100 16917 57140
rect 16875 57091 16917 57100
rect 16204 56512 16340 56552
rect 16396 57056 16436 57065
rect 16107 55124 16149 55133
rect 16107 55084 16108 55124
rect 16148 55084 16149 55124
rect 16107 55075 16149 55084
rect 15915 55040 15957 55049
rect 15915 55000 15916 55040
rect 15956 55000 15957 55040
rect 15915 54991 15957 55000
rect 16107 54956 16149 54965
rect 16107 54916 16108 54956
rect 16148 54916 16149 54956
rect 16107 54907 16149 54916
rect 15916 54858 15956 54867
rect 16108 54822 16148 54907
rect 15916 54293 15956 54818
rect 16011 54452 16053 54461
rect 16011 54412 16012 54452
rect 16052 54412 16053 54452
rect 16011 54403 16053 54412
rect 15915 54284 15957 54293
rect 15915 54244 15916 54284
rect 15956 54244 15957 54284
rect 15915 54235 15957 54244
rect 15916 53360 15956 53369
rect 15916 52529 15956 53320
rect 15915 52520 15957 52529
rect 15915 52480 15916 52520
rect 15956 52480 15957 52520
rect 15915 52471 15957 52480
rect 16012 52109 16052 54403
rect 16107 54032 16149 54041
rect 16107 53992 16108 54032
rect 16148 53992 16149 54032
rect 16107 53983 16149 53992
rect 16108 53898 16148 53983
rect 16204 53621 16244 56512
rect 16300 56384 16340 56393
rect 16300 54461 16340 56344
rect 16396 55460 16436 57016
rect 16491 57056 16533 57065
rect 16491 57016 16492 57056
rect 16532 57016 16533 57056
rect 16491 57007 16533 57016
rect 16684 57056 16724 57065
rect 16876 57056 16916 57091
rect 16972 57065 17012 57150
rect 16724 57016 16820 57056
rect 16684 57007 16724 57016
rect 16492 56922 16532 57007
rect 16588 56888 16628 56897
rect 16780 56888 16820 57016
rect 16876 57005 16916 57016
rect 16971 57056 17013 57065
rect 16971 57016 16972 57056
rect 17012 57016 17013 57056
rect 16971 57007 17013 57016
rect 17068 57056 17108 57184
rect 17068 57007 17108 57016
rect 17259 57056 17301 57065
rect 17259 57016 17260 57056
rect 17300 57016 17301 57056
rect 17259 57007 17301 57016
rect 17356 57056 17396 57184
rect 17356 57007 17396 57016
rect 17548 57056 17588 57065
rect 17164 56888 17204 56897
rect 16780 56848 17164 56888
rect 16588 56393 16628 56848
rect 17164 56839 17204 56848
rect 16779 56720 16821 56729
rect 16779 56680 16780 56720
rect 16820 56680 16821 56720
rect 16779 56671 16821 56680
rect 16587 56384 16629 56393
rect 16587 56344 16588 56384
rect 16628 56344 16629 56384
rect 16587 56335 16629 56344
rect 16780 56384 16820 56671
rect 16971 56636 17013 56645
rect 16971 56596 16972 56636
rect 17012 56596 17013 56636
rect 16971 56587 17013 56596
rect 16972 56552 17012 56587
rect 17260 56552 17300 57007
rect 17548 56972 17588 57016
rect 17548 56932 17684 56972
rect 17452 56888 17492 56897
rect 17492 56848 17588 56888
rect 17452 56839 17492 56848
rect 17452 56552 17492 56561
rect 17260 56512 17452 56552
rect 16972 56501 17012 56512
rect 17452 56503 17492 56512
rect 17164 56384 17204 56393
rect 16780 56379 17164 56384
rect 16820 56344 17164 56379
rect 17548 56384 17588 56848
rect 17644 56645 17684 56932
rect 17643 56636 17685 56645
rect 17643 56596 17644 56636
rect 17684 56596 17685 56636
rect 17643 56587 17685 56596
rect 17644 56384 17684 56393
rect 16780 55460 16820 56339
rect 17164 56335 17204 56344
rect 17260 56342 17300 56351
rect 17163 55964 17205 55973
rect 17260 55964 17300 56302
rect 17356 56342 17396 56351
rect 17548 56344 17644 56384
rect 17644 56335 17684 56344
rect 17740 56309 17780 57184
rect 17836 57056 17876 57595
rect 17931 57560 17973 57569
rect 17931 57520 17932 57560
rect 17972 57520 17973 57560
rect 17931 57511 17973 57520
rect 17836 57007 17876 57016
rect 17932 57056 17972 57511
rect 17835 56384 17877 56393
rect 17835 56344 17836 56384
rect 17876 56344 17877 56384
rect 17835 56335 17877 56344
rect 17356 56225 17396 56302
rect 17739 56300 17781 56309
rect 17739 56260 17740 56300
rect 17780 56260 17781 56300
rect 17739 56251 17781 56260
rect 17836 56250 17876 56335
rect 17355 56216 17397 56225
rect 17355 56176 17356 56216
rect 17396 56176 17397 56216
rect 17355 56167 17397 56176
rect 17643 56132 17685 56141
rect 17643 56092 17644 56132
rect 17684 56092 17685 56132
rect 17643 56083 17685 56092
rect 17644 55998 17684 56083
rect 17163 55924 17164 55964
rect 17204 55924 17300 55964
rect 17163 55915 17205 55924
rect 16971 55628 17013 55637
rect 16971 55588 16972 55628
rect 17012 55588 17013 55628
rect 16971 55579 17013 55588
rect 16396 55420 16532 55460
rect 16492 55049 16532 55420
rect 16588 55420 16820 55460
rect 16491 55040 16533 55049
rect 16491 55000 16492 55040
rect 16532 55000 16533 55040
rect 16491 54991 16533 55000
rect 16396 54872 16436 54881
rect 16588 54872 16628 55420
rect 16436 54832 16628 54872
rect 16684 55000 16916 55040
rect 16684 54872 16724 55000
rect 16396 54823 16436 54832
rect 16684 54823 16724 54832
rect 16780 54872 16820 54881
rect 16299 54452 16341 54461
rect 16299 54412 16300 54452
rect 16340 54412 16341 54452
rect 16299 54403 16341 54412
rect 16491 54452 16533 54461
rect 16491 54412 16492 54452
rect 16532 54412 16533 54452
rect 16491 54403 16533 54412
rect 16299 54284 16341 54293
rect 16299 54244 16300 54284
rect 16340 54244 16341 54284
rect 16299 54235 16341 54244
rect 16300 54150 16340 54235
rect 16203 53612 16245 53621
rect 16203 53572 16204 53612
rect 16244 53572 16245 53612
rect 16203 53563 16245 53572
rect 16107 53276 16149 53285
rect 16107 53236 16108 53276
rect 16148 53236 16149 53276
rect 16107 53227 16149 53236
rect 16108 52277 16148 53227
rect 16107 52268 16149 52277
rect 16107 52228 16108 52268
rect 16148 52228 16149 52268
rect 16107 52219 16149 52228
rect 16011 52100 16053 52109
rect 16011 52060 16012 52100
rect 16052 52060 16053 52100
rect 16011 52051 16053 52060
rect 15820 51976 15956 52016
rect 15723 51932 15765 51941
rect 15723 51892 15724 51932
rect 15764 51892 15765 51932
rect 15723 51883 15765 51892
rect 15820 51848 15860 51859
rect 15820 51773 15860 51808
rect 15819 51764 15861 51773
rect 15819 51724 15820 51764
rect 15860 51724 15861 51764
rect 15819 51715 15861 51724
rect 15628 50959 15668 50968
rect 15723 51008 15765 51017
rect 15723 50968 15724 51008
rect 15764 50968 15765 51008
rect 15723 50959 15765 50968
rect 15724 50874 15764 50959
rect 15723 50756 15765 50765
rect 15723 50716 15724 50756
rect 15764 50716 15765 50756
rect 15723 50707 15765 50716
rect 15051 50588 15093 50597
rect 15051 50548 15052 50588
rect 15092 50548 15093 50588
rect 15051 50539 15093 50548
rect 14860 49540 14996 49580
rect 14524 49505 14564 49514
rect 14564 49465 14804 49496
rect 14524 49456 14804 49465
rect 14764 49412 14804 49456
rect 14860 49412 14900 49421
rect 14380 49372 14516 49412
rect 14764 49372 14860 49412
rect 14379 48824 14421 48833
rect 14379 48784 14380 48824
rect 14420 48784 14421 48824
rect 14476 48824 14516 49372
rect 14860 49363 14900 49372
rect 14668 49328 14708 49337
rect 14668 49001 14708 49288
rect 14763 49244 14805 49253
rect 14763 49204 14764 49244
rect 14804 49204 14805 49244
rect 14763 49195 14805 49204
rect 14667 48992 14709 49001
rect 14667 48952 14668 48992
rect 14708 48952 14709 48992
rect 14667 48943 14709 48952
rect 14476 48784 14708 48824
rect 14379 48775 14421 48784
rect 14380 48656 14420 48775
rect 14380 48616 14516 48656
rect 14283 48572 14325 48581
rect 14283 48532 14284 48572
rect 14324 48532 14325 48572
rect 14283 48523 14325 48532
rect 14284 47998 14324 48523
rect 14379 48068 14421 48077
rect 14379 48028 14380 48068
rect 14420 48028 14421 48068
rect 14379 48019 14421 48028
rect 14284 47949 14324 47958
rect 14380 47900 14420 48019
rect 14476 47984 14516 48616
rect 14571 48572 14613 48581
rect 14571 48532 14572 48572
rect 14612 48532 14613 48572
rect 14571 48523 14613 48532
rect 14572 48438 14612 48523
rect 14668 47984 14708 48784
rect 14476 47944 14612 47984
rect 14380 47860 14516 47900
rect 14476 47816 14516 47860
rect 14476 47767 14516 47776
rect 14187 47312 14229 47321
rect 14187 47272 14188 47312
rect 14228 47272 14229 47312
rect 14187 47263 14229 47272
rect 14475 47312 14517 47321
rect 14475 47272 14476 47312
rect 14516 47272 14517 47312
rect 14475 47263 14517 47272
rect 14188 47178 14228 47263
rect 14380 47060 14420 47069
rect 14284 47020 14380 47060
rect 14284 46640 14324 47020
rect 14380 47011 14420 47020
rect 14188 46600 14324 46640
rect 14188 46486 14228 46600
rect 14188 46437 14228 46446
rect 14380 46388 14420 46397
rect 14476 46388 14516 47263
rect 14572 46640 14612 47944
rect 14668 47935 14708 47944
rect 14572 46600 14708 46640
rect 14420 46348 14516 46388
rect 14380 46339 14420 46348
rect 14091 42776 14133 42785
rect 14091 42736 14092 42776
rect 14132 42736 14133 42776
rect 14091 42727 14133 42736
rect 14379 42776 14421 42785
rect 14379 42736 14380 42776
rect 14420 42736 14421 42776
rect 14379 42727 14421 42736
rect 14380 42642 14420 42727
rect 14572 42524 14612 42533
rect 14572 41950 14612 42484
rect 14092 41936 14132 41945
rect 14132 41896 14516 41936
rect 14572 41901 14612 41910
rect 14092 41887 14132 41896
rect 14283 41768 14325 41777
rect 13900 41728 14132 41768
rect 13995 41600 14037 41609
rect 13995 41560 13996 41600
rect 14036 41560 14037 41600
rect 13995 41551 14037 41560
rect 13707 41432 13749 41441
rect 13707 41392 13708 41432
rect 13748 41392 13749 41432
rect 13707 41383 13749 41392
rect 13804 41264 13844 41273
rect 13652 41224 13748 41264
rect 13612 41215 13652 41224
rect 13419 41012 13461 41021
rect 13419 40972 13420 41012
rect 13460 40972 13461 41012
rect 13419 40963 13461 40972
rect 13612 41012 13652 41021
rect 13228 40888 13364 40928
rect 13131 39920 13173 39929
rect 13131 39880 13132 39920
rect 13172 39880 13173 39920
rect 13131 39871 13173 39880
rect 12940 39677 12980 39712
rect 13131 39752 13173 39761
rect 13131 39712 13132 39752
rect 13172 39712 13173 39752
rect 13131 39703 13173 39712
rect 12939 39668 12981 39677
rect 12939 39628 12940 39668
rect 12980 39628 12981 39668
rect 12939 39619 12981 39628
rect 12652 38863 12692 38872
rect 12748 39040 12884 39080
rect 12651 38324 12693 38333
rect 12651 38284 12652 38324
rect 12692 38284 12693 38324
rect 12651 38275 12693 38284
rect 12652 38240 12692 38275
rect 12652 38189 12692 38200
rect 12748 37820 12788 39040
rect 12843 38912 12885 38921
rect 12843 38872 12844 38912
rect 12884 38872 12885 38912
rect 12843 38863 12885 38872
rect 12940 38912 12980 39619
rect 13035 39500 13077 39509
rect 13035 39460 13036 39500
rect 13076 39460 13077 39500
rect 13035 39451 13077 39460
rect 13036 39366 13076 39451
rect 13132 39248 13172 39703
rect 12940 38863 12980 38872
rect 13036 39208 13172 39248
rect 13036 38912 13076 39208
rect 13228 39005 13268 40888
rect 13420 40878 13460 40963
rect 13612 40844 13652 40972
rect 13708 40937 13748 41224
rect 13707 40928 13749 40937
rect 13707 40888 13708 40928
rect 13748 40888 13749 40928
rect 13707 40879 13749 40888
rect 13611 40804 13652 40844
rect 13324 40685 13364 40770
rect 13611 40760 13651 40804
rect 13611 40720 13652 40760
rect 13323 40676 13365 40685
rect 13323 40636 13324 40676
rect 13364 40636 13365 40676
rect 13323 40627 13365 40636
rect 13515 40592 13557 40601
rect 13515 40552 13516 40592
rect 13556 40552 13557 40592
rect 13515 40543 13557 40552
rect 13324 40424 13364 40433
rect 13324 40340 13364 40384
rect 13516 40424 13556 40543
rect 13516 40375 13556 40384
rect 13612 40424 13652 40720
rect 13612 40375 13652 40384
rect 13324 40300 13460 40340
rect 13323 39752 13365 39761
rect 13323 39712 13324 39752
rect 13364 39712 13365 39752
rect 13323 39703 13365 39712
rect 13227 38996 13269 39005
rect 13227 38956 13228 38996
rect 13268 38956 13269 38996
rect 13227 38947 13269 38956
rect 13036 38863 13076 38872
rect 13132 38912 13172 38921
rect 13324 38912 13364 39703
rect 13420 39593 13460 40300
rect 13707 40256 13749 40265
rect 13707 40216 13708 40256
rect 13748 40216 13749 40256
rect 13707 40207 13749 40216
rect 13611 40172 13653 40181
rect 13611 40132 13612 40172
rect 13652 40132 13653 40172
rect 13611 40123 13653 40132
rect 13515 40004 13557 40013
rect 13515 39964 13516 40004
rect 13556 39964 13557 40004
rect 13515 39955 13557 39964
rect 13419 39584 13461 39593
rect 13419 39544 13420 39584
rect 13460 39544 13461 39584
rect 13419 39535 13461 39544
rect 13420 38912 13460 38921
rect 13324 38872 13420 38912
rect 12844 38778 12884 38863
rect 13132 38753 13172 38872
rect 13420 38863 13460 38872
rect 13227 38828 13269 38837
rect 13227 38788 13228 38828
rect 13268 38788 13269 38828
rect 13227 38779 13269 38788
rect 13131 38744 13173 38753
rect 13131 38704 13132 38744
rect 13172 38704 13173 38744
rect 13131 38695 13173 38704
rect 13132 38585 13172 38695
rect 13131 38576 13173 38585
rect 13131 38536 13132 38576
rect 13172 38536 13173 38576
rect 13131 38527 13173 38536
rect 13131 38156 13173 38165
rect 13131 38116 13132 38156
rect 13172 38116 13173 38156
rect 13131 38107 13173 38116
rect 12748 37780 12980 37820
rect 12748 37400 12788 37409
rect 12748 36896 12788 37360
rect 12844 37400 12884 37411
rect 12844 37325 12884 37360
rect 12843 37316 12885 37325
rect 12843 37276 12844 37316
rect 12884 37276 12885 37316
rect 12843 37267 12885 37276
rect 12748 36856 12884 36896
rect 12747 36728 12789 36737
rect 12747 36688 12748 36728
rect 12788 36688 12789 36728
rect 12747 36679 12789 36688
rect 12844 36728 12884 36856
rect 12748 36594 12788 36679
rect 12844 36653 12884 36688
rect 12843 36644 12885 36653
rect 12843 36604 12844 36644
rect 12884 36604 12885 36644
rect 12843 36595 12885 36604
rect 12652 35888 12692 35897
rect 12267 34880 12309 34889
rect 12267 34840 12268 34880
rect 12308 34840 12309 34880
rect 12267 34831 12309 34840
rect 12555 34880 12597 34889
rect 12555 34840 12556 34880
rect 12596 34840 12597 34880
rect 12555 34831 12597 34840
rect 12076 33328 12212 33368
rect 11979 32192 12021 32201
rect 11979 32152 11980 32192
rect 12020 32152 12021 32192
rect 11979 32143 12021 32152
rect 11980 32058 12020 32143
rect 11979 31352 12021 31361
rect 11979 31312 11980 31352
rect 12020 31312 12021 31352
rect 11979 31303 12021 31312
rect 11980 30605 12020 31303
rect 11979 30596 12021 30605
rect 11979 30556 11980 30596
rect 12020 30556 12021 30596
rect 11979 30547 12021 30556
rect 11884 28960 12020 29000
rect 11980 27824 12020 28960
rect 12076 27917 12116 33328
rect 12268 33209 12308 34831
rect 12555 34712 12597 34721
rect 12555 34672 12556 34712
rect 12596 34672 12597 34712
rect 12555 34663 12597 34672
rect 12363 34376 12405 34385
rect 12363 34336 12364 34376
rect 12404 34336 12405 34376
rect 12363 34327 12405 34336
rect 12364 34242 12404 34327
rect 12460 33690 12500 33699
rect 12267 33200 12309 33209
rect 12267 33160 12268 33200
rect 12308 33160 12309 33200
rect 12267 33151 12309 33160
rect 12460 33116 12500 33650
rect 12460 33067 12500 33076
rect 12267 32948 12309 32957
rect 12267 32908 12268 32948
rect 12308 32908 12309 32948
rect 12267 32899 12309 32908
rect 12268 32864 12308 32899
rect 12268 32813 12308 32824
rect 12171 32276 12213 32285
rect 12171 32236 12172 32276
rect 12212 32236 12213 32276
rect 12171 32227 12213 32236
rect 12459 32276 12501 32285
rect 12459 32236 12460 32276
rect 12500 32236 12501 32276
rect 12459 32227 12501 32236
rect 12172 32142 12212 32227
rect 12460 32192 12500 32227
rect 12460 32141 12500 32152
rect 12556 32192 12596 34663
rect 12652 34049 12692 35848
rect 12843 35720 12885 35729
rect 12843 35680 12844 35720
rect 12884 35680 12885 35720
rect 12843 35671 12885 35680
rect 12844 35586 12884 35671
rect 12747 35132 12789 35141
rect 12747 35092 12748 35132
rect 12788 35092 12789 35132
rect 12747 35083 12789 35092
rect 12844 35132 12884 35143
rect 12748 34721 12788 35083
rect 12844 35057 12884 35092
rect 12843 35048 12885 35057
rect 12843 35008 12844 35048
rect 12884 35008 12885 35048
rect 12843 34999 12885 35008
rect 12747 34712 12789 34721
rect 12747 34672 12748 34712
rect 12788 34672 12789 34712
rect 12747 34663 12789 34672
rect 12651 34040 12693 34049
rect 12651 34000 12652 34040
rect 12692 34000 12693 34040
rect 12651 33991 12693 34000
rect 12651 33872 12693 33881
rect 12940 33872 12980 37780
rect 13035 36560 13077 36569
rect 13035 36520 13036 36560
rect 13076 36520 13077 36560
rect 13035 36511 13077 36520
rect 12651 33832 12652 33872
rect 12692 33832 12693 33872
rect 12651 33823 12693 33832
rect 12748 33832 12980 33872
rect 12652 33738 12692 33823
rect 12556 32117 12596 32152
rect 12555 32108 12597 32117
rect 12555 32068 12556 32108
rect 12596 32068 12597 32108
rect 12555 32059 12597 32068
rect 12651 31352 12693 31361
rect 12651 31312 12652 31352
rect 12692 31312 12693 31352
rect 12651 31303 12693 31312
rect 12652 31218 12692 31303
rect 12748 30680 12788 33832
rect 12940 33704 12980 33713
rect 12651 30596 12693 30605
rect 12651 30556 12652 30596
rect 12692 30556 12693 30596
rect 12651 30547 12693 30556
rect 12267 30428 12309 30437
rect 12267 30388 12268 30428
rect 12308 30388 12309 30428
rect 12267 30379 12309 30388
rect 12268 27917 12308 30379
rect 12652 30269 12692 30547
rect 12651 30260 12693 30269
rect 12651 30220 12652 30260
rect 12692 30220 12693 30260
rect 12651 30211 12693 30220
rect 12748 29882 12788 30640
rect 12844 33664 12940 33704
rect 12844 30260 12884 33664
rect 12940 33655 12980 33664
rect 12940 32108 12980 32119
rect 12940 32033 12980 32068
rect 13036 32108 13076 36511
rect 13132 35477 13172 38107
rect 13228 37493 13268 38779
rect 13227 37484 13269 37493
rect 13227 37444 13228 37484
rect 13268 37444 13269 37484
rect 13227 37435 13269 37444
rect 13323 37400 13365 37409
rect 13323 37360 13324 37400
rect 13364 37360 13460 37400
rect 13323 37351 13365 37360
rect 13227 37316 13269 37325
rect 13227 37276 13228 37316
rect 13268 37276 13269 37316
rect 13227 37267 13269 37276
rect 13228 36644 13268 37267
rect 13324 37266 13364 37351
rect 13324 36653 13364 36738
rect 13131 35468 13173 35477
rect 13131 35428 13132 35468
rect 13172 35428 13173 35468
rect 13131 35419 13173 35428
rect 13131 35048 13173 35057
rect 13228 35048 13268 36604
rect 13323 36644 13365 36653
rect 13323 36604 13324 36644
rect 13364 36604 13365 36644
rect 13323 36595 13365 36604
rect 13420 36476 13460 37360
rect 13324 36436 13460 36476
rect 13324 35216 13364 36436
rect 13420 35888 13460 35897
rect 13420 35477 13460 35848
rect 13419 35468 13461 35477
rect 13419 35428 13420 35468
rect 13460 35428 13461 35468
rect 13419 35419 13461 35428
rect 13324 35167 13364 35176
rect 13131 35008 13132 35048
rect 13172 35008 13268 35048
rect 13131 34999 13173 35008
rect 12939 32024 12981 32033
rect 12939 31984 12940 32024
rect 12980 31984 12981 32024
rect 12939 31975 12981 31984
rect 13036 31025 13076 32068
rect 13132 32033 13172 34999
rect 13420 34964 13460 35419
rect 13228 34924 13460 34964
rect 13131 32024 13173 32033
rect 13131 31984 13132 32024
rect 13172 31984 13173 32024
rect 13131 31975 13173 31984
rect 13228 31361 13268 34924
rect 13516 33881 13556 39955
rect 13612 39779 13652 40123
rect 13708 39836 13748 40207
rect 13708 39787 13748 39796
rect 13612 39730 13652 39739
rect 13804 39509 13844 41224
rect 13900 41264 13940 41273
rect 13803 39500 13845 39509
rect 13803 39460 13804 39500
rect 13844 39460 13845 39500
rect 13803 39451 13845 39460
rect 13707 39332 13749 39341
rect 13707 39292 13708 39332
rect 13748 39292 13749 39332
rect 13707 39283 13749 39292
rect 13708 38912 13748 39283
rect 13900 39164 13940 41224
rect 13996 40424 14036 41551
rect 13996 40088 14036 40384
rect 14092 40349 14132 41728
rect 14283 41728 14284 41768
rect 14324 41728 14325 41768
rect 14283 41719 14325 41728
rect 14187 41516 14229 41525
rect 14187 41476 14188 41516
rect 14228 41476 14229 41516
rect 14187 41467 14229 41476
rect 14188 41264 14228 41467
rect 14091 40340 14133 40349
rect 14091 40300 14092 40340
rect 14132 40300 14133 40340
rect 14091 40291 14133 40300
rect 13996 40048 14132 40088
rect 13996 39500 14036 39509
rect 13996 39341 14036 39460
rect 14092 39416 14132 40048
rect 14188 39929 14228 41224
rect 14187 39920 14229 39929
rect 14187 39880 14188 39920
rect 14228 39880 14229 39920
rect 14187 39871 14229 39880
rect 14284 39845 14324 41719
rect 14379 41348 14421 41357
rect 14379 41308 14380 41348
rect 14420 41308 14421 41348
rect 14379 41299 14421 41308
rect 14380 40853 14420 41299
rect 14476 41180 14516 41896
rect 14668 41357 14708 46600
rect 14764 41852 14804 49195
rect 14956 47489 14996 49540
rect 15052 49496 15092 50539
rect 15724 50336 15764 50707
rect 15916 50345 15956 51976
rect 16492 51941 16532 54403
rect 16587 53444 16629 53453
rect 16587 53404 16588 53444
rect 16628 53404 16629 53444
rect 16587 53395 16629 53404
rect 16012 51932 16052 51941
rect 16491 51932 16533 51941
rect 16052 51892 16148 51932
rect 16012 51883 16052 51892
rect 16108 51773 16148 51892
rect 16491 51892 16492 51932
rect 16532 51892 16533 51932
rect 16588 51932 16628 53395
rect 16683 52100 16725 52109
rect 16683 52060 16684 52100
rect 16724 52060 16725 52100
rect 16683 52051 16725 52060
rect 16588 51892 16629 51932
rect 16491 51883 16533 51892
rect 16589 51859 16629 51892
rect 16204 51848 16244 51857
rect 16107 51764 16149 51773
rect 16107 51724 16108 51764
rect 16148 51724 16149 51764
rect 16107 51715 16149 51724
rect 16107 51596 16149 51605
rect 16107 51556 16108 51596
rect 16148 51556 16149 51596
rect 16107 51547 16149 51556
rect 15627 49748 15669 49757
rect 15627 49708 15628 49748
rect 15668 49708 15669 49748
rect 15627 49699 15669 49708
rect 15052 48833 15092 49456
rect 15051 48824 15093 48833
rect 15051 48784 15052 48824
rect 15092 48784 15093 48824
rect 15051 48775 15093 48784
rect 15531 48824 15573 48833
rect 15531 48784 15532 48824
rect 15572 48784 15573 48824
rect 15531 48775 15573 48784
rect 15628 48824 15668 49699
rect 15532 48690 15572 48775
rect 15628 48488 15668 48784
rect 15724 48749 15764 50296
rect 15915 50336 15957 50345
rect 15915 50296 15916 50336
rect 15956 50296 15957 50336
rect 15915 50287 15957 50296
rect 16108 50336 16148 51547
rect 16204 51269 16244 51808
rect 16396 51848 16436 51857
rect 16589 51810 16629 51819
rect 16299 51764 16341 51773
rect 16299 51724 16300 51764
rect 16340 51724 16341 51764
rect 16299 51715 16341 51724
rect 16300 51630 16340 51715
rect 16396 51596 16436 51808
rect 16588 51596 16628 51605
rect 16396 51556 16588 51596
rect 16588 51547 16628 51556
rect 16203 51260 16245 51269
rect 16203 51220 16204 51260
rect 16244 51220 16245 51260
rect 16203 51211 16245 51220
rect 16300 51101 16340 51132
rect 16299 51092 16341 51101
rect 16299 51052 16300 51092
rect 16340 51052 16341 51092
rect 16299 51043 16341 51052
rect 16300 51008 16340 51043
rect 16300 50933 16340 50968
rect 16299 50924 16341 50933
rect 16299 50884 16300 50924
rect 16340 50884 16341 50924
rect 16299 50875 16341 50884
rect 16587 50420 16629 50429
rect 16587 50380 16588 50420
rect 16628 50380 16629 50420
rect 16587 50371 16629 50380
rect 16108 50177 16148 50296
rect 16203 50336 16245 50345
rect 16203 50296 16204 50336
rect 16244 50296 16245 50336
rect 16203 50287 16245 50296
rect 16107 50168 16149 50177
rect 16107 50128 16108 50168
rect 16148 50128 16149 50168
rect 16107 50119 16149 50128
rect 15916 50084 15956 50093
rect 15916 48833 15956 50044
rect 15915 48824 15957 48833
rect 15915 48784 15916 48824
rect 15956 48784 15957 48824
rect 15915 48775 15957 48784
rect 16108 48824 16148 48833
rect 16204 48824 16244 50287
rect 16395 50168 16437 50177
rect 16395 50128 16396 50168
rect 16436 50128 16437 50168
rect 16395 50119 16437 50128
rect 16299 49580 16341 49589
rect 16299 49540 16300 49580
rect 16340 49540 16341 49580
rect 16299 49531 16341 49540
rect 16300 49496 16340 49531
rect 16300 49445 16340 49456
rect 16396 49169 16436 50119
rect 16588 49505 16628 50371
rect 16587 49496 16629 49505
rect 16587 49456 16588 49496
rect 16628 49456 16629 49496
rect 16587 49447 16629 49456
rect 16395 49160 16437 49169
rect 16395 49120 16396 49160
rect 16436 49120 16437 49160
rect 16395 49111 16437 49120
rect 16491 49076 16533 49085
rect 16491 49036 16492 49076
rect 16532 49036 16533 49076
rect 16491 49027 16533 49036
rect 16148 48784 16244 48824
rect 16108 48775 16148 48784
rect 15723 48740 15765 48749
rect 15723 48700 15724 48740
rect 15764 48700 15765 48740
rect 15723 48691 15765 48700
rect 16012 48740 16052 48751
rect 16012 48665 16052 48700
rect 16011 48656 16053 48665
rect 16011 48616 16012 48656
rect 16052 48616 16053 48656
rect 16011 48607 16053 48616
rect 15532 48448 15668 48488
rect 15435 47816 15477 47825
rect 15435 47776 15436 47816
rect 15476 47776 15477 47816
rect 15435 47767 15477 47776
rect 14955 47480 14997 47489
rect 14955 47440 14956 47480
rect 14996 47440 14997 47480
rect 14955 47431 14997 47440
rect 15436 47312 15476 47767
rect 15436 47263 15476 47272
rect 15532 47312 15572 48448
rect 15916 47993 15956 48078
rect 15915 47984 15957 47993
rect 15915 47944 15916 47984
rect 15956 47944 15957 47984
rect 15915 47935 15957 47944
rect 16012 47732 16052 48607
rect 16108 47825 16148 47910
rect 16107 47816 16149 47825
rect 16107 47776 16108 47816
rect 16148 47776 16149 47816
rect 16107 47767 16149 47776
rect 15916 47692 16052 47732
rect 15916 47312 15956 47692
rect 16204 47648 16244 48784
rect 16492 48572 16532 49027
rect 16587 48824 16629 48833
rect 16587 48784 16588 48824
rect 16628 48784 16629 48824
rect 16587 48775 16629 48784
rect 16588 48690 16628 48775
rect 16492 48532 16628 48572
rect 16491 48404 16533 48413
rect 16491 48364 16492 48404
rect 16532 48364 16533 48404
rect 16491 48355 16533 48364
rect 16492 47993 16532 48355
rect 16588 48077 16628 48532
rect 16587 48068 16629 48077
rect 16587 48028 16588 48068
rect 16628 48028 16629 48068
rect 16587 48019 16629 48028
rect 16491 47984 16533 47993
rect 16491 47944 16492 47984
rect 16532 47944 16533 47984
rect 16491 47935 16533 47944
rect 16492 47850 16532 47935
rect 16299 47816 16341 47825
rect 16299 47776 16300 47816
rect 16340 47776 16341 47816
rect 16299 47767 16341 47776
rect 16300 47682 16340 47767
rect 15532 47263 15572 47272
rect 15628 47272 15916 47312
rect 14955 46472 14997 46481
rect 14955 46432 14956 46472
rect 14996 46432 14997 46472
rect 14955 46423 14997 46432
rect 14956 45800 14996 46423
rect 14956 45751 14996 45760
rect 15148 45548 15188 45557
rect 15052 45508 15148 45548
rect 15052 44297 15092 45508
rect 15148 45499 15188 45508
rect 15436 44960 15476 44969
rect 15436 44372 15476 44920
rect 15340 44332 15476 44372
rect 15532 44960 15572 44969
rect 15628 44960 15668 47272
rect 15916 47263 15956 47272
rect 16012 47608 16244 47648
rect 16012 47312 16052 47608
rect 16299 47396 16341 47405
rect 16299 47356 16300 47396
rect 16340 47356 16341 47396
rect 16299 47347 16341 47356
rect 16012 47144 16052 47272
rect 15916 47104 16052 47144
rect 15724 46472 15764 46483
rect 15724 46397 15764 46432
rect 15723 46388 15765 46397
rect 15723 46348 15724 46388
rect 15764 46348 15860 46388
rect 15723 46339 15765 46348
rect 15820 45800 15860 46348
rect 15820 45751 15860 45760
rect 15572 44920 15668 44960
rect 15916 45044 15956 47104
rect 16203 45380 16245 45389
rect 16203 45340 16204 45380
rect 16244 45340 16245 45380
rect 16203 45331 16245 45340
rect 15051 44288 15093 44297
rect 15051 44248 15052 44288
rect 15092 44248 15093 44288
rect 15051 44239 15093 44248
rect 15148 44213 15188 44298
rect 15147 44204 15189 44213
rect 15147 44164 15148 44204
rect 15188 44164 15189 44204
rect 15147 44155 15189 44164
rect 14955 44120 14997 44129
rect 15340 44120 15380 44332
rect 15532 44288 15572 44920
rect 15436 44269 15476 44278
rect 15532 44239 15572 44248
rect 15916 44288 15956 45004
rect 16011 45044 16053 45053
rect 16011 45004 16012 45044
rect 16052 45004 16053 45044
rect 16011 44995 16053 45004
rect 15916 44239 15956 44248
rect 16012 44288 16052 44995
rect 16204 44297 16244 45331
rect 16012 44239 16052 44248
rect 16203 44288 16245 44297
rect 16203 44248 16204 44288
rect 16244 44248 16245 44288
rect 16203 44239 16245 44248
rect 15436 44213 15476 44229
rect 15435 44204 15477 44213
rect 15435 44164 15436 44204
rect 15476 44164 15477 44204
rect 15435 44155 15477 44164
rect 15436 44134 15476 44155
rect 14955 44080 14956 44120
rect 14996 44080 14997 44120
rect 14955 44071 14997 44080
rect 15244 44080 15380 44120
rect 14956 43986 14996 44071
rect 15244 43700 15284 44080
rect 15244 43651 15284 43660
rect 16204 43457 16244 44239
rect 15052 43448 15092 43457
rect 15243 43448 15285 43457
rect 15092 43408 15244 43448
rect 15284 43408 15285 43448
rect 15052 43399 15092 43408
rect 15243 43399 15285 43408
rect 16203 43448 16245 43457
rect 16203 43408 16204 43448
rect 16244 43408 16245 43448
rect 16203 43399 16245 43408
rect 14956 42692 14996 42701
rect 14764 41803 14804 41812
rect 14860 42652 14956 42692
rect 14860 41525 14900 42652
rect 14956 42643 14996 42652
rect 15147 42608 15189 42617
rect 15147 42568 15148 42608
rect 15188 42568 15189 42608
rect 15147 42559 15189 42568
rect 15148 42474 15188 42559
rect 15147 42188 15189 42197
rect 15147 42148 15148 42188
rect 15188 42148 15189 42188
rect 15147 42139 15189 42148
rect 15148 42054 15188 42139
rect 14956 42020 14996 42029
rect 14956 41609 14996 41980
rect 15244 41936 15284 43399
rect 16108 42692 16148 42701
rect 15148 41896 15284 41936
rect 15724 41936 15764 41945
rect 14955 41600 14997 41609
rect 14955 41560 14956 41600
rect 14996 41560 14997 41600
rect 14955 41551 14997 41560
rect 14859 41516 14901 41525
rect 14859 41476 14860 41516
rect 14900 41476 14901 41516
rect 14859 41467 14901 41476
rect 14667 41348 14709 41357
rect 14667 41308 14668 41348
rect 14708 41308 14709 41348
rect 14667 41299 14709 41308
rect 14476 41140 15092 41180
rect 14667 41012 14709 41021
rect 14667 40972 14668 41012
rect 14708 40972 14709 41012
rect 14667 40963 14709 40972
rect 14379 40844 14421 40853
rect 14379 40804 14380 40844
rect 14420 40804 14421 40844
rect 14379 40795 14421 40804
rect 14475 39920 14517 39929
rect 14475 39880 14476 39920
rect 14516 39880 14517 39920
rect 14475 39871 14517 39880
rect 14283 39836 14325 39845
rect 14283 39796 14284 39836
rect 14324 39796 14325 39836
rect 14283 39787 14325 39796
rect 14187 39752 14229 39761
rect 14187 39712 14188 39752
rect 14228 39712 14229 39752
rect 14187 39703 14229 39712
rect 14284 39752 14324 39787
rect 14476 39786 14516 39871
rect 14188 39618 14228 39703
rect 14284 39702 14324 39712
rect 14380 39752 14420 39763
rect 14380 39677 14420 39712
rect 14668 39752 14708 40963
rect 14859 40928 14901 40937
rect 14859 40888 14860 40928
rect 14900 40888 14901 40928
rect 14859 40879 14901 40888
rect 14763 39920 14805 39929
rect 14763 39880 14764 39920
rect 14804 39880 14805 39920
rect 14763 39871 14805 39880
rect 14668 39703 14708 39712
rect 14764 39752 14804 39871
rect 14764 39703 14804 39712
rect 14860 39752 14900 40879
rect 14860 39703 14900 39712
rect 14956 39752 14996 39761
rect 14379 39668 14421 39677
rect 14379 39628 14380 39668
rect 14420 39628 14421 39668
rect 14379 39619 14421 39628
rect 14475 39584 14517 39593
rect 14475 39544 14476 39584
rect 14516 39544 14517 39584
rect 14475 39535 14517 39544
rect 14667 39584 14709 39593
rect 14667 39544 14668 39584
rect 14708 39544 14709 39584
rect 14667 39535 14709 39544
rect 14379 39500 14421 39509
rect 14379 39460 14380 39500
rect 14420 39460 14421 39500
rect 14379 39451 14421 39460
rect 14092 39376 14228 39416
rect 13995 39332 14037 39341
rect 13995 39292 13996 39332
rect 14036 39292 14037 39332
rect 13995 39283 14037 39292
rect 14092 39164 14132 39173
rect 13900 39124 14092 39164
rect 14092 39115 14132 39124
rect 13708 37820 13748 38872
rect 13804 38828 13844 38837
rect 13804 38669 13844 38788
rect 13803 38660 13845 38669
rect 13803 38620 13804 38660
rect 13844 38620 13845 38660
rect 13803 38611 13845 38620
rect 13995 38324 14037 38333
rect 13995 38284 13996 38324
rect 14036 38284 14037 38324
rect 13995 38275 14037 38284
rect 13899 38240 13941 38249
rect 13899 38200 13900 38240
rect 13940 38200 13941 38240
rect 13899 38191 13941 38200
rect 13900 38106 13940 38191
rect 13803 38072 13845 38081
rect 13803 38032 13804 38072
rect 13844 38032 13845 38072
rect 13803 38023 13845 38032
rect 13612 37780 13748 37820
rect 13612 36737 13652 37780
rect 13804 37414 13844 38023
rect 13804 37365 13844 37374
rect 13996 37316 14036 38275
rect 14091 38072 14133 38081
rect 14091 38032 14092 38072
rect 14132 38032 14133 38072
rect 14091 38023 14133 38032
rect 14092 37938 14132 38023
rect 14188 37820 14228 39376
rect 14283 39332 14325 39341
rect 14283 39292 14284 39332
rect 14324 39292 14325 39332
rect 14283 39283 14325 39292
rect 14284 38912 14324 39283
rect 14284 38863 14324 38872
rect 14380 38912 14420 39451
rect 14380 38863 14420 38872
rect 14476 38828 14516 39535
rect 14572 38921 14612 39006
rect 14571 38912 14613 38921
rect 14571 38872 14572 38912
rect 14612 38872 14613 38912
rect 14571 38863 14613 38872
rect 14476 38779 14516 38788
rect 14668 38744 14708 39535
rect 14859 39164 14901 39173
rect 14859 39124 14860 39164
rect 14900 39124 14901 39164
rect 14859 39115 14901 39124
rect 14572 38704 14708 38744
rect 14188 37780 14324 37820
rect 13996 37267 14036 37276
rect 14284 37400 14324 37780
rect 14475 37652 14517 37661
rect 14475 37612 14476 37652
rect 14516 37612 14517 37652
rect 14475 37603 14517 37612
rect 14284 36821 14324 37360
rect 14476 36896 14516 37603
rect 14476 36847 14516 36856
rect 14572 36821 14612 38704
rect 14667 38240 14709 38249
rect 14667 38200 14668 38240
rect 14708 38200 14709 38240
rect 14667 38191 14709 38200
rect 14283 36812 14325 36821
rect 14283 36772 14284 36812
rect 14324 36772 14325 36812
rect 14283 36763 14325 36772
rect 14571 36812 14613 36821
rect 14571 36772 14572 36812
rect 14612 36772 14613 36812
rect 14571 36763 14613 36772
rect 13611 36728 13653 36737
rect 13804 36728 13844 36737
rect 13611 36688 13612 36728
rect 13652 36688 13653 36728
rect 13611 36679 13653 36688
rect 13708 36688 13804 36728
rect 13612 34553 13652 36679
rect 13611 34544 13653 34553
rect 13611 34504 13612 34544
rect 13652 34504 13653 34544
rect 13611 34495 13653 34504
rect 13612 34376 13652 34385
rect 13612 34049 13652 34336
rect 13708 34301 13748 36688
rect 13804 36679 13844 36688
rect 14332 36686 14372 36695
rect 14091 36644 14133 36653
rect 14091 36604 14092 36644
rect 14132 36604 14133 36644
rect 14332 36644 14372 36646
rect 14332 36604 14516 36644
rect 14091 36595 14133 36604
rect 13996 35300 14036 35309
rect 13900 35260 13996 35300
rect 13804 35202 13844 35211
rect 13804 34628 13844 35162
rect 13804 34579 13844 34588
rect 13803 34460 13845 34469
rect 13803 34420 13804 34460
rect 13844 34420 13845 34460
rect 13803 34411 13845 34420
rect 13707 34292 13749 34301
rect 13707 34252 13708 34292
rect 13748 34252 13749 34292
rect 13707 34243 13749 34252
rect 13611 34040 13653 34049
rect 13611 34000 13612 34040
rect 13652 34000 13653 34040
rect 13611 33991 13653 34000
rect 13515 33872 13557 33881
rect 13515 33832 13516 33872
rect 13556 33832 13557 33872
rect 13515 33823 13557 33832
rect 13323 33704 13365 33713
rect 13708 33704 13748 34243
rect 13323 33664 13324 33704
rect 13364 33664 13365 33704
rect 13323 33655 13365 33664
rect 13516 33664 13748 33704
rect 13227 31352 13269 31361
rect 13227 31312 13228 31352
rect 13268 31312 13269 31352
rect 13227 31303 13269 31312
rect 13324 31025 13364 33655
rect 13419 33620 13461 33629
rect 13419 33580 13420 33620
rect 13460 33580 13461 33620
rect 13419 33571 13461 33580
rect 13420 32957 13460 33571
rect 13419 32948 13461 32957
rect 13419 32908 13420 32948
rect 13460 32908 13461 32948
rect 13419 32899 13461 32908
rect 13035 31016 13077 31025
rect 13035 30976 13036 31016
rect 13076 30976 13077 31016
rect 13035 30967 13077 30976
rect 13323 31016 13365 31025
rect 13323 30976 13324 31016
rect 13364 30976 13365 31016
rect 13323 30967 13365 30976
rect 13227 30848 13269 30857
rect 13227 30808 13228 30848
rect 13268 30808 13269 30848
rect 13227 30799 13269 30808
rect 13131 30680 13173 30689
rect 13131 30640 13132 30680
rect 13172 30640 13173 30680
rect 13131 30631 13173 30640
rect 13228 30680 13268 30799
rect 13228 30631 13268 30640
rect 13324 30680 13364 30689
rect 13132 30546 13172 30631
rect 13324 30512 13364 30640
rect 13420 30680 13460 32899
rect 13516 32192 13556 33664
rect 13516 32143 13556 32152
rect 13515 30848 13557 30857
rect 13515 30808 13516 30848
rect 13556 30808 13557 30848
rect 13515 30799 13557 30808
rect 13420 30631 13460 30640
rect 13228 30472 13460 30512
rect 12940 30428 12980 30437
rect 13228 30428 13268 30472
rect 12980 30388 13268 30428
rect 12940 30379 12980 30388
rect 12844 30220 13364 30260
rect 12939 29924 12981 29933
rect 12844 29882 12884 29891
rect 12556 29842 12844 29882
rect 12939 29884 12940 29924
rect 12980 29884 12981 29924
rect 12939 29875 12981 29884
rect 12363 29168 12405 29177
rect 12363 29128 12364 29168
rect 12404 29128 12405 29168
rect 12363 29119 12405 29128
rect 12556 29168 12596 29842
rect 12844 29833 12884 29842
rect 12940 29756 12980 29875
rect 13035 29840 13077 29849
rect 13035 29800 13036 29840
rect 13076 29800 13077 29840
rect 13035 29791 13077 29800
rect 12748 29716 12980 29756
rect 13036 29756 13076 29791
rect 12748 29336 12788 29716
rect 13036 29705 13076 29716
rect 12939 29588 12981 29597
rect 12939 29548 12940 29588
rect 12980 29548 12981 29588
rect 12939 29539 12981 29548
rect 13131 29588 13173 29597
rect 13131 29548 13132 29588
rect 13172 29548 13173 29588
rect 13131 29539 13173 29548
rect 12748 29287 12788 29296
rect 12651 29252 12693 29261
rect 12651 29212 12652 29252
rect 12692 29212 12693 29252
rect 12651 29203 12693 29212
rect 12364 28580 12404 29119
rect 12459 29084 12501 29093
rect 12459 29044 12460 29084
rect 12500 29044 12501 29084
rect 12459 29035 12501 29044
rect 12364 28531 12404 28540
rect 12460 28328 12500 29035
rect 12460 28279 12500 28288
rect 12556 27917 12596 29128
rect 12652 29009 12692 29203
rect 12940 29179 12980 29539
rect 13132 29177 13172 29539
rect 12940 29130 12980 29139
rect 13131 29168 13173 29177
rect 13131 29128 13132 29168
rect 13172 29128 13173 29168
rect 13131 29119 13173 29128
rect 13132 29034 13172 29119
rect 12651 29000 12693 29009
rect 12651 28960 12652 29000
rect 12692 28960 12693 29000
rect 12651 28951 12693 28960
rect 12940 28916 12980 28925
rect 12843 28748 12885 28757
rect 12843 28708 12844 28748
rect 12884 28708 12885 28748
rect 12843 28699 12885 28708
rect 12747 28328 12789 28337
rect 12747 28288 12748 28328
rect 12788 28288 12789 28328
rect 12747 28279 12789 28288
rect 12844 28328 12884 28699
rect 12844 28279 12884 28288
rect 12940 28328 12980 28876
rect 13035 28916 13077 28925
rect 13324 28916 13364 30220
rect 13420 29840 13460 30472
rect 13516 29933 13556 30799
rect 13612 30680 13652 30691
rect 13612 30605 13652 30640
rect 13611 30596 13653 30605
rect 13611 30556 13612 30596
rect 13652 30556 13653 30596
rect 13611 30547 13653 30556
rect 13804 30512 13844 34411
rect 13900 32621 13940 35260
rect 13996 35251 14036 35260
rect 13996 34208 14036 34217
rect 13996 33713 14036 34168
rect 13995 33704 14037 33713
rect 13995 33664 13996 33704
rect 14036 33664 14037 33704
rect 13995 33655 14037 33664
rect 13899 32612 13941 32621
rect 13899 32572 13900 32612
rect 13940 32572 13941 32612
rect 13899 32563 13941 32572
rect 14092 32453 14132 36595
rect 14476 35729 14516 36604
rect 14475 35720 14517 35729
rect 14475 35680 14476 35720
rect 14516 35680 14517 35720
rect 14475 35671 14517 35680
rect 14475 34796 14517 34805
rect 14475 34756 14476 34796
rect 14516 34756 14517 34796
rect 14475 34747 14517 34756
rect 14187 34376 14229 34385
rect 14187 34336 14188 34376
rect 14228 34336 14229 34376
rect 14187 34327 14229 34336
rect 14188 34242 14228 34327
rect 14187 34040 14229 34049
rect 14187 34000 14188 34040
rect 14228 34000 14229 34040
rect 14187 33991 14229 34000
rect 14188 33704 14228 33991
rect 14228 33664 14324 33704
rect 14188 33655 14228 33664
rect 14091 32444 14133 32453
rect 14091 32404 14092 32444
rect 14132 32404 14133 32444
rect 14091 32395 14133 32404
rect 14188 32276 14228 32285
rect 13899 32192 13941 32201
rect 13899 32152 13900 32192
rect 13940 32152 13941 32192
rect 13899 32143 13941 32152
rect 13996 32178 14036 32187
rect 13900 31352 13940 32143
rect 13996 31772 14036 32138
rect 13996 31732 14132 31772
rect 13995 31604 14037 31613
rect 13995 31564 13996 31604
rect 14036 31564 14037 31604
rect 13995 31555 14037 31564
rect 14092 31604 14132 31732
rect 14092 31555 14132 31564
rect 13900 30689 13940 31312
rect 13899 30680 13941 30689
rect 13899 30640 13900 30680
rect 13940 30640 13941 30680
rect 13899 30631 13941 30640
rect 13804 30472 13847 30512
rect 13807 30428 13847 30472
rect 13804 30388 13847 30428
rect 13804 30344 13844 30388
rect 13612 30304 13844 30344
rect 13515 29924 13557 29933
rect 13515 29884 13516 29924
rect 13556 29884 13557 29924
rect 13515 29875 13557 29884
rect 13420 29765 13460 29800
rect 13419 29756 13461 29765
rect 13612 29756 13652 30304
rect 13996 30260 14036 31555
rect 13804 30220 14036 30260
rect 13707 30008 13749 30017
rect 13707 29968 13708 30008
rect 13748 29968 13749 30008
rect 13707 29959 13749 29968
rect 13419 29716 13420 29756
rect 13460 29716 13461 29756
rect 13419 29707 13461 29716
rect 13516 29716 13652 29756
rect 13708 29840 13748 29959
rect 13420 29168 13460 29707
rect 13420 29093 13460 29128
rect 13419 29084 13461 29093
rect 13419 29044 13420 29084
rect 13460 29044 13461 29084
rect 13419 29035 13461 29044
rect 13035 28876 13036 28916
rect 13076 28876 13077 28916
rect 13035 28867 13077 28876
rect 13132 28876 13364 28916
rect 12940 28279 12980 28288
rect 12748 28194 12788 28279
rect 12651 28160 12693 28169
rect 12651 28120 12652 28160
rect 12692 28120 12693 28160
rect 12651 28111 12693 28120
rect 12652 28026 12692 28111
rect 12075 27908 12117 27917
rect 12075 27868 12076 27908
rect 12116 27868 12117 27908
rect 12075 27859 12117 27868
rect 12267 27908 12309 27917
rect 12267 27868 12268 27908
rect 12308 27868 12309 27908
rect 12267 27859 12309 27868
rect 12555 27908 12597 27917
rect 12555 27868 12556 27908
rect 12596 27868 12597 27908
rect 12555 27859 12597 27868
rect 11980 27775 12020 27784
rect 12844 27824 12884 27833
rect 12844 27665 12884 27784
rect 12939 27824 12981 27833
rect 12939 27784 12940 27824
rect 12980 27784 12981 27824
rect 12939 27775 12981 27784
rect 11979 27656 12021 27665
rect 11822 27641 11862 27650
rect 11979 27616 11980 27656
rect 12020 27616 12021 27656
rect 11979 27607 12021 27616
rect 12076 27656 12116 27665
rect 11822 27497 11862 27601
rect 11980 27522 12020 27607
rect 11499 27448 11500 27488
rect 11540 27448 11541 27488
rect 11499 27439 11541 27448
rect 11596 27448 11732 27488
rect 11821 27488 11863 27497
rect 11821 27448 11822 27488
rect 11862 27448 11863 27488
rect 11500 26069 11540 27439
rect 11499 26060 11541 26069
rect 11499 26020 11500 26060
rect 11540 26020 11541 26060
rect 11499 26011 11541 26020
rect 11500 24641 11540 26011
rect 11499 24632 11541 24641
rect 11499 24592 11500 24632
rect 11540 24592 11541 24632
rect 11499 24583 11541 24592
rect 11499 23960 11541 23969
rect 11499 23920 11500 23960
rect 11540 23920 11541 23960
rect 11499 23911 11541 23920
rect 11500 23288 11540 23911
rect 11596 23801 11636 27448
rect 11821 27439 11863 27448
rect 11883 27320 11925 27329
rect 11788 27280 11884 27320
rect 11924 27280 11925 27320
rect 11691 27068 11733 27077
rect 11691 27028 11692 27068
rect 11732 27028 11733 27068
rect 11691 27019 11733 27028
rect 11692 25061 11732 27019
rect 11691 25052 11733 25061
rect 11691 25012 11692 25052
rect 11732 25012 11733 25052
rect 11691 25003 11733 25012
rect 11692 24641 11732 24726
rect 11691 24632 11733 24641
rect 11691 24592 11692 24632
rect 11732 24592 11733 24632
rect 11691 24583 11733 24592
rect 11788 24464 11828 27280
rect 11883 27271 11925 27280
rect 11979 26900 12021 26909
rect 11979 26860 11980 26900
rect 12020 26860 12021 26900
rect 11979 26851 12021 26860
rect 11884 26816 11924 26825
rect 11884 26657 11924 26776
rect 11883 26648 11925 26657
rect 11883 26608 11884 26648
rect 11924 26608 11925 26648
rect 11883 26599 11925 26608
rect 11884 26144 11924 26599
rect 11884 26095 11924 26104
rect 11980 25304 12020 26851
rect 12076 26825 12116 27616
rect 12267 27656 12309 27665
rect 12267 27616 12268 27656
rect 12308 27616 12309 27656
rect 12267 27607 12309 27616
rect 12364 27656 12404 27665
rect 12556 27656 12596 27665
rect 12404 27616 12500 27656
rect 12364 27607 12404 27616
rect 12268 27522 12308 27607
rect 12171 27488 12213 27497
rect 12171 27448 12172 27488
rect 12212 27448 12213 27488
rect 12171 27439 12213 27448
rect 12172 26984 12212 27439
rect 12363 27404 12405 27413
rect 12363 27364 12364 27404
rect 12404 27364 12405 27404
rect 12363 27355 12405 27364
rect 12364 27270 12404 27355
rect 12460 26984 12500 27616
rect 12556 27413 12596 27616
rect 12652 27656 12692 27665
rect 12652 27497 12692 27616
rect 12843 27656 12885 27665
rect 12843 27616 12844 27656
rect 12884 27616 12885 27656
rect 12843 27607 12885 27616
rect 12651 27488 12693 27497
rect 12651 27448 12652 27488
rect 12692 27448 12693 27488
rect 12651 27439 12693 27448
rect 12555 27404 12597 27413
rect 12555 27364 12556 27404
rect 12596 27364 12597 27404
rect 12555 27355 12597 27364
rect 12940 27320 12980 27775
rect 12172 26944 12404 26984
rect 12075 26816 12117 26825
rect 12075 26776 12076 26816
rect 12116 26776 12117 26816
rect 12075 26767 12117 26776
rect 12076 26648 12116 26657
rect 12172 26648 12212 26944
rect 12267 26816 12309 26825
rect 12267 26776 12268 26816
rect 12308 26776 12309 26816
rect 12267 26767 12309 26776
rect 12364 26816 12404 26944
rect 12460 26935 12500 26944
rect 12652 27280 12980 27320
rect 12364 26767 12404 26776
rect 12555 26816 12597 26825
rect 12555 26776 12556 26816
rect 12596 26776 12597 26816
rect 12555 26767 12597 26776
rect 12116 26608 12212 26648
rect 12076 26599 12116 26608
rect 12076 26312 12116 26321
rect 12268 26312 12308 26767
rect 12556 26682 12596 26767
rect 12116 26272 12308 26312
rect 12076 26263 12116 26272
rect 12171 26144 12213 26153
rect 12171 26104 12172 26144
rect 12212 26104 12213 26144
rect 12171 26095 12213 26104
rect 12076 25304 12116 25313
rect 11980 25264 12076 25304
rect 12076 25255 12116 25264
rect 11883 24968 11925 24977
rect 11883 24928 11884 24968
rect 11924 24928 11925 24968
rect 11883 24919 11925 24928
rect 11884 24800 11924 24919
rect 11884 24751 11924 24760
rect 12172 24548 12212 26095
rect 12652 25313 12692 27280
rect 12843 26564 12885 26573
rect 12843 26524 12844 26564
rect 12884 26524 12885 26564
rect 12843 26515 12885 26524
rect 12556 25304 12596 25313
rect 12268 25220 12308 25229
rect 12556 25220 12596 25264
rect 12651 25304 12693 25313
rect 12651 25264 12652 25304
rect 12692 25264 12693 25304
rect 12651 25255 12693 25264
rect 12308 25180 12596 25220
rect 12268 25171 12308 25180
rect 12652 25170 12692 25255
rect 12267 24968 12309 24977
rect 12267 24928 12268 24968
rect 12308 24928 12309 24968
rect 12267 24919 12309 24928
rect 12268 24644 12308 24919
rect 12268 24595 12308 24604
rect 12363 24632 12405 24641
rect 12363 24592 12364 24632
rect 12404 24592 12405 24632
rect 12363 24583 12405 24592
rect 12460 24632 12500 24641
rect 12172 24508 12308 24548
rect 11692 24424 11828 24464
rect 11595 23792 11637 23801
rect 11595 23752 11596 23792
rect 11636 23752 11637 23792
rect 11595 23743 11637 23752
rect 11692 23624 11732 24424
rect 11884 24380 11924 24389
rect 12076 24380 12116 24389
rect 11500 23239 11540 23248
rect 11596 23584 11732 23624
rect 11788 24340 11884 24380
rect 11596 21701 11636 23584
rect 11691 23456 11733 23465
rect 11691 23416 11692 23456
rect 11732 23416 11733 23456
rect 11691 23407 11733 23416
rect 11595 21692 11637 21701
rect 11595 21652 11596 21692
rect 11636 21652 11637 21692
rect 11595 21643 11637 21652
rect 11596 20768 11636 20777
rect 11596 20189 11636 20728
rect 11595 20180 11637 20189
rect 11404 20140 11540 20180
rect 11307 19928 11349 19937
rect 11307 19888 11308 19928
rect 11348 19888 11349 19928
rect 11307 19879 11349 19888
rect 11308 19349 11348 19879
rect 11403 19592 11445 19601
rect 11403 19552 11404 19592
rect 11444 19552 11445 19592
rect 11403 19543 11445 19552
rect 11307 19340 11349 19349
rect 11307 19300 11308 19340
rect 11348 19300 11349 19340
rect 11307 19291 11349 19300
rect 11308 17417 11348 19291
rect 11307 17408 11349 17417
rect 11307 17368 11308 17408
rect 11348 17368 11349 17408
rect 11307 17359 11349 17368
rect 11307 17072 11349 17081
rect 11307 17032 11308 17072
rect 11348 17032 11349 17072
rect 11307 17023 11349 17032
rect 11308 16938 11348 17023
rect 11308 16232 11348 16243
rect 11308 16157 11348 16192
rect 11307 16148 11349 16157
rect 11307 16108 11308 16148
rect 11348 16108 11349 16148
rect 11307 16099 11349 16108
rect 11116 14428 11252 14468
rect 11307 14468 11349 14477
rect 11307 14428 11308 14468
rect 11348 14428 11349 14468
rect 11116 13376 11156 14428
rect 11307 14419 11349 14428
rect 11211 14048 11253 14057
rect 11211 14008 11212 14048
rect 11252 14008 11253 14048
rect 11211 13999 11253 14008
rect 11308 14048 11348 14419
rect 11308 13999 11348 14008
rect 11212 13914 11252 13999
rect 11307 13796 11349 13805
rect 11307 13756 11308 13796
rect 11348 13756 11349 13796
rect 11307 13747 11349 13756
rect 11116 13336 11252 13376
rect 10636 11320 10868 11360
rect 10924 13252 11060 13292
rect 10539 10940 10581 10949
rect 10539 10900 10540 10940
rect 10580 10900 10581 10940
rect 10539 10891 10581 10900
rect 10540 10361 10580 10891
rect 10539 10352 10581 10361
rect 10539 10312 10540 10352
rect 10580 10312 10581 10352
rect 10539 10303 10581 10312
rect 10540 9512 10580 10303
rect 10540 9463 10580 9472
rect 10347 9260 10389 9269
rect 10347 9220 10348 9260
rect 10388 9220 10389 9260
rect 10347 9211 10389 9220
rect 10347 8924 10389 8933
rect 10347 8884 10348 8924
rect 10388 8884 10389 8924
rect 10347 8875 10389 8884
rect 10251 7496 10293 7505
rect 10251 7456 10252 7496
rect 10292 7456 10293 7496
rect 10251 7447 10293 7456
rect 10252 7160 10292 7447
rect 10252 7111 10292 7120
rect 10155 5984 10197 5993
rect 10155 5944 10156 5984
rect 10196 5944 10197 5984
rect 10155 5935 10197 5944
rect 10251 5732 10293 5741
rect 10251 5692 10252 5732
rect 10292 5692 10293 5732
rect 10251 5683 10293 5692
rect 9964 3844 10100 3884
rect 10156 5648 10196 5657
rect 9867 2792 9909 2801
rect 9867 2752 9868 2792
rect 9908 2752 9909 2792
rect 9867 2743 9909 2752
rect 9868 2658 9908 2743
rect 9867 2456 9909 2465
rect 9867 2416 9868 2456
rect 9908 2416 9909 2456
rect 9867 2407 9909 2416
rect 9771 2372 9813 2381
rect 9771 2332 9772 2372
rect 9812 2332 9813 2372
rect 9771 2323 9813 2332
rect 9868 1952 9908 2407
rect 9772 1912 9868 1952
rect 9484 1660 9620 1700
rect 9676 1700 9716 1709
rect 9387 1028 9429 1037
rect 9387 988 9388 1028
rect 9428 988 9429 1028
rect 9387 979 9429 988
rect 9291 524 9333 533
rect 9291 484 9292 524
rect 9332 484 9333 524
rect 9291 475 9333 484
rect 9292 80 9332 475
rect 9484 80 9524 1660
rect 9579 1532 9621 1541
rect 9579 1492 9580 1532
rect 9620 1492 9621 1532
rect 9579 1483 9621 1492
rect 9580 1112 9620 1483
rect 9676 1289 9716 1660
rect 9772 1457 9812 1912
rect 9868 1903 9908 1912
rect 9964 1784 10004 3844
rect 10156 3641 10196 5608
rect 10252 5598 10292 5683
rect 10251 4808 10293 4817
rect 10251 4768 10252 4808
rect 10292 4768 10293 4808
rect 10251 4759 10293 4768
rect 10252 4136 10292 4759
rect 10348 4220 10388 8875
rect 10444 8168 10484 9388
rect 10636 8672 10676 11320
rect 10924 11192 10964 13252
rect 11116 13208 11156 13217
rect 11116 12965 11156 13168
rect 11115 12956 11157 12965
rect 11115 12916 11116 12956
rect 11156 12916 11157 12956
rect 11115 12907 11157 12916
rect 11115 12536 11157 12545
rect 11115 12496 11116 12536
rect 11156 12496 11157 12536
rect 11115 12487 11157 12496
rect 11116 12368 11156 12487
rect 11116 12319 11156 12328
rect 11212 11789 11252 13336
rect 11308 12452 11348 13747
rect 11308 12403 11348 12412
rect 11019 11780 11061 11789
rect 11019 11740 11020 11780
rect 11060 11740 11061 11780
rect 11019 11731 11061 11740
rect 11211 11780 11253 11789
rect 11211 11740 11212 11780
rect 11252 11740 11253 11780
rect 11211 11731 11253 11740
rect 11020 11360 11060 11731
rect 11020 11320 11348 11360
rect 10924 11152 11060 11192
rect 10732 11068 10964 11108
rect 10732 11024 10772 11068
rect 10732 10975 10772 10984
rect 10827 10940 10869 10949
rect 10827 10900 10828 10940
rect 10868 10900 10869 10940
rect 10827 10891 10869 10900
rect 10828 10806 10868 10891
rect 10924 8765 10964 11068
rect 11020 9689 11060 11152
rect 11308 11024 11348 11320
rect 11308 10975 11348 10984
rect 11320 10193 11360 10212
rect 11308 10184 11360 10193
rect 11404 10184 11444 19543
rect 11500 15401 11540 20140
rect 11595 20140 11596 20180
rect 11636 20140 11637 20180
rect 11595 20131 11637 20140
rect 11596 19181 11636 20131
rect 11595 19172 11637 19181
rect 11595 19132 11596 19172
rect 11636 19132 11637 19172
rect 11595 19123 11637 19132
rect 11595 17072 11637 17081
rect 11595 17032 11596 17072
rect 11636 17032 11637 17072
rect 11595 17023 11637 17032
rect 11499 15392 11541 15401
rect 11499 15352 11500 15392
rect 11540 15352 11541 15392
rect 11499 15343 11541 15352
rect 11499 12536 11541 12545
rect 11499 12496 11500 12536
rect 11540 12496 11541 12536
rect 11499 12487 11541 12496
rect 11500 12402 11540 12487
rect 11596 12377 11636 17023
rect 11692 15653 11732 23407
rect 11788 23120 11828 24340
rect 11884 24331 11924 24340
rect 11980 24340 12076 24380
rect 11883 23792 11925 23801
rect 11883 23752 11884 23792
rect 11924 23752 11925 23792
rect 11883 23743 11925 23752
rect 11884 23465 11924 23743
rect 11883 23456 11925 23465
rect 11883 23416 11884 23456
rect 11924 23416 11925 23456
rect 11883 23407 11925 23416
rect 11788 23071 11828 23080
rect 11883 23120 11925 23129
rect 11883 23080 11884 23120
rect 11924 23080 11925 23120
rect 11883 23071 11925 23080
rect 11980 23120 12020 24340
rect 12076 24331 12116 24340
rect 12171 24380 12213 24389
rect 12171 24340 12172 24380
rect 12212 24340 12213 24380
rect 12171 24331 12213 24340
rect 12172 23960 12212 24331
rect 12076 23920 12212 23960
rect 12076 23288 12116 23920
rect 12172 23792 12212 23801
rect 12268 23792 12308 24508
rect 12364 24221 12404 24583
rect 12363 24212 12405 24221
rect 12363 24172 12364 24212
rect 12404 24172 12405 24212
rect 12363 24163 12405 24172
rect 12460 23969 12500 24592
rect 12748 24632 12788 24641
rect 12748 24473 12788 24592
rect 12747 24464 12789 24473
rect 12747 24424 12748 24464
rect 12788 24424 12789 24464
rect 12747 24415 12789 24424
rect 12844 23969 12884 26515
rect 13036 25556 13076 28867
rect 13132 28328 13172 28876
rect 13516 28832 13556 29716
rect 13708 29672 13748 29800
rect 13132 28001 13172 28288
rect 13324 28792 13556 28832
rect 13612 29632 13748 29672
rect 13804 29840 13844 30220
rect 14188 30017 14228 32236
rect 14284 32117 14324 33664
rect 14380 33452 14420 33461
rect 14380 33041 14420 33412
rect 14476 33209 14516 34747
rect 14572 33536 14612 36763
rect 14668 35888 14708 38191
rect 14763 36140 14805 36149
rect 14763 36100 14764 36140
rect 14804 36100 14805 36140
rect 14763 36091 14805 36100
rect 14668 34385 14708 35848
rect 14764 35468 14804 36091
rect 14860 35972 14900 39115
rect 14956 38921 14996 39712
rect 14955 38912 14997 38921
rect 14955 38872 14956 38912
rect 14996 38872 14997 38912
rect 14955 38863 14997 38872
rect 15052 37820 15092 41140
rect 15148 40256 15188 41896
rect 15531 41432 15573 41441
rect 15531 41392 15532 41432
rect 15572 41392 15573 41432
rect 15531 41383 15573 41392
rect 15628 41432 15668 41441
rect 15724 41432 15764 41896
rect 15819 41936 15861 41945
rect 15819 41896 15820 41936
rect 15860 41896 15861 41936
rect 15819 41887 15861 41896
rect 15820 41802 15860 41887
rect 15915 41516 15957 41525
rect 15915 41476 15916 41516
rect 15956 41476 15957 41516
rect 15915 41467 15957 41476
rect 15668 41392 15764 41432
rect 15628 41383 15668 41392
rect 15436 41264 15476 41275
rect 15436 41189 15476 41224
rect 15243 41180 15285 41189
rect 15243 41140 15244 41180
rect 15284 41140 15285 41180
rect 15243 41131 15285 41140
rect 15435 41180 15477 41189
rect 15435 41140 15436 41180
rect 15476 41140 15477 41180
rect 15435 41131 15477 41140
rect 15244 40424 15284 41131
rect 15435 40676 15477 40685
rect 15435 40636 15436 40676
rect 15476 40636 15477 40676
rect 15435 40627 15477 40636
rect 15339 40592 15381 40601
rect 15339 40552 15340 40592
rect 15380 40552 15381 40592
rect 15339 40543 15381 40552
rect 15244 40375 15284 40384
rect 15148 40216 15284 40256
rect 15147 40004 15189 40013
rect 15147 39964 15148 40004
rect 15188 39964 15189 40004
rect 15147 39955 15189 39964
rect 15148 39752 15188 39955
rect 15244 39929 15284 40216
rect 15243 39920 15285 39929
rect 15243 39880 15244 39920
rect 15284 39880 15285 39920
rect 15340 39920 15380 40543
rect 15436 40542 15476 40627
rect 15436 39920 15476 39929
rect 15340 39880 15436 39920
rect 15243 39871 15285 39880
rect 15436 39871 15476 39880
rect 15148 39703 15188 39712
rect 15244 39752 15284 39761
rect 15147 39584 15189 39593
rect 15147 39544 15148 39584
rect 15188 39544 15189 39584
rect 15147 39535 15189 39544
rect 14956 37780 15092 37820
rect 14956 36149 14996 37780
rect 15148 37577 15188 39535
rect 15244 38837 15284 39712
rect 15340 39752 15380 39761
rect 15340 39089 15380 39712
rect 15435 39752 15477 39761
rect 15435 39712 15436 39752
rect 15476 39712 15477 39752
rect 15435 39703 15477 39712
rect 15339 39080 15381 39089
rect 15339 39040 15340 39080
rect 15380 39040 15381 39080
rect 15339 39031 15381 39040
rect 15436 38912 15476 39703
rect 15532 39593 15572 41383
rect 15916 41264 15956 41467
rect 15916 40760 15956 41224
rect 16108 40937 16148 42652
rect 16300 42608 16340 47347
rect 16491 47312 16533 47321
rect 16491 47272 16492 47312
rect 16532 47272 16533 47312
rect 16491 47263 16533 47272
rect 16492 47178 16532 47263
rect 16588 47060 16628 48019
rect 16396 47020 16628 47060
rect 16396 46640 16436 47020
rect 16587 46808 16629 46817
rect 16587 46768 16588 46808
rect 16628 46768 16629 46808
rect 16587 46759 16629 46768
rect 16396 46600 16532 46640
rect 16492 44960 16532 46600
rect 16492 44288 16532 44920
rect 16492 44239 16532 44248
rect 16588 42860 16628 46759
rect 16684 42944 16724 52051
rect 16780 52025 16820 54832
rect 16876 54200 16916 55000
rect 16972 54284 17012 55579
rect 17067 55544 17109 55553
rect 17067 55504 17068 55544
rect 17108 55504 17109 55544
rect 17067 55495 17109 55504
rect 17068 55410 17108 55495
rect 17067 55040 17109 55049
rect 17067 55000 17068 55040
rect 17108 55000 17109 55040
rect 17067 54991 17109 55000
rect 17068 54704 17108 54991
rect 17068 54655 17108 54664
rect 17164 54461 17204 55915
rect 17451 55712 17493 55721
rect 17451 55672 17452 55712
rect 17492 55672 17493 55712
rect 17451 55663 17493 55672
rect 17452 55544 17492 55663
rect 17452 55495 17492 55504
rect 17260 55460 17300 55469
rect 17260 55217 17300 55420
rect 17259 55208 17301 55217
rect 17259 55168 17260 55208
rect 17300 55168 17301 55208
rect 17259 55159 17301 55168
rect 17835 55208 17877 55217
rect 17835 55168 17836 55208
rect 17876 55168 17877 55208
rect 17835 55159 17877 55168
rect 17836 54872 17876 55159
rect 17836 54823 17876 54832
rect 17932 54872 17972 57016
rect 18124 56384 18164 58108
rect 18124 56057 18164 56344
rect 18123 56048 18165 56057
rect 18123 56008 18124 56048
rect 18164 56008 18165 56048
rect 18123 55999 18165 56008
rect 18123 55712 18165 55721
rect 18123 55672 18124 55712
rect 18164 55672 18165 55712
rect 18123 55663 18165 55672
rect 18124 55460 18164 55663
rect 17163 54452 17205 54461
rect 17163 54412 17164 54452
rect 17204 54412 17205 54452
rect 17163 54403 17205 54412
rect 17835 54368 17877 54377
rect 17835 54328 17836 54368
rect 17876 54328 17877 54368
rect 17835 54319 17877 54328
rect 16972 54244 17204 54284
rect 16876 54160 17108 54200
rect 16971 54032 17013 54041
rect 16971 53992 16972 54032
rect 17012 53992 17013 54032
rect 16971 53983 17013 53992
rect 16875 53024 16917 53033
rect 16875 52984 16876 53024
rect 16916 52984 16917 53024
rect 16875 52975 16917 52984
rect 16779 52016 16821 52025
rect 16779 51976 16780 52016
rect 16820 51976 16821 52016
rect 16779 51967 16821 51976
rect 16780 51848 16820 51857
rect 16780 51689 16820 51808
rect 16779 51680 16821 51689
rect 16779 51640 16780 51680
rect 16820 51640 16821 51680
rect 16779 51631 16821 51640
rect 16876 48152 16916 52975
rect 16972 52520 17012 53983
rect 16972 50345 17012 52480
rect 16971 50336 17013 50345
rect 16971 50296 16972 50336
rect 17012 50296 17013 50336
rect 16971 50287 17013 50296
rect 16972 48413 17012 50287
rect 17068 49085 17108 54160
rect 17164 53360 17204 54244
rect 17739 54200 17781 54209
rect 17739 54160 17740 54200
rect 17780 54160 17781 54200
rect 17739 54151 17781 54160
rect 17836 54200 17876 54319
rect 17836 54151 17876 54160
rect 17643 54116 17685 54125
rect 17643 54076 17644 54116
rect 17684 54076 17685 54116
rect 17643 54067 17685 54076
rect 17644 53982 17684 54067
rect 17204 53320 17300 53360
rect 17164 53311 17204 53320
rect 17163 52436 17205 52445
rect 17163 52396 17164 52436
rect 17204 52396 17205 52436
rect 17163 52387 17205 52396
rect 17164 52302 17204 52387
rect 17163 52016 17205 52025
rect 17163 51976 17164 52016
rect 17204 51976 17205 52016
rect 17163 51967 17205 51976
rect 17164 50429 17204 51967
rect 17260 50756 17300 53320
rect 17356 53108 17396 53117
rect 17356 51848 17396 53068
rect 17643 52940 17685 52949
rect 17643 52900 17644 52940
rect 17684 52900 17685 52940
rect 17643 52891 17685 52900
rect 17547 52856 17589 52865
rect 17547 52816 17548 52856
rect 17588 52816 17589 52856
rect 17547 52807 17589 52816
rect 17452 52520 17492 52531
rect 17452 52445 17492 52480
rect 17548 52520 17588 52807
rect 17451 52436 17493 52445
rect 17451 52396 17452 52436
rect 17492 52396 17493 52436
rect 17451 52387 17493 52396
rect 17356 51799 17396 51808
rect 17452 51848 17492 51857
rect 17548 51848 17588 52480
rect 17492 51808 17588 51848
rect 17452 51799 17492 51808
rect 17547 51008 17589 51017
rect 17547 50968 17548 51008
rect 17588 50968 17589 51008
rect 17547 50959 17589 50968
rect 17548 50765 17588 50959
rect 17355 50756 17397 50765
rect 17260 50716 17356 50756
rect 17396 50716 17397 50756
rect 17355 50707 17397 50716
rect 17547 50756 17589 50765
rect 17547 50716 17548 50756
rect 17588 50716 17589 50756
rect 17547 50707 17589 50716
rect 17163 50420 17205 50429
rect 17163 50380 17164 50420
rect 17204 50380 17205 50420
rect 17163 50371 17205 50380
rect 17356 50315 17396 50707
rect 17644 50429 17684 52891
rect 17740 51680 17780 54151
rect 17932 52604 17972 54832
rect 18028 55420 18164 55460
rect 18028 54032 18068 55420
rect 18028 53983 18068 53992
rect 18027 53696 18069 53705
rect 18027 53656 18028 53696
rect 18068 53656 18069 53696
rect 18027 53647 18069 53656
rect 17836 52564 17932 52604
rect 17836 51848 17876 52564
rect 17932 52555 17972 52564
rect 18028 52604 18068 53647
rect 17836 51799 17876 51808
rect 17932 51848 17972 51857
rect 18028 51848 18068 52564
rect 17972 51808 18068 51848
rect 17932 51799 17972 51808
rect 17740 51640 17876 51680
rect 17740 50840 17780 50849
rect 17740 50513 17780 50800
rect 17739 50504 17781 50513
rect 17739 50464 17740 50504
rect 17780 50464 17781 50504
rect 17739 50455 17781 50464
rect 17643 50420 17685 50429
rect 17643 50380 17644 50420
rect 17684 50380 17685 50420
rect 17643 50371 17685 50380
rect 17356 50266 17396 50275
rect 17836 50252 17876 51640
rect 18027 50504 18069 50513
rect 18027 50464 18028 50504
rect 18068 50464 18069 50504
rect 18027 50455 18069 50464
rect 17931 50336 17973 50345
rect 17931 50296 17932 50336
rect 17972 50296 17973 50336
rect 17931 50287 17973 50296
rect 17644 50212 17876 50252
rect 17548 50084 17588 50093
rect 17164 50044 17548 50084
rect 17067 49076 17109 49085
rect 17067 49036 17068 49076
rect 17108 49036 17109 49076
rect 17067 49027 17109 49036
rect 17164 48824 17204 50044
rect 17548 50035 17588 50044
rect 17116 48814 17204 48824
rect 17156 48784 17204 48814
rect 17260 48908 17300 48917
rect 17116 48765 17156 48774
rect 16971 48404 17013 48413
rect 16971 48364 16972 48404
rect 17012 48364 17013 48404
rect 16971 48355 17013 48364
rect 17260 48329 17300 48868
rect 17259 48320 17301 48329
rect 17259 48280 17260 48320
rect 17300 48280 17301 48320
rect 17259 48271 17301 48280
rect 16876 48112 17396 48152
rect 17259 47984 17301 47993
rect 17259 47944 17260 47984
rect 17300 47944 17301 47984
rect 17259 47935 17301 47944
rect 16971 47816 17013 47825
rect 16971 47776 16972 47816
rect 17012 47776 17013 47816
rect 16971 47767 17013 47776
rect 16972 47307 17012 47767
rect 16972 47258 17012 47267
rect 17164 47396 17204 47405
rect 17164 46817 17204 47356
rect 17163 46808 17205 46817
rect 17163 46768 17164 46808
rect 17204 46768 17205 46808
rect 17163 46759 17205 46768
rect 16972 46481 17012 46566
rect 16971 46472 17013 46481
rect 16971 46432 16972 46472
rect 17012 46432 17013 46472
rect 16971 46423 17013 46432
rect 17164 46304 17204 46313
rect 16876 46264 17164 46304
rect 16876 44876 16916 46264
rect 17164 46255 17204 46264
rect 17068 45800 17108 45809
rect 17260 45800 17300 47935
rect 17356 46640 17396 48112
rect 17356 46600 17588 46640
rect 17355 46472 17397 46481
rect 17355 46432 17356 46472
rect 17396 46432 17397 46472
rect 17355 46423 17397 46432
rect 17356 45809 17396 46423
rect 17451 46052 17493 46061
rect 17451 46012 17452 46052
rect 17492 46012 17493 46052
rect 17451 46003 17493 46012
rect 16972 45760 17068 45800
rect 17108 45760 17300 45800
rect 17355 45800 17397 45809
rect 17355 45760 17356 45800
rect 17396 45760 17397 45800
rect 16972 45389 17012 45760
rect 17068 45751 17108 45760
rect 17355 45751 17397 45760
rect 17452 45800 17492 46003
rect 17452 45751 17492 45760
rect 17355 45632 17397 45641
rect 17355 45592 17356 45632
rect 17396 45592 17397 45632
rect 17355 45583 17397 45592
rect 17260 45548 17300 45557
rect 17068 45508 17260 45548
rect 16971 45380 17013 45389
rect 16971 45340 16972 45380
rect 17012 45340 17013 45380
rect 16971 45331 17013 45340
rect 17068 45044 17108 45508
rect 17260 45499 17300 45508
rect 17020 45004 17108 45044
rect 17020 45002 17060 45004
rect 17020 44953 17060 44962
rect 16876 44836 17012 44876
rect 16972 44283 17012 44836
rect 17164 44792 17204 44801
rect 16972 44234 17012 44243
rect 17068 44752 17164 44792
rect 16684 42904 16916 42944
rect 16588 42820 16724 42860
rect 16300 42559 16340 42568
rect 16588 42692 16628 42701
rect 16204 41936 16244 41945
rect 16107 40928 16149 40937
rect 16107 40888 16108 40928
rect 16148 40888 16149 40928
rect 16107 40879 16149 40888
rect 15628 40720 15956 40760
rect 15531 39584 15573 39593
rect 15531 39544 15532 39584
rect 15572 39544 15573 39584
rect 15531 39535 15573 39544
rect 15340 38872 15476 38912
rect 15243 38828 15285 38837
rect 15243 38788 15244 38828
rect 15284 38788 15285 38828
rect 15243 38779 15285 38788
rect 15243 38408 15285 38417
rect 15243 38368 15244 38408
rect 15284 38368 15285 38408
rect 15243 38359 15285 38368
rect 15147 37568 15189 37577
rect 15147 37528 15148 37568
rect 15188 37528 15189 37568
rect 15147 37519 15189 37528
rect 15148 37232 15188 37519
rect 15244 37409 15284 38359
rect 15340 37652 15380 38872
rect 15628 38576 15668 40720
rect 16107 40676 16149 40685
rect 16204 40676 16244 41896
rect 16107 40636 16108 40676
rect 16148 40636 16244 40676
rect 16300 41936 16340 41945
rect 16107 40627 16149 40636
rect 15723 40592 15765 40601
rect 16300 40592 16340 41896
rect 16395 41768 16437 41777
rect 16395 41728 16396 41768
rect 16436 41728 16437 41768
rect 16395 41719 16437 41728
rect 15723 40552 15724 40592
rect 15764 40552 15765 40592
rect 15723 40543 15765 40552
rect 16204 40552 16340 40592
rect 15724 40424 15764 40543
rect 15819 40508 15861 40517
rect 15819 40468 15820 40508
rect 15860 40468 15861 40508
rect 15819 40459 15861 40468
rect 16204 40508 16244 40552
rect 15724 40375 15764 40384
rect 15820 40424 15860 40459
rect 15723 40004 15765 40013
rect 15723 39964 15724 40004
rect 15764 39964 15765 40004
rect 15723 39955 15765 39964
rect 15436 38536 15668 38576
rect 15724 39752 15764 39955
rect 15436 37913 15476 38536
rect 15724 38417 15764 39712
rect 15723 38408 15765 38417
rect 15723 38368 15724 38408
rect 15764 38368 15765 38408
rect 15723 38359 15765 38368
rect 15532 38240 15572 38249
rect 15435 37904 15477 37913
rect 15435 37864 15436 37904
rect 15476 37864 15477 37904
rect 15435 37855 15477 37864
rect 15436 37736 15476 37855
rect 15532 37820 15572 38200
rect 15628 38240 15668 38249
rect 15820 38240 15860 40384
rect 16107 40340 16149 40349
rect 16107 40300 16108 40340
rect 16148 40300 16149 40340
rect 16107 40291 16149 40300
rect 15668 38200 15860 38240
rect 15628 38191 15668 38200
rect 15532 37780 15764 37820
rect 15436 37696 15668 37736
rect 15340 37612 15572 37652
rect 15243 37400 15285 37409
rect 15243 37360 15244 37400
rect 15284 37360 15285 37400
rect 15243 37351 15285 37360
rect 15532 37400 15572 37612
rect 15148 37192 15284 37232
rect 15051 36896 15093 36905
rect 15051 36856 15052 36896
rect 15092 36856 15093 36896
rect 15051 36847 15093 36856
rect 14955 36140 14997 36149
rect 14955 36100 14956 36140
rect 14996 36100 14997 36140
rect 14955 36091 14997 36100
rect 15052 36056 15092 36847
rect 15052 36016 15188 36056
rect 14860 35932 15092 35972
rect 15052 35888 15092 35932
rect 15052 35839 15092 35848
rect 14859 35720 14901 35729
rect 15148 35720 15188 36016
rect 14859 35680 14860 35720
rect 14900 35680 14901 35720
rect 14859 35671 14901 35680
rect 15052 35680 15188 35720
rect 14860 35586 14900 35671
rect 14764 35428 14996 35468
rect 14667 34376 14709 34385
rect 14667 34336 14668 34376
rect 14708 34336 14709 34376
rect 14667 34327 14709 34336
rect 14668 33713 14708 33798
rect 14667 33704 14709 33713
rect 14667 33664 14668 33704
rect 14708 33664 14709 33704
rect 14667 33655 14709 33664
rect 14764 33704 14804 33713
rect 14804 33664 14900 33704
rect 14764 33655 14804 33664
rect 14572 33496 14708 33536
rect 14475 33200 14517 33209
rect 14475 33160 14476 33200
rect 14516 33160 14517 33200
rect 14475 33151 14517 33160
rect 14379 33032 14421 33041
rect 14379 32992 14380 33032
rect 14420 32992 14421 33032
rect 14379 32983 14421 32992
rect 14571 32696 14613 32705
rect 14571 32656 14572 32696
rect 14612 32656 14613 32696
rect 14571 32647 14613 32656
rect 14283 32108 14325 32117
rect 14283 32068 14284 32108
rect 14324 32068 14325 32108
rect 14283 32059 14325 32068
rect 14380 31352 14420 31361
rect 14420 31312 14516 31352
rect 14380 31303 14420 31312
rect 14284 31184 14324 31193
rect 14092 30008 14132 30017
rect 13131 27992 13173 28001
rect 13131 27952 13132 27992
rect 13172 27952 13173 27992
rect 13131 27943 13173 27952
rect 13132 26153 13172 27943
rect 13324 27833 13364 28792
rect 13515 28664 13557 28673
rect 13515 28624 13516 28664
rect 13556 28624 13557 28664
rect 13515 28615 13557 28624
rect 13516 28001 13556 28615
rect 13515 27992 13557 28001
rect 13515 27952 13516 27992
rect 13556 27952 13557 27992
rect 13515 27943 13557 27952
rect 13323 27824 13365 27833
rect 13612 27824 13652 29632
rect 13707 29504 13749 29513
rect 13707 29464 13708 29504
rect 13748 29464 13749 29504
rect 13707 29455 13749 29464
rect 13708 29168 13748 29455
rect 13804 29345 13844 29800
rect 13996 29968 14092 30008
rect 13803 29336 13845 29345
rect 13803 29296 13804 29336
rect 13844 29296 13845 29336
rect 13803 29287 13845 29296
rect 13708 29119 13748 29128
rect 13804 29168 13844 29179
rect 13804 29093 13844 29128
rect 13803 29084 13845 29093
rect 13803 29044 13804 29084
rect 13844 29044 13845 29084
rect 13803 29035 13845 29044
rect 13899 29000 13941 29009
rect 13899 28960 13900 29000
rect 13940 28960 13941 29000
rect 13899 28951 13941 28960
rect 13803 28916 13845 28925
rect 13803 28876 13804 28916
rect 13844 28876 13845 28916
rect 13803 28867 13845 28876
rect 13707 28664 13749 28673
rect 13707 28624 13708 28664
rect 13748 28624 13749 28664
rect 13707 28615 13749 28624
rect 13708 28421 13748 28615
rect 13707 28412 13749 28421
rect 13707 28372 13708 28412
rect 13748 28372 13749 28412
rect 13707 28363 13749 28372
rect 13707 28160 13749 28169
rect 13707 28120 13708 28160
rect 13748 28120 13749 28160
rect 13707 28111 13749 28120
rect 13323 27784 13324 27824
rect 13364 27784 13365 27824
rect 13323 27775 13365 27784
rect 13420 27784 13652 27824
rect 13227 27740 13269 27749
rect 13227 27700 13228 27740
rect 13268 27700 13269 27740
rect 13227 27691 13269 27700
rect 13228 27656 13268 27691
rect 13228 27605 13268 27616
rect 13323 27656 13365 27665
rect 13323 27616 13324 27656
rect 13364 27616 13365 27656
rect 13323 27607 13365 27616
rect 13324 27522 13364 27607
rect 13227 27488 13269 27497
rect 13227 27448 13228 27488
rect 13268 27448 13269 27488
rect 13227 27439 13269 27448
rect 13131 26144 13173 26153
rect 13131 26104 13132 26144
rect 13172 26104 13173 26144
rect 13131 26095 13173 26104
rect 12940 25516 13076 25556
rect 12459 23960 12501 23969
rect 12459 23920 12460 23960
rect 12500 23920 12501 23960
rect 12459 23911 12501 23920
rect 12843 23960 12885 23969
rect 12843 23920 12844 23960
rect 12884 23920 12885 23960
rect 12843 23911 12885 23920
rect 12212 23752 12308 23792
rect 12172 23743 12212 23752
rect 12076 23239 12116 23248
rect 12268 23129 12308 23752
rect 12652 23792 12692 23801
rect 12364 23708 12404 23717
rect 12652 23708 12692 23752
rect 12404 23668 12692 23708
rect 12748 23792 12788 23801
rect 12364 23659 12404 23668
rect 12748 23549 12788 23752
rect 12843 23792 12885 23801
rect 12843 23752 12844 23792
rect 12884 23752 12885 23792
rect 12843 23743 12885 23752
rect 12747 23540 12789 23549
rect 12747 23500 12748 23540
rect 12788 23500 12789 23540
rect 12747 23491 12789 23500
rect 11980 23071 12020 23080
rect 12267 23120 12309 23129
rect 12267 23080 12268 23120
rect 12308 23080 12309 23120
rect 12267 23071 12309 23080
rect 11884 22986 11924 23071
rect 12555 23036 12597 23045
rect 12555 22996 12556 23036
rect 12596 22996 12597 23036
rect 12555 22987 12597 22996
rect 12556 22625 12596 22987
rect 12651 22700 12693 22709
rect 12651 22660 12652 22700
rect 12692 22660 12693 22700
rect 12651 22651 12693 22660
rect 11883 22616 11925 22625
rect 11883 22576 11884 22616
rect 11924 22576 11925 22616
rect 11883 22567 11925 22576
rect 12555 22616 12597 22625
rect 12555 22576 12556 22616
rect 12596 22576 12597 22616
rect 12555 22567 12597 22576
rect 11788 22280 11828 22289
rect 11788 21533 11828 22240
rect 11787 21524 11829 21533
rect 11787 21484 11788 21524
rect 11828 21484 11829 21524
rect 11787 21475 11829 21484
rect 11884 17081 11924 22567
rect 12363 22448 12405 22457
rect 12363 22408 12364 22448
rect 12404 22408 12405 22448
rect 12363 22399 12405 22408
rect 12268 22280 12308 22289
rect 11980 22196 12020 22205
rect 12268 22196 12308 22240
rect 12020 22156 12308 22196
rect 12364 22280 12404 22399
rect 11980 22147 12020 22156
rect 12364 21953 12404 22240
rect 12363 21944 12405 21953
rect 12363 21904 12364 21944
rect 12404 21904 12405 21944
rect 12363 21895 12405 21904
rect 11979 21692 12021 21701
rect 11979 21652 11980 21692
rect 12020 21652 12021 21692
rect 11979 21643 12021 21652
rect 11980 20096 12020 21643
rect 12268 21608 12308 21617
rect 12268 21449 12308 21568
rect 12267 21440 12309 21449
rect 12267 21400 12268 21440
rect 12308 21400 12309 21440
rect 12267 21391 12309 21400
rect 12124 20777 12164 20786
rect 12164 20737 12212 20768
rect 12124 20728 12212 20737
rect 12172 20264 12212 20728
rect 12268 20600 12308 20609
rect 12308 20560 12404 20600
rect 12268 20551 12308 20560
rect 12268 20264 12308 20273
rect 12172 20224 12268 20264
rect 12268 20215 12308 20224
rect 12076 20096 12116 20124
rect 11980 20056 12076 20096
rect 11980 19769 12020 20056
rect 12076 20047 12116 20056
rect 11979 19760 12021 19769
rect 11979 19720 11980 19760
rect 12020 19720 12021 19760
rect 11979 19711 12021 19720
rect 11980 18929 12020 19711
rect 12075 19676 12117 19685
rect 12075 19636 12076 19676
rect 12116 19636 12117 19676
rect 12075 19627 12117 19636
rect 12076 19256 12116 19627
rect 12364 19340 12404 20560
rect 11979 18920 12021 18929
rect 11979 18880 11980 18920
rect 12020 18880 12021 18920
rect 11979 18871 12021 18880
rect 12076 18845 12116 19216
rect 12172 19300 12404 19340
rect 12075 18836 12117 18845
rect 12075 18796 12076 18836
rect 12116 18796 12117 18836
rect 12075 18787 12117 18796
rect 11883 17072 11925 17081
rect 11883 17032 11884 17072
rect 11924 17032 11925 17072
rect 11883 17023 11925 17032
rect 11836 16241 11876 16250
rect 11876 16201 11924 16232
rect 11836 16192 11924 16201
rect 11691 15644 11733 15653
rect 11691 15604 11692 15644
rect 11732 15604 11733 15644
rect 11691 15595 11733 15604
rect 11691 15476 11733 15485
rect 11691 15436 11692 15476
rect 11732 15436 11733 15476
rect 11691 15427 11733 15436
rect 11692 14552 11732 15427
rect 11787 15392 11829 15401
rect 11787 15352 11788 15392
rect 11828 15352 11829 15392
rect 11787 15343 11829 15352
rect 11788 14720 11828 15343
rect 11884 14972 11924 16192
rect 12172 16073 12212 19300
rect 12556 19256 12596 19265
rect 12268 19172 12308 19181
rect 12556 19172 12596 19216
rect 12652 19256 12692 22651
rect 12748 22457 12788 23491
rect 12844 23465 12884 23743
rect 12843 23456 12885 23465
rect 12843 23416 12844 23456
rect 12884 23416 12885 23456
rect 12843 23407 12885 23416
rect 12747 22448 12789 22457
rect 12747 22408 12748 22448
rect 12788 22408 12789 22448
rect 12747 22399 12789 22408
rect 12844 22364 12884 23407
rect 12844 22315 12884 22324
rect 12940 23120 12980 25516
rect 13035 25388 13077 25397
rect 13035 25348 13036 25388
rect 13076 25348 13077 25388
rect 13035 25339 13077 25348
rect 13036 25254 13076 25339
rect 13131 25304 13173 25313
rect 13131 25264 13132 25304
rect 13172 25264 13173 25304
rect 13131 25255 13173 25264
rect 13132 25170 13172 25255
rect 13228 25052 13268 27439
rect 13323 27152 13365 27161
rect 13323 27112 13324 27152
rect 13364 27112 13365 27152
rect 13323 27103 13365 27112
rect 12747 22280 12789 22289
rect 12747 22240 12748 22280
rect 12788 22240 12789 22280
rect 12747 22231 12789 22240
rect 12748 22146 12788 22231
rect 12843 21356 12885 21365
rect 12843 21316 12844 21356
rect 12884 21316 12885 21356
rect 12843 21307 12885 21316
rect 12844 20096 12884 21307
rect 12844 20021 12884 20056
rect 12843 20012 12885 20021
rect 12843 19972 12844 20012
rect 12884 19972 12885 20012
rect 12843 19963 12885 19972
rect 12692 19216 12884 19256
rect 12652 19207 12692 19216
rect 12308 19132 12596 19172
rect 12268 19123 12308 19132
rect 12363 18920 12405 18929
rect 12363 18880 12364 18920
rect 12404 18880 12405 18920
rect 12363 18871 12405 18880
rect 12267 18836 12309 18845
rect 12267 18796 12268 18836
rect 12308 18796 12309 18836
rect 12267 18787 12309 18796
rect 12268 18593 12308 18787
rect 12267 18584 12309 18593
rect 12267 18544 12268 18584
rect 12308 18544 12309 18584
rect 12267 18535 12309 18544
rect 11980 16064 12020 16073
rect 12171 16064 12213 16073
rect 12020 16024 12116 16064
rect 11980 16015 12020 16024
rect 11980 14972 12020 14981
rect 11884 14932 11980 14972
rect 11980 14923 12020 14932
rect 11788 14636 11828 14680
rect 11788 14596 12020 14636
rect 11692 14512 11828 14552
rect 11788 14048 11828 14512
rect 11883 14132 11925 14141
rect 11883 14092 11884 14132
rect 11924 14092 11925 14132
rect 11883 14083 11925 14092
rect 11788 13999 11828 14008
rect 11692 13964 11732 13975
rect 11692 13889 11732 13924
rect 11691 13880 11733 13889
rect 11691 13840 11692 13880
rect 11732 13840 11733 13880
rect 11691 13831 11733 13840
rect 11884 12704 11924 14083
rect 11980 13628 12020 14596
rect 12076 13805 12116 16024
rect 12171 16024 12172 16064
rect 12212 16024 12213 16064
rect 12171 16015 12213 16024
rect 12268 15812 12308 18535
rect 12364 15812 12404 18871
rect 12460 18668 12500 18677
rect 12500 18628 12788 18668
rect 12460 18619 12500 18628
rect 12748 18584 12788 18628
rect 12748 18535 12788 18544
rect 12844 18584 12884 19216
rect 12459 17828 12501 17837
rect 12459 17788 12460 17828
rect 12500 17788 12501 17828
rect 12459 17779 12501 17788
rect 12460 17669 12500 17779
rect 12459 17660 12501 17669
rect 12459 17620 12460 17660
rect 12500 17620 12501 17660
rect 12459 17611 12501 17620
rect 12555 17240 12597 17249
rect 12555 17200 12556 17240
rect 12596 17200 12597 17240
rect 12555 17191 12597 17200
rect 12556 17072 12596 17191
rect 12556 17023 12596 17032
rect 12748 16820 12788 16829
rect 12748 16232 12788 16780
rect 12748 16183 12788 16192
rect 12844 16232 12884 18544
rect 12268 15772 12311 15812
rect 12271 15728 12311 15772
rect 12267 15688 12311 15728
rect 12353 15772 12404 15812
rect 12267 15644 12307 15688
rect 12267 15604 12308 15644
rect 12268 15560 12308 15604
rect 12353 15560 12393 15772
rect 12460 15644 12500 15653
rect 12500 15604 12788 15644
rect 12460 15595 12500 15604
rect 12748 15560 12788 15604
rect 12353 15520 12404 15560
rect 12268 15511 12308 15520
rect 12267 15224 12309 15233
rect 12267 15184 12268 15224
rect 12308 15184 12309 15224
rect 12267 15175 12309 15184
rect 12268 14048 12308 15175
rect 12268 13999 12308 14008
rect 12075 13796 12117 13805
rect 12075 13756 12076 13796
rect 12116 13756 12117 13796
rect 12075 13747 12117 13756
rect 11980 13588 12116 13628
rect 11692 12664 11924 12704
rect 11595 12368 11637 12377
rect 11595 12328 11596 12368
rect 11636 12328 11637 12368
rect 11595 12319 11637 12328
rect 11595 12200 11637 12209
rect 11595 12160 11596 12200
rect 11636 12160 11637 12200
rect 11595 12151 11637 12160
rect 11348 10144 11444 10184
rect 11308 10135 11348 10144
rect 11404 10025 11444 10144
rect 11596 10109 11636 12151
rect 11595 10100 11637 10109
rect 11595 10060 11596 10100
rect 11636 10060 11637 10100
rect 11595 10051 11637 10060
rect 11403 10016 11445 10025
rect 11403 9976 11404 10016
rect 11444 9976 11445 10016
rect 11403 9967 11445 9976
rect 11692 9764 11732 12664
rect 11787 12368 11829 12377
rect 11787 12328 11788 12368
rect 11828 12328 11829 12368
rect 11787 12319 11829 12328
rect 11788 11696 11828 12319
rect 11788 11453 11828 11656
rect 11980 11528 12020 11537
rect 11787 11444 11829 11453
rect 11787 11404 11788 11444
rect 11828 11404 11829 11444
rect 11787 11395 11829 11404
rect 11980 11360 12020 11488
rect 11884 11320 12020 11360
rect 11884 11024 11924 11320
rect 11979 11192 12021 11201
rect 11979 11152 11980 11192
rect 12020 11152 12021 11192
rect 11979 11143 12021 11152
rect 11980 11058 12020 11143
rect 11836 11014 11924 11024
rect 11876 10984 11924 11014
rect 11836 10965 11876 10974
rect 12076 10184 12116 13588
rect 12171 13544 12213 13553
rect 12171 13504 12172 13544
rect 12212 13504 12213 13544
rect 12171 13495 12213 13504
rect 12172 11948 12212 13495
rect 12364 13217 12404 15520
rect 12748 15511 12788 15520
rect 12844 15560 12884 16192
rect 12844 14477 12884 15520
rect 12940 15317 12980 23080
rect 13036 25012 13268 25052
rect 13324 26816 13364 27103
rect 13036 20180 13076 25012
rect 13227 23960 13269 23969
rect 13227 23920 13228 23960
rect 13268 23920 13269 23960
rect 13227 23911 13269 23920
rect 13228 23876 13268 23911
rect 13131 23792 13173 23801
rect 13131 23752 13132 23792
rect 13172 23752 13173 23792
rect 13131 23743 13173 23752
rect 13132 23658 13172 23743
rect 13228 23045 13268 23836
rect 13324 23381 13364 26776
rect 13323 23372 13365 23381
rect 13323 23332 13324 23372
rect 13364 23332 13365 23372
rect 13323 23323 13365 23332
rect 13227 23036 13269 23045
rect 13227 22996 13228 23036
rect 13268 22996 13269 23036
rect 13227 22987 13269 22996
rect 13131 22784 13173 22793
rect 13131 22744 13132 22784
rect 13172 22744 13173 22784
rect 13131 22735 13173 22744
rect 13132 22289 13172 22735
rect 13227 22532 13269 22541
rect 13227 22492 13228 22532
rect 13268 22492 13269 22532
rect 13227 22483 13269 22492
rect 13131 22280 13173 22289
rect 13131 22240 13132 22280
rect 13172 22240 13173 22280
rect 13131 22231 13173 22240
rect 13228 20525 13268 22483
rect 13323 22280 13365 22289
rect 13323 22240 13324 22280
rect 13364 22240 13365 22280
rect 13323 22231 13365 22240
rect 13324 22146 13364 22231
rect 13227 20516 13269 20525
rect 13227 20476 13228 20516
rect 13268 20476 13269 20516
rect 13227 20467 13269 20476
rect 13036 20140 13172 20180
rect 13036 19256 13076 19265
rect 13036 18500 13076 19216
rect 13132 19256 13172 20140
rect 13132 18668 13172 19216
rect 13420 19013 13460 27784
rect 13516 27656 13556 27665
rect 13708 27656 13748 28111
rect 13556 27616 13652 27656
rect 13516 27607 13556 27616
rect 13612 27488 13652 27616
rect 13708 27607 13748 27616
rect 13708 27488 13748 27497
rect 13612 27448 13708 27488
rect 13708 27439 13748 27448
rect 13515 27404 13557 27413
rect 13515 27364 13516 27404
rect 13556 27364 13557 27404
rect 13515 27355 13557 27364
rect 13516 27270 13556 27355
rect 13707 27320 13749 27329
rect 13707 27280 13708 27320
rect 13748 27280 13749 27320
rect 13707 27271 13749 27280
rect 13611 26144 13653 26153
rect 13611 26104 13612 26144
rect 13652 26104 13653 26144
rect 13611 26095 13653 26104
rect 13612 26010 13652 26095
rect 13612 25304 13652 25313
rect 13708 25304 13748 27271
rect 13652 25264 13748 25304
rect 13612 25255 13652 25264
rect 13708 23792 13748 23801
rect 13708 23204 13748 23752
rect 13516 23164 13748 23204
rect 13516 22289 13556 23164
rect 13804 23120 13844 28867
rect 13900 27656 13940 28951
rect 13900 27607 13940 27616
rect 13996 27656 14036 29968
rect 14092 29959 14132 29968
rect 14187 30008 14229 30017
rect 14187 29968 14188 30008
rect 14228 29968 14229 30008
rect 14187 29959 14229 29968
rect 14187 29756 14229 29765
rect 14187 29716 14188 29756
rect 14228 29716 14229 29756
rect 14187 29707 14229 29716
rect 14091 29420 14133 29429
rect 14091 29380 14092 29420
rect 14132 29380 14133 29420
rect 14091 29371 14133 29380
rect 14092 29000 14132 29371
rect 14188 29168 14228 29707
rect 14284 29513 14324 31144
rect 14379 30092 14421 30101
rect 14379 30052 14380 30092
rect 14420 30052 14421 30092
rect 14379 30043 14421 30052
rect 14380 29840 14420 30043
rect 14476 29933 14516 31312
rect 14572 30101 14612 32647
rect 14571 30092 14613 30101
rect 14571 30052 14572 30092
rect 14612 30052 14613 30092
rect 14571 30043 14613 30052
rect 14475 29924 14517 29933
rect 14475 29884 14476 29924
rect 14516 29884 14517 29924
rect 14475 29875 14517 29884
rect 14380 29791 14420 29800
rect 14283 29504 14325 29513
rect 14283 29464 14284 29504
rect 14324 29464 14325 29504
rect 14283 29455 14325 29464
rect 14284 29345 14324 29455
rect 14283 29336 14325 29345
rect 14283 29296 14284 29336
rect 14324 29296 14325 29336
rect 14283 29287 14325 29296
rect 14284 29189 14324 29198
rect 14188 29149 14284 29168
rect 14476 29189 14516 29875
rect 14188 29128 14324 29149
rect 14380 29168 14420 29177
rect 14476 29140 14516 29149
rect 14572 29168 14612 29177
rect 14380 29084 14420 29128
rect 14475 29084 14517 29093
rect 14380 29044 14476 29084
rect 14516 29044 14517 29084
rect 14475 29035 14517 29044
rect 14092 28951 14132 28960
rect 14572 28757 14612 29128
rect 14571 28748 14613 28757
rect 14571 28708 14572 28748
rect 14612 28708 14613 28748
rect 14571 28699 14613 28708
rect 14374 28664 14416 28673
rect 14475 28664 14517 28673
rect 14374 28624 14375 28664
rect 14415 28624 14420 28664
rect 14374 28615 14420 28624
rect 14475 28624 14476 28664
rect 14516 28624 14517 28664
rect 14475 28615 14517 28624
rect 14091 28412 14133 28421
rect 14091 28372 14092 28412
rect 14132 28372 14133 28412
rect 14091 28363 14133 28372
rect 13996 27607 14036 27616
rect 14092 27488 14132 28363
rect 14380 28328 14420 28615
rect 14380 28279 14420 28288
rect 14379 28160 14421 28169
rect 14379 28120 14380 28160
rect 14420 28120 14421 28160
rect 14379 28111 14421 28120
rect 14283 27656 14325 27665
rect 14283 27616 14284 27656
rect 14324 27616 14325 27656
rect 14283 27607 14325 27616
rect 13900 27448 14132 27488
rect 13900 25313 13940 27448
rect 14187 27236 14229 27245
rect 14187 27196 14188 27236
rect 14228 27196 14229 27236
rect 14187 27187 14229 27196
rect 14188 25472 14228 27187
rect 13996 25432 14228 25472
rect 13899 25304 13941 25313
rect 13899 25264 13900 25304
rect 13940 25264 13941 25304
rect 13899 25255 13941 25264
rect 13612 23080 13844 23120
rect 13515 22280 13557 22289
rect 13515 22240 13516 22280
rect 13556 22240 13557 22280
rect 13515 22231 13557 22240
rect 13516 21608 13556 21619
rect 13516 21533 13556 21568
rect 13515 21524 13557 21533
rect 13515 21484 13516 21524
rect 13556 21484 13557 21524
rect 13515 21475 13557 21484
rect 13612 20180 13652 23080
rect 13804 22285 13844 22294
rect 13708 21776 13748 21785
rect 13804 21776 13844 22245
rect 13900 21869 13940 25255
rect 13996 24800 14036 25432
rect 14140 25313 14180 25322
rect 14284 25304 14324 27607
rect 14380 25388 14420 28111
rect 14476 27824 14516 28615
rect 14668 28421 14708 33496
rect 14763 33032 14805 33041
rect 14763 32992 14764 33032
rect 14804 32992 14805 33032
rect 14763 32983 14805 32992
rect 14764 32864 14804 32983
rect 14764 32815 14804 32824
rect 14860 32864 14900 33664
rect 14764 31352 14804 31361
rect 14764 31193 14804 31312
rect 14860 31352 14900 32824
rect 14763 31184 14805 31193
rect 14763 31144 14764 31184
rect 14804 31144 14805 31184
rect 14763 31135 14805 31144
rect 14860 31016 14900 31312
rect 14764 30976 14900 31016
rect 14764 30176 14804 30976
rect 14859 30680 14901 30689
rect 14859 30640 14860 30680
rect 14900 30640 14901 30680
rect 14859 30631 14901 30640
rect 14860 30546 14900 30631
rect 14859 30176 14901 30185
rect 14764 30136 14860 30176
rect 14900 30136 14901 30176
rect 14859 30127 14901 30136
rect 14763 29588 14805 29597
rect 14763 29548 14764 29588
rect 14804 29548 14805 29588
rect 14763 29539 14805 29548
rect 14764 29168 14804 29539
rect 14860 29345 14900 30127
rect 14956 29588 14996 35428
rect 15052 32369 15092 35680
rect 15244 34376 15284 37192
rect 15435 36980 15477 36989
rect 15435 36940 15436 36980
rect 15476 36940 15477 36980
rect 15435 36931 15477 36940
rect 15436 35216 15476 36931
rect 15532 36569 15572 37360
rect 15628 36989 15668 37696
rect 15724 37652 15764 37780
rect 15724 37603 15764 37612
rect 15627 36980 15669 36989
rect 15627 36940 15628 36980
rect 15668 36940 15669 36980
rect 15627 36931 15669 36940
rect 15628 36728 15668 36737
rect 15531 36560 15573 36569
rect 15531 36520 15532 36560
rect 15572 36520 15573 36560
rect 15531 36511 15573 36520
rect 15628 35729 15668 36688
rect 15723 36728 15765 36737
rect 15723 36688 15724 36728
rect 15764 36688 15765 36728
rect 15723 36679 15765 36688
rect 15724 36594 15764 36679
rect 15820 36653 15860 38200
rect 16108 38240 16148 40291
rect 16108 38191 16148 38200
rect 16012 38156 16052 38165
rect 16012 38072 16052 38116
rect 16204 38072 16244 40468
rect 16300 40424 16340 40435
rect 16300 40349 16340 40384
rect 16299 40340 16341 40349
rect 16299 40300 16300 40340
rect 16340 40300 16341 40340
rect 16299 40291 16341 40300
rect 16299 39080 16341 39089
rect 16299 39040 16300 39080
rect 16340 39040 16341 39080
rect 16299 39031 16341 39040
rect 16012 38032 16244 38072
rect 16011 37484 16053 37493
rect 16011 37444 16012 37484
rect 16052 37444 16053 37484
rect 16011 37435 16053 37444
rect 15915 37400 15957 37409
rect 15915 37360 15916 37400
rect 15956 37360 15957 37400
rect 15915 37351 15957 37360
rect 15916 37266 15956 37351
rect 15819 36644 15861 36653
rect 15819 36604 15820 36644
rect 15860 36604 15861 36644
rect 15819 36595 15861 36604
rect 16012 36476 16052 37435
rect 16108 36653 16148 36738
rect 16107 36644 16149 36653
rect 16107 36604 16108 36644
rect 16148 36604 16149 36644
rect 16107 36595 16149 36604
rect 16204 36644 16244 38032
rect 16300 38912 16340 39031
rect 16300 37829 16340 38872
rect 16299 37820 16341 37829
rect 16299 37780 16300 37820
rect 16340 37780 16341 37820
rect 16299 37771 16341 37780
rect 16012 36436 16148 36476
rect 15627 35720 15669 35729
rect 15627 35680 15628 35720
rect 15668 35680 15669 35720
rect 15627 35671 15669 35680
rect 15628 35216 15668 35225
rect 15436 35176 15628 35216
rect 15628 35167 15668 35176
rect 15436 34376 15476 34385
rect 15244 34336 15436 34376
rect 15436 34040 15476 34336
rect 15819 34376 15861 34385
rect 15819 34336 15820 34376
rect 15860 34336 15861 34376
rect 15819 34327 15861 34336
rect 15820 34242 15860 34327
rect 15628 34208 15668 34217
rect 15668 34168 15764 34208
rect 15628 34159 15668 34168
rect 15436 34000 15668 34040
rect 15148 33620 15188 33629
rect 15148 32864 15188 33580
rect 15244 33620 15284 33629
rect 15244 33041 15284 33580
rect 15243 33032 15285 33041
rect 15243 32992 15244 33032
rect 15284 32992 15285 33032
rect 15243 32983 15285 32992
rect 15244 32864 15284 32873
rect 15148 32824 15244 32864
rect 15051 32360 15093 32369
rect 15051 32320 15052 32360
rect 15092 32320 15093 32360
rect 15051 32311 15093 32320
rect 15051 32192 15093 32201
rect 15051 32152 15052 32192
rect 15092 32152 15093 32192
rect 15051 32143 15093 32152
rect 15052 32058 15092 32143
rect 15244 31352 15284 32824
rect 15340 32864 15380 32873
rect 15380 32824 15572 32864
rect 15340 32815 15380 32824
rect 15339 31688 15381 31697
rect 15339 31648 15340 31688
rect 15380 31648 15381 31688
rect 15339 31639 15381 31648
rect 15340 31436 15380 31639
rect 15340 31387 15380 31396
rect 15244 31268 15284 31312
rect 15244 31228 15380 31268
rect 15147 31184 15189 31193
rect 15147 31144 15148 31184
rect 15188 31144 15189 31184
rect 15147 31135 15189 31144
rect 15148 30932 15188 31135
rect 15052 30892 15188 30932
rect 15052 30848 15092 30892
rect 15052 30799 15092 30808
rect 15243 30680 15285 30689
rect 15243 30640 15244 30680
rect 15284 30640 15285 30680
rect 15243 30631 15285 30640
rect 15244 30546 15284 30631
rect 15243 29840 15285 29849
rect 15243 29800 15244 29840
rect 15284 29800 15285 29840
rect 15243 29791 15285 29800
rect 14956 29548 15092 29588
rect 14859 29336 14901 29345
rect 14859 29296 14860 29336
rect 14900 29296 14901 29336
rect 15052 29336 15092 29548
rect 15052 29296 15188 29336
rect 14859 29287 14901 29296
rect 14955 29252 14997 29261
rect 14955 29212 14956 29252
rect 14996 29212 14997 29252
rect 14955 29203 14997 29212
rect 14764 29119 14804 29128
rect 14860 29168 14900 29177
rect 14860 28757 14900 29128
rect 14956 29168 14996 29203
rect 14956 29117 14996 29128
rect 15052 29168 15092 29177
rect 14955 29000 14997 29009
rect 14955 28960 14956 29000
rect 14996 28960 14997 29000
rect 14955 28951 14997 28960
rect 14859 28748 14901 28757
rect 14859 28708 14860 28748
rect 14900 28708 14901 28748
rect 14859 28699 14901 28708
rect 14667 28412 14709 28421
rect 14667 28372 14668 28412
rect 14708 28372 14709 28412
rect 14667 28363 14709 28372
rect 14860 28328 14900 28337
rect 14572 28244 14612 28253
rect 14860 28244 14900 28288
rect 14956 28328 14996 28951
rect 15052 28337 15092 29128
rect 15148 28673 15188 29296
rect 15244 29168 15284 29791
rect 15244 29119 15284 29128
rect 15244 28925 15284 29010
rect 15243 28916 15285 28925
rect 15243 28876 15244 28916
rect 15284 28876 15285 28916
rect 15243 28867 15285 28876
rect 15340 28748 15380 31228
rect 15532 29588 15572 32824
rect 15628 30605 15668 34000
rect 15724 33881 15764 34168
rect 15819 34040 15861 34049
rect 15819 34000 15820 34040
rect 15860 34000 15861 34040
rect 15819 33991 15861 34000
rect 15723 33872 15765 33881
rect 15723 33832 15724 33872
rect 15764 33832 15765 33872
rect 15723 33823 15765 33832
rect 15724 33704 15764 33713
rect 15724 31613 15764 33664
rect 15820 32864 15860 33991
rect 16011 32864 16053 32873
rect 15860 32824 15956 32864
rect 15820 32815 15860 32824
rect 15723 31604 15765 31613
rect 15723 31564 15724 31604
rect 15764 31564 15765 31604
rect 15723 31555 15765 31564
rect 15724 31352 15764 31555
rect 15820 31352 15860 31361
rect 15724 31312 15820 31352
rect 15820 31303 15860 31312
rect 15916 31184 15956 32824
rect 16011 32824 16012 32864
rect 16052 32824 16053 32864
rect 16011 32815 16053 32824
rect 15724 31144 15956 31184
rect 15627 30596 15669 30605
rect 15627 30556 15628 30596
rect 15668 30556 15669 30596
rect 15627 30547 15669 30556
rect 15628 29849 15668 29934
rect 15627 29840 15669 29849
rect 15627 29800 15628 29840
rect 15668 29800 15669 29840
rect 15627 29791 15669 29800
rect 15532 29548 15668 29588
rect 15435 29504 15477 29513
rect 15435 29464 15436 29504
rect 15476 29464 15477 29504
rect 15435 29455 15477 29464
rect 15436 29168 15476 29455
rect 15531 29420 15573 29429
rect 15531 29380 15532 29420
rect 15572 29380 15573 29420
rect 15531 29371 15573 29380
rect 15436 29119 15476 29128
rect 15532 29168 15572 29371
rect 15532 29119 15572 29128
rect 15244 28708 15380 28748
rect 15147 28664 15189 28673
rect 15147 28624 15148 28664
rect 15188 28624 15189 28664
rect 15147 28615 15189 28624
rect 15244 28580 15284 28708
rect 15237 28540 15284 28580
rect 15237 28412 15277 28540
rect 15237 28372 15284 28412
rect 14956 28279 14996 28288
rect 15051 28328 15093 28337
rect 15051 28288 15052 28328
rect 15092 28288 15093 28328
rect 15244 28328 15284 28372
rect 15340 28328 15380 28337
rect 15244 28288 15340 28328
rect 15051 28279 15093 28288
rect 14612 28204 14900 28244
rect 14572 28195 14612 28204
rect 14955 28160 14997 28169
rect 14476 27775 14516 27784
rect 14764 28120 14956 28160
rect 14996 28120 14997 28160
rect 14471 27656 14511 27665
rect 14572 27656 14612 27665
rect 14511 27616 14516 27656
rect 14471 27607 14516 27616
rect 14476 26489 14516 27607
rect 14572 26993 14612 27616
rect 14668 27656 14708 27665
rect 14668 27068 14708 27616
rect 14764 27236 14804 28120
rect 14955 28111 14997 28120
rect 14859 27656 14901 27665
rect 14859 27616 14860 27656
rect 14900 27616 14901 27656
rect 14859 27607 14901 27616
rect 14956 27656 14996 27665
rect 15148 27656 15188 27665
rect 14996 27616 15092 27656
rect 14956 27607 14996 27616
rect 14860 27522 14900 27607
rect 14956 27404 14996 27415
rect 14956 27329 14996 27364
rect 14955 27320 14997 27329
rect 14955 27280 14956 27320
rect 14996 27280 14997 27320
rect 14955 27271 14997 27280
rect 14764 27196 14900 27236
rect 14763 27068 14805 27077
rect 14668 27028 14764 27068
rect 14804 27028 14805 27068
rect 14763 27019 14805 27028
rect 14571 26984 14613 26993
rect 14571 26944 14572 26984
rect 14612 26944 14613 26984
rect 14571 26935 14613 26944
rect 14764 26934 14804 27019
rect 14572 26816 14612 26825
rect 14860 26816 14900 27196
rect 14955 27068 14997 27077
rect 14955 27028 14956 27068
rect 14996 27028 14997 27068
rect 14955 27019 14997 27028
rect 14572 26657 14612 26776
rect 14764 26776 14900 26816
rect 14956 26816 14996 27019
rect 15052 26984 15092 27616
rect 15148 27161 15188 27616
rect 15147 27152 15189 27161
rect 15147 27112 15148 27152
rect 15188 27112 15189 27152
rect 15147 27103 15189 27112
rect 15052 26935 15092 26944
rect 14571 26648 14613 26657
rect 14571 26608 14572 26648
rect 14612 26608 14613 26648
rect 14571 26599 14613 26608
rect 14475 26480 14517 26489
rect 14475 26440 14476 26480
rect 14516 26440 14517 26480
rect 14475 26431 14517 26440
rect 14380 25348 14516 25388
rect 14180 25273 14228 25304
rect 14140 25264 14228 25273
rect 14284 25264 14420 25304
rect 14188 24800 14228 25264
rect 14284 25136 14324 25145
rect 14284 24977 14324 25096
rect 14283 24968 14325 24977
rect 14283 24928 14284 24968
rect 14324 24928 14325 24968
rect 14283 24919 14325 24928
rect 13996 24760 14132 24800
rect 13996 24632 14036 24643
rect 13996 24557 14036 24592
rect 13995 24548 14037 24557
rect 13995 24508 13996 24548
rect 14036 24508 14037 24548
rect 13995 24499 14037 24508
rect 14092 24128 14132 24760
rect 14188 24751 14228 24760
rect 13996 24088 14132 24128
rect 13996 23297 14036 24088
rect 14091 23960 14133 23969
rect 14091 23920 14092 23960
rect 14132 23920 14133 23960
rect 14091 23911 14133 23920
rect 13995 23288 14037 23297
rect 13995 23248 13996 23288
rect 14036 23248 14037 23288
rect 13995 23239 14037 23248
rect 13995 23120 14037 23129
rect 13995 23080 13996 23120
rect 14036 23080 14037 23120
rect 13995 23071 14037 23080
rect 13996 22280 14036 23071
rect 14092 22709 14132 23911
rect 14380 23885 14420 25264
rect 14379 23876 14421 23885
rect 14379 23836 14380 23876
rect 14420 23836 14421 23876
rect 14379 23827 14421 23836
rect 14236 23801 14276 23810
rect 14236 23624 14276 23761
rect 14379 23708 14421 23717
rect 14379 23668 14380 23708
rect 14420 23668 14421 23708
rect 14379 23659 14421 23668
rect 14236 23584 14324 23624
rect 14284 23372 14324 23584
rect 14380 23574 14420 23659
rect 14284 23332 14420 23372
rect 14380 23288 14420 23332
rect 14380 23239 14420 23248
rect 14187 23120 14229 23129
rect 14187 23080 14188 23120
rect 14228 23080 14229 23120
rect 14187 23071 14229 23080
rect 14188 22986 14228 23071
rect 14091 22700 14133 22709
rect 14091 22660 14092 22700
rect 14132 22660 14133 22700
rect 14091 22651 14133 22660
rect 14283 22700 14325 22709
rect 14283 22660 14284 22700
rect 14324 22660 14325 22700
rect 14283 22651 14325 22660
rect 13996 22240 14132 22280
rect 13996 22112 14036 22121
rect 13899 21860 13941 21869
rect 13899 21820 13900 21860
rect 13940 21820 13941 21860
rect 13899 21811 13941 21820
rect 13748 21736 13844 21776
rect 13708 21727 13748 21736
rect 13707 21608 13749 21617
rect 13707 21568 13708 21608
rect 13748 21568 13749 21608
rect 13707 21559 13749 21568
rect 13899 21608 13941 21617
rect 13899 21568 13900 21608
rect 13940 21568 13941 21608
rect 13899 21559 13941 21568
rect 13516 20140 13652 20180
rect 13708 20768 13748 21559
rect 13900 21474 13940 21559
rect 13996 21113 14036 22072
rect 14092 21944 14132 22240
rect 14092 21904 14228 21944
rect 13995 21104 14037 21113
rect 13995 21064 13996 21104
rect 14036 21064 14037 21104
rect 13995 21055 14037 21064
rect 13419 19004 13461 19013
rect 13419 18964 13420 19004
rect 13460 18964 13461 19004
rect 13419 18955 13461 18964
rect 13516 18677 13556 20140
rect 13611 19256 13653 19265
rect 13611 19216 13612 19256
rect 13652 19216 13653 19256
rect 13611 19207 13653 19216
rect 13612 19122 13652 19207
rect 13515 18668 13557 18677
rect 13132 18628 13364 18668
rect 13228 18500 13268 18509
rect 13036 18460 13228 18500
rect 13228 16232 13268 18460
rect 13324 18500 13364 18628
rect 13515 18628 13516 18668
rect 13556 18628 13557 18668
rect 13515 18619 13557 18628
rect 13324 17240 13364 18460
rect 13420 17744 13460 17755
rect 13420 17585 13460 17704
rect 13419 17576 13461 17585
rect 13419 17536 13420 17576
rect 13460 17536 13461 17576
rect 13419 17527 13461 17536
rect 13324 17200 13460 17240
rect 13323 17072 13365 17081
rect 13323 17032 13324 17072
rect 13364 17032 13365 17072
rect 13323 17023 13365 17032
rect 13324 16938 13364 17023
rect 13131 15644 13173 15653
rect 13131 15604 13132 15644
rect 13172 15604 13173 15644
rect 13131 15595 13173 15604
rect 12939 15308 12981 15317
rect 12939 15268 12940 15308
rect 12980 15268 12981 15308
rect 12939 15259 12981 15268
rect 13132 14720 13172 15595
rect 13228 15569 13268 16192
rect 13324 16232 13364 16241
rect 13420 16232 13460 17200
rect 13364 16192 13460 16232
rect 13227 15560 13269 15569
rect 13227 15520 13228 15560
rect 13268 15520 13269 15560
rect 13227 15511 13269 15520
rect 13228 15426 13268 15511
rect 13324 15485 13364 16192
rect 13708 15728 13748 20728
rect 13995 20768 14037 20777
rect 13995 20728 13996 20768
rect 14036 20728 14037 20768
rect 13995 20719 14037 20728
rect 13899 19424 13941 19433
rect 13899 19384 13900 19424
rect 13940 19384 13941 19424
rect 13899 19375 13941 19384
rect 13803 19256 13845 19265
rect 13803 19216 13804 19256
rect 13844 19216 13845 19256
rect 13803 19207 13845 19216
rect 13804 18584 13844 19207
rect 13804 16241 13844 18544
rect 13803 16232 13845 16241
rect 13803 16192 13804 16232
rect 13844 16192 13845 16232
rect 13803 16183 13845 16192
rect 13420 15688 13748 15728
rect 13323 15476 13365 15485
rect 13323 15436 13324 15476
rect 13364 15436 13365 15476
rect 13323 15427 13365 15436
rect 13324 15342 13364 15427
rect 13227 15308 13269 15317
rect 13227 15268 13228 15308
rect 13268 15268 13269 15308
rect 13227 15259 13269 15268
rect 12940 14680 13132 14720
rect 12843 14468 12885 14477
rect 12843 14428 12844 14468
rect 12884 14428 12885 14468
rect 12843 14419 12885 14428
rect 12940 14300 12980 14680
rect 13132 14671 13172 14680
rect 13228 14552 13268 15259
rect 12844 14260 12980 14300
rect 13132 14512 13268 14552
rect 12748 14034 12788 14043
rect 12556 13460 12596 13469
rect 12748 13460 12788 13994
rect 12596 13420 12788 13460
rect 12556 13411 12596 13420
rect 12651 13292 12693 13301
rect 12651 13252 12652 13292
rect 12692 13252 12693 13292
rect 12651 13243 12693 13252
rect 12363 13208 12405 13217
rect 12363 13168 12364 13208
rect 12404 13168 12405 13208
rect 12363 13159 12405 13168
rect 12364 13074 12404 13159
rect 12172 11899 12212 11908
rect 12652 11864 12692 13243
rect 12747 13208 12789 13217
rect 12747 13168 12748 13208
rect 12788 13168 12789 13208
rect 12747 13159 12789 13168
rect 12748 12536 12788 13159
rect 12844 12545 12884 14260
rect 13035 14216 13077 14225
rect 13035 14176 13036 14216
rect 13076 14176 13077 14216
rect 13035 14167 13077 14176
rect 12939 14132 12981 14141
rect 12939 14092 12940 14132
rect 12980 14092 12981 14132
rect 12939 14083 12981 14092
rect 12940 13998 12980 14083
rect 12940 12620 12980 12629
rect 13036 12620 13076 14167
rect 12980 12580 13076 12620
rect 13132 13208 13172 14512
rect 13227 14216 13269 14225
rect 13227 14176 13228 14216
rect 13268 14176 13269 14216
rect 13227 14167 13269 14176
rect 13228 14048 13268 14167
rect 13228 13999 13268 14008
rect 13323 14048 13365 14057
rect 13323 14008 13324 14048
rect 13364 14008 13365 14048
rect 13323 13999 13365 14008
rect 13227 13796 13269 13805
rect 13227 13756 13228 13796
rect 13268 13756 13269 13796
rect 13227 13747 13269 13756
rect 12940 12571 12980 12580
rect 12748 12377 12788 12496
rect 12843 12536 12885 12545
rect 12843 12496 12844 12536
rect 12884 12496 12885 12536
rect 12843 12487 12885 12496
rect 12747 12368 12789 12377
rect 12747 12328 12748 12368
rect 12788 12328 12789 12368
rect 12747 12319 12789 12328
rect 12652 11824 12788 11864
rect 12364 11780 12404 11789
rect 12364 11201 12404 11740
rect 12652 11696 12692 11707
rect 12652 11621 12692 11656
rect 12651 11612 12693 11621
rect 12651 11572 12652 11612
rect 12692 11572 12693 11612
rect 12651 11563 12693 11572
rect 12748 11360 12788 11824
rect 12652 11320 12788 11360
rect 12363 11192 12405 11201
rect 12363 11152 12364 11192
rect 12404 11152 12405 11192
rect 12363 11143 12405 11152
rect 12556 11024 12596 11033
rect 12556 10445 12596 10984
rect 12652 11024 12692 11320
rect 12555 10436 12597 10445
rect 12555 10396 12556 10436
rect 12596 10396 12597 10436
rect 12555 10387 12597 10396
rect 12556 10184 12596 10193
rect 12076 10144 12556 10184
rect 11787 10016 11829 10025
rect 11787 9976 11788 10016
rect 11828 9976 11829 10016
rect 11787 9967 11829 9976
rect 11979 10016 12021 10025
rect 11979 9976 11980 10016
rect 12020 9976 12021 10016
rect 11979 9967 12021 9976
rect 11404 9724 11732 9764
rect 11019 9680 11061 9689
rect 11019 9640 11020 9680
rect 11060 9640 11061 9680
rect 11019 9631 11061 9640
rect 11020 9512 11060 9521
rect 11060 9472 11348 9512
rect 11020 9463 11060 9472
rect 10923 8756 10965 8765
rect 10923 8716 10924 8756
rect 10964 8716 10965 8756
rect 10923 8707 10965 8716
rect 10676 8632 10772 8672
rect 10636 8623 10676 8632
rect 10444 8128 10676 8168
rect 10443 8000 10485 8009
rect 10443 7960 10444 8000
rect 10484 7960 10485 8000
rect 10443 7951 10485 7960
rect 10540 8000 10580 8009
rect 10444 6320 10484 7951
rect 10540 7505 10580 7960
rect 10636 7832 10676 8128
rect 10732 8009 10772 8632
rect 10731 8000 10773 8009
rect 10731 7960 10732 8000
rect 10772 7960 10773 8000
rect 10924 8000 10964 8707
rect 11020 8000 11060 8009
rect 10924 7960 11020 8000
rect 10731 7951 10773 7960
rect 11020 7951 11060 7960
rect 11116 7916 11156 7925
rect 11156 7876 11252 7916
rect 11116 7832 11156 7876
rect 10636 7792 11156 7832
rect 10539 7496 10581 7505
rect 10539 7456 10540 7496
rect 10580 7456 10581 7496
rect 10539 7447 10581 7456
rect 10540 7169 10580 7447
rect 10827 7328 10869 7337
rect 10827 7288 10828 7328
rect 10868 7288 10869 7328
rect 10827 7279 10869 7288
rect 10539 7160 10581 7169
rect 10731 7160 10773 7169
rect 10539 7120 10540 7160
rect 10580 7120 10581 7160
rect 10539 7111 10581 7120
rect 10636 7120 10732 7160
rect 10772 7120 10773 7160
rect 10540 6488 10580 6497
rect 10636 6488 10676 7120
rect 10731 7111 10773 7120
rect 10731 6656 10773 6665
rect 10731 6616 10732 6656
rect 10772 6616 10773 6656
rect 10731 6607 10773 6616
rect 10732 6522 10772 6607
rect 10580 6448 10676 6488
rect 10540 6439 10580 6448
rect 10444 6280 10580 6320
rect 10540 5060 10580 6280
rect 10828 6068 10868 7279
rect 11115 6992 11157 7001
rect 11115 6952 11116 6992
rect 11156 6952 11157 6992
rect 11115 6943 11157 6952
rect 11116 6404 11156 6943
rect 11116 6355 11156 6364
rect 10923 6320 10965 6329
rect 10923 6280 10924 6320
rect 10964 6280 10965 6320
rect 10923 6271 10965 6280
rect 10924 6186 10964 6271
rect 11212 6236 11252 7876
rect 11308 6320 11348 9472
rect 11404 6992 11444 9724
rect 11499 9596 11541 9605
rect 11499 9556 11500 9596
rect 11540 9556 11541 9596
rect 11499 9547 11541 9556
rect 11692 9596 11732 9605
rect 11500 9507 11540 9547
rect 11500 9458 11540 9467
rect 11499 9260 11541 9269
rect 11499 9220 11500 9260
rect 11540 9220 11541 9260
rect 11499 9211 11541 9220
rect 11500 8000 11540 9211
rect 11692 8429 11732 9556
rect 11691 8420 11733 8429
rect 11691 8380 11692 8420
rect 11732 8380 11733 8420
rect 11691 8371 11733 8380
rect 11500 7951 11540 7960
rect 11596 8000 11636 8009
rect 11500 7169 11540 7254
rect 11499 7160 11541 7169
rect 11499 7120 11500 7160
rect 11540 7120 11541 7160
rect 11499 7111 11541 7120
rect 11404 6952 11540 6992
rect 11403 6320 11445 6329
rect 11308 6280 11404 6320
rect 11444 6280 11445 6320
rect 11403 6271 11445 6280
rect 11212 6196 11348 6236
rect 11115 6068 11157 6077
rect 10828 6028 10964 6068
rect 10731 5648 10773 5657
rect 10731 5608 10732 5648
rect 10772 5608 10773 5648
rect 10731 5599 10773 5608
rect 10732 5514 10772 5599
rect 10540 5020 10868 5060
rect 10443 4976 10485 4985
rect 10443 4936 10444 4976
rect 10484 4936 10485 4976
rect 10443 4927 10485 4936
rect 10828 4976 10868 5020
rect 10444 4842 10484 4927
rect 10636 4724 10676 4733
rect 10636 4481 10676 4684
rect 10828 4565 10868 4936
rect 10827 4556 10869 4565
rect 10827 4516 10828 4556
rect 10868 4516 10869 4556
rect 10827 4507 10869 4516
rect 10635 4472 10677 4481
rect 10635 4432 10636 4472
rect 10676 4432 10677 4472
rect 10635 4423 10677 4432
rect 10827 4220 10869 4229
rect 10348 4180 10484 4220
rect 10155 3632 10197 3641
rect 10155 3592 10156 3632
rect 10196 3592 10197 3632
rect 10155 3583 10197 3592
rect 10252 3557 10292 4096
rect 10348 4116 10388 4125
rect 10348 3977 10388 4076
rect 10347 3968 10389 3977
rect 10347 3928 10348 3968
rect 10388 3928 10389 3968
rect 10347 3919 10389 3928
rect 10444 3716 10484 4180
rect 10827 4180 10828 4220
rect 10868 4180 10869 4220
rect 10827 4171 10869 4180
rect 10828 4086 10868 4171
rect 10348 3676 10484 3716
rect 10636 3968 10676 3977
rect 10348 3632 10388 3676
rect 10348 3583 10388 3592
rect 10251 3548 10293 3557
rect 10251 3508 10252 3548
rect 10292 3508 10293 3548
rect 10251 3499 10293 3508
rect 10204 3422 10244 3431
rect 10059 3380 10101 3389
rect 10059 3340 10060 3380
rect 10100 3340 10101 3380
rect 10540 3389 10580 3474
rect 10204 3380 10244 3382
rect 10539 3380 10581 3389
rect 10204 3340 10388 3380
rect 10059 3331 10101 3340
rect 10060 2624 10100 3331
rect 10060 2575 10100 2584
rect 10155 2624 10197 2633
rect 10155 2584 10156 2624
rect 10196 2584 10197 2624
rect 10155 2575 10197 2584
rect 10059 2204 10101 2213
rect 10059 2164 10060 2204
rect 10100 2164 10101 2204
rect 10059 2155 10101 2164
rect 9868 1744 10004 1784
rect 9771 1448 9813 1457
rect 9771 1408 9772 1448
rect 9812 1408 9813 1448
rect 9771 1399 9813 1408
rect 9675 1280 9717 1289
rect 9675 1240 9676 1280
rect 9716 1240 9717 1280
rect 9675 1231 9717 1240
rect 9580 1072 9716 1112
rect 9676 80 9716 1072
rect 9868 80 9908 1744
rect 10060 1112 10100 2155
rect 10060 1063 10100 1072
rect 10156 1028 10196 2575
rect 10348 2204 10388 3340
rect 10539 3340 10540 3380
rect 10580 3340 10581 3380
rect 10539 3331 10581 3340
rect 10539 3212 10581 3221
rect 10539 3172 10540 3212
rect 10580 3172 10581 3212
rect 10539 3163 10581 3172
rect 10252 2164 10388 2204
rect 10252 1280 10292 2164
rect 10347 2036 10389 2045
rect 10347 1996 10348 2036
rect 10388 1996 10389 2036
rect 10347 1987 10389 1996
rect 10252 1231 10292 1240
rect 10156 988 10292 1028
rect 10059 608 10101 617
rect 10059 568 10060 608
rect 10100 568 10101 608
rect 10059 559 10101 568
rect 10060 80 10100 559
rect 10252 80 10292 988
rect 10348 617 10388 1987
rect 10443 944 10485 953
rect 10443 904 10444 944
rect 10484 904 10485 944
rect 10443 895 10485 904
rect 10444 810 10484 895
rect 10540 692 10580 3163
rect 10636 2045 10676 3928
rect 10924 3380 10964 6028
rect 11115 6028 11116 6068
rect 11156 6028 11157 6068
rect 11115 6019 11157 6028
rect 10924 3331 10964 3340
rect 11020 3968 11060 3977
rect 11020 3305 11060 3928
rect 11116 3548 11156 6019
rect 11212 5653 11252 5662
rect 11212 4481 11252 5613
rect 11211 4472 11253 4481
rect 11211 4432 11212 4472
rect 11252 4432 11253 4472
rect 11211 4423 11253 4432
rect 11211 4220 11253 4229
rect 11211 4180 11212 4220
rect 11252 4180 11253 4220
rect 11211 4171 11253 4180
rect 11212 4086 11252 4171
rect 11308 4145 11348 6196
rect 11404 5564 11444 6271
rect 11404 5069 11444 5524
rect 11403 5060 11445 5069
rect 11403 5020 11404 5060
rect 11444 5020 11445 5060
rect 11403 5011 11445 5020
rect 11500 4220 11540 6952
rect 11596 6665 11636 7960
rect 11691 7412 11733 7421
rect 11691 7372 11692 7412
rect 11732 7372 11733 7412
rect 11691 7363 11733 7372
rect 11692 7278 11732 7363
rect 11595 6656 11637 6665
rect 11595 6616 11596 6656
rect 11636 6616 11637 6656
rect 11595 6607 11637 6616
rect 11788 5993 11828 9967
rect 11883 9596 11925 9605
rect 11883 9556 11884 9596
rect 11924 9556 11925 9596
rect 11883 9547 11925 9556
rect 11884 9462 11924 9547
rect 11883 8672 11925 8681
rect 11883 8632 11884 8672
rect 11924 8632 11925 8672
rect 11883 8623 11925 8632
rect 11884 8538 11924 8623
rect 11980 8336 12020 9967
rect 12268 9521 12308 10144
rect 12556 10135 12596 10144
rect 12652 10025 12692 10984
rect 12748 10445 12788 10530
rect 12747 10436 12789 10445
rect 12747 10396 12748 10436
rect 12788 10396 12789 10436
rect 12747 10387 12789 10396
rect 12651 10016 12693 10025
rect 12651 9976 12652 10016
rect 12692 9976 12693 10016
rect 12651 9967 12693 9976
rect 12555 9848 12597 9857
rect 12555 9808 12556 9848
rect 12596 9808 12597 9848
rect 12555 9799 12597 9808
rect 12075 9512 12117 9521
rect 12075 9472 12076 9512
rect 12116 9472 12117 9512
rect 12075 9463 12117 9472
rect 12267 9512 12309 9521
rect 12267 9472 12268 9512
rect 12308 9472 12309 9512
rect 12267 9463 12309 9472
rect 12076 9378 12116 9463
rect 12364 8672 12404 8681
rect 12076 8588 12116 8597
rect 12364 8588 12404 8632
rect 12460 8672 12500 8683
rect 12460 8597 12500 8632
rect 12116 8548 12404 8588
rect 12459 8588 12501 8597
rect 12459 8548 12460 8588
rect 12500 8548 12501 8588
rect 12076 8539 12116 8548
rect 12459 8539 12501 8548
rect 11980 8296 12212 8336
rect 12076 6488 12116 6497
rect 11787 5984 11829 5993
rect 11787 5944 11788 5984
rect 11828 5944 11829 5984
rect 11787 5935 11829 5944
rect 11595 5900 11637 5909
rect 11595 5860 11596 5900
rect 11636 5860 11637 5900
rect 11595 5851 11637 5860
rect 11596 5766 11636 5851
rect 11691 5816 11733 5825
rect 11691 5776 11692 5816
rect 11732 5776 11828 5816
rect 11691 5767 11733 5776
rect 11788 5743 11828 5776
rect 11788 5694 11828 5703
rect 11595 5648 11637 5657
rect 11595 5608 11596 5648
rect 11636 5608 11637 5648
rect 11595 5599 11637 5608
rect 11596 4817 11636 5599
rect 11980 5480 12020 5489
rect 11980 5321 12020 5440
rect 11979 5312 12021 5321
rect 11979 5272 11980 5312
rect 12020 5272 12021 5312
rect 11979 5263 12021 5272
rect 12076 5153 12116 6448
rect 12172 6488 12212 8296
rect 12460 8000 12500 8009
rect 12556 8000 12596 9799
rect 12844 9521 12884 12487
rect 13132 11360 13172 13168
rect 12940 11320 13172 11360
rect 12940 10016 12980 11320
rect 13132 11024 13172 11033
rect 13228 11024 13268 13747
rect 13324 13385 13364 13999
rect 13323 13376 13365 13385
rect 13323 13336 13324 13376
rect 13364 13336 13365 13376
rect 13323 13327 13365 13336
rect 13172 10984 13268 11024
rect 13132 10975 13172 10984
rect 13036 10940 13076 10949
rect 13036 10697 13076 10900
rect 13420 10856 13460 15688
rect 13804 15560 13844 16183
rect 13804 15511 13844 15520
rect 13611 14972 13653 14981
rect 13611 14932 13612 14972
rect 13652 14932 13653 14972
rect 13611 14923 13653 14932
rect 13132 10816 13460 10856
rect 13612 11024 13652 14923
rect 13803 14216 13845 14225
rect 13803 14176 13804 14216
rect 13844 14176 13845 14216
rect 13803 14167 13845 14176
rect 13708 13964 13748 13973
rect 13708 11453 13748 13924
rect 13804 13964 13844 14167
rect 13804 13805 13844 13924
rect 13803 13796 13845 13805
rect 13803 13756 13804 13796
rect 13844 13756 13845 13796
rect 13803 13747 13845 13756
rect 13900 12200 13940 19375
rect 13996 17249 14036 20719
rect 14092 20096 14132 20105
rect 14092 19685 14132 20056
rect 14091 19676 14133 19685
rect 14091 19636 14092 19676
rect 14132 19636 14133 19676
rect 14091 19627 14133 19636
rect 14188 19433 14228 21904
rect 14284 20105 14324 22651
rect 14379 22448 14421 22457
rect 14375 22408 14380 22448
rect 14420 22408 14421 22448
rect 14375 22399 14421 22408
rect 14375 22293 14415 22399
rect 14375 22244 14415 22253
rect 14476 22280 14516 25348
rect 14668 24632 14708 24641
rect 14668 24221 14708 24592
rect 14667 24212 14709 24221
rect 14667 24172 14668 24212
rect 14708 24172 14709 24212
rect 14667 24163 14709 24172
rect 14764 23885 14804 26776
rect 14956 26767 14996 26776
rect 15052 26816 15092 26825
rect 14859 26648 14901 26657
rect 14859 26608 14860 26648
rect 14900 26608 14901 26648
rect 14859 26599 14901 26608
rect 14860 26153 14900 26599
rect 15052 26489 15092 26776
rect 15243 26816 15285 26825
rect 15243 26776 15244 26816
rect 15284 26776 15285 26816
rect 15243 26767 15285 26776
rect 15244 26682 15284 26767
rect 15051 26480 15093 26489
rect 15051 26440 15052 26480
rect 15092 26440 15093 26480
rect 15051 26431 15093 26440
rect 15052 26312 15092 26431
rect 15092 26272 15284 26312
rect 15052 26263 15092 26272
rect 14859 26144 14901 26153
rect 14859 26104 14860 26144
rect 14900 26104 14901 26144
rect 14859 26095 14901 26104
rect 15244 26144 15284 26272
rect 15340 26228 15380 28288
rect 15436 28328 15476 28337
rect 15628 28328 15668 29548
rect 15724 28757 15764 31144
rect 15915 30092 15957 30101
rect 15915 30052 15916 30092
rect 15956 30052 15957 30092
rect 15915 30043 15957 30052
rect 15820 29672 15860 29681
rect 15820 29177 15860 29632
rect 15819 29168 15861 29177
rect 15819 29128 15820 29168
rect 15860 29128 15861 29168
rect 15916 29168 15956 30043
rect 16012 29840 16052 32815
rect 16012 29791 16052 29800
rect 16012 29168 16052 29177
rect 15916 29128 16012 29168
rect 15819 29119 15861 29128
rect 16012 29119 16052 29128
rect 15723 28748 15765 28757
rect 15723 28708 15724 28748
rect 15764 28708 15765 28748
rect 15723 28699 15765 28708
rect 15915 28748 15957 28757
rect 15915 28708 15916 28748
rect 15956 28708 15957 28748
rect 15915 28699 15957 28708
rect 15476 28288 15668 28328
rect 15916 28328 15956 28699
rect 15436 28085 15476 28288
rect 15916 28279 15956 28288
rect 15435 28076 15477 28085
rect 15435 28036 15436 28076
rect 15476 28036 15477 28076
rect 15435 28027 15477 28036
rect 15915 27992 15957 28001
rect 15915 27952 15916 27992
rect 15956 27952 15957 27992
rect 15915 27943 15957 27952
rect 15819 27740 15861 27749
rect 15819 27700 15820 27740
rect 15860 27700 15861 27740
rect 15819 27691 15861 27700
rect 15435 27656 15477 27665
rect 15435 27616 15436 27656
rect 15476 27616 15477 27656
rect 15435 27607 15477 27616
rect 15436 26312 15476 27607
rect 15723 26984 15765 26993
rect 15723 26944 15724 26984
rect 15764 26944 15765 26984
rect 15723 26935 15765 26944
rect 15532 26816 15572 26825
rect 15572 26776 15668 26816
rect 15532 26767 15572 26776
rect 15532 26312 15572 26321
rect 15436 26272 15532 26312
rect 15532 26263 15572 26272
rect 15340 26188 15476 26228
rect 15244 26095 15284 26104
rect 15345 26134 15385 26143
rect 14860 26010 14900 26095
rect 15345 26069 15385 26094
rect 15339 26060 15385 26069
rect 15339 26020 15340 26060
rect 15380 26020 15385 26060
rect 15339 26011 15381 26020
rect 15340 26004 15380 26011
rect 15436 25985 15476 26188
rect 15435 25976 15477 25985
rect 15435 25936 15436 25976
rect 15476 25936 15477 25976
rect 15435 25927 15477 25936
rect 15628 25733 15668 26776
rect 15724 26312 15764 26935
rect 15820 26489 15860 27691
rect 15819 26480 15861 26489
rect 15819 26440 15820 26480
rect 15860 26440 15861 26480
rect 15819 26431 15861 26440
rect 15724 26263 15764 26272
rect 15820 26144 15860 26153
rect 15916 26134 15956 27943
rect 16108 26489 16148 36436
rect 16204 34460 16244 36604
rect 16299 36560 16341 36569
rect 16299 36520 16300 36560
rect 16340 36520 16341 36560
rect 16299 36511 16341 36520
rect 16300 35888 16340 36511
rect 16300 35477 16340 35848
rect 16299 35468 16341 35477
rect 16299 35428 16300 35468
rect 16340 35428 16341 35468
rect 16299 35419 16341 35428
rect 16204 34420 16340 34460
rect 16203 33872 16245 33881
rect 16203 33832 16204 33872
rect 16244 33832 16245 33872
rect 16203 33823 16245 33832
rect 16204 33699 16244 33823
rect 16204 33650 16244 33659
rect 16300 33536 16340 34420
rect 16396 33872 16436 41719
rect 16588 41525 16628 42652
rect 16587 41516 16629 41525
rect 16587 41476 16588 41516
rect 16628 41476 16629 41516
rect 16587 41467 16629 41476
rect 16587 40172 16629 40181
rect 16587 40132 16588 40172
rect 16628 40132 16629 40172
rect 16587 40123 16629 40132
rect 16491 38744 16533 38753
rect 16491 38704 16492 38744
rect 16532 38704 16533 38744
rect 16491 38695 16533 38704
rect 16492 35897 16532 38695
rect 16588 38240 16628 40123
rect 16588 36056 16628 38200
rect 16684 37577 16724 42820
rect 16779 42608 16821 42617
rect 16779 42568 16780 42608
rect 16820 42568 16821 42608
rect 16779 42559 16821 42568
rect 16780 42474 16820 42559
rect 16779 41936 16821 41945
rect 16779 41896 16780 41936
rect 16820 41896 16821 41936
rect 16779 41887 16821 41896
rect 16780 41802 16820 41887
rect 16876 41609 16916 42904
rect 16875 41600 16917 41609
rect 16875 41560 16876 41600
rect 16916 41560 16917 41600
rect 16875 41551 16917 41560
rect 16971 41180 17013 41189
rect 16971 41140 16972 41180
rect 17012 41140 17013 41180
rect 16971 41131 17013 41140
rect 16780 40424 16820 40433
rect 16780 40181 16820 40384
rect 16779 40172 16821 40181
rect 16779 40132 16780 40172
rect 16820 40132 16821 40172
rect 16779 40123 16821 40132
rect 16972 39752 17012 41131
rect 17068 40181 17108 44752
rect 17164 44743 17204 44752
rect 17164 44456 17204 44465
rect 17356 44456 17396 45583
rect 17204 44416 17396 44456
rect 17164 44407 17204 44416
rect 17355 44120 17397 44129
rect 17355 44080 17356 44120
rect 17396 44080 17397 44120
rect 17355 44071 17397 44080
rect 17356 42944 17396 44071
rect 17548 43961 17588 46600
rect 17547 43952 17589 43961
rect 17547 43912 17548 43952
rect 17588 43912 17589 43952
rect 17547 43903 17589 43912
rect 17547 43532 17589 43541
rect 17547 43492 17548 43532
rect 17588 43492 17589 43532
rect 17547 43483 17589 43492
rect 17451 43448 17493 43457
rect 17451 43408 17452 43448
rect 17492 43408 17493 43448
rect 17451 43399 17493 43408
rect 17356 42895 17396 42904
rect 17163 42692 17205 42701
rect 17355 42692 17397 42701
rect 17163 42652 17164 42692
rect 17204 42652 17205 42692
rect 17163 42643 17205 42652
rect 17260 42652 17356 42692
rect 17396 42652 17397 42692
rect 17164 42558 17204 42643
rect 17260 42449 17300 42652
rect 17355 42643 17397 42652
rect 17259 42440 17301 42449
rect 17259 42400 17260 42440
rect 17300 42400 17301 42440
rect 17259 42391 17301 42400
rect 17308 41945 17348 41954
rect 17348 41905 17396 41936
rect 17308 41896 17396 41905
rect 17356 41432 17396 41896
rect 17452 41852 17492 43399
rect 17452 41803 17492 41812
rect 17356 41383 17396 41392
rect 17548 41348 17588 43483
rect 17644 42449 17684 50212
rect 17932 50202 17972 50287
rect 17740 50084 17780 50093
rect 17780 50044 17972 50084
rect 17740 50035 17780 50044
rect 17739 49160 17781 49169
rect 17739 49120 17740 49160
rect 17780 49120 17781 49160
rect 17739 49111 17781 49120
rect 17740 47984 17780 49111
rect 17932 48824 17972 50044
rect 18028 49496 18068 50455
rect 18028 49447 18068 49456
rect 18124 49496 18164 49507
rect 18124 49421 18164 49456
rect 18123 49412 18165 49421
rect 18123 49372 18124 49412
rect 18164 49372 18165 49412
rect 18123 49363 18165 49372
rect 18124 49169 18164 49363
rect 18123 49160 18165 49169
rect 18123 49120 18124 49160
rect 18164 49120 18165 49160
rect 18123 49111 18165 49120
rect 18028 48824 18068 48833
rect 17932 48784 18028 48824
rect 18028 48775 18068 48784
rect 18124 48824 18164 49111
rect 18124 48775 18164 48784
rect 18123 48404 18165 48413
rect 18123 48364 18124 48404
rect 18164 48364 18165 48404
rect 18123 48355 18165 48364
rect 17740 47935 17780 47944
rect 17835 47984 17877 47993
rect 17835 47944 17836 47984
rect 17876 47944 17877 47984
rect 17835 47935 17877 47944
rect 18124 47984 18164 48355
rect 18124 47935 18164 47944
rect 17836 46061 17876 47935
rect 17932 47816 17972 47825
rect 17932 47321 17972 47776
rect 17931 47312 17973 47321
rect 17931 47272 17932 47312
rect 17972 47272 17973 47312
rect 17931 47263 17973 47272
rect 18220 46640 18260 59359
rect 18316 57056 18356 57065
rect 18316 54788 18356 57016
rect 18412 57056 18452 57065
rect 18412 54881 18452 57016
rect 18411 54872 18453 54881
rect 18411 54832 18412 54872
rect 18452 54832 18453 54872
rect 18411 54823 18453 54832
rect 18316 53705 18356 54748
rect 18412 54738 18452 54823
rect 18315 53696 18357 53705
rect 18315 53656 18316 53696
rect 18356 53656 18357 53696
rect 18315 53647 18357 53656
rect 18316 53360 18356 53369
rect 18508 53360 18548 60787
rect 18604 58745 18644 63559
rect 18699 63524 18741 63533
rect 18699 63484 18700 63524
rect 18740 63484 18741 63524
rect 18699 63475 18741 63484
rect 18808 63524 19176 63533
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 18808 63475 19176 63484
rect 18603 58736 18645 58745
rect 18603 58696 18604 58736
rect 18644 58696 18645 58736
rect 18603 58687 18645 58696
rect 18700 58064 18740 63475
rect 18987 63104 19029 63113
rect 18987 63064 18988 63104
rect 19028 63064 19029 63104
rect 18987 63055 19029 63064
rect 18988 62432 19028 63055
rect 19276 63020 19316 64072
rect 19372 63944 19412 63955
rect 19372 63869 19412 63904
rect 19371 63860 19413 63869
rect 19371 63820 19372 63860
rect 19412 63820 19413 63860
rect 19371 63811 19413 63820
rect 19564 63188 19604 65920
rect 19756 65911 19796 65920
rect 19755 65708 19797 65717
rect 19755 65668 19756 65708
rect 19796 65668 19797 65708
rect 19755 65659 19797 65668
rect 19659 64448 19701 64457
rect 19659 64408 19660 64448
rect 19700 64408 19701 64448
rect 19659 64399 19701 64408
rect 19516 63148 19604 63188
rect 19516 63146 19556 63148
rect 19516 63097 19556 63106
rect 19660 63104 19700 64399
rect 19756 64280 19796 65659
rect 19852 64877 19892 67171
rect 20524 66809 20564 69103
rect 20619 68144 20661 68153
rect 20619 68104 20620 68144
rect 20660 68104 20661 68144
rect 20619 68095 20661 68104
rect 20523 66800 20565 66809
rect 20523 66760 20524 66800
rect 20564 66760 20565 66800
rect 20523 66751 20565 66760
rect 20523 66128 20565 66137
rect 20523 66088 20524 66128
rect 20564 66088 20565 66128
rect 20523 66079 20565 66088
rect 20048 65792 20416 65801
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20048 65743 20416 65752
rect 20524 64961 20564 66079
rect 20620 65045 20660 68095
rect 20716 68060 20756 72472
rect 21099 72472 21100 72512
rect 21140 72472 21141 72512
rect 21099 72463 21141 72472
rect 20716 68020 20852 68060
rect 20715 67136 20757 67145
rect 20715 67096 20716 67136
rect 20756 67096 20757 67136
rect 20715 67087 20757 67096
rect 20619 65036 20661 65045
rect 20619 64996 20620 65036
rect 20660 64996 20661 65036
rect 20619 64987 20661 64996
rect 20523 64952 20565 64961
rect 20523 64912 20524 64952
rect 20564 64912 20565 64952
rect 20523 64903 20565 64912
rect 19851 64868 19893 64877
rect 19851 64828 19852 64868
rect 19892 64828 19893 64868
rect 19851 64819 19893 64828
rect 19852 64700 19892 64711
rect 19852 64625 19892 64660
rect 19851 64616 19893 64625
rect 19851 64576 19852 64616
rect 19892 64576 19893 64616
rect 19851 64567 19893 64576
rect 20044 64457 20084 64542
rect 20043 64448 20085 64457
rect 20043 64408 20044 64448
rect 20084 64408 20085 64448
rect 20043 64399 20085 64408
rect 20619 64448 20661 64457
rect 20619 64408 20620 64448
rect 20660 64408 20661 64448
rect 20619 64399 20661 64408
rect 20048 64280 20416 64289
rect 19756 64240 19892 64280
rect 19756 63860 19796 63869
rect 19756 63365 19796 63820
rect 19755 63356 19797 63365
rect 19755 63316 19756 63356
rect 19796 63316 19797 63356
rect 19755 63307 19797 63316
rect 19852 63188 19892 64240
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20048 64231 20416 64240
rect 19947 63692 19989 63701
rect 19947 63652 19948 63692
rect 19988 63652 19989 63692
rect 19947 63643 19989 63652
rect 19948 63558 19988 63643
rect 19852 63139 19892 63148
rect 19660 63064 19796 63104
rect 19276 62980 19508 63020
rect 18988 62383 19028 62392
rect 19468 62427 19508 62980
rect 19660 62936 19700 62945
rect 19468 62378 19508 62387
rect 19564 62896 19660 62936
rect 18808 62012 19176 62021
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 18808 61963 19176 61972
rect 19372 61592 19412 61603
rect 19564 61601 19604 62896
rect 19660 62887 19700 62896
rect 19659 62684 19701 62693
rect 19659 62644 19660 62684
rect 19700 62644 19701 62684
rect 19659 62635 19701 62644
rect 19660 62600 19700 62635
rect 19660 62549 19700 62560
rect 19756 62432 19796 63064
rect 20044 62936 20084 62945
rect 19660 62392 19796 62432
rect 19948 62896 20044 62936
rect 19372 61517 19412 61552
rect 19563 61592 19605 61601
rect 19563 61552 19564 61592
rect 19604 61552 19605 61592
rect 19563 61543 19605 61552
rect 19371 61508 19413 61517
rect 19371 61468 19372 61508
rect 19412 61468 19413 61508
rect 19660 61508 19700 62392
rect 19851 62348 19893 62357
rect 19851 62308 19852 62348
rect 19892 62308 19893 62348
rect 19851 62299 19893 62308
rect 19852 62214 19892 62299
rect 19756 61685 19796 61770
rect 19755 61676 19797 61685
rect 19755 61636 19756 61676
rect 19796 61636 19797 61676
rect 19755 61627 19797 61636
rect 19948 61592 19988 62896
rect 20044 62887 20084 62896
rect 20048 62768 20416 62777
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20048 62719 20416 62728
rect 20523 62768 20565 62777
rect 20523 62728 20524 62768
rect 20564 62728 20565 62768
rect 20523 62719 20565 62728
rect 19852 61552 19988 61592
rect 20044 62180 20084 62189
rect 19660 61468 19796 61508
rect 19371 61459 19413 61468
rect 19564 61424 19604 61433
rect 19604 61384 19700 61424
rect 19564 61375 19604 61384
rect 19275 60920 19317 60929
rect 19372 60920 19412 60929
rect 19275 60880 19276 60920
rect 19316 60880 19372 60920
rect 19275 60871 19317 60880
rect 19372 60871 19412 60880
rect 18808 60500 19176 60509
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 18808 60451 19176 60460
rect 18891 60332 18933 60341
rect 18891 60292 18892 60332
rect 18932 60292 18933 60332
rect 18891 60283 18933 60292
rect 18892 60080 18932 60283
rect 18892 59408 18932 60040
rect 18892 59359 18932 59368
rect 18808 58988 19176 58997
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 18808 58939 19176 58948
rect 19276 58568 19316 60871
rect 19564 60668 19604 60677
rect 19468 60628 19564 60668
rect 19468 60164 19508 60628
rect 19564 60619 19604 60628
rect 19420 60124 19508 60164
rect 19420 60122 19460 60124
rect 19420 60073 19460 60082
rect 19563 59912 19605 59921
rect 19563 59872 19564 59912
rect 19604 59872 19605 59912
rect 19563 59863 19605 59872
rect 19564 59778 19604 59863
rect 19660 59660 19700 61384
rect 19756 61097 19796 61468
rect 19755 61088 19797 61097
rect 19755 61048 19756 61088
rect 19796 61048 19797 61088
rect 19755 61039 19797 61048
rect 19756 60164 19796 60173
rect 19756 59669 19796 60124
rect 19468 59620 19700 59660
rect 19755 59660 19797 59669
rect 19755 59620 19756 59660
rect 19796 59620 19797 59660
rect 19468 59408 19508 59620
rect 19755 59611 19797 59620
rect 19563 59492 19605 59501
rect 19563 59452 19564 59492
rect 19604 59452 19605 59492
rect 19563 59443 19605 59452
rect 19420 59398 19508 59408
rect 19460 59368 19508 59398
rect 19564 59358 19604 59443
rect 19420 59349 19460 59358
rect 19756 59333 19796 59418
rect 19755 59324 19797 59333
rect 19755 59284 19756 59324
rect 19796 59284 19797 59324
rect 19755 59275 19797 59284
rect 19755 59156 19797 59165
rect 19755 59116 19756 59156
rect 19796 59116 19797 59156
rect 19755 59107 19797 59116
rect 19659 58652 19701 58661
rect 19659 58612 19660 58652
rect 19700 58612 19701 58652
rect 19659 58603 19701 58612
rect 18700 58024 18932 58064
rect 18796 57896 18836 57905
rect 18796 57812 18836 57856
rect 18604 57772 18836 57812
rect 18604 55805 18644 57772
rect 18892 57728 18932 58024
rect 19276 57989 19316 58528
rect 19660 58518 19700 58603
rect 19468 58400 19508 58409
rect 19372 58360 19468 58400
rect 19275 57980 19317 57989
rect 19275 57940 19276 57980
rect 19316 57940 19317 57980
rect 19275 57931 19317 57940
rect 19083 57896 19125 57905
rect 19083 57856 19084 57896
rect 19124 57856 19125 57896
rect 19083 57847 19125 57856
rect 19084 57762 19124 57847
rect 18700 57688 18932 57728
rect 18700 56225 18740 57688
rect 18808 57476 19176 57485
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 18808 57427 19176 57436
rect 19372 57070 19412 58360
rect 19468 58351 19508 58360
rect 19564 57644 19604 57653
rect 18892 57056 18932 57065
rect 18932 57016 19316 57056
rect 19372 57021 19412 57030
rect 19468 57604 19564 57644
rect 18892 57007 18932 57016
rect 18699 56216 18741 56225
rect 18699 56176 18700 56216
rect 18740 56176 18741 56216
rect 18699 56167 18741 56176
rect 18808 55964 19176 55973
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 18808 55915 19176 55924
rect 18603 55796 18645 55805
rect 18603 55756 18604 55796
rect 18644 55756 18645 55796
rect 18603 55747 18645 55756
rect 18699 55628 18741 55637
rect 18699 55588 18700 55628
rect 18740 55588 18741 55628
rect 18699 55579 18741 55588
rect 18700 55544 18740 55579
rect 18700 55493 18740 55504
rect 18892 55376 18932 55385
rect 18356 53320 18548 53360
rect 18700 55336 18892 55376
rect 18316 51008 18356 53320
rect 18700 52772 18740 55336
rect 18892 55327 18932 55336
rect 19276 55133 19316 57016
rect 19372 56393 19412 56478
rect 19371 56384 19413 56393
rect 19371 56344 19372 56384
rect 19412 56344 19413 56384
rect 19371 56335 19413 56344
rect 19371 56216 19413 56225
rect 19371 56176 19372 56216
rect 19412 56176 19413 56216
rect 19371 56167 19413 56176
rect 19372 55628 19412 56167
rect 19372 55579 19412 55588
rect 19371 55460 19413 55469
rect 19371 55420 19372 55460
rect 19412 55420 19413 55460
rect 19371 55411 19413 55420
rect 18891 55124 18933 55133
rect 18891 55084 18892 55124
rect 18932 55084 18933 55124
rect 18891 55075 18933 55084
rect 19275 55124 19317 55133
rect 19275 55084 19276 55124
rect 19316 55084 19317 55124
rect 19275 55075 19317 55084
rect 18892 54872 18932 55075
rect 19275 54956 19317 54965
rect 19275 54916 19276 54956
rect 19316 54916 19317 54956
rect 19275 54907 19317 54916
rect 18892 54713 18932 54832
rect 18891 54704 18933 54713
rect 18891 54664 18892 54704
rect 18932 54664 18933 54704
rect 18891 54655 18933 54664
rect 18808 54452 19176 54461
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 18808 54403 19176 54412
rect 19276 54284 19316 54907
rect 19372 54867 19412 55411
rect 19372 54818 19412 54827
rect 19180 54244 19316 54284
rect 19083 54032 19125 54041
rect 19083 53992 19084 54032
rect 19124 53992 19125 54032
rect 19083 53983 19125 53992
rect 18891 53864 18933 53873
rect 18891 53824 18892 53864
rect 18932 53824 18933 53864
rect 18891 53815 18933 53824
rect 18892 53117 18932 53815
rect 19084 53369 19124 53983
rect 19180 53537 19220 54244
rect 19276 54041 19316 54126
rect 19275 54032 19317 54041
rect 19468 54032 19508 57604
rect 19564 57595 19604 57604
rect 19756 57560 19796 59107
rect 19852 58745 19892 61552
rect 20044 61517 20084 62140
rect 20524 61937 20564 62719
rect 20523 61928 20565 61937
rect 20523 61888 20524 61928
rect 20564 61888 20565 61928
rect 20523 61879 20565 61888
rect 20043 61508 20085 61517
rect 20043 61468 20044 61508
rect 20084 61468 20085 61508
rect 20043 61459 20085 61468
rect 19947 61424 19989 61433
rect 19947 61384 19948 61424
rect 19988 61384 19989 61424
rect 19947 61375 19989 61384
rect 19948 61290 19988 61375
rect 20048 61256 20416 61265
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20048 61207 20416 61216
rect 20043 60836 20085 60845
rect 20043 60796 20044 60836
rect 20084 60796 20085 60836
rect 20043 60787 20085 60796
rect 20044 60702 20084 60787
rect 20235 60668 20277 60677
rect 20235 60628 20236 60668
rect 20276 60628 20277 60668
rect 20235 60619 20277 60628
rect 20236 60534 20276 60619
rect 19948 59912 19988 59921
rect 19948 59324 19988 59872
rect 20048 59744 20416 59753
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20048 59695 20416 59704
rect 19948 59284 20084 59324
rect 19947 59156 19989 59165
rect 19947 59116 19948 59156
rect 19988 59116 19989 59156
rect 19947 59107 19989 59116
rect 19948 59022 19988 59107
rect 20044 58820 20084 59284
rect 19948 58780 20084 58820
rect 19851 58736 19893 58745
rect 19851 58696 19852 58736
rect 19892 58696 19893 58736
rect 19851 58687 19893 58696
rect 19660 57520 19796 57560
rect 19852 58400 19892 58409
rect 19563 56888 19605 56897
rect 19563 56848 19564 56888
rect 19604 56848 19605 56888
rect 19563 56839 19605 56848
rect 19564 56754 19604 56839
rect 19564 56132 19604 56141
rect 19564 55553 19604 56092
rect 19660 56057 19700 57520
rect 19755 57308 19797 57317
rect 19755 57268 19756 57308
rect 19796 57268 19797 57308
rect 19755 57259 19797 57268
rect 19756 57140 19796 57259
rect 19756 57091 19796 57100
rect 19755 56972 19797 56981
rect 19755 56932 19756 56972
rect 19796 56932 19797 56972
rect 19755 56923 19797 56932
rect 19756 56477 19796 56923
rect 19852 56813 19892 58360
rect 19948 57065 19988 58780
rect 20043 58652 20085 58661
rect 20043 58612 20044 58652
rect 20084 58612 20085 58652
rect 20043 58603 20085 58612
rect 20044 58518 20084 58603
rect 20236 58400 20276 58409
rect 20276 58360 20564 58400
rect 20236 58351 20276 58360
rect 20048 58232 20416 58241
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20048 58183 20416 58192
rect 19947 57056 19989 57065
rect 19947 57016 19948 57056
rect 19988 57016 19989 57056
rect 19947 57007 19989 57016
rect 19948 56888 19988 56897
rect 19851 56804 19893 56813
rect 19851 56764 19852 56804
rect 19892 56764 19893 56804
rect 19851 56755 19893 56764
rect 19755 56468 19797 56477
rect 19755 56428 19756 56468
rect 19796 56428 19797 56468
rect 19755 56419 19797 56428
rect 19756 56300 19796 56309
rect 19948 56300 19988 56848
rect 20048 56720 20416 56729
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20048 56671 20416 56680
rect 19948 56260 20084 56300
rect 19756 56141 19796 56260
rect 19755 56132 19797 56141
rect 19755 56092 19756 56132
rect 19796 56092 19797 56132
rect 19755 56083 19797 56092
rect 19947 56132 19989 56141
rect 19947 56092 19948 56132
rect 19988 56092 19989 56132
rect 19947 56083 19989 56092
rect 19659 56048 19701 56057
rect 19659 56008 19660 56048
rect 19700 56008 19701 56048
rect 19659 55999 19701 56008
rect 19948 55998 19988 56083
rect 19755 55796 19797 55805
rect 19755 55756 19756 55796
rect 19796 55756 19797 55796
rect 19755 55747 19797 55756
rect 19756 55628 19796 55747
rect 19756 55579 19796 55588
rect 20044 55553 20084 56260
rect 20524 55721 20564 58360
rect 20523 55712 20565 55721
rect 20523 55672 20524 55712
rect 20564 55672 20565 55712
rect 20523 55663 20565 55672
rect 19563 55544 19605 55553
rect 19563 55504 19564 55544
rect 19604 55504 19605 55544
rect 19563 55495 19605 55504
rect 20043 55544 20085 55553
rect 20043 55504 20044 55544
rect 20084 55504 20085 55544
rect 20043 55495 20085 55504
rect 19564 55376 19604 55385
rect 19948 55376 19988 55385
rect 19604 55336 19700 55376
rect 19564 55327 19604 55336
rect 19563 54956 19605 54965
rect 19563 54916 19564 54956
rect 19604 54916 19605 54956
rect 19563 54907 19605 54916
rect 19564 54822 19604 54907
rect 19660 54620 19700 55336
rect 19756 54797 19796 54882
rect 19948 54797 19988 55336
rect 20048 55208 20416 55217
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20048 55159 20416 55168
rect 19755 54788 19797 54797
rect 19755 54748 19756 54788
rect 19796 54748 19797 54788
rect 19755 54739 19797 54748
rect 19947 54788 19989 54797
rect 19947 54748 19948 54788
rect 19988 54748 19989 54788
rect 19947 54739 19989 54748
rect 19948 54620 19988 54629
rect 19660 54580 19796 54620
rect 19563 54200 19605 54209
rect 19563 54160 19564 54200
rect 19604 54160 19605 54200
rect 19563 54151 19605 54160
rect 19275 53992 19276 54032
rect 19316 53992 19317 54032
rect 19275 53983 19317 53992
rect 19372 53992 19508 54032
rect 19372 53864 19412 53992
rect 19564 53948 19604 54151
rect 19660 54125 19700 54210
rect 19659 54116 19701 54125
rect 19659 54076 19660 54116
rect 19700 54076 19701 54116
rect 19659 54067 19701 54076
rect 19564 53908 19700 53948
rect 19276 53824 19412 53864
rect 19468 53864 19508 53873
rect 19179 53528 19221 53537
rect 19179 53488 19180 53528
rect 19220 53488 19221 53528
rect 19179 53479 19221 53488
rect 19083 53360 19125 53369
rect 19083 53320 19084 53360
rect 19124 53320 19125 53360
rect 19083 53311 19125 53320
rect 18891 53108 18933 53117
rect 18891 53068 18892 53108
rect 18932 53068 18933 53108
rect 18891 53059 18933 53068
rect 18808 52940 19176 52949
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 18808 52891 19176 52900
rect 18700 52732 18932 52772
rect 18508 52520 18548 52529
rect 18412 52480 18508 52520
rect 18412 51857 18452 52480
rect 18508 52471 18548 52480
rect 18411 51848 18453 51857
rect 18411 51808 18412 51848
rect 18452 51808 18453 51848
rect 18411 51799 18453 51808
rect 18892 51843 18932 52732
rect 18987 52688 19029 52697
rect 18987 52648 18988 52688
rect 19028 52648 19029 52688
rect 18987 52639 19029 52648
rect 18988 52534 19028 52639
rect 18988 52485 19028 52494
rect 19179 52352 19221 52361
rect 19179 52312 19180 52352
rect 19220 52312 19221 52352
rect 19179 52303 19221 52312
rect 19180 52218 19220 52303
rect 19083 51932 19125 51941
rect 19083 51892 19084 51932
rect 19124 51892 19125 51932
rect 19083 51883 19125 51892
rect 18412 51714 18452 51799
rect 18892 51794 18932 51803
rect 19084 51798 19124 51883
rect 18808 51428 19176 51437
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 18808 51379 19176 51388
rect 18316 50849 18356 50968
rect 18315 50840 18357 50849
rect 18315 50800 18316 50840
rect 18356 50800 18357 50840
rect 18315 50791 18357 50800
rect 19179 50336 19221 50345
rect 19179 50296 19180 50336
rect 19220 50296 19221 50336
rect 19179 50287 19221 50296
rect 19180 50202 19220 50287
rect 19276 50252 19316 53824
rect 19468 52697 19508 53824
rect 19563 53360 19605 53369
rect 19563 53320 19564 53360
rect 19604 53320 19605 53360
rect 19563 53311 19605 53320
rect 19564 53226 19604 53311
rect 19660 52949 19700 53908
rect 19756 53789 19796 54580
rect 19852 53864 19892 53873
rect 19755 53780 19797 53789
rect 19755 53740 19756 53780
rect 19796 53740 19797 53780
rect 19755 53731 19797 53740
rect 19756 53108 19796 53117
rect 19659 52940 19701 52949
rect 19659 52900 19660 52940
rect 19700 52900 19701 52940
rect 19659 52891 19701 52900
rect 19756 52772 19796 53068
rect 19852 53033 19892 53824
rect 19948 53453 19988 54580
rect 20044 54116 20084 54125
rect 20044 53873 20084 54076
rect 20235 54032 20277 54041
rect 20235 53992 20236 54032
rect 20276 53992 20277 54032
rect 20235 53983 20277 53992
rect 20043 53864 20085 53873
rect 20043 53824 20044 53864
rect 20084 53824 20085 53864
rect 20043 53815 20085 53824
rect 20236 53864 20276 53983
rect 20236 53815 20276 53824
rect 20048 53696 20416 53705
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20048 53647 20416 53656
rect 19947 53444 19989 53453
rect 19947 53404 19948 53444
rect 19988 53404 19989 53444
rect 19947 53395 19989 53404
rect 19947 53276 19989 53285
rect 19947 53236 19948 53276
rect 19988 53236 19989 53276
rect 19947 53227 19989 53236
rect 19948 53142 19988 53227
rect 20140 53108 20180 53117
rect 19851 53024 19893 53033
rect 19851 52984 19852 53024
rect 19892 52984 19893 53024
rect 19851 52975 19893 52984
rect 19756 52732 19892 52772
rect 19467 52688 19509 52697
rect 19467 52648 19468 52688
rect 19508 52648 19509 52688
rect 19467 52639 19509 52648
rect 19372 52604 19412 52613
rect 19372 52193 19412 52564
rect 19755 52604 19797 52613
rect 19755 52564 19756 52604
rect 19796 52564 19797 52604
rect 19755 52555 19797 52564
rect 19756 52470 19796 52555
rect 19564 52352 19604 52361
rect 19371 52184 19413 52193
rect 19371 52144 19372 52184
rect 19412 52144 19413 52184
rect 19371 52135 19413 52144
rect 19564 52025 19604 52312
rect 19563 52016 19605 52025
rect 19563 51976 19564 52016
rect 19604 51976 19605 52016
rect 19563 51967 19605 51976
rect 19372 51764 19412 51773
rect 19755 51764 19797 51773
rect 19412 51724 19508 51764
rect 19372 51715 19412 51724
rect 19372 50252 19412 50261
rect 19276 50212 19372 50252
rect 19372 50203 19412 50212
rect 18603 50084 18645 50093
rect 19468 50084 19508 51724
rect 19755 51724 19756 51764
rect 19796 51724 19797 51764
rect 19755 51715 19797 51724
rect 19563 51680 19605 51689
rect 19563 51640 19564 51680
rect 19604 51640 19605 51680
rect 19563 51631 19605 51640
rect 19564 51546 19604 51631
rect 19756 51630 19796 51715
rect 19563 51008 19605 51017
rect 19563 50968 19564 51008
rect 19604 50968 19605 51008
rect 19563 50959 19605 50968
rect 19564 50874 19604 50959
rect 19756 50840 19796 50849
rect 19563 50336 19605 50345
rect 19563 50296 19564 50336
rect 19604 50296 19605 50336
rect 19563 50287 19605 50296
rect 19564 50168 19604 50287
rect 19564 50119 19604 50128
rect 18603 50044 18604 50084
rect 18644 50044 18645 50084
rect 18603 50035 18645 50044
rect 19372 50044 19508 50084
rect 18604 49580 18644 50035
rect 18808 49916 19176 49925
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 18808 49867 19176 49876
rect 18508 49496 18548 49507
rect 18508 49421 18548 49456
rect 18507 49412 18549 49421
rect 18507 49372 18508 49412
rect 18548 49372 18549 49412
rect 18507 49363 18549 49372
rect 18411 49160 18453 49169
rect 18411 49120 18412 49160
rect 18452 49120 18453 49160
rect 18411 49111 18453 49120
rect 18315 48992 18357 49001
rect 18315 48952 18316 48992
rect 18356 48952 18357 48992
rect 18315 48943 18357 48952
rect 18316 47573 18356 48943
rect 18315 47564 18357 47573
rect 18315 47524 18316 47564
rect 18356 47524 18357 47564
rect 18315 47515 18357 47524
rect 18315 47312 18357 47321
rect 18315 47272 18316 47312
rect 18356 47272 18357 47312
rect 18315 47263 18357 47272
rect 18412 47312 18452 49111
rect 18508 48824 18548 49363
rect 18508 47321 18548 48784
rect 18604 48824 18644 49540
rect 19083 49496 19125 49505
rect 19083 49456 19084 49496
rect 19124 49456 19125 49496
rect 19083 49447 19125 49456
rect 18604 48775 18644 48784
rect 19084 48824 19124 49447
rect 19084 48775 19124 48784
rect 18808 48404 19176 48413
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 18808 48355 19176 48364
rect 19275 48236 19317 48245
rect 19275 48196 19276 48236
rect 19316 48196 19317 48236
rect 19275 48187 19317 48196
rect 18891 47480 18933 47489
rect 18891 47440 18892 47480
rect 18932 47440 18933 47480
rect 18891 47431 18933 47440
rect 18316 47178 18356 47263
rect 18028 46600 18260 46640
rect 18412 46640 18452 47272
rect 18507 47312 18549 47321
rect 18795 47312 18837 47321
rect 18507 47272 18508 47312
rect 18548 47272 18549 47312
rect 18507 47263 18549 47272
rect 18700 47272 18796 47312
rect 18836 47272 18837 47312
rect 18700 46724 18740 47272
rect 18795 47263 18837 47272
rect 18892 47312 18932 47431
rect 18796 47178 18836 47263
rect 18892 47069 18932 47272
rect 18891 47060 18933 47069
rect 18891 47020 18892 47060
rect 18932 47020 18933 47060
rect 18891 47011 18933 47020
rect 18808 46892 19176 46901
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 18808 46843 19176 46852
rect 18987 46724 19029 46733
rect 18700 46684 18932 46724
rect 18412 46600 18548 46640
rect 17835 46052 17877 46061
rect 17835 46012 17836 46052
rect 17876 46012 17877 46052
rect 17835 46003 17877 46012
rect 17931 44708 17973 44717
rect 17931 44668 17932 44708
rect 17972 44668 17973 44708
rect 17931 44659 17973 44668
rect 17932 44456 17972 44659
rect 17932 44407 17972 44416
rect 17740 44204 17780 44213
rect 17780 44164 17876 44204
rect 17740 44155 17780 44164
rect 17739 43700 17781 43709
rect 17739 43660 17740 43700
rect 17780 43660 17781 43700
rect 17739 43651 17781 43660
rect 17740 43566 17780 43651
rect 17740 42692 17780 42701
rect 17643 42440 17685 42449
rect 17643 42400 17644 42440
rect 17684 42400 17685 42440
rect 17643 42391 17685 42400
rect 17644 42020 17684 42029
rect 17644 41357 17684 41980
rect 17740 41525 17780 42652
rect 17836 42356 17876 44164
rect 18028 44036 18068 46600
rect 18412 46472 18452 46481
rect 18412 45977 18452 46432
rect 18508 46472 18548 46600
rect 18892 46556 18932 46684
rect 18987 46684 18988 46724
rect 19028 46684 19029 46724
rect 18987 46675 19029 46684
rect 18892 46507 18932 46516
rect 18988 46556 19028 46675
rect 18988 46507 19028 46516
rect 18508 46423 18548 46432
rect 18411 45968 18453 45977
rect 18411 45928 18412 45968
rect 18452 45928 18453 45968
rect 18411 45919 18453 45928
rect 18795 45968 18837 45977
rect 18892 45968 18932 45977
rect 18795 45928 18796 45968
rect 18836 45928 18892 45968
rect 18795 45919 18837 45928
rect 18892 45919 18932 45928
rect 18699 45800 18741 45809
rect 18699 45760 18700 45800
rect 18740 45760 18741 45800
rect 18699 45751 18741 45760
rect 18700 45473 18740 45751
rect 18699 45464 18741 45473
rect 18699 45424 18700 45464
rect 18740 45424 18741 45464
rect 18699 45415 18741 45424
rect 18808 45380 19176 45389
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 18808 45331 19176 45340
rect 18315 45212 18357 45221
rect 18315 45172 18316 45212
rect 18356 45172 18357 45212
rect 18315 45163 18357 45172
rect 18316 45078 18356 45163
rect 18124 45044 18164 45053
rect 18124 44708 18164 45004
rect 18507 44960 18549 44969
rect 18507 44920 18508 44960
rect 18548 44920 18549 44960
rect 18507 44911 18549 44920
rect 18124 44668 18452 44708
rect 18315 44540 18357 44549
rect 18315 44500 18316 44540
rect 18356 44500 18357 44540
rect 18315 44491 18357 44500
rect 18123 44456 18165 44465
rect 18123 44416 18124 44456
rect 18164 44416 18165 44456
rect 18123 44407 18165 44416
rect 18316 44456 18356 44491
rect 18124 44204 18164 44407
rect 18316 44405 18356 44416
rect 18124 44155 18164 44164
rect 18028 43996 18356 44036
rect 17932 43532 17972 43541
rect 17932 42785 17972 43492
rect 18124 43280 18164 43289
rect 18124 42953 18164 43240
rect 18123 42944 18165 42953
rect 18123 42904 18124 42944
rect 18164 42904 18165 42944
rect 18123 42895 18165 42904
rect 17931 42776 17973 42785
rect 17931 42736 17932 42776
rect 17972 42736 17973 42776
rect 17931 42727 17973 42736
rect 18124 42692 18164 42701
rect 17931 42608 17973 42617
rect 17931 42568 17932 42608
rect 17972 42568 17973 42608
rect 17931 42559 17973 42568
rect 17932 42474 17972 42559
rect 17836 42316 17972 42356
rect 17835 42188 17877 42197
rect 17835 42148 17836 42188
rect 17876 42148 17877 42188
rect 17835 42139 17877 42148
rect 17836 42054 17876 42139
rect 17835 41600 17877 41609
rect 17835 41560 17836 41600
rect 17876 41560 17877 41600
rect 17835 41551 17877 41560
rect 17739 41516 17781 41525
rect 17739 41476 17740 41516
rect 17780 41476 17781 41516
rect 17739 41467 17781 41476
rect 17452 41308 17588 41348
rect 17643 41348 17685 41357
rect 17643 41308 17644 41348
rect 17684 41308 17685 41348
rect 17164 41264 17204 41275
rect 17164 41189 17204 41224
rect 17163 41180 17205 41189
rect 17163 41140 17164 41180
rect 17204 41140 17205 41180
rect 17163 41131 17205 41140
rect 17452 41096 17492 41308
rect 17643 41299 17685 41308
rect 17356 41056 17492 41096
rect 17548 41180 17588 41189
rect 17260 40429 17300 40438
rect 17067 40172 17109 40181
rect 17067 40132 17068 40172
rect 17108 40132 17109 40172
rect 17067 40123 17109 40132
rect 17164 39920 17204 39929
rect 17260 39920 17300 40389
rect 17204 39880 17300 39920
rect 17164 39871 17204 39880
rect 16972 38921 17012 39712
rect 16971 38912 17013 38921
rect 16971 38872 16972 38912
rect 17012 38872 17013 38912
rect 16971 38863 17013 38872
rect 17260 38324 17300 38333
rect 16780 38284 17260 38324
rect 16683 37568 16725 37577
rect 16683 37528 16684 37568
rect 16724 37528 16725 37568
rect 16683 37519 16725 37528
rect 16683 36812 16725 36821
rect 16683 36772 16684 36812
rect 16724 36772 16725 36812
rect 16683 36763 16725 36772
rect 16684 36728 16724 36763
rect 16684 36677 16724 36688
rect 16588 36016 16724 36056
rect 16492 35857 16628 35897
rect 16492 35729 16532 35814
rect 16491 35720 16533 35729
rect 16491 35680 16492 35720
rect 16532 35680 16533 35720
rect 16491 35671 16533 35680
rect 16588 35552 16628 35857
rect 16396 33823 16436 33832
rect 16492 35512 16628 35552
rect 16204 33496 16340 33536
rect 16204 27833 16244 33496
rect 16348 32873 16388 32882
rect 16388 32833 16436 32864
rect 16348 32824 16436 32833
rect 16396 32360 16436 32824
rect 16492 32780 16532 35512
rect 16587 33704 16629 33713
rect 16587 33664 16588 33704
rect 16628 33664 16629 33704
rect 16587 33655 16629 33664
rect 16588 33377 16628 33655
rect 16684 33461 16724 36016
rect 16683 33452 16725 33461
rect 16683 33412 16684 33452
rect 16724 33412 16725 33452
rect 16683 33403 16725 33412
rect 16587 33368 16629 33377
rect 16587 33328 16588 33368
rect 16628 33328 16629 33368
rect 16587 33319 16629 33328
rect 16492 32731 16532 32740
rect 16492 32360 16532 32369
rect 16396 32320 16492 32360
rect 16492 32311 16532 32320
rect 16300 32192 16340 32203
rect 16300 32117 16340 32152
rect 16299 32108 16341 32117
rect 16299 32068 16300 32108
rect 16340 32068 16436 32108
rect 16299 32059 16341 32068
rect 16300 31357 16340 31366
rect 16300 31025 16340 31317
rect 16299 31016 16341 31025
rect 16299 30976 16300 31016
rect 16340 30976 16341 31016
rect 16299 30967 16341 30976
rect 16396 30680 16436 32068
rect 16588 31352 16628 33319
rect 16684 31352 16724 31361
rect 16588 31312 16684 31352
rect 16684 31303 16724 31312
rect 16492 31184 16532 31193
rect 16492 30857 16532 31144
rect 16683 31016 16725 31025
rect 16683 30976 16684 31016
rect 16724 30976 16725 31016
rect 16683 30967 16725 30976
rect 16491 30848 16533 30857
rect 16491 30808 16492 30848
rect 16532 30808 16533 30848
rect 16491 30799 16533 30808
rect 16684 30848 16724 30967
rect 16684 30799 16724 30808
rect 16491 30680 16533 30689
rect 16396 30640 16492 30680
rect 16532 30640 16533 30680
rect 16491 30631 16533 30640
rect 16492 30546 16532 30631
rect 16395 30512 16437 30521
rect 16395 30472 16396 30512
rect 16436 30472 16437 30512
rect 16395 30463 16437 30472
rect 16396 29000 16436 30463
rect 16780 30185 16820 38284
rect 17260 38275 17300 38284
rect 17356 38240 17396 41056
rect 17451 40676 17493 40685
rect 17451 40636 17452 40676
rect 17492 40636 17493 40676
rect 17451 40627 17493 40636
rect 17452 40340 17492 40627
rect 17452 40291 17492 40300
rect 17451 40172 17493 40181
rect 17451 40132 17452 40172
rect 17492 40132 17493 40172
rect 17451 40123 17493 40132
rect 17452 38744 17492 40123
rect 17548 39173 17588 41140
rect 17739 41012 17781 41021
rect 17739 40972 17740 41012
rect 17780 40972 17781 41012
rect 17739 40963 17781 40972
rect 17740 40878 17780 40963
rect 17836 40769 17876 41551
rect 17932 41432 17972 42316
rect 18124 42113 18164 42652
rect 18316 42608 18356 43996
rect 18316 42559 18356 42568
rect 18219 42356 18261 42365
rect 18219 42316 18220 42356
rect 18260 42316 18261 42356
rect 18219 42307 18261 42316
rect 18220 42188 18260 42307
rect 18412 42188 18452 44668
rect 18508 44288 18548 44911
rect 18604 44288 18644 44297
rect 18508 44248 18604 44288
rect 18604 44239 18644 44248
rect 18808 43868 19176 43877
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 18808 43819 19176 43828
rect 18795 43700 18837 43709
rect 19276 43700 19316 48187
rect 19372 47993 19412 50044
rect 19756 49580 19796 50800
rect 19612 49540 19796 49580
rect 19612 49538 19652 49540
rect 19612 49489 19652 49498
rect 19852 49496 19892 52732
rect 20140 52697 20180 53068
rect 20139 52688 20181 52697
rect 20139 52648 20140 52688
rect 20180 52648 20181 52688
rect 20139 52639 20181 52648
rect 19947 52352 19989 52361
rect 19947 52312 19948 52352
rect 19988 52312 19989 52352
rect 19947 52303 19989 52312
rect 19948 52218 19988 52303
rect 20048 52184 20416 52193
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20048 52135 20416 52144
rect 19948 51680 19988 51689
rect 20139 51680 20181 51689
rect 19988 51640 20140 51680
rect 20180 51640 20181 51680
rect 19948 51631 19988 51640
rect 20139 51631 20181 51640
rect 20139 51008 20181 51017
rect 20139 50968 20140 51008
rect 20180 50968 20181 51008
rect 20139 50959 20181 50968
rect 20140 50882 20180 50959
rect 20140 50833 20180 50842
rect 20048 50672 20416 50681
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20048 50623 20416 50632
rect 19947 50588 19989 50597
rect 19947 50548 19948 50588
rect 19988 50548 19989 50588
rect 19947 50539 19989 50548
rect 19948 50168 19988 50539
rect 19948 50119 19988 50128
rect 19756 49456 19892 49496
rect 19756 49412 19796 49456
rect 19660 49372 19796 49412
rect 19660 48824 19700 49372
rect 19756 49286 19796 49295
rect 19756 49076 19796 49246
rect 20048 49160 20416 49169
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20048 49111 20416 49120
rect 19756 49036 19988 49076
rect 19612 48814 19700 48824
rect 19652 48784 19700 48814
rect 19756 48908 19796 48917
rect 19612 48765 19652 48774
rect 19371 47984 19413 47993
rect 19371 47944 19372 47984
rect 19412 47944 19413 47984
rect 19371 47935 19413 47944
rect 19372 47850 19412 47935
rect 19371 47564 19413 47573
rect 19371 47524 19372 47564
rect 19412 47524 19413 47564
rect 19371 47515 19413 47524
rect 19372 47312 19412 47515
rect 19563 47312 19605 47321
rect 19412 47272 19508 47312
rect 19372 47263 19412 47272
rect 19468 46472 19508 47272
rect 19563 47272 19564 47312
rect 19604 47272 19605 47312
rect 19563 47263 19605 47272
rect 19468 46423 19508 46432
rect 19371 46136 19413 46145
rect 19371 46096 19372 46136
rect 19412 46096 19413 46136
rect 19371 46087 19413 46096
rect 19372 45716 19412 46087
rect 19467 45884 19509 45893
rect 19467 45844 19468 45884
rect 19508 45844 19509 45884
rect 19467 45835 19509 45844
rect 19372 45667 19412 45676
rect 18795 43660 18796 43700
rect 18836 43660 18837 43700
rect 18795 43651 18837 43660
rect 18892 43660 19316 43700
rect 18796 43566 18836 43651
rect 18604 43532 18644 43541
rect 18604 43373 18644 43492
rect 18603 43364 18645 43373
rect 18603 43324 18604 43364
rect 18644 43324 18645 43364
rect 18603 43315 18645 43324
rect 18796 42701 18836 42786
rect 18795 42692 18837 42701
rect 18795 42652 18796 42692
rect 18836 42652 18837 42692
rect 18795 42643 18837 42652
rect 18892 42524 18932 43660
rect 18988 43532 19028 43541
rect 19372 43532 19412 43541
rect 19028 43492 19316 43532
rect 18988 43483 19028 43492
rect 19179 43280 19221 43289
rect 19179 43240 19180 43280
rect 19220 43240 19221 43280
rect 19179 43231 19221 43240
rect 19180 43146 19220 43231
rect 18987 42860 19029 42869
rect 18987 42820 18988 42860
rect 19028 42820 19029 42860
rect 18987 42811 19029 42820
rect 18988 42608 19028 42811
rect 18988 42559 19028 42568
rect 18700 42484 18932 42524
rect 18603 42440 18645 42449
rect 18603 42400 18604 42440
rect 18644 42400 18645 42440
rect 18603 42391 18645 42400
rect 18220 42139 18260 42148
rect 18316 42148 18452 42188
rect 18604 42188 18644 42391
rect 18123 42104 18165 42113
rect 18123 42064 18124 42104
rect 18164 42064 18165 42104
rect 18123 42055 18165 42064
rect 18028 42020 18068 42029
rect 18028 41516 18068 41980
rect 18028 41476 18164 41516
rect 17932 41392 18068 41432
rect 17932 41264 17972 41273
rect 17932 41189 17972 41224
rect 17931 41180 17973 41189
rect 17931 41140 17932 41180
rect 17972 41140 17973 41180
rect 17931 41131 17973 41140
rect 17835 40760 17877 40769
rect 17835 40720 17836 40760
rect 17876 40720 17877 40760
rect 17835 40711 17877 40720
rect 17739 39836 17781 39845
rect 17739 39796 17740 39836
rect 17780 39796 17781 39836
rect 17739 39787 17781 39796
rect 17547 39164 17589 39173
rect 17547 39124 17548 39164
rect 17588 39124 17589 39164
rect 17547 39115 17589 39124
rect 17740 39164 17780 39787
rect 17740 39115 17780 39124
rect 17835 39080 17877 39089
rect 17835 39040 17836 39080
rect 17876 39040 17877 39080
rect 17835 39031 17877 39040
rect 17548 38912 17588 38921
rect 17588 38872 17674 38912
rect 17548 38863 17588 38872
rect 17634 38837 17674 38872
rect 17634 38828 17685 38837
rect 17634 38788 17644 38828
rect 17684 38788 17685 38828
rect 17643 38779 17685 38788
rect 17452 38704 17588 38744
rect 17452 38240 17492 38249
rect 17116 38198 17156 38207
rect 17356 38200 17452 38240
rect 17116 38156 17156 38158
rect 17116 38116 17396 38156
rect 16875 37736 16917 37745
rect 16875 37696 16876 37736
rect 16916 37696 16917 37736
rect 16875 37687 16917 37696
rect 16876 35888 16916 37687
rect 17356 37652 17396 38116
rect 17356 37603 17396 37612
rect 17164 37400 17204 37409
rect 17204 37360 17300 37400
rect 17164 37351 17204 37360
rect 17067 36896 17109 36905
rect 17067 36856 17068 36896
rect 17108 36856 17109 36896
rect 17067 36847 17109 36856
rect 16971 36308 17013 36317
rect 16971 36268 16972 36308
rect 17012 36268 17013 36308
rect 16971 36259 17013 36268
rect 16876 35645 16916 35848
rect 16875 35636 16917 35645
rect 16875 35596 16876 35636
rect 16916 35596 16917 35636
rect 16875 35587 16917 35596
rect 16875 35468 16917 35477
rect 16875 35428 16876 35468
rect 16916 35428 16917 35468
rect 16875 35419 16917 35428
rect 16876 35216 16916 35419
rect 16876 35167 16916 35176
rect 16875 35048 16917 35057
rect 16875 35008 16876 35048
rect 16916 35008 16917 35048
rect 16875 34999 16917 35008
rect 16876 30680 16916 34999
rect 16779 30176 16821 30185
rect 16779 30136 16780 30176
rect 16820 30136 16821 30176
rect 16779 30127 16821 30136
rect 16876 29093 16916 30640
rect 16972 30521 17012 36259
rect 17068 35225 17108 36847
rect 17164 36714 17204 36723
rect 17067 35216 17109 35225
rect 17067 35176 17068 35216
rect 17108 35176 17109 35216
rect 17067 35167 17109 35176
rect 17068 34964 17108 34973
rect 17164 34964 17204 36674
rect 17260 35477 17300 37360
rect 17356 36812 17396 36821
rect 17356 36653 17396 36772
rect 17355 36644 17397 36653
rect 17355 36604 17356 36644
rect 17396 36604 17397 36644
rect 17355 36595 17397 36604
rect 17452 36569 17492 38200
rect 17451 36560 17493 36569
rect 17451 36520 17452 36560
rect 17492 36520 17493 36560
rect 17451 36511 17493 36520
rect 17548 36317 17588 38704
rect 17836 38501 17876 39031
rect 17835 38492 17877 38501
rect 17835 38452 17836 38492
rect 17876 38452 17877 38492
rect 17835 38443 17877 38452
rect 17835 38240 17877 38249
rect 17835 38200 17836 38240
rect 17876 38200 17877 38240
rect 17835 38191 17877 38200
rect 17547 36308 17589 36317
rect 17547 36268 17548 36308
rect 17588 36268 17589 36308
rect 17547 36259 17589 36268
rect 17259 35468 17301 35477
rect 17259 35428 17260 35468
rect 17300 35428 17301 35468
rect 17259 35419 17301 35428
rect 17451 35468 17493 35477
rect 17451 35428 17452 35468
rect 17492 35428 17493 35468
rect 17451 35419 17493 35428
rect 17260 35216 17300 35227
rect 17260 35141 17300 35176
rect 17355 35216 17397 35225
rect 17355 35176 17356 35216
rect 17396 35176 17397 35216
rect 17355 35167 17397 35176
rect 17259 35132 17301 35141
rect 17259 35092 17260 35132
rect 17300 35092 17301 35132
rect 17259 35083 17301 35092
rect 17108 34924 17204 34964
rect 17068 34915 17108 34924
rect 17067 34796 17109 34805
rect 17067 34756 17068 34796
rect 17108 34756 17109 34796
rect 17067 34747 17109 34756
rect 17068 34376 17108 34747
rect 17068 34327 17108 34336
rect 17356 33620 17396 35167
rect 17164 33580 17396 33620
rect 16971 30512 17013 30521
rect 16971 30472 16972 30512
rect 17012 30472 17013 30512
rect 16971 30463 17013 30472
rect 16875 29084 16917 29093
rect 16875 29044 16876 29084
rect 16916 29044 16917 29084
rect 16875 29035 16917 29044
rect 16396 28960 16724 29000
rect 16444 28337 16484 28346
rect 16484 28297 16532 28328
rect 16444 28288 16532 28297
rect 16395 28160 16437 28169
rect 16395 28120 16396 28160
rect 16436 28120 16437 28160
rect 16395 28111 16437 28120
rect 16203 27824 16245 27833
rect 16203 27784 16204 27824
rect 16244 27784 16245 27824
rect 16203 27775 16245 27784
rect 16396 27656 16436 28111
rect 16492 27824 16532 28288
rect 16587 28160 16629 28169
rect 16587 28120 16588 28160
rect 16628 28120 16629 28160
rect 16587 28111 16629 28120
rect 16588 28026 16628 28111
rect 16588 27824 16628 27833
rect 16492 27784 16588 27824
rect 16588 27775 16628 27784
rect 16396 26825 16436 27616
rect 16587 27656 16629 27665
rect 16587 27616 16588 27656
rect 16628 27616 16629 27656
rect 16587 27607 16629 27616
rect 16395 26816 16437 26825
rect 16395 26776 16396 26816
rect 16436 26776 16437 26816
rect 16395 26767 16437 26776
rect 16107 26480 16149 26489
rect 16107 26440 16108 26480
rect 16148 26440 16149 26480
rect 16107 26431 16149 26440
rect 16108 26228 16148 26237
rect 15860 26104 15956 26134
rect 15820 26094 15956 26104
rect 16012 26144 16052 26153
rect 16012 25976 16052 26104
rect 15820 25936 16052 25976
rect 15627 25724 15669 25733
rect 15627 25684 15628 25724
rect 15668 25684 15669 25724
rect 15627 25675 15669 25684
rect 15147 25304 15189 25313
rect 14956 25264 15148 25304
rect 15188 25264 15189 25304
rect 14763 23876 14805 23885
rect 14763 23836 14764 23876
rect 14804 23836 14805 23876
rect 14763 23827 14805 23836
rect 14572 23792 14612 23801
rect 14572 23633 14612 23752
rect 14668 23771 14708 23780
rect 14571 23624 14613 23633
rect 14571 23584 14572 23624
rect 14612 23584 14613 23624
rect 14571 23575 14613 23584
rect 14572 22793 14612 23575
rect 14668 23120 14708 23731
rect 14764 23771 14804 23780
rect 14764 23297 14804 23731
rect 14859 23624 14901 23633
rect 14859 23584 14860 23624
rect 14900 23584 14901 23624
rect 14859 23575 14901 23584
rect 14860 23490 14900 23575
rect 14763 23288 14805 23297
rect 14763 23248 14764 23288
rect 14804 23248 14805 23288
rect 14763 23239 14805 23248
rect 14860 23288 14900 23297
rect 14956 23288 14996 25264
rect 15147 25255 15189 25264
rect 15340 25304 15380 25313
rect 15148 25170 15188 25255
rect 15243 25220 15285 25229
rect 15243 25180 15244 25220
rect 15284 25180 15285 25220
rect 15243 25171 15285 25180
rect 15244 25086 15284 25171
rect 15340 24641 15380 25264
rect 15532 25304 15572 25315
rect 15532 25229 15572 25264
rect 15628 25304 15668 25313
rect 15531 25220 15573 25229
rect 15531 25180 15532 25220
rect 15572 25180 15573 25220
rect 15531 25171 15573 25180
rect 15339 24632 15381 24641
rect 15339 24592 15340 24632
rect 15380 24592 15381 24632
rect 15339 24583 15381 24592
rect 15243 24548 15285 24557
rect 15243 24508 15244 24548
rect 15284 24508 15285 24548
rect 15243 24499 15285 24508
rect 15147 23792 15189 23801
rect 15147 23752 15148 23792
rect 15188 23752 15189 23792
rect 15147 23743 15189 23752
rect 14900 23248 14996 23288
rect 15051 23288 15093 23297
rect 15051 23248 15052 23288
rect 15092 23248 15093 23288
rect 14860 23239 14900 23248
rect 15051 23239 15093 23248
rect 15052 23154 15092 23239
rect 15148 23129 15188 23743
rect 14763 23120 14805 23129
rect 14668 23080 14764 23120
rect 14804 23080 14805 23120
rect 14763 23071 14805 23080
rect 15147 23120 15189 23129
rect 15147 23080 15148 23120
rect 15188 23080 15189 23120
rect 15147 23071 15189 23080
rect 15244 23120 15284 24499
rect 15435 23876 15477 23885
rect 15435 23836 15436 23876
rect 15476 23836 15477 23876
rect 15435 23827 15477 23836
rect 15436 23792 15476 23827
rect 15436 23741 15476 23752
rect 15531 23708 15573 23717
rect 15531 23668 15532 23708
rect 15572 23668 15573 23708
rect 15531 23659 15573 23668
rect 14764 22986 14804 23071
rect 14571 22784 14613 22793
rect 14571 22744 14572 22784
rect 14612 22744 14613 22784
rect 14571 22735 14613 22744
rect 15051 22784 15093 22793
rect 15051 22744 15052 22784
rect 15092 22744 15093 22784
rect 15051 22735 15093 22744
rect 14668 22280 14708 22289
rect 14476 22240 14612 22280
rect 14476 22112 14516 22121
rect 14476 22037 14516 22072
rect 14470 22028 14516 22037
rect 14470 21988 14471 22028
rect 14511 21988 14516 22028
rect 14470 21979 14512 21988
rect 14475 21860 14517 21869
rect 14475 21820 14476 21860
rect 14516 21820 14517 21860
rect 14475 21811 14517 21820
rect 14283 20096 14325 20105
rect 14283 20056 14284 20096
rect 14324 20056 14325 20096
rect 14283 20047 14325 20056
rect 14284 19844 14324 19853
rect 14187 19424 14229 19433
rect 14187 19384 14188 19424
rect 14228 19384 14229 19424
rect 14187 19375 14229 19384
rect 14140 19265 14180 19274
rect 14284 19256 14324 19804
rect 14180 19225 14324 19256
rect 14140 19216 14324 19225
rect 14091 19088 14133 19097
rect 14091 19048 14092 19088
rect 14132 19048 14133 19088
rect 14091 19039 14133 19048
rect 14284 19088 14324 19099
rect 13995 17240 14037 17249
rect 13995 17200 13996 17240
rect 14036 17200 14037 17240
rect 13995 17191 14037 17200
rect 14092 16073 14132 19039
rect 14284 19013 14324 19048
rect 14476 19013 14516 21811
rect 14283 19004 14325 19013
rect 14283 18964 14284 19004
rect 14324 18964 14325 19004
rect 14283 18955 14325 18964
rect 14475 19004 14517 19013
rect 14475 18964 14476 19004
rect 14516 18964 14517 19004
rect 14475 18955 14517 18964
rect 14572 18761 14612 22240
rect 14668 19424 14708 22240
rect 14860 22280 14900 22289
rect 14764 22112 14804 22121
rect 14764 21617 14804 22072
rect 14763 21608 14805 21617
rect 14763 21568 14764 21608
rect 14804 21568 14805 21608
rect 14763 21559 14805 21568
rect 14763 21440 14805 21449
rect 14763 21400 14764 21440
rect 14804 21400 14805 21440
rect 14860 21440 14900 22240
rect 14956 22280 14996 22289
rect 14956 21785 14996 22240
rect 14955 21776 14997 21785
rect 14955 21736 14956 21776
rect 14996 21736 14997 21776
rect 14955 21727 14997 21736
rect 15052 21692 15092 22735
rect 15148 22532 15188 23071
rect 15148 22483 15188 22492
rect 15244 22280 15284 23080
rect 15532 22961 15572 23659
rect 15628 23381 15668 25264
rect 15724 25304 15764 25313
rect 15724 24389 15764 25264
rect 15820 25304 15860 25936
rect 16108 25565 16148 26188
rect 16204 26153 16244 26238
rect 16203 26144 16245 26153
rect 16203 26104 16204 26144
rect 16244 26104 16245 26144
rect 16203 26095 16245 26104
rect 16300 26144 16340 26153
rect 16203 25976 16245 25985
rect 16300 25976 16340 26104
rect 16396 25985 16436 26767
rect 16588 26489 16628 27607
rect 16684 26648 16724 28960
rect 16780 28337 16820 28422
rect 16779 28328 16821 28337
rect 16779 28288 16780 28328
rect 16820 28288 16821 28328
rect 16779 28279 16821 28288
rect 16780 27656 16820 27667
rect 16780 27581 16820 27616
rect 16779 27572 16821 27581
rect 16779 27532 16780 27572
rect 16820 27532 16821 27572
rect 16779 27523 16821 27532
rect 17067 27572 17109 27581
rect 17067 27532 17068 27572
rect 17108 27532 17109 27572
rect 17067 27523 17109 27532
rect 16971 26984 17013 26993
rect 16971 26944 16972 26984
rect 17012 26944 17013 26984
rect 16971 26935 17013 26944
rect 16780 26825 16820 26910
rect 16972 26850 17012 26935
rect 16779 26816 16821 26825
rect 16779 26776 16780 26816
rect 16820 26776 16821 26816
rect 16779 26767 16821 26776
rect 16971 26648 17013 26657
rect 16684 26608 16820 26648
rect 16587 26480 16629 26489
rect 16587 26440 16588 26480
rect 16628 26440 16629 26480
rect 16587 26431 16629 26440
rect 16491 26312 16533 26321
rect 16491 26272 16492 26312
rect 16532 26272 16533 26312
rect 16491 26263 16533 26272
rect 16492 26144 16532 26263
rect 16532 26104 16628 26144
rect 16492 26095 16532 26104
rect 16203 25936 16204 25976
rect 16244 25936 16340 25976
rect 16395 25976 16437 25985
rect 16395 25936 16396 25976
rect 16436 25936 16437 25976
rect 16203 25927 16245 25936
rect 16395 25927 16437 25936
rect 16107 25556 16149 25565
rect 16107 25516 16108 25556
rect 16148 25516 16149 25556
rect 16107 25507 16149 25516
rect 16107 25388 16149 25397
rect 16107 25348 16108 25388
rect 16148 25348 16149 25388
rect 16107 25339 16149 25348
rect 15820 25255 15860 25264
rect 16011 25304 16053 25313
rect 16011 25264 16012 25304
rect 16052 25264 16053 25304
rect 16011 25255 16053 25264
rect 16108 25304 16148 25339
rect 16300 25313 16340 25398
rect 16012 25170 16052 25255
rect 16108 25253 16148 25264
rect 16204 25304 16244 25313
rect 16204 25136 16244 25264
rect 16299 25304 16341 25313
rect 16299 25264 16300 25304
rect 16340 25264 16341 25304
rect 16299 25255 16341 25264
rect 16491 25304 16533 25313
rect 16491 25264 16492 25304
rect 16532 25264 16533 25304
rect 16491 25255 16533 25264
rect 16108 25096 16244 25136
rect 15916 24632 15956 24643
rect 15916 24557 15956 24592
rect 16108 24557 16148 25096
rect 16203 24968 16245 24977
rect 16203 24928 16204 24968
rect 16244 24928 16245 24968
rect 16203 24919 16245 24928
rect 15915 24548 15957 24557
rect 15915 24508 15916 24548
rect 15956 24508 15957 24548
rect 15915 24499 15957 24508
rect 16107 24548 16149 24557
rect 16107 24508 16108 24548
rect 16148 24508 16149 24548
rect 16107 24499 16149 24508
rect 15723 24380 15765 24389
rect 15723 24340 15724 24380
rect 15764 24340 15765 24380
rect 15723 24331 15765 24340
rect 16107 24380 16149 24389
rect 16107 24340 16108 24380
rect 16148 24340 16149 24380
rect 16107 24331 16149 24340
rect 16108 24246 16148 24331
rect 16012 24044 16052 24053
rect 16204 24044 16244 24919
rect 16395 24884 16437 24893
rect 16395 24844 16396 24884
rect 16436 24844 16437 24884
rect 16395 24835 16437 24844
rect 16396 24800 16436 24835
rect 16396 24749 16436 24760
rect 16299 24632 16341 24641
rect 16299 24592 16300 24632
rect 16340 24592 16341 24632
rect 16299 24583 16341 24592
rect 16492 24632 16532 25255
rect 16588 25229 16628 26104
rect 16683 25724 16725 25733
rect 16683 25684 16684 25724
rect 16724 25684 16725 25724
rect 16683 25675 16725 25684
rect 16684 25304 16724 25675
rect 16780 25481 16820 26608
rect 16971 26608 16972 26648
rect 17012 26608 17013 26648
rect 16971 26599 17013 26608
rect 16875 26144 16917 26153
rect 16875 26104 16876 26144
rect 16916 26104 16917 26144
rect 16875 26095 16917 26104
rect 16779 25472 16821 25481
rect 16779 25432 16780 25472
rect 16820 25432 16821 25472
rect 16779 25423 16821 25432
rect 16684 25255 16724 25264
rect 16587 25220 16629 25229
rect 16587 25180 16588 25220
rect 16628 25180 16629 25220
rect 16587 25171 16629 25180
rect 16492 24583 16532 24592
rect 16588 24632 16628 24641
rect 16780 24632 16820 24641
rect 16300 24498 16340 24583
rect 16491 24128 16533 24137
rect 16491 24088 16492 24128
rect 16532 24088 16533 24128
rect 16491 24079 16533 24088
rect 16052 24004 16244 24044
rect 16012 23995 16052 24004
rect 15820 23960 15860 23969
rect 15723 23876 15765 23885
rect 15723 23836 15724 23876
rect 15764 23836 15765 23876
rect 15723 23827 15765 23836
rect 15724 23549 15764 23827
rect 15723 23540 15765 23549
rect 15723 23500 15724 23540
rect 15764 23500 15765 23540
rect 15723 23491 15765 23500
rect 15627 23372 15669 23381
rect 15627 23332 15628 23372
rect 15668 23332 15669 23372
rect 15627 23323 15669 23332
rect 15531 22952 15573 22961
rect 15531 22912 15532 22952
rect 15572 22912 15573 22952
rect 15531 22903 15573 22912
rect 15724 22793 15764 23491
rect 15820 23129 15860 23920
rect 16299 23876 16341 23885
rect 16299 23836 16300 23876
rect 16340 23836 16341 23876
rect 16299 23827 16341 23836
rect 16300 23792 16340 23827
rect 16300 23741 16340 23752
rect 16396 23792 16436 23801
rect 16203 23204 16245 23213
rect 16203 23164 16204 23204
rect 16244 23164 16245 23204
rect 16203 23155 16245 23164
rect 15819 23120 15861 23129
rect 15819 23080 15820 23120
rect 15860 23080 15861 23120
rect 15819 23071 15861 23080
rect 15723 22784 15765 22793
rect 15723 22744 15724 22784
rect 15764 22744 15765 22784
rect 15723 22735 15765 22744
rect 15340 22280 15380 22289
rect 15244 22240 15340 22280
rect 15052 21652 15188 21692
rect 15053 21524 15093 21652
rect 15148 21608 15188 21652
rect 15148 21559 15188 21568
rect 15244 21533 15284 22240
rect 15340 22231 15380 22240
rect 15723 22280 15765 22289
rect 15723 22240 15724 22280
rect 15764 22240 15765 22280
rect 15723 22231 15765 22240
rect 15339 21776 15381 21785
rect 15339 21736 15340 21776
rect 15380 21736 15381 21776
rect 15339 21727 15381 21736
rect 15724 21776 15764 22231
rect 15915 22028 15957 22037
rect 15915 21988 15916 22028
rect 15956 21988 15957 22028
rect 15915 21979 15957 21988
rect 15724 21727 15764 21736
rect 15819 21776 15861 21785
rect 15819 21736 15820 21776
rect 15860 21736 15861 21776
rect 15819 21727 15861 21736
rect 15340 21642 15380 21727
rect 15532 21617 15572 21702
rect 15531 21608 15573 21617
rect 15531 21568 15532 21608
rect 15572 21568 15573 21608
rect 15531 21559 15573 21568
rect 15628 21608 15668 21617
rect 15052 21484 15093 21524
rect 15243 21524 15285 21533
rect 15243 21484 15244 21524
rect 15284 21484 15285 21524
rect 14955 21440 14997 21449
rect 14860 21400 14956 21440
rect 14996 21400 14997 21440
rect 14763 21391 14805 21400
rect 14955 21391 14997 21400
rect 14764 20180 14804 21391
rect 14955 20768 14997 20777
rect 15052 20768 15092 21484
rect 15243 21475 15285 21484
rect 15147 21440 15189 21449
rect 15147 21400 15148 21440
rect 15188 21400 15189 21440
rect 15147 21391 15189 21400
rect 15148 21020 15188 21391
rect 15148 20971 15188 20980
rect 14955 20728 14956 20768
rect 14996 20728 15092 20768
rect 14955 20719 14997 20728
rect 14956 20634 14996 20719
rect 15244 20273 15284 21475
rect 15339 21440 15381 21449
rect 15339 21400 15340 21440
rect 15380 21400 15381 21440
rect 15339 21391 15381 21400
rect 15340 20768 15380 21391
rect 15340 20719 15380 20728
rect 15435 20768 15477 20777
rect 15435 20728 15436 20768
rect 15476 20728 15477 20768
rect 15435 20719 15477 20728
rect 15436 20634 15476 20719
rect 15339 20600 15381 20609
rect 15339 20560 15340 20600
rect 15380 20560 15381 20600
rect 15339 20551 15381 20560
rect 15628 20600 15668 21568
rect 15820 21608 15860 21727
rect 15820 21559 15860 21568
rect 15916 21608 15956 21979
rect 15916 21559 15956 21568
rect 16017 21608 16057 21617
rect 15723 21524 15765 21533
rect 15723 21484 15724 21524
rect 15764 21484 15765 21524
rect 15723 21475 15765 21484
rect 15724 21029 15764 21475
rect 16017 21449 16057 21568
rect 16016 21440 16058 21449
rect 16016 21400 16017 21440
rect 16057 21400 16058 21440
rect 16016 21391 16058 21400
rect 15723 21020 15765 21029
rect 15723 20980 15724 21020
rect 15764 20980 15765 21020
rect 15723 20971 15765 20980
rect 16107 20768 16149 20777
rect 16107 20728 16108 20768
rect 16148 20728 16149 20768
rect 16107 20719 16149 20728
rect 16108 20634 16148 20719
rect 16012 20600 16052 20609
rect 15628 20551 15668 20560
rect 15820 20560 16012 20600
rect 15243 20264 15285 20273
rect 15243 20224 15244 20264
rect 15284 20224 15285 20264
rect 15243 20215 15285 20224
rect 14764 20140 14900 20180
rect 14860 20096 14900 20140
rect 14860 19601 14900 20056
rect 15051 19844 15093 19853
rect 15051 19804 15052 19844
rect 15092 19804 15093 19844
rect 15051 19795 15093 19804
rect 14859 19592 14901 19601
rect 14859 19552 14860 19592
rect 14900 19552 14901 19592
rect 14859 19543 14901 19552
rect 14668 19384 14996 19424
rect 14668 19256 14708 19265
rect 14668 19181 14708 19216
rect 14860 19256 14900 19267
rect 14860 19181 14900 19216
rect 14667 19172 14709 19181
rect 14667 19132 14668 19172
rect 14708 19132 14709 19172
rect 14667 19123 14709 19132
rect 14859 19172 14901 19181
rect 14859 19132 14860 19172
rect 14900 19132 14901 19172
rect 14859 19123 14901 19132
rect 14668 18929 14708 19123
rect 14763 19088 14805 19097
rect 14763 19048 14764 19088
rect 14804 19048 14805 19088
rect 14763 19039 14805 19048
rect 14764 18954 14804 19039
rect 14667 18920 14709 18929
rect 14667 18880 14668 18920
rect 14708 18880 14709 18920
rect 14667 18871 14709 18880
rect 14187 18752 14229 18761
rect 14187 18712 14188 18752
rect 14228 18712 14229 18752
rect 14187 18703 14229 18712
rect 14571 18752 14613 18761
rect 14571 18712 14572 18752
rect 14612 18712 14613 18752
rect 14571 18703 14613 18712
rect 14763 18752 14805 18761
rect 14763 18712 14764 18752
rect 14804 18712 14805 18752
rect 14763 18703 14805 18712
rect 14091 16064 14133 16073
rect 14091 16024 14092 16064
rect 14132 16024 14133 16064
rect 14091 16015 14133 16024
rect 13995 13460 14037 13469
rect 13995 13420 13996 13460
rect 14036 13420 14037 13460
rect 13995 13411 14037 13420
rect 13996 12368 14036 13411
rect 14092 12797 14132 16015
rect 14188 15644 14228 18703
rect 14475 18668 14517 18677
rect 14475 18628 14476 18668
rect 14516 18628 14517 18668
rect 14475 18619 14517 18628
rect 14284 18570 14324 18579
rect 14476 18534 14516 18619
rect 14667 18584 14709 18593
rect 14667 18544 14668 18584
rect 14708 18544 14709 18584
rect 14667 18535 14709 18544
rect 14284 18005 14324 18530
rect 14475 18248 14517 18257
rect 14475 18208 14476 18248
rect 14516 18208 14517 18248
rect 14475 18199 14517 18208
rect 14283 17996 14325 18005
rect 14283 17956 14284 17996
rect 14324 17956 14325 17996
rect 14283 17947 14325 17956
rect 14283 16820 14325 16829
rect 14283 16780 14284 16820
rect 14324 16780 14325 16820
rect 14283 16771 14325 16780
rect 14284 16246 14324 16771
rect 14284 16197 14324 16206
rect 14476 16232 14516 18199
rect 14668 17744 14708 18535
rect 14764 17828 14804 18703
rect 14956 18416 14996 19384
rect 15052 19256 15092 19795
rect 15052 19207 15092 19216
rect 15148 19256 15188 19265
rect 15148 19013 15188 19216
rect 15340 19256 15380 20551
rect 15435 19760 15477 19769
rect 15435 19720 15436 19760
rect 15476 19720 15477 19760
rect 15435 19711 15477 19720
rect 15340 19207 15380 19216
rect 15244 19088 15284 19097
rect 15147 19004 15189 19013
rect 15147 18964 15148 19004
rect 15188 18964 15189 19004
rect 15147 18955 15189 18964
rect 15052 18593 15092 18678
rect 15051 18584 15093 18593
rect 15051 18544 15052 18584
rect 15092 18544 15188 18584
rect 15051 18535 15093 18544
rect 14956 18376 15092 18416
rect 14860 18005 14900 18090
rect 14859 17996 14901 18005
rect 14859 17956 14860 17996
rect 14900 17956 14901 17996
rect 14859 17947 14901 17956
rect 14764 17788 14900 17828
rect 14571 17240 14613 17249
rect 14571 17200 14572 17240
rect 14612 17200 14613 17240
rect 14571 17191 14613 17200
rect 14572 17072 14612 17191
rect 14572 16997 14612 17032
rect 14571 16988 14613 16997
rect 14571 16948 14572 16988
rect 14612 16948 14613 16988
rect 14571 16939 14613 16948
rect 14476 16192 14612 16232
rect 14475 16064 14517 16073
rect 14475 16024 14476 16064
rect 14516 16024 14517 16064
rect 14475 16015 14517 16024
rect 14476 15930 14516 16015
rect 14476 15644 14516 15653
rect 14188 15604 14476 15644
rect 14188 14393 14228 15604
rect 14476 15595 14516 15604
rect 14332 15550 14372 15559
rect 14372 15510 14516 15550
rect 14332 15501 14372 15510
rect 14476 14972 14516 15510
rect 14572 15140 14612 16192
rect 14668 15728 14708 17704
rect 14763 16820 14805 16829
rect 14763 16780 14764 16820
rect 14804 16780 14805 16820
rect 14763 16771 14805 16780
rect 14764 16686 14804 16771
rect 14668 15688 14804 15728
rect 14667 15560 14709 15569
rect 14667 15520 14668 15560
rect 14708 15520 14709 15560
rect 14667 15511 14709 15520
rect 14668 15426 14708 15511
rect 14572 15100 14708 15140
rect 14572 14972 14612 14981
rect 14476 14932 14572 14972
rect 14572 14923 14612 14932
rect 14379 14804 14421 14813
rect 14379 14764 14380 14804
rect 14420 14764 14421 14804
rect 14379 14755 14421 14764
rect 14380 14720 14420 14755
rect 14380 14669 14420 14680
rect 14668 14552 14708 15100
rect 14764 14813 14804 15688
rect 14763 14804 14805 14813
rect 14763 14764 14764 14804
rect 14804 14764 14805 14804
rect 14763 14755 14805 14764
rect 14284 14512 14708 14552
rect 14187 14384 14229 14393
rect 14187 14344 14188 14384
rect 14228 14344 14229 14384
rect 14187 14335 14229 14344
rect 14284 14048 14324 14512
rect 14860 14468 14900 17788
rect 14955 15140 14997 15149
rect 14955 15100 14956 15140
rect 14996 15100 14997 15140
rect 14955 15091 14997 15100
rect 14956 14477 14996 15091
rect 14188 14008 14284 14048
rect 14091 12788 14133 12797
rect 14091 12748 14092 12788
rect 14132 12748 14133 12788
rect 14091 12739 14133 12748
rect 14188 12620 14228 14008
rect 14284 13999 14324 14008
rect 14380 14428 14900 14468
rect 14955 14468 14997 14477
rect 14955 14428 14956 14468
rect 14996 14428 14997 14468
rect 14380 13880 14420 14428
rect 14955 14419 14997 14428
rect 14956 14132 14996 14141
rect 14284 13840 14420 13880
rect 14476 14092 14956 14132
rect 14284 12881 14324 13840
rect 14379 13208 14421 13217
rect 14379 13168 14380 13208
rect 14420 13168 14421 13208
rect 14379 13159 14421 13168
rect 14380 13074 14420 13159
rect 14283 12872 14325 12881
rect 14283 12832 14284 12872
rect 14324 12832 14325 12872
rect 14283 12823 14325 12832
rect 13996 12319 14036 12328
rect 14092 12580 14228 12620
rect 14092 12284 14132 12580
rect 14188 12452 14228 12461
rect 14476 12452 14516 14092
rect 14956 14083 14996 14092
rect 14764 14034 14804 14043
rect 15052 14034 15092 18376
rect 15148 17081 15188 18544
rect 15244 17669 15284 19048
rect 15436 18593 15476 19711
rect 15723 19424 15765 19433
rect 15723 19384 15724 19424
rect 15764 19384 15765 19424
rect 15723 19375 15765 19384
rect 15627 19256 15669 19265
rect 15627 19216 15628 19256
rect 15668 19216 15669 19256
rect 15627 19207 15669 19216
rect 15724 19256 15764 19375
rect 15628 19122 15668 19207
rect 15532 19088 15572 19099
rect 15532 19013 15572 19048
rect 15531 19004 15573 19013
rect 15531 18964 15532 19004
rect 15572 18964 15573 19004
rect 15531 18955 15573 18964
rect 15627 18920 15669 18929
rect 15627 18880 15628 18920
rect 15668 18880 15669 18920
rect 15627 18871 15669 18880
rect 15435 18584 15477 18593
rect 15435 18544 15436 18584
rect 15476 18544 15477 18584
rect 15435 18535 15477 18544
rect 15436 17837 15476 17868
rect 15435 17828 15477 17837
rect 15435 17788 15436 17828
rect 15476 17788 15477 17828
rect 15435 17779 15477 17788
rect 15436 17744 15476 17779
rect 15243 17660 15285 17669
rect 15243 17620 15244 17660
rect 15284 17620 15285 17660
rect 15243 17611 15285 17620
rect 15147 17072 15189 17081
rect 15147 17032 15148 17072
rect 15188 17032 15189 17072
rect 15147 17023 15189 17032
rect 15243 16988 15285 16997
rect 15243 16948 15244 16988
rect 15284 16948 15285 16988
rect 15243 16939 15285 16948
rect 15244 15065 15284 16939
rect 15436 15569 15476 17704
rect 15628 16820 15668 18871
rect 15724 17249 15764 19216
rect 15820 19256 15860 20560
rect 16012 20551 16052 20560
rect 15915 20096 15957 20105
rect 15915 20056 15916 20096
rect 15956 20056 15957 20096
rect 15915 20047 15957 20056
rect 16108 20096 16148 20105
rect 15820 19181 15860 19216
rect 15819 19172 15861 19181
rect 15819 19132 15820 19172
rect 15860 19132 15861 19172
rect 15819 19123 15861 19132
rect 15820 19092 15860 19123
rect 15916 19004 15956 20047
rect 16108 19769 16148 20056
rect 16107 19760 16149 19769
rect 16107 19720 16108 19760
rect 16148 19720 16149 19760
rect 16107 19711 16149 19720
rect 16011 19592 16053 19601
rect 16011 19552 16012 19592
rect 16052 19552 16053 19592
rect 16011 19543 16053 19552
rect 15820 18964 15956 19004
rect 15723 17240 15765 17249
rect 15723 17200 15724 17240
rect 15764 17200 15765 17240
rect 15723 17191 15765 17200
rect 15723 17072 15765 17081
rect 15723 17032 15724 17072
rect 15764 17032 15765 17072
rect 15723 17023 15765 17032
rect 15724 16938 15764 17023
rect 15628 16780 15764 16820
rect 15724 16241 15764 16780
rect 15532 16232 15572 16241
rect 15532 16073 15572 16192
rect 15628 16232 15668 16241
rect 15531 16064 15573 16073
rect 15531 16024 15532 16064
rect 15572 16024 15573 16064
rect 15531 16015 15573 16024
rect 15628 15728 15668 16192
rect 15723 16232 15765 16241
rect 15723 16192 15724 16232
rect 15764 16192 15765 16232
rect 15723 16183 15765 16192
rect 15723 16064 15765 16073
rect 15723 16024 15724 16064
rect 15764 16024 15765 16064
rect 15723 16015 15765 16024
rect 15724 15737 15764 16015
rect 15532 15688 15668 15728
rect 15723 15728 15765 15737
rect 15723 15688 15724 15728
rect 15764 15688 15765 15728
rect 15435 15560 15477 15569
rect 15435 15520 15436 15560
rect 15476 15520 15477 15560
rect 15435 15511 15477 15520
rect 15339 15476 15381 15485
rect 15339 15436 15340 15476
rect 15380 15436 15381 15476
rect 15339 15427 15381 15436
rect 15243 15056 15285 15065
rect 15243 15016 15244 15056
rect 15284 15016 15285 15056
rect 15243 15007 15285 15016
rect 15243 14804 15285 14813
rect 15243 14764 15244 14804
rect 15284 14764 15285 14804
rect 15243 14755 15285 14764
rect 15148 14720 15188 14729
rect 15148 14216 15188 14680
rect 15244 14720 15284 14755
rect 15244 14669 15284 14680
rect 15340 14300 15380 15427
rect 15532 15149 15572 15688
rect 15723 15679 15765 15688
rect 15627 15560 15669 15569
rect 15627 15520 15628 15560
rect 15668 15520 15669 15560
rect 15627 15511 15669 15520
rect 15531 15140 15573 15149
rect 15531 15100 15532 15140
rect 15572 15100 15573 15140
rect 15531 15091 15573 15100
rect 15628 14888 15668 15511
rect 15820 15392 15860 18964
rect 16012 18920 16052 19543
rect 16108 19256 16148 19267
rect 16108 19181 16148 19216
rect 16107 19172 16149 19181
rect 16107 19132 16108 19172
rect 16148 19132 16149 19172
rect 16107 19123 16149 19132
rect 15916 18880 16052 18920
rect 15916 16157 15956 18880
rect 16107 18668 16149 18677
rect 16107 18628 16108 18668
rect 16148 18628 16149 18668
rect 16107 18619 16149 18628
rect 16012 16232 16052 16241
rect 15915 16148 15957 16157
rect 15915 16108 15916 16148
rect 15956 16108 15957 16148
rect 15915 16099 15957 16108
rect 16012 16073 16052 16192
rect 16108 16232 16148 18619
rect 16204 17837 16244 23155
rect 16396 22625 16436 23752
rect 16492 23456 16532 24079
rect 16588 23624 16628 24592
rect 16684 24592 16780 24632
rect 16684 24053 16724 24592
rect 16780 24583 16820 24592
rect 16683 24044 16725 24053
rect 16683 24004 16684 24044
rect 16724 24004 16725 24044
rect 16683 23995 16725 24004
rect 16684 23801 16724 23886
rect 16683 23792 16725 23801
rect 16683 23752 16684 23792
rect 16724 23752 16725 23792
rect 16683 23743 16725 23752
rect 16588 23584 16724 23624
rect 16492 23416 16628 23456
rect 16492 23078 16532 23131
rect 16491 23038 16492 23045
rect 16532 23038 16533 23045
rect 16491 23036 16533 23038
rect 16491 22996 16492 23036
rect 16532 22996 16533 23036
rect 16491 22987 16533 22996
rect 16395 22616 16437 22625
rect 16395 22576 16396 22616
rect 16436 22576 16437 22616
rect 16395 22567 16437 22576
rect 16588 22541 16628 23416
rect 16684 23288 16724 23584
rect 16780 23288 16820 23297
rect 16684 23248 16780 23288
rect 16780 23239 16820 23248
rect 16876 23213 16916 26095
rect 16972 25313 17012 26599
rect 16971 25304 17013 25313
rect 16971 25264 16972 25304
rect 17012 25264 17013 25304
rect 16971 25255 17013 25264
rect 17068 24800 17108 27523
rect 16972 24760 17108 24800
rect 16972 24137 17012 24760
rect 17067 24212 17109 24221
rect 17067 24172 17068 24212
rect 17108 24172 17109 24212
rect 17067 24163 17109 24172
rect 16971 24128 17013 24137
rect 16971 24088 16972 24128
rect 17012 24088 17013 24128
rect 16971 24079 17013 24088
rect 17068 23771 17108 24163
rect 17164 23969 17204 33580
rect 17355 33452 17397 33461
rect 17355 33412 17356 33452
rect 17396 33412 17397 33452
rect 17355 33403 17397 33412
rect 17259 31436 17301 31445
rect 17259 31396 17260 31436
rect 17300 31396 17301 31436
rect 17259 31387 17301 31396
rect 17260 30689 17300 31387
rect 17259 30680 17301 30689
rect 17259 30640 17260 30680
rect 17300 30640 17301 30680
rect 17259 30631 17301 30640
rect 17260 29840 17300 30631
rect 17260 29168 17300 29800
rect 17260 28925 17300 29128
rect 17356 29000 17396 33403
rect 17452 31445 17492 35419
rect 17739 35216 17781 35225
rect 17739 35176 17740 35216
rect 17780 35176 17781 35216
rect 17739 35167 17781 35176
rect 17740 34385 17780 35167
rect 17836 35141 17876 38191
rect 17932 36569 17972 41131
rect 18028 37820 18068 41392
rect 18124 40013 18164 41476
rect 18316 41441 18356 42148
rect 18604 42139 18644 42148
rect 18412 42020 18452 42029
rect 18315 41432 18357 41441
rect 18315 41392 18316 41432
rect 18356 41392 18357 41432
rect 18315 41383 18357 41392
rect 18219 40676 18261 40685
rect 18219 40636 18220 40676
rect 18260 40636 18261 40676
rect 18219 40627 18261 40636
rect 18220 40424 18260 40627
rect 18260 40384 18356 40424
rect 18220 40375 18260 40384
rect 18123 40004 18165 40013
rect 18123 39964 18124 40004
rect 18164 39964 18165 40004
rect 18123 39955 18165 39964
rect 18114 39845 18154 39857
rect 18113 39836 18155 39845
rect 18113 39796 18114 39836
rect 18154 39796 18164 39836
rect 18113 39787 18164 39796
rect 18124 39772 18164 39787
rect 18124 39723 18164 39732
rect 18220 39752 18260 39761
rect 18220 39668 18260 39712
rect 18124 39628 18260 39668
rect 18124 38669 18164 39628
rect 18316 39584 18356 40384
rect 18412 39929 18452 41980
rect 18507 41348 18549 41357
rect 18507 41308 18508 41348
rect 18548 41308 18549 41348
rect 18507 41299 18549 41308
rect 18411 39920 18453 39929
rect 18411 39880 18412 39920
rect 18452 39880 18453 39920
rect 18411 39871 18453 39880
rect 18220 39544 18356 39584
rect 18123 38660 18165 38669
rect 18123 38620 18124 38660
rect 18164 38620 18165 38660
rect 18123 38611 18165 38620
rect 18028 37780 18164 37820
rect 18124 36905 18164 37780
rect 18123 36896 18165 36905
rect 18123 36856 18124 36896
rect 18164 36856 18165 36896
rect 18123 36847 18165 36856
rect 17931 36560 17973 36569
rect 17931 36520 17932 36560
rect 17972 36520 17973 36560
rect 17931 36511 17973 36520
rect 17932 35309 17972 36511
rect 18124 35888 18164 35897
rect 18124 35729 18164 35848
rect 18220 35813 18260 39544
rect 18508 39089 18548 41299
rect 18700 40676 18740 42484
rect 18808 42356 19176 42365
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 18808 42307 19176 42316
rect 18987 42188 19029 42197
rect 18987 42148 18988 42188
rect 19028 42148 19029 42188
rect 18987 42139 19029 42148
rect 18988 42054 19028 42139
rect 18796 42020 18836 42029
rect 18796 41189 18836 41980
rect 19179 42020 19221 42029
rect 19179 41980 19180 42020
rect 19220 41980 19221 42020
rect 19179 41971 19221 41980
rect 19180 41886 19220 41971
rect 19180 41264 19220 41273
rect 18795 41180 18837 41189
rect 18795 41140 18796 41180
rect 18836 41140 18837 41180
rect 18795 41131 18837 41140
rect 19180 41021 19220 41224
rect 19179 41012 19221 41021
rect 19179 40972 19180 41012
rect 19220 40972 19221 41012
rect 19179 40963 19221 40972
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 19276 40685 19316 43492
rect 19372 43205 19412 43492
rect 19371 43196 19413 43205
rect 19371 43156 19372 43196
rect 19412 43156 19413 43196
rect 19371 43147 19413 43156
rect 19372 42692 19412 42701
rect 19372 42533 19412 42652
rect 19371 42524 19413 42533
rect 19371 42484 19372 42524
rect 19412 42484 19413 42524
rect 19371 42475 19413 42484
rect 19371 42188 19413 42197
rect 19371 42148 19372 42188
rect 19412 42148 19413 42188
rect 19371 42139 19413 42148
rect 19372 42054 19412 42139
rect 19371 41012 19413 41021
rect 19371 40972 19372 41012
rect 19412 40972 19413 41012
rect 19371 40963 19413 40972
rect 19372 40878 19412 40963
rect 19275 40676 19317 40685
rect 18700 40636 18932 40676
rect 18892 40340 18932 40636
rect 19275 40636 19276 40676
rect 19316 40636 19317 40676
rect 19275 40627 19317 40636
rect 19468 40592 19508 45835
rect 19564 45716 19604 47263
rect 19756 45893 19796 48868
rect 19852 47298 19892 47307
rect 19755 45884 19797 45893
rect 19755 45844 19756 45884
rect 19796 45844 19797 45884
rect 19755 45835 19797 45844
rect 19755 45716 19797 45725
rect 19564 45676 19700 45716
rect 19563 45548 19605 45557
rect 19563 45508 19564 45548
rect 19604 45508 19605 45548
rect 19563 45499 19605 45508
rect 19564 45414 19604 45499
rect 19563 44120 19605 44129
rect 19563 44080 19564 44120
rect 19604 44080 19605 44120
rect 19563 44071 19605 44080
rect 19564 43700 19604 44071
rect 19564 43651 19604 43660
rect 19563 42776 19605 42785
rect 19563 42736 19564 42776
rect 19604 42736 19605 42776
rect 19563 42727 19605 42736
rect 19564 42608 19604 42727
rect 19564 42559 19604 42568
rect 19564 42020 19604 42029
rect 19564 41777 19604 41980
rect 19563 41768 19605 41777
rect 19563 41728 19564 41768
rect 19604 41728 19605 41768
rect 19563 41719 19605 41728
rect 19660 41516 19700 45676
rect 19755 45676 19756 45716
rect 19796 45676 19797 45716
rect 19755 45667 19797 45676
rect 19756 45582 19796 45667
rect 19755 45464 19797 45473
rect 19755 45424 19756 45464
rect 19796 45424 19797 45464
rect 19755 45415 19797 45424
rect 19756 44960 19796 45415
rect 19756 44045 19796 44920
rect 19852 44456 19892 47258
rect 19948 46985 19988 49036
rect 20048 47648 20416 47657
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20048 47599 20416 47608
rect 20043 47396 20085 47405
rect 20043 47356 20044 47396
rect 20084 47356 20085 47396
rect 20043 47347 20085 47356
rect 20044 47262 20084 47347
rect 19947 46976 19989 46985
rect 19947 46936 19948 46976
rect 19988 46936 19989 46976
rect 19947 46927 19989 46936
rect 19948 46477 19988 46486
rect 19948 45716 19988 46437
rect 20140 46304 20180 46313
rect 20180 46264 20564 46304
rect 20140 46255 20180 46264
rect 20048 46136 20416 46145
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20048 46087 20416 46096
rect 19948 45676 20084 45716
rect 19947 45548 19989 45557
rect 19947 45508 19948 45548
rect 19988 45508 19989 45548
rect 19947 45499 19989 45508
rect 19948 45414 19988 45499
rect 19948 45212 19988 45221
rect 20044 45212 20084 45676
rect 19988 45172 20084 45212
rect 19948 45163 19988 45172
rect 20048 44624 20416 44633
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20048 44575 20416 44584
rect 20044 44456 20084 44465
rect 19852 44416 20044 44456
rect 20044 44407 20084 44416
rect 20524 44297 20564 46264
rect 19851 44288 19893 44297
rect 19851 44248 19852 44288
rect 19892 44248 19893 44288
rect 19851 44239 19893 44248
rect 20523 44288 20565 44297
rect 20523 44248 20524 44288
rect 20564 44248 20565 44288
rect 20523 44239 20565 44248
rect 19852 44154 19892 44239
rect 20620 44129 20660 64399
rect 20716 63785 20756 67087
rect 20812 66053 20852 68020
rect 20907 67808 20949 67817
rect 20907 67768 20908 67808
rect 20948 67768 20949 67808
rect 20907 67759 20949 67768
rect 20811 66044 20853 66053
rect 20811 66004 20812 66044
rect 20852 66004 20853 66044
rect 20811 65995 20853 66004
rect 20811 65792 20853 65801
rect 20811 65752 20812 65792
rect 20852 65752 20853 65792
rect 20811 65743 20853 65752
rect 20812 64205 20852 65743
rect 20811 64196 20853 64205
rect 20811 64156 20812 64196
rect 20852 64156 20853 64196
rect 20811 64147 20853 64156
rect 20908 63869 20948 67759
rect 21003 66800 21045 66809
rect 21003 66760 21004 66800
rect 21044 66760 21045 66800
rect 21003 66751 21045 66760
rect 21004 64709 21044 66751
rect 21003 64700 21045 64709
rect 21003 64660 21004 64700
rect 21044 64660 21045 64700
rect 21003 64651 21045 64660
rect 20907 63860 20949 63869
rect 20907 63820 20908 63860
rect 20948 63820 20949 63860
rect 20907 63811 20949 63820
rect 20715 63776 20757 63785
rect 20715 63736 20716 63776
rect 20756 63736 20757 63776
rect 20715 63727 20757 63736
rect 20811 63692 20853 63701
rect 20811 63652 20812 63692
rect 20852 63652 20853 63692
rect 20811 63643 20853 63652
rect 20715 60668 20757 60677
rect 20715 60628 20716 60668
rect 20756 60628 20757 60668
rect 20715 60619 20757 60628
rect 20716 57065 20756 60619
rect 20812 59753 20852 63643
rect 21003 63104 21045 63113
rect 21003 63064 21004 63104
rect 21044 63064 21045 63104
rect 21003 63055 21045 63064
rect 20907 59912 20949 59921
rect 20907 59872 20908 59912
rect 20948 59872 20949 59912
rect 20907 59863 20949 59872
rect 20811 59744 20853 59753
rect 20811 59704 20812 59744
rect 20852 59704 20853 59744
rect 20811 59695 20853 59704
rect 20715 57056 20757 57065
rect 20715 57016 20716 57056
rect 20756 57016 20757 57056
rect 20715 57007 20757 57016
rect 20811 56888 20853 56897
rect 20811 56848 20812 56888
rect 20852 56848 20853 56888
rect 20811 56839 20853 56848
rect 20715 52856 20757 52865
rect 20715 52816 20716 52856
rect 20756 52816 20757 52856
rect 20715 52807 20757 52816
rect 20716 44633 20756 52807
rect 20812 45977 20852 56839
rect 20908 47321 20948 59863
rect 20907 47312 20949 47321
rect 20907 47272 20908 47312
rect 20948 47272 20949 47312
rect 20907 47263 20949 47272
rect 20811 45968 20853 45977
rect 20811 45928 20812 45968
rect 20852 45928 20853 45968
rect 20811 45919 20853 45928
rect 20715 44624 20757 44633
rect 20715 44584 20716 44624
rect 20756 44584 20757 44624
rect 20715 44575 20757 44584
rect 20619 44120 20661 44129
rect 20619 44080 20620 44120
rect 20660 44080 20661 44120
rect 20619 44071 20661 44080
rect 19755 44036 19797 44045
rect 19755 43996 19756 44036
rect 19796 43996 19797 44036
rect 19755 43987 19797 43996
rect 19755 43784 19797 43793
rect 19755 43744 19756 43784
rect 19796 43744 19797 43784
rect 19755 43735 19797 43744
rect 19756 43532 19796 43735
rect 19947 43700 19989 43709
rect 19947 43660 19948 43700
rect 19988 43660 19989 43700
rect 19947 43651 19989 43660
rect 19948 43566 19988 43651
rect 19756 43483 19796 43492
rect 20048 43112 20416 43121
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20048 43063 20416 43072
rect 20907 42944 20949 42953
rect 20907 42904 20908 42944
rect 20948 42904 20949 42944
rect 20907 42895 20949 42904
rect 19756 42692 19796 42701
rect 19756 42113 19796 42652
rect 19947 42524 19989 42533
rect 19947 42484 19948 42524
rect 19988 42484 19989 42524
rect 19947 42475 19989 42484
rect 19948 42390 19988 42475
rect 20139 42188 20181 42197
rect 20139 42148 20140 42188
rect 20180 42148 20181 42188
rect 20139 42139 20181 42148
rect 19755 42104 19797 42113
rect 19755 42064 19756 42104
rect 19796 42064 19797 42104
rect 19755 42055 19797 42064
rect 20140 42054 20180 42139
rect 19948 42020 19988 42029
rect 19755 41768 19797 41777
rect 19755 41728 19756 41768
rect 19796 41728 19797 41768
rect 19755 41719 19797 41728
rect 19756 41634 19796 41719
rect 19948 41609 19988 41980
rect 19947 41600 19989 41609
rect 19947 41560 19948 41600
rect 19988 41560 19989 41600
rect 19947 41551 19989 41560
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 19660 41476 19796 41516
rect 19756 41432 19796 41476
rect 19756 41383 19796 41392
rect 20235 41432 20277 41441
rect 20235 41392 20236 41432
rect 20276 41392 20277 41432
rect 20235 41383 20277 41392
rect 20236 41298 20276 41383
rect 19563 41264 19605 41273
rect 19563 41224 19564 41264
rect 19604 41224 19605 41264
rect 19852 41264 19892 41273
rect 19563 41215 19605 41224
rect 19660 41250 19700 41259
rect 19564 41130 19604 41215
rect 19660 41021 19700 41210
rect 19659 41012 19701 41021
rect 19659 40972 19660 41012
rect 19700 40972 19796 41012
rect 19659 40963 19701 40972
rect 19372 40552 19508 40592
rect 18892 40300 19316 40340
rect 19179 40172 19221 40181
rect 19179 40132 19180 40172
rect 19220 40132 19221 40172
rect 19179 40123 19221 40132
rect 19180 39752 19220 40123
rect 18604 39668 18644 39677
rect 18507 39080 18549 39089
rect 18507 39040 18508 39080
rect 18548 39040 18549 39080
rect 18507 39031 18549 39040
rect 18411 38912 18453 38921
rect 18411 38872 18412 38912
rect 18452 38872 18453 38912
rect 18411 38863 18453 38872
rect 18508 38912 18548 38921
rect 18412 38778 18452 38863
rect 18508 38669 18548 38872
rect 18604 38837 18644 39628
rect 18700 39668 18740 39677
rect 18603 38828 18645 38837
rect 18603 38788 18604 38828
rect 18644 38788 18645 38828
rect 18603 38779 18645 38788
rect 18315 38660 18357 38669
rect 18315 38620 18316 38660
rect 18356 38620 18357 38660
rect 18315 38611 18357 38620
rect 18507 38660 18549 38669
rect 18507 38620 18508 38660
rect 18548 38620 18549 38660
rect 18507 38611 18549 38620
rect 18316 38408 18356 38611
rect 18700 38585 18740 39628
rect 19180 39509 19220 39712
rect 19179 39500 19221 39509
rect 19179 39460 19180 39500
rect 19220 39460 19221 39500
rect 19179 39451 19221 39460
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19083 39164 19125 39173
rect 19083 39124 19084 39164
rect 19124 39124 19125 39164
rect 19083 39115 19125 39124
rect 18795 38912 18837 38921
rect 18795 38872 18796 38912
rect 18836 38872 18837 38912
rect 18795 38863 18837 38872
rect 18892 38912 18932 38923
rect 18699 38576 18741 38585
rect 18699 38536 18700 38576
rect 18740 38536 18741 38576
rect 18699 38527 18741 38536
rect 18700 38408 18740 38527
rect 18316 38368 18452 38408
rect 18315 38240 18357 38249
rect 18315 38200 18316 38240
rect 18356 38200 18357 38240
rect 18315 38191 18357 38200
rect 18316 37241 18356 38191
rect 18315 37232 18357 37241
rect 18315 37192 18316 37232
rect 18356 37192 18357 37232
rect 18315 37183 18357 37192
rect 18316 36728 18356 36737
rect 18316 36140 18356 36688
rect 18316 36091 18356 36100
rect 18412 36728 18452 38368
rect 18604 38368 18740 38408
rect 18796 38408 18836 38863
rect 18892 38837 18932 38872
rect 18987 38912 19029 38921
rect 18987 38872 18988 38912
rect 19028 38872 19029 38912
rect 18987 38863 19029 38872
rect 18891 38828 18933 38837
rect 18891 38788 18892 38828
rect 18932 38788 18933 38828
rect 18891 38779 18933 38788
rect 18988 38778 19028 38863
rect 18892 38408 18932 38417
rect 18796 38368 18892 38408
rect 18604 38249 18644 38368
rect 18892 38359 18932 38368
rect 18603 38240 18645 38249
rect 18603 38200 18604 38240
rect 18644 38200 18645 38240
rect 18603 38191 18645 38200
rect 18700 38240 18740 38249
rect 19084 38240 19124 39115
rect 18740 38200 19124 38240
rect 18700 37409 18740 38200
rect 19276 37913 19316 40300
rect 19372 38744 19412 40552
rect 19468 40424 19508 40435
rect 19756 40424 19796 40972
rect 19852 40760 19892 41224
rect 20043 41180 20085 41189
rect 20043 41140 20044 41180
rect 20084 41140 20085 41180
rect 20043 41131 20085 41140
rect 20044 41046 20084 41131
rect 19852 40720 20180 40760
rect 19948 40433 19988 40518
rect 19852 40424 19892 40433
rect 19756 40384 19852 40424
rect 19468 40349 19508 40384
rect 19852 40375 19892 40384
rect 19947 40424 19989 40433
rect 19947 40384 19948 40424
rect 19988 40384 19989 40424
rect 19947 40375 19989 40384
rect 20044 40424 20084 40433
rect 19467 40340 19509 40349
rect 19467 40300 19468 40340
rect 19508 40300 19509 40340
rect 19467 40291 19509 40300
rect 19468 39173 19508 40291
rect 19660 40256 19700 40265
rect 20044 40256 20084 40384
rect 20140 40424 20180 40720
rect 20140 40375 20180 40384
rect 19660 39747 19700 40216
rect 19660 39698 19700 39707
rect 19756 40216 20084 40256
rect 20523 40256 20565 40265
rect 20523 40216 20524 40256
rect 20564 40216 20565 40256
rect 19467 39164 19509 39173
rect 19467 39124 19468 39164
rect 19508 39124 19509 39164
rect 19467 39115 19509 39124
rect 19756 39080 19796 40216
rect 20523 40207 20565 40216
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 19851 39920 19893 39929
rect 19851 39880 19852 39920
rect 19892 39880 19893 39920
rect 19851 39871 19893 39880
rect 19852 39786 19892 39871
rect 20139 39584 20181 39593
rect 20139 39544 20140 39584
rect 20180 39544 20181 39584
rect 20139 39535 20181 39544
rect 19660 39040 19796 39080
rect 19467 38996 19509 39005
rect 19467 38956 19468 38996
rect 19508 38956 19509 38996
rect 19467 38947 19509 38956
rect 19468 38912 19508 38947
rect 19468 38861 19508 38872
rect 19372 38704 19508 38744
rect 19372 38156 19412 38165
rect 19372 37997 19412 38116
rect 19371 37988 19413 37997
rect 19371 37948 19372 37988
rect 19412 37948 19413 37988
rect 19371 37939 19413 37948
rect 19275 37904 19317 37913
rect 19275 37864 19276 37904
rect 19316 37864 19317 37904
rect 19275 37855 19317 37864
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 18219 35804 18261 35813
rect 18219 35764 18220 35804
rect 18260 35764 18261 35804
rect 18219 35755 18261 35764
rect 18123 35720 18165 35729
rect 18123 35680 18124 35720
rect 18164 35680 18165 35720
rect 18123 35671 18165 35680
rect 18124 35477 18164 35671
rect 18123 35468 18165 35477
rect 18123 35428 18124 35468
rect 18164 35428 18165 35468
rect 18123 35419 18165 35428
rect 17931 35300 17973 35309
rect 17931 35260 17932 35300
rect 17972 35260 17973 35300
rect 17931 35251 17973 35260
rect 17835 35132 17877 35141
rect 17835 35092 17836 35132
rect 17876 35092 17877 35132
rect 17835 35083 17877 35092
rect 18412 34544 18452 36688
rect 18508 37400 18548 37409
rect 18508 36569 18548 37360
rect 18699 37400 18741 37409
rect 18699 37360 18700 37400
rect 18740 37360 18741 37400
rect 18699 37351 18741 37360
rect 18891 37232 18933 37241
rect 18891 37192 18892 37232
rect 18932 37192 18933 37232
rect 18891 37183 18933 37192
rect 18892 36728 18932 37183
rect 18892 36679 18932 36688
rect 19371 36728 19413 36737
rect 19371 36688 19372 36728
rect 19412 36688 19413 36728
rect 19371 36679 19413 36688
rect 18796 36644 18836 36655
rect 18796 36569 18836 36604
rect 19372 36594 19412 36679
rect 18507 36560 18549 36569
rect 18507 36520 18508 36560
rect 18548 36520 18549 36560
rect 18507 36511 18549 36520
rect 18795 36560 18837 36569
rect 18795 36520 18796 36560
rect 18836 36520 18837 36560
rect 18795 36511 18837 36520
rect 19468 36317 19508 38704
rect 19563 38408 19605 38417
rect 19563 38368 19564 38408
rect 19604 38368 19605 38408
rect 19563 38359 19605 38368
rect 19564 38274 19604 38359
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 19467 36308 19509 36317
rect 19467 36268 19468 36308
rect 19508 36268 19509 36308
rect 19467 36259 19509 36268
rect 18508 35888 18548 35899
rect 18508 35813 18548 35848
rect 18507 35804 18549 35813
rect 18507 35764 18508 35804
rect 18548 35764 18549 35804
rect 18507 35755 18549 35764
rect 18507 35216 18549 35225
rect 18507 35176 18508 35216
rect 18548 35176 18549 35216
rect 18507 35167 18549 35176
rect 18508 35082 18548 35167
rect 18700 34964 18740 34973
rect 17836 34504 18068 34544
rect 17739 34376 17781 34385
rect 17739 34336 17740 34376
rect 17780 34336 17781 34376
rect 17739 34327 17781 34336
rect 17836 34376 17876 34504
rect 17836 34327 17876 34336
rect 17932 34376 17972 34385
rect 17643 34040 17685 34049
rect 17643 34000 17644 34040
rect 17684 34000 17685 34040
rect 17643 33991 17685 34000
rect 17644 33797 17684 33991
rect 17643 33788 17685 33797
rect 17643 33748 17644 33788
rect 17684 33748 17685 33788
rect 17643 33739 17685 33748
rect 17644 33452 17684 33739
rect 17740 33704 17780 34327
rect 17932 34049 17972 34336
rect 17931 34040 17973 34049
rect 17931 34000 17932 34040
rect 17972 34000 17973 34040
rect 17931 33991 17973 34000
rect 18028 33872 18068 34504
rect 18028 33823 18068 33832
rect 18124 34504 18452 34544
rect 18508 34924 18700 34964
rect 17836 33704 17876 33713
rect 17740 33664 17836 33704
rect 17876 33664 17972 33704
rect 17836 33655 17876 33664
rect 17644 33412 17876 33452
rect 17740 32192 17780 32201
rect 17740 31688 17780 32152
rect 17836 32192 17876 33412
rect 17932 33125 17972 33664
rect 17931 33116 17973 33125
rect 17931 33076 17932 33116
rect 17972 33076 17973 33116
rect 17931 33067 17973 33076
rect 17931 32864 17973 32873
rect 17931 32824 17932 32864
rect 17972 32824 17973 32864
rect 17931 32815 17973 32824
rect 17932 32730 17972 32815
rect 17836 32143 17876 32152
rect 18124 31940 18164 34504
rect 18316 34376 18356 34385
rect 18316 33536 18356 34336
rect 18412 34376 18452 34385
rect 18412 34049 18452 34336
rect 18411 34040 18453 34049
rect 18411 34000 18412 34040
rect 18452 34000 18453 34040
rect 18411 33991 18453 34000
rect 18508 33704 18548 34924
rect 18700 34915 18740 34924
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18892 34376 18932 34385
rect 18699 34040 18741 34049
rect 18699 34000 18700 34040
rect 18740 34000 18741 34040
rect 18699 33991 18741 34000
rect 18508 33655 18548 33664
rect 18604 33704 18644 33713
rect 18604 33536 18644 33664
rect 18316 33496 18644 33536
rect 18604 32276 18644 33496
rect 18220 32236 18644 32276
rect 18700 33620 18740 33991
rect 18892 33797 18932 34336
rect 19372 34381 19412 34390
rect 19660 34385 19700 39040
rect 19948 38917 19988 38926
rect 19948 38408 19988 38877
rect 20140 38828 20180 39535
rect 20140 38779 20180 38788
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 19852 38368 19988 38408
rect 19755 38156 19797 38165
rect 19755 38116 19756 38156
rect 19796 38116 19797 38156
rect 19755 38107 19797 38116
rect 19756 38022 19796 38107
rect 19852 37652 19892 38368
rect 19947 38072 19989 38081
rect 19947 38032 19948 38072
rect 19988 38032 19989 38072
rect 19947 38023 19989 38032
rect 19948 37938 19988 38023
rect 19948 37652 19988 37661
rect 19852 37612 19948 37652
rect 19948 37603 19988 37612
rect 19755 37400 19797 37409
rect 19755 37360 19756 37400
rect 19796 37360 19797 37400
rect 19755 37351 19797 37360
rect 19756 36056 19796 37351
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 20044 36812 20084 36821
rect 19852 36714 19892 36723
rect 19852 36140 19892 36674
rect 19948 36140 19988 36149
rect 19852 36100 19948 36140
rect 19948 36091 19988 36100
rect 19756 36016 19892 36056
rect 19756 35888 19796 35899
rect 19756 35813 19796 35848
rect 19755 35804 19797 35813
rect 19755 35764 19756 35804
rect 19796 35764 19797 35804
rect 19755 35755 19797 35764
rect 19852 35636 19892 36016
rect 20044 35720 20084 36772
rect 19756 35596 19892 35636
rect 19948 35680 20084 35720
rect 19756 35225 19796 35596
rect 19851 35300 19893 35309
rect 19851 35260 19852 35300
rect 19892 35260 19893 35300
rect 19851 35251 19893 35260
rect 19755 35216 19797 35225
rect 19755 35176 19756 35216
rect 19796 35176 19797 35216
rect 19755 35167 19797 35176
rect 18891 33788 18933 33797
rect 18891 33748 18892 33788
rect 18932 33748 18933 33788
rect 18891 33739 18933 33748
rect 18988 33620 19028 33629
rect 18700 33580 18988 33620
rect 18220 32192 18260 32236
rect 18220 32143 18260 32152
rect 18315 32108 18357 32117
rect 18315 32068 18316 32108
rect 18356 32068 18357 32108
rect 18315 32059 18357 32068
rect 18316 31974 18356 32059
rect 18124 31900 18260 31940
rect 17740 31648 18164 31688
rect 18124 31604 18164 31648
rect 18124 31555 18164 31564
rect 17451 31436 17493 31445
rect 17451 31396 17452 31436
rect 17492 31396 17493 31436
rect 17451 31387 17493 31396
rect 17931 31352 17973 31361
rect 17931 31312 17932 31352
rect 17972 31312 17973 31352
rect 17931 31303 17973 31312
rect 18123 31352 18165 31361
rect 18123 31312 18124 31352
rect 18164 31312 18165 31352
rect 18123 31303 18165 31312
rect 17932 31218 17972 31303
rect 17451 30764 17493 30773
rect 17451 30724 17452 30764
rect 17492 30724 17493 30764
rect 17451 30715 17493 30724
rect 17452 30092 17492 30715
rect 18124 30680 18164 31303
rect 18124 30631 18164 30640
rect 18220 30512 18260 31900
rect 18412 31352 18452 31361
rect 18316 30848 18356 30857
rect 18412 30848 18452 31312
rect 18508 31352 18548 32236
rect 18603 32108 18645 32117
rect 18700 32108 18740 33580
rect 18988 33571 19028 33580
rect 19084 33620 19124 33631
rect 19084 33545 19124 33580
rect 19083 33536 19125 33545
rect 19083 33496 19084 33536
rect 19124 33496 19125 33536
rect 19083 33487 19125 33496
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 19179 33116 19221 33125
rect 19179 33076 19180 33116
rect 19220 33076 19221 33116
rect 19179 33067 19221 33076
rect 19372 33116 19412 34341
rect 19659 34376 19701 34385
rect 19659 34336 19660 34376
rect 19700 34336 19701 34376
rect 19659 34327 19701 34336
rect 19563 34292 19605 34301
rect 19563 34252 19564 34292
rect 19604 34252 19605 34292
rect 19563 34243 19605 34252
rect 19564 34158 19604 34243
rect 19467 33788 19509 33797
rect 19467 33748 19468 33788
rect 19508 33748 19509 33788
rect 19467 33739 19509 33748
rect 19372 33067 19412 33076
rect 19180 32864 19220 33067
rect 18795 32780 18837 32789
rect 18795 32740 18796 32780
rect 18836 32740 18837 32780
rect 18795 32731 18837 32740
rect 18796 32192 18836 32731
rect 19180 32276 19220 32824
rect 19468 32789 19508 33739
rect 19564 33704 19604 33715
rect 19564 33629 19604 33664
rect 19563 33620 19605 33629
rect 19563 33580 19564 33620
rect 19604 33580 19605 33620
rect 19563 33571 19605 33580
rect 19467 32780 19509 32789
rect 19467 32740 19468 32780
rect 19508 32740 19509 32780
rect 19467 32731 19509 32740
rect 19467 32276 19509 32285
rect 19180 32236 19412 32276
rect 18796 32143 18836 32152
rect 19276 32178 19316 32187
rect 18603 32068 18604 32108
rect 18644 32068 18740 32108
rect 18603 32059 18645 32068
rect 18508 31277 18548 31312
rect 18507 31268 18549 31277
rect 18507 31228 18508 31268
rect 18548 31228 18549 31268
rect 18507 31219 18549 31228
rect 18604 31268 18644 32059
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18987 31436 19029 31445
rect 18987 31396 18988 31436
rect 19028 31396 19029 31436
rect 18987 31387 19029 31396
rect 18892 31352 18932 31361
rect 18892 31268 18932 31312
rect 18988 31302 19028 31387
rect 18604 31228 18932 31268
rect 18356 30808 18452 30848
rect 18316 30799 18356 30808
rect 17452 30043 17492 30052
rect 18124 30472 18260 30512
rect 17740 29840 17780 29849
rect 17548 29800 17740 29840
rect 17452 29336 17492 29345
rect 17548 29336 17588 29800
rect 17740 29791 17780 29800
rect 17836 29840 17876 29849
rect 17876 29800 18068 29840
rect 17836 29791 17876 29800
rect 17835 29672 17877 29681
rect 17835 29632 17836 29672
rect 17876 29632 17877 29672
rect 17835 29623 17877 29632
rect 17492 29296 17588 29336
rect 17452 29287 17492 29296
rect 17643 29252 17685 29261
rect 17643 29212 17644 29252
rect 17684 29212 17685 29252
rect 17643 29203 17685 29212
rect 17547 29084 17589 29093
rect 17547 29044 17548 29084
rect 17588 29044 17589 29084
rect 17547 29035 17589 29044
rect 17356 28960 17492 29000
rect 17259 28916 17301 28925
rect 17259 28876 17260 28916
rect 17300 28876 17301 28916
rect 17259 28867 17301 28876
rect 17355 27488 17397 27497
rect 17355 27448 17356 27488
rect 17396 27448 17397 27488
rect 17355 27439 17397 27448
rect 17259 26984 17301 26993
rect 17259 26944 17260 26984
rect 17300 26944 17301 26984
rect 17259 26935 17301 26944
rect 17260 26816 17300 26935
rect 17260 26767 17300 26776
rect 17356 26816 17396 27439
rect 17356 26153 17396 26776
rect 17355 26144 17397 26153
rect 17355 26104 17356 26144
rect 17396 26104 17397 26144
rect 17355 26095 17397 26104
rect 17163 23960 17205 23969
rect 17163 23920 17164 23960
rect 17204 23920 17205 23960
rect 17163 23911 17205 23920
rect 17164 23792 17204 23801
rect 17068 23752 17164 23771
rect 17068 23731 17204 23752
rect 17259 23792 17301 23801
rect 17259 23752 17260 23792
rect 17300 23752 17301 23792
rect 17259 23743 17301 23752
rect 16875 23204 16917 23213
rect 16875 23164 16876 23204
rect 16916 23164 16917 23204
rect 16875 23155 16917 23164
rect 16684 23120 16724 23129
rect 16684 22877 16724 23080
rect 16876 23120 16916 23155
rect 16876 23070 16916 23080
rect 16971 23120 17013 23129
rect 16971 23080 16972 23120
rect 17012 23080 17013 23120
rect 16971 23071 17013 23080
rect 16972 22986 17012 23071
rect 16683 22868 16725 22877
rect 16683 22828 16684 22868
rect 16724 22828 16725 22868
rect 16683 22819 16725 22828
rect 16779 22700 16821 22709
rect 16779 22660 16780 22700
rect 16820 22660 16821 22700
rect 16779 22651 16821 22660
rect 16587 22532 16629 22541
rect 16587 22492 16588 22532
rect 16628 22492 16629 22532
rect 16587 22483 16629 22492
rect 16588 22280 16628 22483
rect 16588 22231 16628 22240
rect 16780 22280 16820 22651
rect 16780 22231 16820 22240
rect 16684 21608 16724 21617
rect 16299 21356 16341 21365
rect 16299 21316 16300 21356
rect 16340 21316 16341 21356
rect 16299 21307 16341 21316
rect 16300 20768 16340 21307
rect 16300 20719 16340 20728
rect 16395 20768 16437 20777
rect 16395 20728 16396 20768
rect 16436 20728 16437 20768
rect 16395 20719 16437 20728
rect 16492 20768 16532 20777
rect 16396 20096 16436 20719
rect 16492 20264 16532 20728
rect 16684 20693 16724 21568
rect 17068 21533 17108 23731
rect 17260 23624 17300 23743
rect 17356 23717 17396 26095
rect 17452 23876 17492 28960
rect 17548 24137 17588 29035
rect 17547 24128 17589 24137
rect 17547 24088 17548 24128
rect 17588 24088 17589 24128
rect 17547 24079 17589 24088
rect 17644 23885 17684 29203
rect 17739 29084 17781 29093
rect 17739 29044 17740 29084
rect 17780 29044 17781 29084
rect 17739 29035 17781 29044
rect 17740 26909 17780 29035
rect 17836 28337 17876 29623
rect 17931 29168 17973 29177
rect 17931 29128 17932 29168
rect 17972 29128 17973 29168
rect 17931 29119 17973 29128
rect 18028 29168 18068 29800
rect 18124 29681 18164 30472
rect 18220 29840 18260 29849
rect 18123 29672 18165 29681
rect 18123 29632 18124 29672
rect 18164 29632 18165 29672
rect 18123 29623 18165 29632
rect 18220 29588 18260 29800
rect 18316 29840 18356 29849
rect 18356 29800 18548 29840
rect 18316 29791 18356 29800
rect 18220 29548 18356 29588
rect 18219 29420 18261 29429
rect 18219 29380 18220 29420
rect 18260 29380 18261 29420
rect 18219 29371 18261 29380
rect 18068 29128 18164 29168
rect 18028 29119 18068 29128
rect 17932 29034 17972 29119
rect 18027 28916 18069 28925
rect 18027 28876 18028 28916
rect 18068 28876 18069 28916
rect 18027 28867 18069 28876
rect 17931 28664 17973 28673
rect 17931 28624 17932 28664
rect 17972 28624 17973 28664
rect 17931 28615 17973 28624
rect 17835 28328 17877 28337
rect 17835 28288 17836 28328
rect 17876 28288 17877 28328
rect 17835 28279 17877 28288
rect 17836 27917 17876 28279
rect 17932 28085 17972 28615
rect 18028 28328 18068 28867
rect 17931 28076 17973 28085
rect 17931 28036 17932 28076
rect 17972 28036 17973 28076
rect 17931 28027 17973 28036
rect 17835 27908 17877 27917
rect 17835 27868 17836 27908
rect 17876 27868 17877 27908
rect 17835 27859 17877 27868
rect 17931 27740 17973 27749
rect 17931 27700 17932 27740
rect 17972 27700 17973 27740
rect 17931 27691 17973 27700
rect 17739 26900 17781 26909
rect 17739 26860 17740 26900
rect 17780 26860 17781 26900
rect 17739 26851 17781 26860
rect 17740 26766 17780 26851
rect 17836 26816 17876 26825
rect 17836 26564 17876 26776
rect 17740 26524 17876 26564
rect 17740 26405 17780 26524
rect 17932 26480 17972 27691
rect 18028 27665 18068 28288
rect 18027 27656 18069 27665
rect 18027 27616 18028 27656
rect 18068 27616 18069 27656
rect 18027 27607 18069 27616
rect 17836 26440 17972 26480
rect 17739 26396 17781 26405
rect 17739 26356 17740 26396
rect 17780 26356 17781 26396
rect 17739 26347 17781 26356
rect 17740 26144 17780 26153
rect 17740 25985 17780 26104
rect 17739 25976 17781 25985
rect 17739 25936 17740 25976
rect 17780 25936 17781 25976
rect 17739 25927 17781 25936
rect 17739 24548 17781 24557
rect 17739 24508 17740 24548
rect 17780 24508 17781 24548
rect 17739 24499 17781 24508
rect 17643 23876 17685 23885
rect 17452 23836 17588 23876
rect 17355 23708 17397 23717
rect 17355 23668 17356 23708
rect 17396 23668 17397 23708
rect 17355 23659 17397 23668
rect 17164 23584 17300 23624
rect 17164 23120 17204 23584
rect 17259 23456 17301 23465
rect 17259 23416 17260 23456
rect 17300 23416 17301 23456
rect 17259 23407 17301 23416
rect 17164 23071 17204 23080
rect 17260 23120 17300 23407
rect 17451 23372 17493 23381
rect 17451 23332 17452 23372
rect 17492 23332 17493 23372
rect 17451 23323 17493 23332
rect 17355 23288 17397 23297
rect 17355 23248 17356 23288
rect 17396 23248 17397 23288
rect 17355 23239 17397 23248
rect 17452 23288 17492 23323
rect 17260 23071 17300 23080
rect 17356 23120 17396 23239
rect 17452 23237 17492 23248
rect 17356 23071 17396 23080
rect 17451 23120 17493 23129
rect 17451 23080 17452 23120
rect 17492 23080 17493 23120
rect 17451 23071 17493 23080
rect 17067 21524 17109 21533
rect 17067 21484 17068 21524
rect 17108 21484 17109 21524
rect 17067 21475 17109 21484
rect 16780 20768 16820 20777
rect 16683 20684 16725 20693
rect 16683 20644 16684 20684
rect 16724 20644 16725 20684
rect 16683 20635 16725 20644
rect 16588 20600 16628 20609
rect 16588 20441 16628 20560
rect 16587 20432 16629 20441
rect 16587 20392 16588 20432
rect 16628 20392 16629 20432
rect 16587 20383 16629 20392
rect 16492 20224 16724 20264
rect 16588 20096 16628 20105
rect 16396 20056 16588 20096
rect 16300 19844 16340 19853
rect 16396 19844 16436 20056
rect 16588 20047 16628 20056
rect 16340 19804 16436 19844
rect 16300 19181 16340 19804
rect 16491 19424 16533 19433
rect 16491 19384 16492 19424
rect 16532 19384 16533 19424
rect 16396 19349 16436 19380
rect 16491 19375 16533 19384
rect 16395 19340 16437 19349
rect 16395 19300 16396 19340
rect 16436 19300 16437 19340
rect 16395 19291 16437 19300
rect 16396 19256 16436 19291
rect 16299 19172 16341 19181
rect 16299 19132 16300 19172
rect 16340 19132 16341 19172
rect 16299 19123 16341 19132
rect 16299 18584 16341 18593
rect 16299 18544 16300 18584
rect 16340 18544 16341 18584
rect 16299 18535 16341 18544
rect 16300 18005 16340 18535
rect 16299 17996 16341 18005
rect 16299 17956 16300 17996
rect 16340 17956 16341 17996
rect 16299 17947 16341 17956
rect 16203 17828 16245 17837
rect 16203 17788 16204 17828
rect 16244 17788 16245 17828
rect 16203 17779 16245 17788
rect 16396 17240 16436 19216
rect 16492 19256 16532 19375
rect 16684 19340 16724 20224
rect 16780 19508 16820 20728
rect 16875 20768 16917 20777
rect 16875 20728 16876 20768
rect 16916 20728 16917 20768
rect 16875 20719 16917 20728
rect 17068 20768 17108 20777
rect 16876 20634 16916 20719
rect 16971 20600 17013 20609
rect 16971 20560 16972 20600
rect 17012 20560 17013 20600
rect 16971 20551 17013 20560
rect 16972 20466 17012 20551
rect 17068 20357 17108 20728
rect 17259 20600 17301 20609
rect 17259 20560 17260 20600
rect 17300 20560 17301 20600
rect 17259 20551 17301 20560
rect 16875 20348 16917 20357
rect 16875 20308 16876 20348
rect 16916 20308 16917 20348
rect 16875 20299 16917 20308
rect 17067 20348 17109 20357
rect 17067 20308 17068 20348
rect 17108 20308 17109 20348
rect 17067 20299 17109 20308
rect 16876 20096 16916 20299
rect 16971 20180 17013 20189
rect 16971 20140 16972 20180
rect 17012 20140 17013 20180
rect 16971 20131 17013 20140
rect 16876 20047 16916 20056
rect 16972 20046 17012 20131
rect 17260 20096 17300 20551
rect 17355 20348 17397 20357
rect 17355 20308 17356 20348
rect 17396 20308 17397 20348
rect 17355 20299 17397 20308
rect 17164 20056 17300 20096
rect 16971 19928 17013 19937
rect 16971 19888 16972 19928
rect 17012 19888 17013 19928
rect 16971 19879 17013 19888
rect 16780 19459 16820 19468
rect 16492 19207 16532 19216
rect 16588 19300 16724 19340
rect 16492 18752 16532 18761
rect 16588 18752 16628 19300
rect 16972 19256 17012 19879
rect 17164 19349 17204 20056
rect 17259 19928 17301 19937
rect 17259 19888 17260 19928
rect 17300 19888 17301 19928
rect 17259 19879 17301 19888
rect 17260 19794 17300 19879
rect 17163 19340 17205 19349
rect 17163 19300 17164 19340
rect 17204 19300 17205 19340
rect 17163 19291 17205 19300
rect 16972 19207 17012 19216
rect 16683 19172 16725 19181
rect 16683 19132 16684 19172
rect 16724 19132 16725 19172
rect 16683 19123 16725 19132
rect 16532 18712 16628 18752
rect 16492 18703 16532 18712
rect 16588 18593 16628 18712
rect 16587 18584 16629 18593
rect 16587 18544 16588 18584
rect 16628 18544 16629 18584
rect 16587 18535 16629 18544
rect 16684 18584 16724 19123
rect 17163 19088 17205 19097
rect 17163 19048 17164 19088
rect 17204 19048 17205 19088
rect 17163 19039 17205 19048
rect 16779 18836 16821 18845
rect 16779 18796 16780 18836
rect 16820 18796 16821 18836
rect 16779 18787 16821 18796
rect 16684 18535 16724 18544
rect 16780 18584 16820 18787
rect 16876 18593 16916 18678
rect 17164 18605 17204 19039
rect 17356 18752 17396 20299
rect 17452 20273 17492 23071
rect 17548 20609 17588 23836
rect 17643 23836 17644 23876
rect 17684 23836 17685 23876
rect 17643 23827 17685 23836
rect 17643 23624 17685 23633
rect 17643 23584 17644 23624
rect 17684 23584 17685 23624
rect 17643 23575 17685 23584
rect 17644 23120 17684 23575
rect 17740 23288 17780 24499
rect 17740 23239 17780 23248
rect 17644 23071 17684 23080
rect 17643 20768 17685 20777
rect 17643 20728 17644 20768
rect 17684 20728 17685 20768
rect 17643 20719 17685 20728
rect 17547 20600 17589 20609
rect 17547 20560 17548 20600
rect 17588 20560 17589 20600
rect 17547 20551 17589 20560
rect 17451 20264 17493 20273
rect 17451 20224 17452 20264
rect 17492 20224 17493 20264
rect 17451 20215 17493 20224
rect 17452 20096 17492 20105
rect 17644 20096 17684 20719
rect 17492 20056 17588 20096
rect 17452 20047 17492 20056
rect 17451 19844 17493 19853
rect 17451 19804 17452 19844
rect 17492 19804 17493 19844
rect 17451 19795 17493 19804
rect 17452 19710 17492 19795
rect 17452 18752 17492 18761
rect 17356 18712 17452 18752
rect 17452 18703 17492 18712
rect 16683 17996 16725 18005
rect 16683 17956 16684 17996
rect 16724 17956 16725 17996
rect 16683 17947 16725 17956
rect 16684 17837 16724 17947
rect 16683 17828 16725 17837
rect 16683 17788 16684 17828
rect 16724 17788 16725 17828
rect 16780 17828 16820 18544
rect 16875 18584 16917 18593
rect 16875 18544 16876 18584
rect 16916 18544 16917 18584
rect 16875 18535 16917 18544
rect 16972 18584 17012 18593
rect 17164 18556 17204 18565
rect 17260 18584 17300 18593
rect 16972 18500 17012 18544
rect 17260 18500 17300 18544
rect 16972 18460 17300 18500
rect 17356 18584 17396 18593
rect 17548 18584 17588 20056
rect 17644 18752 17684 20056
rect 17740 20096 17780 20105
rect 17740 19937 17780 20056
rect 17739 19928 17781 19937
rect 17739 19888 17740 19928
rect 17780 19888 17781 19928
rect 17739 19879 17781 19888
rect 17740 18752 17780 18761
rect 17644 18712 17740 18752
rect 17740 18703 17780 18712
rect 17396 18544 17588 18584
rect 17643 18584 17685 18593
rect 17643 18544 17644 18584
rect 17684 18544 17685 18584
rect 17356 18416 17396 18544
rect 17643 18535 17685 18544
rect 17644 18450 17684 18535
rect 16876 18376 17396 18416
rect 17451 18416 17493 18425
rect 17451 18376 17452 18416
rect 17492 18376 17493 18416
rect 16876 17996 16916 18376
rect 17451 18367 17493 18376
rect 16876 17947 16916 17956
rect 16780 17788 16916 17828
rect 16683 17779 16725 17788
rect 16684 17744 16724 17779
rect 16684 17694 16724 17704
rect 16779 17660 16821 17669
rect 16779 17620 16780 17660
rect 16820 17620 16821 17660
rect 16779 17611 16821 17620
rect 16396 17200 16532 17240
rect 16395 17072 16437 17081
rect 16395 17032 16396 17072
rect 16436 17032 16437 17072
rect 16395 17023 16437 17032
rect 16011 16064 16053 16073
rect 16011 16024 16012 16064
rect 16052 16024 16053 16064
rect 16011 16015 16053 16024
rect 16108 15821 16148 16192
rect 16299 16064 16341 16073
rect 16299 16024 16300 16064
rect 16340 16024 16341 16064
rect 16299 16015 16341 16024
rect 16203 15980 16245 15989
rect 16203 15940 16204 15980
rect 16244 15940 16245 15980
rect 16203 15931 16245 15940
rect 16107 15812 16149 15821
rect 16107 15772 16108 15812
rect 16148 15772 16149 15812
rect 16107 15763 16149 15772
rect 16011 15728 16053 15737
rect 16011 15688 16012 15728
rect 16052 15688 16053 15728
rect 16011 15679 16053 15688
rect 15916 15560 15956 15569
rect 16012 15560 16052 15679
rect 16108 15644 16148 15653
rect 16108 15560 16148 15604
rect 16012 15520 16148 15560
rect 15916 15476 15956 15520
rect 15916 15436 16052 15476
rect 15820 15352 15956 15392
rect 15723 15140 15765 15149
rect 15723 15100 15724 15140
rect 15764 15100 15765 15140
rect 15723 15091 15765 15100
rect 15148 14167 15188 14176
rect 15244 14260 15380 14300
rect 15436 14848 15668 14888
rect 14572 13994 14764 14034
rect 14572 13460 14612 13994
rect 14764 13985 14804 13994
rect 14860 13994 15092 14034
rect 14667 13880 14709 13889
rect 14667 13840 14668 13880
rect 14708 13840 14709 13880
rect 14667 13831 14709 13840
rect 14572 13411 14612 13420
rect 14571 12536 14613 12545
rect 14571 12496 14572 12536
rect 14612 12496 14613 12536
rect 14571 12487 14613 12496
rect 14228 12412 14516 12452
rect 14188 12403 14228 12412
rect 14092 12244 14228 12284
rect 13900 12160 14036 12200
rect 13900 11696 13940 11705
rect 13707 11444 13749 11453
rect 13707 11404 13708 11444
rect 13748 11404 13749 11444
rect 13707 11395 13749 11404
rect 13035 10688 13077 10697
rect 13035 10648 13036 10688
rect 13076 10648 13077 10688
rect 13035 10639 13077 10648
rect 13036 10184 13076 10193
rect 13132 10184 13172 10816
rect 13227 10688 13269 10697
rect 13227 10648 13228 10688
rect 13268 10648 13269 10688
rect 13227 10639 13269 10648
rect 13076 10144 13172 10184
rect 13036 10135 13076 10144
rect 12940 9976 13076 10016
rect 12843 9512 12885 9521
rect 12843 9472 12844 9512
rect 12884 9472 12885 9512
rect 12843 9463 12885 9472
rect 12651 8840 12693 8849
rect 12651 8800 12652 8840
rect 12692 8800 12693 8840
rect 12651 8791 12693 8800
rect 12172 5657 12212 6448
rect 12268 7960 12460 8000
rect 12500 7960 12596 8000
rect 12171 5648 12213 5657
rect 12171 5608 12172 5648
rect 12212 5608 12213 5648
rect 12171 5599 12213 5608
rect 12268 5648 12308 7960
rect 12460 7951 12500 7960
rect 12459 7496 12501 7505
rect 12459 7456 12460 7496
rect 12500 7456 12501 7496
rect 12459 7447 12501 7456
rect 12363 6404 12405 6413
rect 12363 6364 12364 6404
rect 12404 6364 12405 6404
rect 12363 6355 12405 6364
rect 12268 5396 12308 5608
rect 12172 5356 12308 5396
rect 12075 5144 12117 5153
rect 12075 5104 12076 5144
rect 12116 5104 12117 5144
rect 12075 5095 12117 5104
rect 12075 4976 12117 4985
rect 12075 4936 12076 4976
rect 12116 4936 12117 4976
rect 12075 4927 12117 4936
rect 12076 4842 12116 4927
rect 11595 4808 11637 4817
rect 11595 4768 11596 4808
rect 11636 4768 11637 4808
rect 11595 4759 11637 4768
rect 12172 4733 12212 5356
rect 12268 5069 12308 5154
rect 12267 5060 12309 5069
rect 12267 5020 12268 5060
rect 12308 5020 12309 5060
rect 12267 5011 12309 5020
rect 12364 4892 12404 6355
rect 12268 4852 12404 4892
rect 12171 4724 12213 4733
rect 12171 4684 12172 4724
rect 12212 4684 12213 4724
rect 12171 4675 12213 4684
rect 11883 4304 11925 4313
rect 11883 4264 11884 4304
rect 11924 4264 11925 4304
rect 11883 4255 11925 4264
rect 11596 4220 11636 4229
rect 11500 4180 11596 4220
rect 11596 4171 11636 4180
rect 11307 4136 11349 4145
rect 11307 4096 11308 4136
rect 11348 4096 11349 4136
rect 11307 4087 11349 4096
rect 11884 4136 11924 4255
rect 11884 4087 11924 4096
rect 11403 3968 11445 3977
rect 11403 3928 11404 3968
rect 11444 3928 11445 3968
rect 11403 3919 11445 3928
rect 11979 3968 12021 3977
rect 11979 3928 11980 3968
rect 12020 3928 12021 3968
rect 11979 3919 12021 3928
rect 11404 3834 11444 3919
rect 11883 3548 11925 3557
rect 11116 3508 11444 3548
rect 11019 3296 11061 3305
rect 11019 3256 11020 3296
rect 11060 3256 11061 3296
rect 11019 3247 11061 3256
rect 10732 3212 10772 3221
rect 10732 2633 10772 3172
rect 11116 3212 11156 3221
rect 11308 3212 11348 3221
rect 11116 2885 11156 3172
rect 11212 3172 11308 3212
rect 10827 2876 10869 2885
rect 10827 2836 10828 2876
rect 10868 2836 10869 2876
rect 10827 2827 10869 2836
rect 11115 2876 11157 2885
rect 11115 2836 11116 2876
rect 11156 2836 11157 2876
rect 11115 2827 11157 2836
rect 10731 2624 10773 2633
rect 10731 2584 10732 2624
rect 10772 2584 10773 2624
rect 10731 2575 10773 2584
rect 10635 2036 10677 2045
rect 10635 1996 10636 2036
rect 10676 1996 10677 2036
rect 10635 1987 10677 1996
rect 10828 1784 10868 2827
rect 11115 2372 11157 2381
rect 11115 2332 11116 2372
rect 11156 2332 11157 2372
rect 11115 2323 11157 2332
rect 11116 2213 11156 2323
rect 11115 2204 11157 2213
rect 11115 2164 11116 2204
rect 11156 2164 11157 2204
rect 11115 2155 11157 2164
rect 11116 1952 11156 2155
rect 11116 1903 11156 1912
rect 10732 1744 10868 1784
rect 10635 1448 10677 1457
rect 10635 1408 10636 1448
rect 10676 1408 10677 1448
rect 10635 1399 10677 1408
rect 10636 1112 10676 1399
rect 10636 1063 10676 1072
rect 10732 944 10772 1744
rect 11212 1196 11252 3172
rect 11308 3163 11348 3172
rect 11308 2624 11348 2633
rect 11308 2381 11348 2584
rect 11307 2372 11349 2381
rect 11307 2332 11308 2372
rect 11348 2332 11349 2372
rect 11307 2323 11349 2332
rect 11307 2120 11349 2129
rect 11307 2080 11308 2120
rect 11348 2080 11349 2120
rect 11307 2071 11349 2080
rect 11308 1986 11348 2071
rect 10444 652 10580 692
rect 10636 904 10772 944
rect 11020 1156 11252 1196
rect 10347 608 10389 617
rect 10347 568 10348 608
rect 10388 568 10389 608
rect 10347 559 10389 568
rect 10444 80 10484 652
rect 10636 80 10676 904
rect 11020 608 11060 1156
rect 11211 1028 11253 1037
rect 11211 988 11212 1028
rect 11252 988 11253 1028
rect 11211 979 11253 988
rect 10828 568 11060 608
rect 10828 80 10868 568
rect 11019 272 11061 281
rect 11019 232 11020 272
rect 11060 232 11061 272
rect 11019 223 11061 232
rect 11020 80 11060 223
rect 11212 80 11252 979
rect 11404 80 11444 3508
rect 11883 3508 11884 3548
rect 11924 3508 11925 3548
rect 11883 3499 11925 3508
rect 11788 3464 11828 3473
rect 11787 3459 11788 3464
rect 11692 3424 11788 3459
rect 11692 3419 11828 3424
rect 11499 3380 11541 3389
rect 11499 3340 11500 3380
rect 11540 3340 11541 3380
rect 11499 3331 11541 3340
rect 11500 3246 11540 3331
rect 11500 2876 11540 2885
rect 11692 2876 11732 3419
rect 11788 3415 11828 3419
rect 11884 3464 11924 3499
rect 11540 2836 11732 2876
rect 11500 2827 11540 2836
rect 11691 2624 11733 2633
rect 11691 2584 11692 2624
rect 11732 2584 11733 2624
rect 11691 2575 11733 2584
rect 11788 2624 11828 2633
rect 11595 2204 11637 2213
rect 11595 2164 11596 2204
rect 11636 2164 11637 2204
rect 11595 2155 11637 2164
rect 11500 1952 11540 1961
rect 11500 1793 11540 1912
rect 11499 1784 11541 1793
rect 11499 1744 11500 1784
rect 11540 1744 11541 1784
rect 11499 1735 11541 1744
rect 11500 1373 11540 1735
rect 11499 1364 11541 1373
rect 11499 1324 11500 1364
rect 11540 1324 11541 1364
rect 11499 1315 11541 1324
rect 11596 80 11636 2155
rect 11692 1616 11732 2575
rect 11788 2129 11828 2584
rect 11884 2624 11924 3424
rect 11884 2575 11924 2584
rect 11787 2120 11829 2129
rect 11787 2080 11788 2120
rect 11828 2080 11829 2120
rect 11787 2071 11829 2080
rect 11980 1961 12020 3919
rect 12268 3548 12308 4852
rect 12076 3508 12308 3548
rect 11979 1952 12021 1961
rect 11979 1912 11980 1952
rect 12020 1912 12021 1952
rect 11979 1903 12021 1912
rect 11979 1700 12021 1709
rect 11979 1660 11980 1700
rect 12020 1660 12021 1700
rect 11979 1651 12021 1660
rect 11692 1576 11828 1616
rect 11788 80 11828 1576
rect 11883 1196 11925 1205
rect 11883 1156 11884 1196
rect 11924 1156 11925 1196
rect 11883 1147 11925 1156
rect 11884 1112 11924 1147
rect 11884 869 11924 1072
rect 11883 860 11925 869
rect 11883 820 11884 860
rect 11924 820 11925 860
rect 11883 811 11925 820
rect 11980 80 12020 1651
rect 12076 1280 12116 3508
rect 12364 3464 12404 3473
rect 12460 3464 12500 7447
rect 12555 7076 12597 7085
rect 12555 7036 12556 7076
rect 12596 7036 12597 7076
rect 12555 7027 12597 7036
rect 12556 6497 12596 7027
rect 12555 6488 12597 6497
rect 12555 6448 12556 6488
rect 12596 6448 12597 6488
rect 12555 6439 12597 6448
rect 12652 6488 12692 8791
rect 12940 8765 12980 8796
rect 12939 8756 12981 8765
rect 12939 8716 12940 8756
rect 12980 8716 12981 8756
rect 12939 8707 12981 8716
rect 12843 8672 12885 8681
rect 12843 8632 12844 8672
rect 12884 8632 12885 8672
rect 12843 8623 12885 8632
rect 12940 8672 12980 8707
rect 12844 7841 12884 8623
rect 12940 8429 12980 8632
rect 12939 8420 12981 8429
rect 12939 8380 12940 8420
rect 12980 8380 12981 8420
rect 12939 8371 12981 8380
rect 13036 8261 13076 9976
rect 13035 8252 13077 8261
rect 13035 8212 13036 8252
rect 13076 8212 13077 8252
rect 13035 8203 13077 8212
rect 12843 7832 12885 7841
rect 12843 7792 12844 7832
rect 12884 7792 12885 7832
rect 12843 7783 12885 7792
rect 12844 7160 12884 7169
rect 12844 6917 12884 7120
rect 12843 6908 12885 6917
rect 12843 6868 12844 6908
rect 12884 6868 12885 6908
rect 12843 6859 12885 6868
rect 12652 6439 12692 6448
rect 12556 6354 12596 6439
rect 12651 6152 12693 6161
rect 12651 6112 12652 6152
rect 12692 6112 12693 6152
rect 12651 6103 12693 6112
rect 12556 4976 12596 4985
rect 12556 4817 12596 4936
rect 12555 4808 12597 4817
rect 12555 4768 12556 4808
rect 12596 4768 12597 4808
rect 12555 4759 12597 4768
rect 12556 3893 12596 4759
rect 12555 3884 12597 3893
rect 12555 3844 12556 3884
rect 12596 3844 12597 3884
rect 12555 3835 12597 3844
rect 12404 3424 12500 3464
rect 12268 3380 12308 3389
rect 12171 2876 12213 2885
rect 12171 2836 12172 2876
rect 12212 2836 12213 2876
rect 12171 2827 12213 2836
rect 12076 1231 12116 1240
rect 12172 80 12212 2827
rect 12268 2801 12308 3340
rect 12267 2792 12309 2801
rect 12267 2752 12268 2792
rect 12308 2752 12309 2792
rect 12267 2743 12309 2752
rect 12268 2708 12308 2743
rect 12268 2657 12308 2668
rect 12364 2708 12404 3424
rect 12364 2659 12404 2668
rect 12267 2372 12309 2381
rect 12267 2332 12268 2372
rect 12308 2332 12309 2372
rect 12267 2323 12309 2332
rect 12268 1961 12308 2323
rect 12267 1952 12309 1961
rect 12267 1912 12268 1952
rect 12308 1912 12309 1952
rect 12267 1903 12309 1912
rect 12268 1112 12308 1903
rect 12363 1280 12405 1289
rect 12363 1240 12364 1280
rect 12404 1240 12405 1280
rect 12363 1231 12405 1240
rect 12268 1063 12308 1072
rect 12364 80 12404 1231
rect 12652 1205 12692 6103
rect 12747 4388 12789 4397
rect 12747 4348 12748 4388
rect 12788 4348 12789 4388
rect 12747 4339 12789 4348
rect 12748 1961 12788 4339
rect 12844 3464 12884 3473
rect 12844 3137 12884 3424
rect 12843 3128 12885 3137
rect 12843 3088 12844 3128
rect 12884 3088 12885 3128
rect 12843 3079 12885 3088
rect 12844 2624 12884 3079
rect 12844 2575 12884 2584
rect 12939 2624 12981 2633
rect 12939 2584 12940 2624
rect 12980 2584 12981 2624
rect 12939 2575 12981 2584
rect 12940 2120 12980 2575
rect 13036 2381 13076 8203
rect 13132 6917 13172 10144
rect 13131 6908 13173 6917
rect 13131 6868 13132 6908
rect 13172 6868 13173 6908
rect 13131 6859 13173 6868
rect 13228 6497 13268 10639
rect 13419 10268 13461 10277
rect 13419 10228 13420 10268
rect 13460 10228 13461 10268
rect 13419 10219 13461 10228
rect 13323 9512 13365 9521
rect 13323 9472 13324 9512
rect 13364 9472 13365 9512
rect 13323 9463 13365 9472
rect 13132 6488 13172 6497
rect 13132 6329 13172 6448
rect 13227 6488 13269 6497
rect 13227 6448 13228 6488
rect 13268 6448 13269 6488
rect 13227 6439 13269 6448
rect 13131 6320 13173 6329
rect 13131 6280 13132 6320
rect 13172 6280 13173 6320
rect 13131 6271 13173 6280
rect 13324 6161 13364 9463
rect 13420 8840 13460 10219
rect 13515 10100 13557 10109
rect 13515 10060 13516 10100
rect 13556 10060 13557 10100
rect 13515 10051 13557 10060
rect 13516 9680 13556 10051
rect 13516 9631 13556 9640
rect 13420 8800 13556 8840
rect 13419 8672 13461 8681
rect 13419 8632 13420 8672
rect 13460 8632 13461 8672
rect 13419 8623 13461 8632
rect 13420 8538 13460 8623
rect 13516 6656 13556 8800
rect 13612 7505 13652 10984
rect 13900 10277 13940 11656
rect 13899 10268 13941 10277
rect 13899 10228 13900 10268
rect 13940 10228 13941 10268
rect 13899 10219 13941 10228
rect 13708 9428 13748 9437
rect 13708 8597 13748 9388
rect 13900 8677 13940 8686
rect 13707 8588 13749 8597
rect 13707 8548 13708 8588
rect 13748 8548 13749 8588
rect 13707 8539 13749 8548
rect 13900 8168 13940 8637
rect 13900 8119 13940 8128
rect 13707 8000 13749 8009
rect 13707 7960 13708 8000
rect 13748 7960 13749 8000
rect 13707 7951 13749 7960
rect 13611 7496 13653 7505
rect 13611 7456 13612 7496
rect 13652 7456 13653 7496
rect 13611 7447 13653 7456
rect 13420 6616 13556 6656
rect 13323 6152 13365 6161
rect 13323 6112 13324 6152
rect 13364 6112 13365 6152
rect 13323 6103 13365 6112
rect 13227 4892 13269 4901
rect 13227 4852 13228 4892
rect 13268 4852 13269 4892
rect 13227 4843 13269 4852
rect 13131 4388 13173 4397
rect 13131 4348 13132 4388
rect 13172 4348 13173 4388
rect 13131 4339 13173 4348
rect 13132 4136 13172 4339
rect 13132 4087 13172 4096
rect 13131 3632 13173 3641
rect 13131 3592 13132 3632
rect 13172 3592 13173 3632
rect 13131 3583 13173 3592
rect 13132 3305 13172 3583
rect 13131 3296 13173 3305
rect 13131 3256 13132 3296
rect 13172 3256 13173 3296
rect 13131 3247 13173 3256
rect 13131 2876 13173 2885
rect 13131 2836 13132 2876
rect 13172 2836 13173 2876
rect 13131 2827 13173 2836
rect 13035 2372 13077 2381
rect 13035 2332 13036 2372
rect 13076 2332 13077 2372
rect 13035 2323 13077 2332
rect 12940 2071 12980 2080
rect 12747 1952 12789 1961
rect 12747 1912 12748 1952
rect 12788 1912 12789 1952
rect 12747 1903 12789 1912
rect 13132 1952 13172 2827
rect 13228 2036 13268 4843
rect 13324 3968 13364 3977
rect 13324 3459 13364 3928
rect 13324 3410 13364 3419
rect 13324 2629 13364 2638
rect 13324 2465 13364 2589
rect 13420 2540 13460 6616
rect 13515 6488 13557 6497
rect 13515 6448 13516 6488
rect 13556 6448 13557 6488
rect 13708 6488 13748 7951
rect 13803 7916 13845 7925
rect 13803 7876 13804 7916
rect 13844 7876 13845 7916
rect 13803 7867 13845 7876
rect 13804 6656 13844 7867
rect 13996 6992 14036 12160
rect 14092 11528 14132 11537
rect 14092 11019 14132 11488
rect 14092 10970 14132 10979
rect 14091 8588 14133 8597
rect 14091 8548 14092 8588
rect 14132 8548 14133 8588
rect 14091 8539 14133 8548
rect 14092 8454 14132 8539
rect 14188 8261 14228 12244
rect 14572 12041 14612 12487
rect 14571 12032 14613 12041
rect 14571 11992 14572 12032
rect 14612 11992 14613 12032
rect 14571 11983 14613 11992
rect 14668 11864 14708 13831
rect 14763 12872 14805 12881
rect 14763 12832 14764 12872
rect 14804 12832 14805 12872
rect 14763 12823 14805 12832
rect 14764 12125 14804 12823
rect 14763 12116 14805 12125
rect 14763 12076 14764 12116
rect 14804 12076 14805 12116
rect 14763 12067 14805 12076
rect 14380 11824 14708 11864
rect 14283 11528 14325 11537
rect 14283 11488 14284 11528
rect 14324 11488 14325 11528
rect 14283 11479 14325 11488
rect 14284 11192 14324 11479
rect 14284 11143 14324 11152
rect 14283 10268 14325 10277
rect 14283 10228 14284 10268
rect 14324 10228 14325 10268
rect 14283 10219 14325 10228
rect 14284 10184 14324 10219
rect 14284 10109 14324 10144
rect 14283 10100 14325 10109
rect 14283 10060 14284 10100
rect 14324 10060 14325 10100
rect 14283 10051 14325 10060
rect 14284 10020 14324 10051
rect 14380 9848 14420 11824
rect 14572 11696 14612 11705
rect 14475 11528 14517 11537
rect 14475 11488 14476 11528
rect 14516 11488 14517 11528
rect 14475 11479 14517 11488
rect 14476 11201 14516 11479
rect 14475 11192 14517 11201
rect 14475 11152 14476 11192
rect 14516 11152 14517 11192
rect 14475 11143 14517 11152
rect 14475 10856 14517 10865
rect 14475 10816 14476 10856
rect 14516 10816 14517 10856
rect 14475 10807 14517 10816
rect 14476 10722 14516 10807
rect 14476 10436 14516 10445
rect 14572 10436 14612 11656
rect 14668 11696 14708 11824
rect 14668 11647 14708 11656
rect 14667 11192 14709 11201
rect 14667 11152 14668 11192
rect 14708 11152 14709 11192
rect 14667 11143 14709 11152
rect 14668 10940 14708 11143
rect 14668 10891 14708 10900
rect 14516 10396 14612 10436
rect 14476 10387 14516 10396
rect 14763 10268 14805 10277
rect 14763 10228 14764 10268
rect 14804 10228 14805 10268
rect 14763 10219 14805 10228
rect 14284 9808 14420 9848
rect 14764 10184 14804 10219
rect 14187 8252 14229 8261
rect 14187 8212 14188 8252
rect 14228 8212 14229 8252
rect 14187 8203 14229 8212
rect 14284 8177 14324 9808
rect 14379 9680 14421 9689
rect 14379 9640 14380 9680
rect 14420 9640 14421 9680
rect 14379 9631 14421 9640
rect 14380 9512 14420 9631
rect 14380 9463 14420 9472
rect 14764 8681 14804 10144
rect 14860 9185 14900 13994
rect 15244 13880 15284 14260
rect 15339 14048 15381 14057
rect 15339 14008 15340 14048
rect 15380 14008 15381 14048
rect 15339 13999 15381 14008
rect 15052 13840 15284 13880
rect 15052 11873 15092 13840
rect 15340 13796 15380 13999
rect 15244 13756 15380 13796
rect 15147 13544 15189 13553
rect 15147 13504 15148 13544
rect 15188 13504 15189 13544
rect 15147 13495 15189 13504
rect 15051 11864 15093 11873
rect 15051 11824 15052 11864
rect 15092 11824 15093 11864
rect 15051 11815 15093 11824
rect 15052 11780 15092 11815
rect 15052 11730 15092 11740
rect 15148 11696 15188 13495
rect 15244 13217 15284 13756
rect 15436 13712 15476 14848
rect 15628 14804 15668 14848
rect 15628 14755 15668 14764
rect 15724 14804 15764 15091
rect 15627 14636 15669 14645
rect 15627 14596 15628 14636
rect 15668 14596 15669 14636
rect 15627 14587 15669 14596
rect 15340 13672 15476 13712
rect 15243 13208 15285 13217
rect 15243 13168 15244 13208
rect 15284 13168 15285 13208
rect 15243 13159 15285 13168
rect 15243 11780 15285 11789
rect 15243 11740 15244 11780
rect 15284 11740 15285 11780
rect 15243 11731 15285 11740
rect 14955 10016 14997 10025
rect 14955 9976 14956 10016
rect 14996 9976 14997 10016
rect 14955 9967 14997 9976
rect 14859 9176 14901 9185
rect 14859 9136 14860 9176
rect 14900 9136 14901 9176
rect 14859 9127 14901 9136
rect 14763 8672 14805 8681
rect 14763 8632 14764 8672
rect 14804 8632 14805 8672
rect 14763 8623 14805 8632
rect 14283 8168 14325 8177
rect 14283 8128 14284 8168
rect 14324 8128 14325 8168
rect 14283 8119 14325 8128
rect 14091 8000 14133 8009
rect 14091 7960 14092 8000
rect 14132 7960 14133 8000
rect 14091 7951 14133 7960
rect 14092 7866 14132 7951
rect 14187 7580 14229 7589
rect 14187 7540 14188 7580
rect 14228 7540 14229 7580
rect 14187 7531 14229 7540
rect 13804 6607 13844 6616
rect 13900 6952 14036 6992
rect 14092 7160 14132 7169
rect 13515 6439 13557 6448
rect 13612 6474 13652 6483
rect 13516 5648 13556 6439
rect 13708 6448 13844 6488
rect 13612 5900 13652 6434
rect 13708 5900 13748 5909
rect 13612 5860 13708 5900
rect 13708 5851 13748 5860
rect 13516 4985 13556 5608
rect 13804 4985 13844 6448
rect 13515 4976 13557 4985
rect 13515 4936 13516 4976
rect 13556 4936 13557 4976
rect 13515 4927 13557 4936
rect 13803 4976 13845 4985
rect 13803 4936 13804 4976
rect 13844 4936 13845 4976
rect 13803 4927 13845 4936
rect 13516 4397 13556 4927
rect 13804 4842 13844 4927
rect 13515 4388 13557 4397
rect 13515 4348 13516 4388
rect 13556 4348 13557 4388
rect 13515 4339 13557 4348
rect 13515 4220 13557 4229
rect 13515 4180 13516 4220
rect 13556 4180 13557 4220
rect 13515 4171 13557 4180
rect 13516 3632 13556 4171
rect 13707 4136 13749 4145
rect 13707 4096 13708 4136
rect 13748 4096 13749 4136
rect 13707 4087 13749 4096
rect 13708 4002 13748 4087
rect 13516 3583 13556 3592
rect 13707 3380 13749 3389
rect 13900 3380 13940 6952
rect 14092 6497 14132 7120
rect 14091 6488 14133 6497
rect 14091 6448 14092 6488
rect 14132 6448 14133 6488
rect 14091 6439 14133 6448
rect 13996 5648 14036 5657
rect 13996 5144 14036 5608
rect 14091 5648 14133 5657
rect 14091 5608 14092 5648
rect 14132 5608 14133 5648
rect 14091 5599 14133 5608
rect 13996 5095 14036 5104
rect 14092 3557 14132 5599
rect 14188 5405 14228 7531
rect 14667 7496 14709 7505
rect 14667 7456 14668 7496
rect 14708 7456 14709 7496
rect 14667 7447 14709 7456
rect 14572 7160 14612 7171
rect 14572 7085 14612 7120
rect 14668 7160 14708 7447
rect 14764 7421 14804 8623
rect 14860 8504 14900 8513
rect 14860 7589 14900 8464
rect 14859 7580 14901 7589
rect 14859 7540 14860 7580
rect 14900 7540 14901 7580
rect 14859 7531 14901 7540
rect 14763 7412 14805 7421
rect 14763 7372 14764 7412
rect 14804 7372 14805 7412
rect 14763 7363 14805 7372
rect 14956 7244 14996 9967
rect 15052 8677 15092 8686
rect 15052 8177 15092 8637
rect 15051 8168 15093 8177
rect 15051 8128 15052 8168
rect 15092 8128 15093 8168
rect 15051 8119 15093 8128
rect 15148 7832 15188 11656
rect 15244 8597 15284 11731
rect 15243 8588 15285 8597
rect 15243 8548 15244 8588
rect 15284 8548 15285 8588
rect 15243 8539 15285 8548
rect 15340 8345 15380 13672
rect 15628 13628 15668 14587
rect 15436 13588 15668 13628
rect 15436 8765 15476 13588
rect 15724 13469 15764 14764
rect 15531 13460 15573 13469
rect 15531 13420 15532 13460
rect 15572 13420 15573 13460
rect 15531 13411 15573 13420
rect 15723 13460 15765 13469
rect 15723 13420 15724 13460
rect 15764 13420 15765 13460
rect 15723 13411 15765 13420
rect 15532 8840 15572 13411
rect 15723 13292 15765 13301
rect 15723 13252 15724 13292
rect 15764 13252 15765 13292
rect 15723 13243 15765 13252
rect 15627 11780 15669 11789
rect 15627 11740 15628 11780
rect 15668 11740 15669 11780
rect 15627 11731 15669 11740
rect 15628 11696 15668 11731
rect 15628 11645 15668 11656
rect 15724 11360 15764 13243
rect 15819 13208 15861 13217
rect 15819 13168 15820 13208
rect 15860 13168 15861 13208
rect 15819 13159 15861 13168
rect 15820 12713 15860 13159
rect 15819 12704 15861 12713
rect 15819 12664 15820 12704
rect 15860 12664 15861 12704
rect 15819 12655 15861 12664
rect 15820 12536 15860 12655
rect 15820 12487 15860 12496
rect 15628 11320 15764 11360
rect 15628 9521 15668 11320
rect 15724 11024 15764 11033
rect 15724 9680 15764 10984
rect 15819 11024 15861 11033
rect 15819 10984 15820 11024
rect 15860 10984 15861 11024
rect 15819 10975 15861 10984
rect 15820 10890 15860 10975
rect 15916 10529 15956 15352
rect 16012 15317 16052 15436
rect 16204 15401 16244 15931
rect 16300 15569 16340 16015
rect 16299 15560 16341 15569
rect 16299 15520 16300 15560
rect 16340 15520 16341 15560
rect 16299 15511 16341 15520
rect 16203 15392 16245 15401
rect 16203 15352 16204 15392
rect 16244 15352 16245 15392
rect 16203 15343 16245 15352
rect 16011 15308 16053 15317
rect 16011 15268 16012 15308
rect 16052 15268 16053 15308
rect 16011 15259 16053 15268
rect 16299 15308 16341 15317
rect 16299 15268 16300 15308
rect 16340 15268 16341 15308
rect 16299 15259 16341 15268
rect 16012 14057 16052 15259
rect 16300 15174 16340 15259
rect 16203 14972 16245 14981
rect 16203 14932 16204 14972
rect 16244 14932 16245 14972
rect 16203 14923 16245 14932
rect 16204 14720 16244 14923
rect 16204 14671 16244 14680
rect 16011 14048 16053 14057
rect 16011 14008 16012 14048
rect 16052 14008 16053 14048
rect 16011 13999 16053 14008
rect 16203 13460 16245 13469
rect 16203 13420 16204 13460
rect 16244 13420 16245 13460
rect 16203 13411 16245 13420
rect 16012 13208 16052 13217
rect 16012 12704 16052 13168
rect 16107 13208 16149 13217
rect 16107 13168 16108 13208
rect 16148 13168 16149 13208
rect 16107 13159 16149 13168
rect 16108 13074 16148 13159
rect 16012 12655 16052 12664
rect 16204 12536 16244 13411
rect 16300 12545 16340 12630
rect 16012 12496 16244 12536
rect 16299 12536 16341 12545
rect 16299 12496 16300 12536
rect 16340 12496 16341 12536
rect 15915 10520 15957 10529
rect 15915 10480 15916 10520
rect 15956 10480 15957 10520
rect 15915 10471 15957 10480
rect 16012 10352 16052 12496
rect 16299 12487 16341 12496
rect 16299 12368 16341 12377
rect 16299 12328 16300 12368
rect 16340 12328 16341 12368
rect 16299 12319 16341 12328
rect 16108 11701 16148 11710
rect 16108 10436 16148 11661
rect 16300 11612 16340 12319
rect 16300 11563 16340 11572
rect 16396 11360 16436 17023
rect 16492 16073 16532 17200
rect 16587 16232 16629 16241
rect 16587 16192 16588 16232
rect 16628 16192 16629 16232
rect 16587 16183 16629 16192
rect 16588 16098 16628 16183
rect 16491 16064 16533 16073
rect 16491 16024 16492 16064
rect 16532 16024 16533 16064
rect 16491 16015 16533 16024
rect 16587 15728 16629 15737
rect 16587 15688 16588 15728
rect 16628 15688 16629 15728
rect 16587 15679 16629 15688
rect 16491 15644 16533 15653
rect 16491 15604 16492 15644
rect 16532 15604 16533 15644
rect 16491 15595 16533 15604
rect 16492 15560 16532 15595
rect 16492 15509 16532 15520
rect 16491 15392 16533 15401
rect 16491 15352 16492 15392
rect 16532 15352 16533 15392
rect 16491 15343 16533 15352
rect 16492 14048 16532 15343
rect 16588 14813 16628 15679
rect 16683 15308 16725 15317
rect 16683 15268 16684 15308
rect 16724 15268 16725 15308
rect 16683 15259 16725 15268
rect 16587 14804 16629 14813
rect 16587 14764 16588 14804
rect 16628 14764 16629 14804
rect 16587 14755 16629 14764
rect 16588 14216 16628 14755
rect 16684 14734 16724 15259
rect 16684 14685 16724 14694
rect 16588 14176 16724 14216
rect 16587 14048 16629 14057
rect 16492 14008 16588 14048
rect 16628 14008 16629 14048
rect 16587 13999 16629 14008
rect 16588 13914 16628 13999
rect 16491 13880 16533 13889
rect 16491 13840 16492 13880
rect 16532 13840 16533 13880
rect 16491 13831 16533 13840
rect 16492 13301 16532 13831
rect 16587 13460 16629 13469
rect 16587 13420 16588 13460
rect 16628 13420 16629 13460
rect 16587 13411 16629 13420
rect 16491 13292 16533 13301
rect 16491 13252 16492 13292
rect 16532 13252 16533 13292
rect 16491 13243 16533 13252
rect 16588 13292 16628 13411
rect 16588 13243 16628 13252
rect 16492 13158 16532 13243
rect 16684 13040 16724 14176
rect 16588 13000 16724 13040
rect 16396 11320 16532 11360
rect 16299 11192 16341 11201
rect 16299 11152 16300 11192
rect 16340 11152 16341 11192
rect 16299 11143 16341 11152
rect 16300 11024 16340 11143
rect 16300 10975 16340 10984
rect 16203 10940 16245 10949
rect 16203 10900 16204 10940
rect 16244 10900 16245 10940
rect 16203 10891 16245 10900
rect 16204 10806 16244 10891
rect 16204 10436 16244 10445
rect 16108 10396 16204 10436
rect 16204 10387 16244 10396
rect 15916 10312 16052 10352
rect 15820 9680 15860 9689
rect 15724 9640 15820 9680
rect 15820 9631 15860 9640
rect 15627 9512 15669 9521
rect 15627 9472 15628 9512
rect 15668 9472 15669 9512
rect 15627 9463 15669 9472
rect 15628 9378 15668 9463
rect 15532 8800 15668 8840
rect 15435 8756 15477 8765
rect 15435 8716 15436 8756
rect 15476 8716 15477 8756
rect 15435 8707 15477 8716
rect 15532 8672 15572 8683
rect 15532 8597 15572 8632
rect 15531 8588 15573 8597
rect 15531 8548 15532 8588
rect 15572 8548 15573 8588
rect 15531 8539 15573 8548
rect 15339 8336 15381 8345
rect 15339 8296 15340 8336
rect 15380 8296 15381 8336
rect 15339 8287 15381 8296
rect 15243 8252 15285 8261
rect 15243 8212 15244 8252
rect 15284 8212 15285 8252
rect 15243 8203 15285 8212
rect 15531 8252 15573 8261
rect 15531 8212 15532 8252
rect 15572 8212 15573 8252
rect 15531 8203 15573 8212
rect 15244 8084 15284 8203
rect 15532 8168 15572 8203
rect 15532 8117 15572 8128
rect 15244 8044 15380 8084
rect 15340 8000 15380 8044
rect 15340 7951 15380 7960
rect 15148 7792 15476 7832
rect 15243 7664 15285 7673
rect 15243 7624 15244 7664
rect 15284 7624 15285 7664
rect 15243 7615 15285 7624
rect 15052 7244 15092 7253
rect 14283 7076 14325 7085
rect 14283 7036 14284 7076
rect 14324 7036 14325 7076
rect 14283 7027 14325 7036
rect 14571 7076 14613 7085
rect 14571 7036 14572 7076
rect 14612 7036 14613 7076
rect 14571 7027 14613 7036
rect 14284 6942 14324 7027
rect 14379 6404 14421 6413
rect 14379 6364 14380 6404
rect 14420 6364 14421 6404
rect 14379 6355 14421 6364
rect 14187 5396 14229 5405
rect 14187 5356 14188 5396
rect 14228 5356 14229 5396
rect 14187 5347 14229 5356
rect 14284 4976 14324 4985
rect 14380 4976 14420 6355
rect 14475 5816 14517 5825
rect 14475 5776 14476 5816
rect 14516 5776 14517 5816
rect 14475 5767 14517 5776
rect 14476 5732 14516 5767
rect 14476 5681 14516 5692
rect 14571 5732 14613 5741
rect 14571 5692 14572 5732
rect 14612 5692 14613 5732
rect 14571 5683 14613 5692
rect 14572 5598 14612 5683
rect 14324 4936 14420 4976
rect 14284 4313 14324 4936
rect 14283 4304 14325 4313
rect 14283 4264 14284 4304
rect 14324 4264 14325 4304
rect 14283 4255 14325 4264
rect 14091 3548 14133 3557
rect 14091 3508 14092 3548
rect 14132 3508 14133 3548
rect 14091 3499 14133 3508
rect 13707 3340 13708 3380
rect 13748 3340 13749 3380
rect 13707 3331 13749 3340
rect 13804 3340 13940 3380
rect 14476 3464 14516 3473
rect 13611 2960 13653 2969
rect 13611 2920 13612 2960
rect 13652 2920 13653 2960
rect 13611 2911 13653 2920
rect 13516 2540 13556 2549
rect 13420 2500 13516 2540
rect 13516 2491 13556 2500
rect 13323 2456 13365 2465
rect 13323 2416 13324 2456
rect 13364 2416 13365 2456
rect 13323 2407 13365 2416
rect 13228 1996 13460 2036
rect 13132 1903 13172 1912
rect 12748 1818 12788 1903
rect 12747 1280 12789 1289
rect 12747 1240 12748 1280
rect 12788 1240 12789 1280
rect 12747 1231 12789 1240
rect 13323 1280 13365 1289
rect 13323 1240 13324 1280
rect 13364 1240 13365 1280
rect 13323 1231 13365 1240
rect 12651 1196 12693 1205
rect 12651 1156 12652 1196
rect 12692 1156 12693 1196
rect 12651 1147 12693 1156
rect 12555 944 12597 953
rect 12555 904 12556 944
rect 12596 904 12597 944
rect 12555 895 12597 904
rect 12556 80 12596 895
rect 12748 80 12788 1231
rect 13131 1196 13173 1205
rect 13131 1156 13132 1196
rect 13172 1156 13173 1196
rect 13131 1147 13173 1156
rect 12939 944 12981 953
rect 12939 904 12940 944
rect 12980 904 12981 944
rect 12939 895 12981 904
rect 12940 80 12980 895
rect 13132 80 13172 1147
rect 13324 80 13364 1231
rect 13420 1112 13460 1996
rect 13612 1280 13652 2911
rect 13708 2792 13748 3331
rect 13804 3044 13844 3340
rect 13900 3212 13940 3221
rect 13940 3172 14132 3212
rect 13900 3163 13940 3172
rect 13804 3004 13940 3044
rect 13708 2743 13748 2752
rect 13900 1373 13940 3004
rect 13996 2456 14036 2465
rect 13899 1364 13941 1373
rect 13899 1324 13900 1364
rect 13940 1324 13941 1364
rect 13899 1315 13941 1324
rect 13708 1280 13748 1289
rect 13612 1240 13708 1280
rect 13708 1231 13748 1240
rect 13899 1196 13941 1205
rect 13899 1156 13900 1196
rect 13940 1156 13941 1196
rect 13899 1147 13941 1156
rect 13516 1112 13556 1121
rect 13420 1072 13516 1112
rect 13516 1063 13556 1072
rect 13900 1112 13940 1147
rect 13996 1121 14036 2416
rect 13900 1061 13940 1072
rect 13995 1112 14037 1121
rect 13995 1072 13996 1112
rect 14036 1072 14037 1112
rect 13995 1063 14037 1072
rect 13899 944 13941 953
rect 13899 904 13900 944
rect 13940 904 13941 944
rect 13899 895 13941 904
rect 13515 860 13557 869
rect 13515 820 13516 860
rect 13556 820 13557 860
rect 13515 811 13557 820
rect 13516 80 13556 811
rect 13707 776 13749 785
rect 13707 736 13708 776
rect 13748 736 13749 776
rect 13707 727 13749 736
rect 13708 80 13748 727
rect 13900 80 13940 895
rect 14092 80 14132 3172
rect 14283 2876 14325 2885
rect 14283 2836 14284 2876
rect 14324 2836 14325 2876
rect 14283 2827 14325 2836
rect 14187 2708 14229 2717
rect 14187 2668 14188 2708
rect 14228 2668 14229 2708
rect 14187 2659 14229 2668
rect 14188 2574 14228 2659
rect 14187 2456 14229 2465
rect 14187 2416 14188 2456
rect 14228 2416 14229 2456
rect 14187 2407 14229 2416
rect 14188 533 14228 2407
rect 14284 1784 14324 2827
rect 14379 2456 14421 2465
rect 14379 2416 14380 2456
rect 14420 2416 14421 2456
rect 14379 2407 14421 2416
rect 14380 2322 14420 2407
rect 14476 2120 14516 3424
rect 14572 3464 14612 3473
rect 14668 3464 14708 7120
rect 14764 7204 15052 7244
rect 14764 5825 14804 7204
rect 15052 7195 15092 7204
rect 15148 7160 15188 7169
rect 15244 7160 15284 7615
rect 15339 7580 15381 7589
rect 15339 7540 15340 7580
rect 15380 7540 15381 7580
rect 15339 7531 15381 7540
rect 15188 7120 15284 7160
rect 15148 7111 15188 7120
rect 14859 7076 14901 7085
rect 15051 7076 15093 7085
rect 14859 7036 14860 7076
rect 14900 7036 14901 7076
rect 14859 7027 14901 7036
rect 14956 7036 15052 7076
rect 15092 7036 15093 7076
rect 14860 6581 14900 7027
rect 14859 6572 14901 6581
rect 14859 6532 14860 6572
rect 14900 6532 14901 6572
rect 14859 6523 14901 6532
rect 14860 6488 14900 6523
rect 14860 6438 14900 6448
rect 14763 5816 14805 5825
rect 14763 5776 14764 5816
rect 14804 5776 14900 5816
rect 14763 5767 14805 5776
rect 14612 3424 14708 3464
rect 14860 3464 14900 5776
rect 14956 4901 14996 7036
rect 15051 7027 15093 7036
rect 15051 5648 15093 5657
rect 15051 5608 15052 5648
rect 15092 5608 15093 5648
rect 15051 5599 15093 5608
rect 15052 5514 15092 5599
rect 14955 4892 14997 4901
rect 14955 4852 14956 4892
rect 14996 4852 14997 4892
rect 14955 4843 14997 4852
rect 14955 4136 14997 4145
rect 14955 4096 14956 4136
rect 14996 4096 14997 4136
rect 14955 4087 14997 4096
rect 14956 4002 14996 4087
rect 15148 3968 15188 3977
rect 15052 3473 15092 3558
rect 14956 3464 14996 3473
rect 14860 3424 14956 3464
rect 14572 3415 14612 3424
rect 14571 2708 14613 2717
rect 14571 2668 14572 2708
rect 14612 2668 14613 2708
rect 14571 2659 14613 2668
rect 14572 2574 14612 2659
rect 14668 2633 14708 3424
rect 14956 3415 14996 3424
rect 15051 3464 15093 3473
rect 15051 3424 15052 3464
rect 15092 3424 15093 3464
rect 15051 3415 15093 3424
rect 15051 3212 15093 3221
rect 15051 3172 15052 3212
rect 15092 3172 15093 3212
rect 15051 3163 15093 3172
rect 14667 2624 14709 2633
rect 14667 2584 14668 2624
rect 14708 2584 14709 2624
rect 14667 2575 14709 2584
rect 14572 2120 14612 2129
rect 14476 2080 14572 2120
rect 14572 2071 14612 2080
rect 14380 1961 14420 2046
rect 14379 1952 14421 1961
rect 14379 1912 14380 1952
rect 14420 1912 14421 1952
rect 14379 1903 14421 1912
rect 14763 1952 14805 1961
rect 14763 1912 14764 1952
rect 14804 1912 14805 1952
rect 14763 1903 14805 1912
rect 14764 1818 14804 1903
rect 14284 1744 14516 1784
rect 14283 944 14325 953
rect 14283 904 14284 944
rect 14324 904 14325 944
rect 14283 895 14325 904
rect 14187 524 14229 533
rect 14187 484 14188 524
rect 14228 484 14229 524
rect 14187 475 14229 484
rect 14284 80 14324 895
rect 14476 80 14516 1744
rect 14859 524 14901 533
rect 14859 484 14860 524
rect 14900 484 14901 524
rect 14859 475 14901 484
rect 14667 356 14709 365
rect 14667 316 14668 356
rect 14708 316 14709 356
rect 14667 307 14709 316
rect 14668 80 14708 307
rect 14860 80 14900 475
rect 15052 80 15092 3163
rect 15148 2624 15188 3928
rect 15244 3473 15284 7120
rect 15340 4136 15380 7531
rect 15436 6245 15476 7792
rect 15628 7160 15668 8800
rect 15916 8672 15956 10312
rect 16012 10184 16052 10193
rect 16012 10025 16052 10144
rect 16395 10184 16437 10193
rect 16395 10144 16396 10184
rect 16436 10144 16437 10184
rect 16395 10135 16437 10144
rect 16396 10050 16436 10135
rect 16011 10016 16053 10025
rect 16011 9976 16012 10016
rect 16052 9976 16053 10016
rect 16011 9967 16053 9976
rect 16203 10016 16245 10025
rect 16203 9976 16204 10016
rect 16244 9976 16245 10016
rect 16203 9967 16245 9976
rect 16107 8756 16149 8765
rect 16107 8716 16108 8756
rect 16148 8716 16149 8756
rect 16107 8707 16149 8716
rect 16012 8672 16052 8681
rect 15916 8632 16012 8672
rect 15819 8336 15861 8345
rect 15819 8296 15820 8336
rect 15860 8296 15861 8336
rect 15819 8287 15861 8296
rect 15723 8168 15765 8177
rect 15723 8128 15724 8168
rect 15764 8128 15765 8168
rect 15723 8119 15765 8128
rect 15724 8034 15764 8119
rect 15628 6329 15668 7120
rect 15627 6320 15669 6329
rect 15627 6280 15628 6320
rect 15668 6280 15669 6320
rect 15627 6271 15669 6280
rect 15435 6236 15477 6245
rect 15435 6196 15436 6236
rect 15476 6196 15477 6236
rect 15435 6187 15477 6196
rect 15580 5657 15620 5666
rect 15620 5617 15668 5648
rect 15580 5608 15668 5617
rect 15628 5144 15668 5608
rect 15820 5564 15860 8287
rect 16012 8177 16052 8632
rect 16011 8168 16053 8177
rect 16011 8128 16012 8168
rect 16052 8128 16053 8168
rect 16011 8119 16053 8128
rect 15916 8000 15956 8011
rect 15916 7925 15956 7960
rect 15915 7916 15957 7925
rect 15915 7876 15916 7916
rect 15956 7876 15957 7916
rect 15915 7867 15957 7876
rect 16108 7328 16148 8707
rect 16204 7925 16244 9967
rect 16492 9689 16532 11320
rect 16491 9680 16533 9689
rect 16491 9640 16492 9680
rect 16532 9640 16533 9680
rect 16491 9631 16533 9640
rect 16492 9512 16532 9521
rect 16492 9101 16532 9472
rect 16491 9092 16533 9101
rect 16491 9052 16492 9092
rect 16532 9052 16533 9092
rect 16491 9043 16533 9052
rect 16395 9008 16437 9017
rect 16395 8968 16396 9008
rect 16436 8968 16437 9008
rect 16395 8959 16437 8968
rect 16203 7916 16245 7925
rect 16203 7876 16204 7916
rect 16244 7876 16245 7916
rect 16203 7867 16245 7876
rect 16012 7288 16148 7328
rect 16012 5648 16052 7288
rect 16156 7169 16196 7178
rect 16196 7129 16244 7160
rect 16156 7120 16244 7129
rect 16204 6656 16244 7120
rect 16299 6992 16341 7001
rect 16299 6952 16300 6992
rect 16340 6952 16341 6992
rect 16299 6943 16341 6952
rect 16300 6858 16340 6943
rect 16396 6740 16436 8959
rect 16588 8840 16628 13000
rect 16780 11360 16820 17611
rect 16876 15653 16916 17788
rect 16972 17072 17012 17081
rect 16972 15821 17012 17032
rect 17355 17072 17397 17081
rect 17452 17072 17492 18367
rect 17547 18332 17589 18341
rect 17547 18292 17548 18332
rect 17588 18292 17589 18332
rect 17547 18283 17589 18292
rect 17355 17032 17356 17072
rect 17396 17032 17492 17072
rect 17355 17023 17397 17032
rect 17356 16938 17396 17023
rect 17164 16820 17204 16829
rect 17068 16780 17164 16820
rect 17068 16246 17108 16780
rect 17164 16771 17204 16780
rect 17259 16316 17301 16325
rect 17259 16276 17260 16316
rect 17300 16276 17301 16316
rect 17259 16267 17301 16276
rect 17068 16197 17108 16206
rect 17260 16148 17300 16267
rect 17260 16099 17300 16108
rect 17163 16064 17205 16073
rect 17163 16024 17164 16064
rect 17204 16024 17205 16064
rect 17163 16015 17205 16024
rect 17452 16064 17492 16073
rect 16971 15812 17013 15821
rect 16971 15772 16972 15812
rect 17012 15772 17013 15812
rect 16971 15763 17013 15772
rect 16875 15644 16917 15653
rect 16875 15604 16876 15644
rect 16916 15604 16917 15644
rect 16875 15595 16917 15604
rect 16971 15308 17013 15317
rect 16971 15268 16972 15308
rect 17012 15268 17013 15308
rect 16971 15259 17013 15268
rect 16875 14804 16917 14813
rect 16875 14764 16876 14804
rect 16916 14764 16917 14804
rect 16875 14755 16917 14764
rect 16876 14636 16916 14755
rect 16876 14587 16916 14596
rect 16972 14468 17012 15259
rect 17067 14552 17109 14561
rect 17067 14512 17068 14552
rect 17108 14512 17109 14552
rect 17067 14503 17109 14512
rect 16492 8800 16628 8840
rect 16684 11320 16820 11360
rect 16876 14428 17012 14468
rect 16492 8672 16532 8800
rect 16492 7505 16532 8632
rect 16588 8672 16628 8681
rect 16588 8261 16628 8632
rect 16587 8252 16629 8261
rect 16587 8212 16588 8252
rect 16628 8212 16629 8252
rect 16587 8203 16629 8212
rect 16491 7496 16533 7505
rect 16491 7456 16492 7496
rect 16532 7456 16533 7496
rect 16491 7447 16533 7456
rect 16587 7328 16629 7337
rect 16587 7288 16588 7328
rect 16628 7288 16629 7328
rect 16587 7279 16629 7288
rect 16588 7160 16628 7279
rect 16588 6917 16628 7120
rect 16587 6908 16629 6917
rect 16587 6868 16588 6908
rect 16628 6868 16629 6908
rect 16587 6859 16629 6868
rect 16396 6700 16628 6740
rect 16300 6656 16340 6665
rect 16204 6616 16300 6656
rect 16300 6607 16340 6616
rect 16492 6497 16532 6582
rect 16107 6488 16149 6497
rect 16107 6448 16108 6488
rect 16148 6448 16149 6488
rect 16107 6439 16149 6448
rect 16491 6488 16533 6497
rect 16491 6448 16492 6488
rect 16532 6448 16533 6488
rect 16491 6439 16533 6448
rect 16108 6354 16148 6439
rect 16203 6320 16245 6329
rect 16203 6280 16204 6320
rect 16244 6280 16245 6320
rect 16203 6271 16245 6280
rect 16491 6320 16533 6329
rect 16491 6280 16492 6320
rect 16532 6280 16533 6320
rect 16491 6271 16533 6280
rect 16012 5608 16148 5648
rect 15820 5524 16052 5564
rect 15724 5480 15764 5489
rect 15764 5440 15860 5480
rect 15724 5431 15764 5440
rect 15724 5144 15764 5153
rect 15628 5104 15724 5144
rect 15724 5095 15764 5104
rect 15531 4976 15573 4985
rect 15531 4936 15532 4976
rect 15572 4936 15573 4976
rect 15531 4927 15573 4936
rect 15723 4976 15765 4985
rect 15723 4936 15724 4976
rect 15764 4936 15765 4976
rect 15723 4927 15765 4936
rect 15532 4145 15572 4927
rect 15340 3893 15380 4096
rect 15531 4136 15573 4145
rect 15531 4096 15532 4136
rect 15572 4096 15573 4136
rect 15531 4087 15573 4096
rect 15724 3968 15764 4927
rect 15820 4061 15860 5440
rect 15916 4976 15956 4987
rect 15916 4901 15956 4936
rect 15915 4892 15957 4901
rect 15915 4852 15916 4892
rect 15956 4852 15957 4892
rect 15915 4843 15957 4852
rect 15819 4052 15861 4061
rect 15819 4012 15820 4052
rect 15860 4012 15861 4052
rect 15819 4003 15861 4012
rect 15532 3928 15764 3968
rect 15339 3884 15381 3893
rect 15339 3844 15340 3884
rect 15380 3844 15381 3884
rect 15339 3835 15381 3844
rect 15243 3464 15285 3473
rect 15243 3424 15244 3464
rect 15284 3424 15285 3464
rect 15243 3415 15285 3424
rect 15532 3464 15572 3928
rect 15819 3884 15861 3893
rect 15819 3844 15820 3884
rect 15860 3844 15861 3884
rect 15819 3835 15861 3844
rect 15627 3716 15669 3725
rect 15627 3676 15628 3716
rect 15668 3676 15669 3716
rect 15627 3667 15669 3676
rect 15532 3415 15572 3424
rect 15628 2801 15668 3667
rect 15723 3548 15765 3557
rect 15723 3508 15724 3548
rect 15764 3508 15765 3548
rect 15723 3499 15765 3508
rect 15627 2792 15669 2801
rect 15627 2752 15628 2792
rect 15668 2752 15669 2792
rect 15627 2743 15669 2752
rect 15244 2633 15284 2718
rect 15628 2708 15668 2743
rect 15628 2658 15668 2668
rect 15724 2708 15764 3499
rect 15724 2659 15764 2668
rect 15148 2575 15188 2584
rect 15243 2624 15285 2633
rect 15243 2584 15244 2624
rect 15284 2584 15285 2624
rect 15243 2575 15285 2584
rect 15147 2120 15189 2129
rect 15147 2080 15148 2120
rect 15188 2080 15189 2120
rect 15147 2071 15189 2080
rect 15148 1112 15188 2071
rect 15820 1961 15860 3835
rect 16012 3557 16052 5524
rect 16108 3725 16148 5608
rect 16204 5069 16244 6271
rect 16203 5060 16245 5069
rect 16203 5020 16204 5060
rect 16244 5020 16245 5060
rect 16203 5011 16245 5020
rect 16299 4976 16341 4985
rect 16299 4936 16300 4976
rect 16340 4936 16341 4976
rect 16299 4927 16341 4936
rect 16107 3716 16149 3725
rect 16107 3676 16108 3716
rect 16148 3676 16149 3716
rect 16107 3667 16149 3676
rect 16203 3632 16245 3641
rect 16203 3592 16204 3632
rect 16244 3592 16245 3632
rect 16203 3583 16245 3592
rect 16011 3548 16053 3557
rect 16011 3508 16012 3548
rect 16052 3508 16053 3548
rect 16011 3499 16053 3508
rect 16204 3498 16244 3583
rect 16060 3422 16100 3431
rect 16060 3380 16100 3382
rect 16060 3340 16148 3380
rect 16108 2120 16148 3340
rect 16203 3128 16245 3137
rect 16203 3088 16204 3128
rect 16244 3088 16245 3128
rect 16203 3079 16245 3088
rect 16204 2624 16244 3079
rect 16204 2575 16244 2584
rect 16204 2120 16244 2129
rect 16108 2080 16204 2120
rect 16204 2071 16244 2080
rect 15243 1952 15285 1961
rect 15243 1912 15244 1952
rect 15284 1912 15285 1952
rect 15243 1903 15285 1912
rect 15819 1952 15861 1961
rect 15819 1912 15820 1952
rect 15860 1912 15861 1952
rect 15819 1903 15861 1912
rect 16011 1952 16053 1961
rect 16011 1912 16012 1952
rect 16052 1912 16053 1952
rect 16011 1903 16053 1912
rect 15244 1373 15284 1903
rect 16012 1818 16052 1903
rect 16203 1700 16245 1709
rect 16203 1660 16204 1700
rect 16244 1660 16245 1700
rect 16203 1651 16245 1660
rect 15339 1616 15381 1625
rect 15339 1576 15340 1616
rect 15380 1576 15381 1616
rect 15339 1567 15381 1576
rect 15243 1364 15285 1373
rect 15243 1324 15244 1364
rect 15284 1324 15285 1364
rect 15243 1315 15285 1324
rect 15340 1280 15380 1567
rect 15435 1532 15477 1541
rect 15435 1492 15436 1532
rect 15476 1492 15477 1532
rect 15435 1483 15477 1492
rect 15340 1231 15380 1240
rect 15148 1063 15188 1072
rect 15243 272 15285 281
rect 15243 232 15244 272
rect 15284 232 15285 272
rect 15243 223 15285 232
rect 15244 80 15284 223
rect 15436 80 15476 1483
rect 15531 1112 15573 1121
rect 15531 1072 15532 1112
rect 15572 1072 15573 1112
rect 15531 1063 15573 1072
rect 15819 1112 15861 1121
rect 15819 1072 15820 1112
rect 15860 1072 15861 1112
rect 15819 1063 15861 1072
rect 15532 978 15572 1063
rect 15627 776 15669 785
rect 15627 736 15628 776
rect 15668 736 15669 776
rect 15627 727 15669 736
rect 15628 80 15668 727
rect 15820 80 15860 1063
rect 16011 860 16053 869
rect 16011 820 16012 860
rect 16052 820 16053 860
rect 16011 811 16053 820
rect 16012 80 16052 811
rect 16204 80 16244 1651
rect 16300 1121 16340 4927
rect 16395 3212 16437 3221
rect 16395 3172 16396 3212
rect 16436 3172 16437 3212
rect 16395 3163 16437 3172
rect 16396 3078 16436 3163
rect 16492 2540 16532 6271
rect 16588 5060 16628 6700
rect 16684 5573 16724 11320
rect 16779 11024 16821 11033
rect 16779 10984 16780 11024
rect 16820 10984 16821 11024
rect 16779 10975 16821 10984
rect 16780 10890 16820 10975
rect 16876 8840 16916 14428
rect 17068 14418 17108 14503
rect 16971 14048 17013 14057
rect 16971 14008 16972 14048
rect 17012 14008 17013 14048
rect 16971 13999 17013 14008
rect 16972 12956 17012 13999
rect 17068 13208 17108 13219
rect 17068 13133 17108 13168
rect 17067 13124 17109 13133
rect 17067 13084 17068 13124
rect 17108 13084 17109 13124
rect 17067 13075 17109 13084
rect 16972 12916 17108 12956
rect 16971 12536 17013 12545
rect 16971 12496 16972 12536
rect 17012 12496 17013 12536
rect 16971 12487 17013 12496
rect 16972 10193 17012 12487
rect 16971 10184 17013 10193
rect 16971 10144 16972 10184
rect 17012 10144 17013 10184
rect 16971 10135 17013 10144
rect 16780 8800 16916 8840
rect 16780 6329 16820 8800
rect 16875 8672 16917 8681
rect 16875 8632 16876 8672
rect 16916 8632 16917 8672
rect 16875 8623 16917 8632
rect 16876 8538 16916 8623
rect 17068 8009 17108 12916
rect 17164 11453 17204 16015
rect 17452 15905 17492 16024
rect 17451 15896 17493 15905
rect 17451 15856 17452 15896
rect 17492 15856 17493 15896
rect 17451 15847 17493 15856
rect 17451 15644 17493 15653
rect 17451 15604 17452 15644
rect 17492 15604 17493 15644
rect 17451 15595 17493 15604
rect 17259 14804 17301 14813
rect 17259 14764 17260 14804
rect 17300 14764 17301 14804
rect 17259 14755 17301 14764
rect 17260 14670 17300 14755
rect 17452 14216 17492 15595
rect 17548 15317 17588 18283
rect 17643 17996 17685 18005
rect 17643 17956 17644 17996
rect 17684 17956 17685 17996
rect 17643 17947 17685 17956
rect 17644 17862 17684 17947
rect 17740 17744 17780 17753
rect 17740 17249 17780 17704
rect 17836 17744 17876 26440
rect 17931 26312 17973 26321
rect 17931 26272 17932 26312
rect 17972 26272 17973 26312
rect 17931 26263 17973 26272
rect 17932 26178 17972 26263
rect 17932 25304 17972 25313
rect 18028 25304 18068 27607
rect 18124 27497 18164 29128
rect 18220 28580 18260 29371
rect 18316 29084 18356 29548
rect 18412 29093 18452 29178
rect 18508 29168 18548 29800
rect 18604 29765 18644 31228
rect 19276 30773 19316 32138
rect 19275 30764 19317 30773
rect 19275 30724 19276 30764
rect 19316 30724 19317 30764
rect 19275 30715 19317 30724
rect 18795 30680 18837 30689
rect 18700 30640 18796 30680
rect 18836 30640 18837 30680
rect 18603 29756 18645 29765
rect 18603 29716 18604 29756
rect 18644 29716 18645 29756
rect 18603 29707 18645 29716
rect 18411 29084 18453 29093
rect 18316 29044 18412 29084
rect 18452 29044 18453 29084
rect 18411 29035 18453 29044
rect 18508 28673 18548 29128
rect 18507 28664 18549 28673
rect 18507 28624 18508 28664
rect 18548 28624 18549 28664
rect 18507 28615 18549 28624
rect 18700 28580 18740 30640
rect 18795 30631 18837 30640
rect 18796 30546 18836 30631
rect 19372 30605 19412 32236
rect 19467 32236 19468 32276
rect 19508 32236 19509 32276
rect 19467 32227 19509 32236
rect 19468 32142 19508 32227
rect 19468 31352 19508 31361
rect 19564 31352 19604 33571
rect 19508 31312 19604 31352
rect 19468 31303 19508 31312
rect 19659 30680 19701 30689
rect 19659 30640 19660 30680
rect 19700 30640 19701 30680
rect 19659 30631 19701 30640
rect 19371 30596 19413 30605
rect 19371 30556 19372 30596
rect 19412 30556 19413 30596
rect 19371 30547 19413 30556
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 18796 29840 18836 29849
rect 18796 29261 18836 29800
rect 19276 29845 19316 29854
rect 19372 29849 19412 30547
rect 19467 30512 19509 30521
rect 19467 30472 19468 30512
rect 19508 30472 19509 30512
rect 19467 30463 19509 30472
rect 19276 29429 19316 29805
rect 19371 29840 19413 29849
rect 19371 29800 19372 29840
rect 19412 29800 19413 29840
rect 19371 29791 19413 29800
rect 19275 29420 19317 29429
rect 19275 29380 19276 29420
rect 19316 29380 19317 29420
rect 19275 29371 19317 29380
rect 18795 29252 18837 29261
rect 18795 29212 18796 29252
rect 18836 29212 18837 29252
rect 18795 29203 18837 29212
rect 18987 29252 19029 29261
rect 18987 29212 18988 29252
rect 19028 29212 19029 29252
rect 18987 29203 19029 29212
rect 18988 29168 19028 29203
rect 18988 29117 19028 29128
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 18700 28540 18836 28580
rect 18220 28531 18260 28540
rect 18508 28328 18548 28337
rect 18220 28288 18508 28328
rect 18220 27824 18260 28288
rect 18508 28279 18548 28288
rect 18603 28328 18645 28337
rect 18603 28288 18604 28328
rect 18644 28288 18645 28328
rect 18603 28279 18645 28288
rect 18604 28194 18644 28279
rect 18220 27775 18260 27784
rect 18796 27749 18836 28540
rect 18987 28328 19029 28337
rect 18987 28288 18988 28328
rect 19028 28288 19029 28328
rect 18987 28279 19029 28288
rect 19084 28328 19124 28337
rect 18988 28194 19028 28279
rect 19084 28001 19124 28288
rect 19083 27992 19125 28001
rect 19083 27952 19084 27992
rect 19124 27952 19125 27992
rect 19083 27943 19125 27952
rect 19275 27824 19317 27833
rect 19275 27784 19276 27824
rect 19316 27784 19317 27824
rect 19275 27775 19317 27784
rect 18795 27740 18837 27749
rect 18795 27700 18796 27740
rect 18836 27700 18837 27740
rect 18795 27698 18837 27700
rect 18795 27691 18796 27698
rect 18836 27691 18837 27698
rect 18796 27649 18836 27658
rect 18123 27488 18165 27497
rect 18123 27448 18124 27488
rect 18164 27448 18165 27488
rect 18123 27439 18165 27448
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 18316 26816 18356 26825
rect 18316 26657 18356 26776
rect 18796 26821 18836 26830
rect 18315 26648 18357 26657
rect 18315 26608 18316 26648
rect 18356 26608 18357 26648
rect 18315 26599 18357 26608
rect 18507 26396 18549 26405
rect 18507 26356 18508 26396
rect 18548 26356 18549 26396
rect 18507 26347 18549 26356
rect 18508 26153 18548 26347
rect 18699 26312 18741 26321
rect 18796 26312 18836 26781
rect 18988 26732 19028 26741
rect 19276 26732 19316 27775
rect 19028 26692 19316 26732
rect 18988 26683 19028 26692
rect 19275 26480 19317 26489
rect 19275 26440 19276 26480
rect 19316 26440 19317 26480
rect 19372 26480 19412 29791
rect 19468 29756 19508 30463
rect 19468 29707 19508 29716
rect 19660 29336 19700 30631
rect 19660 29287 19700 29296
rect 19516 29158 19700 29168
rect 19556 29128 19700 29158
rect 19516 29109 19556 29118
rect 19564 28328 19604 28339
rect 19564 28253 19604 28288
rect 19563 28244 19605 28253
rect 19563 28204 19564 28244
rect 19604 28204 19605 28244
rect 19563 28195 19605 28204
rect 19372 26440 19508 26480
rect 19275 26431 19317 26440
rect 18699 26272 18700 26312
rect 18740 26272 18836 26312
rect 18699 26263 18741 26272
rect 18220 26144 18260 26153
rect 18124 25556 18164 25565
rect 18220 25556 18260 26104
rect 18315 26144 18357 26153
rect 18315 26104 18316 26144
rect 18356 26104 18357 26144
rect 18315 26095 18357 26104
rect 18507 26144 18549 26153
rect 18700 26144 18740 26153
rect 18507 26104 18508 26144
rect 18548 26104 18549 26144
rect 18507 26095 18549 26104
rect 18604 26104 18700 26144
rect 18316 26010 18356 26095
rect 18604 25649 18644 26104
rect 18700 26095 18740 26104
rect 18795 26144 18837 26153
rect 18795 26104 18796 26144
rect 18836 26104 18837 26144
rect 18795 26095 18837 26104
rect 19276 26144 19316 26431
rect 18796 26010 18836 26095
rect 19276 25901 19316 26104
rect 18699 25892 18741 25901
rect 18699 25852 18700 25892
rect 18740 25852 18741 25892
rect 18699 25843 18741 25852
rect 19275 25892 19317 25901
rect 19275 25852 19276 25892
rect 19316 25852 19317 25892
rect 19275 25843 19317 25852
rect 18603 25640 18645 25649
rect 18603 25600 18604 25640
rect 18644 25600 18645 25640
rect 18603 25591 18645 25600
rect 18164 25516 18260 25556
rect 18124 25507 18164 25516
rect 18700 25397 18740 25843
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18699 25388 18741 25397
rect 18699 25348 18700 25388
rect 18740 25348 18741 25388
rect 18699 25339 18741 25348
rect 17972 25264 18068 25304
rect 17932 25255 17972 25264
rect 18028 24632 18068 25264
rect 18315 25304 18357 25313
rect 18315 25264 18316 25304
rect 18356 25264 18357 25304
rect 18315 25255 18357 25264
rect 18123 25220 18165 25229
rect 18123 25180 18124 25220
rect 18164 25180 18165 25220
rect 18123 25171 18165 25180
rect 18028 23801 18068 24592
rect 18124 24044 18164 25171
rect 18316 25170 18356 25255
rect 18220 24716 18260 24725
rect 18260 24676 18548 24716
rect 18220 24667 18260 24676
rect 18508 24632 18548 24676
rect 18508 24583 18548 24592
rect 18604 24632 18644 24641
rect 18604 24305 18644 24592
rect 18603 24296 18645 24305
rect 18508 24256 18604 24296
rect 18644 24256 18645 24296
rect 18124 24004 18260 24044
rect 18123 23876 18165 23885
rect 18123 23836 18124 23876
rect 18164 23836 18165 23876
rect 18123 23827 18165 23836
rect 18027 23792 18069 23801
rect 18027 23752 18028 23792
rect 18068 23752 18069 23792
rect 18027 23743 18069 23752
rect 17931 23288 17973 23297
rect 17931 23248 17932 23288
rect 17972 23248 17973 23288
rect 17931 23239 17973 23248
rect 17932 23120 17972 23239
rect 18027 23204 18069 23213
rect 18027 23164 18028 23204
rect 18068 23164 18069 23204
rect 18027 23155 18069 23164
rect 17932 23071 17972 23080
rect 18028 23070 18068 23155
rect 17931 22700 17973 22709
rect 17931 22660 17932 22700
rect 17972 22660 17973 22700
rect 17931 22651 17973 22660
rect 17932 21608 17972 22651
rect 17932 21365 17972 21568
rect 18028 22280 18068 22289
rect 17931 21356 17973 21365
rect 17931 21316 17932 21356
rect 17972 21316 17973 21356
rect 17931 21307 17973 21316
rect 17931 20432 17973 20441
rect 17931 20392 17932 20432
rect 17972 20392 17973 20432
rect 17931 20383 17973 20392
rect 17932 20096 17972 20383
rect 18028 20189 18068 22240
rect 18124 22028 18164 23827
rect 18220 23129 18260 24004
rect 18411 23792 18453 23801
rect 18411 23752 18412 23792
rect 18452 23752 18453 23792
rect 18411 23743 18453 23752
rect 18219 23120 18261 23129
rect 18219 23080 18220 23120
rect 18260 23080 18261 23120
rect 18219 23071 18261 23080
rect 18315 22784 18357 22793
rect 18315 22744 18316 22784
rect 18356 22744 18357 22784
rect 18315 22735 18357 22744
rect 18219 22448 18261 22457
rect 18219 22408 18220 22448
rect 18260 22408 18261 22448
rect 18219 22399 18261 22408
rect 18220 22314 18260 22399
rect 18316 22112 18356 22735
rect 18412 22709 18452 23743
rect 18411 22700 18453 22709
rect 18411 22660 18412 22700
rect 18452 22660 18453 22700
rect 18411 22651 18453 22660
rect 18508 22616 18548 24256
rect 18603 24247 18645 24256
rect 18603 23960 18645 23969
rect 18603 23920 18604 23960
rect 18644 23920 18645 23960
rect 18603 23911 18645 23920
rect 18604 23826 18644 23911
rect 18700 23708 18740 25339
rect 19468 25304 19508 26440
rect 19660 25556 19700 29128
rect 19852 26312 19892 35251
rect 19948 34721 19988 35680
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 19947 34712 19989 34721
rect 19947 34672 19948 34712
rect 19988 34672 19989 34712
rect 19947 34663 19989 34672
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 20236 33872 20276 33881
rect 20524 33872 20564 40207
rect 20619 39836 20661 39845
rect 20619 39796 20620 39836
rect 20660 39796 20661 39836
rect 20619 39787 20661 39796
rect 20276 33832 20564 33872
rect 20236 33823 20276 33832
rect 20044 33690 20084 33699
rect 20044 33293 20084 33650
rect 20043 33284 20085 33293
rect 20043 33244 20044 33284
rect 20084 33244 20085 33284
rect 20043 33235 20085 33244
rect 20523 33284 20565 33293
rect 20523 33244 20524 33284
rect 20564 33244 20565 33284
rect 20523 33235 20565 33244
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 19948 31357 19988 31366
rect 19948 27824 19988 31317
rect 20140 31193 20180 31278
rect 20139 31184 20181 31193
rect 20139 31144 20140 31184
rect 20180 31144 20181 31184
rect 20139 31135 20181 31144
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 20236 30848 20276 30857
rect 20524 30848 20564 33235
rect 20276 30808 20564 30848
rect 20236 30799 20276 30808
rect 20044 30680 20084 30691
rect 20044 30605 20084 30640
rect 20043 30596 20085 30605
rect 20043 30556 20044 30596
rect 20084 30556 20085 30596
rect 20043 30547 20085 30556
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 20235 28832 20277 28841
rect 20235 28792 20236 28832
rect 20276 28792 20277 28832
rect 20235 28783 20277 28792
rect 20044 28337 20084 28342
rect 20043 28333 20085 28337
rect 20043 28288 20044 28333
rect 20084 28288 20085 28333
rect 20043 28279 20085 28288
rect 20044 28198 20084 28279
rect 20236 28244 20276 28783
rect 20523 28328 20565 28337
rect 20523 28288 20524 28328
rect 20564 28288 20565 28328
rect 20523 28279 20565 28288
rect 20236 28195 20276 28204
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 19948 27784 20180 27824
rect 20140 27740 20180 27784
rect 20236 27740 20276 27749
rect 20140 27700 20236 27740
rect 20236 27691 20276 27700
rect 20043 27656 20085 27665
rect 20043 27616 20044 27656
rect 20084 27616 20085 27656
rect 20043 27607 20085 27616
rect 20044 27522 20084 27607
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 19948 26312 19988 26321
rect 19852 26272 19948 26312
rect 19948 26263 19988 26272
rect 19804 26134 19988 26144
rect 19844 26104 19988 26134
rect 19804 26085 19844 26094
rect 19756 25556 19796 25565
rect 19660 25516 19756 25556
rect 19756 25507 19796 25516
rect 19564 25304 19604 25313
rect 19468 25264 19564 25304
rect 19604 25264 19796 25304
rect 19564 25255 19604 25264
rect 18987 24716 19029 24725
rect 18987 24676 18988 24716
rect 19028 24676 19029 24716
rect 18987 24667 19029 24676
rect 19371 24716 19413 24725
rect 19371 24676 19372 24716
rect 19412 24676 19413 24716
rect 19371 24667 19413 24676
rect 18988 24632 19028 24667
rect 18988 24581 19028 24592
rect 19084 24548 19124 24557
rect 19124 24508 19316 24548
rect 19084 24499 19124 24508
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 18604 23668 18740 23708
rect 18796 23792 18836 23801
rect 18604 22952 18644 23668
rect 18700 23129 18740 23214
rect 18699 23120 18741 23129
rect 18699 23080 18700 23120
rect 18740 23080 18741 23120
rect 18699 23071 18741 23080
rect 18796 23045 18836 23752
rect 18795 23036 18837 23045
rect 18795 22996 18796 23036
rect 18836 22996 18837 23036
rect 18795 22987 18837 22996
rect 19276 22961 19316 24508
rect 19275 22952 19317 22961
rect 18604 22912 18740 22952
rect 18508 22576 18644 22616
rect 18507 22448 18549 22457
rect 18507 22408 18508 22448
rect 18548 22408 18549 22448
rect 18507 22399 18549 22408
rect 18508 22280 18548 22399
rect 18604 22289 18644 22576
rect 18508 22231 18548 22240
rect 18603 22280 18645 22289
rect 18603 22240 18604 22280
rect 18644 22240 18645 22280
rect 18603 22231 18645 22240
rect 18604 22146 18644 22231
rect 18316 22072 18548 22112
rect 18124 21988 18356 22028
rect 18124 21701 18164 21786
rect 18123 21692 18165 21701
rect 18123 21652 18124 21692
rect 18164 21652 18165 21692
rect 18123 21643 18165 21652
rect 18316 21608 18356 21988
rect 18411 21692 18453 21701
rect 18411 21652 18412 21692
rect 18452 21652 18453 21692
rect 18411 21643 18453 21652
rect 18220 21568 18356 21608
rect 18412 21608 18452 21643
rect 18220 21524 18260 21568
rect 18412 21557 18452 21568
rect 18508 21608 18548 22072
rect 18548 21568 18644 21608
rect 18508 21559 18548 21568
rect 18124 21484 18260 21524
rect 18027 20180 18069 20189
rect 18027 20140 18028 20180
rect 18068 20140 18069 20180
rect 18027 20131 18069 20140
rect 17932 20047 17972 20056
rect 18028 19844 18068 19853
rect 18028 19265 18068 19804
rect 18027 19256 18069 19265
rect 18027 19216 18028 19256
rect 18068 19216 18069 19256
rect 18027 19207 18069 19216
rect 17932 17744 17972 17753
rect 17836 17704 17932 17744
rect 17739 17240 17781 17249
rect 17739 17200 17740 17240
rect 17780 17200 17781 17240
rect 17739 17191 17781 17200
rect 17836 17072 17876 17704
rect 17932 17695 17972 17704
rect 17931 17576 17973 17585
rect 17931 17536 17932 17576
rect 17972 17536 17973 17576
rect 17931 17527 17973 17536
rect 17740 17032 17876 17072
rect 17643 16316 17685 16325
rect 17643 16276 17644 16316
rect 17684 16276 17685 16316
rect 17643 16267 17685 16276
rect 17644 16182 17684 16267
rect 17740 16064 17780 17032
rect 17644 16024 17780 16064
rect 17836 16232 17876 16241
rect 17547 15308 17589 15317
rect 17547 15268 17548 15308
rect 17588 15268 17589 15308
rect 17547 15259 17589 15268
rect 17547 14720 17589 14729
rect 17547 14680 17548 14720
rect 17588 14680 17589 14720
rect 17547 14671 17589 14680
rect 17548 14586 17588 14671
rect 17356 14176 17492 14216
rect 17259 11696 17301 11705
rect 17259 11656 17260 11696
rect 17300 11656 17301 11696
rect 17259 11647 17301 11656
rect 17260 11562 17300 11647
rect 17163 11444 17205 11453
rect 17163 11404 17164 11444
rect 17204 11404 17205 11444
rect 17163 11395 17205 11404
rect 17163 11276 17205 11285
rect 17163 11236 17164 11276
rect 17204 11236 17205 11276
rect 17163 11227 17205 11236
rect 17164 10361 17204 11227
rect 17356 11108 17396 14176
rect 17644 13376 17684 16024
rect 17739 15560 17781 15569
rect 17739 15520 17740 15560
rect 17780 15520 17781 15560
rect 17739 15511 17781 15520
rect 17740 15426 17780 15511
rect 17836 15401 17876 16192
rect 17932 16232 17972 17527
rect 18124 16400 18164 21484
rect 18315 21356 18357 21365
rect 18315 21316 18316 21356
rect 18356 21316 18357 21356
rect 18315 21307 18357 21316
rect 18507 21356 18549 21365
rect 18507 21316 18508 21356
rect 18548 21316 18549 21356
rect 18507 21307 18549 21316
rect 18219 20180 18261 20189
rect 18219 20140 18220 20180
rect 18260 20140 18261 20180
rect 18219 20131 18261 20140
rect 18220 19601 18260 20131
rect 18219 19592 18261 19601
rect 18219 19552 18220 19592
rect 18260 19552 18261 19592
rect 18219 19543 18261 19552
rect 18220 19256 18260 19543
rect 18316 19265 18356 21307
rect 18508 20768 18548 21307
rect 18508 20719 18548 20728
rect 18508 20096 18548 20105
rect 18412 19508 18452 19517
rect 18508 19508 18548 20056
rect 18604 20096 18644 21568
rect 18700 20180 18740 22912
rect 19275 22912 19276 22952
rect 19316 22912 19317 22952
rect 19275 22903 19317 22912
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 19275 22616 19317 22625
rect 19275 22576 19276 22616
rect 19316 22576 19317 22616
rect 19275 22567 19317 22576
rect 19083 22532 19125 22541
rect 19083 22492 19084 22532
rect 19124 22492 19125 22532
rect 19083 22483 19125 22492
rect 18987 22448 19029 22457
rect 18987 22408 18988 22448
rect 19028 22408 19029 22448
rect 18987 22399 19029 22408
rect 18988 22364 19028 22399
rect 18891 22280 18933 22289
rect 18891 22240 18892 22280
rect 18932 22240 18933 22280
rect 18891 22231 18933 22240
rect 18892 21608 18932 22231
rect 18988 21617 19028 22324
rect 19084 22364 19124 22483
rect 19084 22315 19124 22324
rect 18892 21559 18932 21568
rect 18987 21608 19029 21617
rect 18987 21568 18988 21608
rect 19028 21568 19029 21608
rect 18987 21559 19029 21568
rect 18988 21474 19028 21559
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 18987 20180 19029 20189
rect 18700 20140 18836 20180
rect 18644 20056 18740 20096
rect 18604 20047 18644 20056
rect 18603 19928 18645 19937
rect 18603 19888 18604 19928
rect 18644 19888 18645 19928
rect 18603 19879 18645 19888
rect 18452 19468 18548 19508
rect 18412 19459 18452 19468
rect 18604 19424 18644 19879
rect 18508 19384 18644 19424
rect 18220 19207 18260 19216
rect 18315 19256 18357 19265
rect 18315 19216 18316 19256
rect 18356 19216 18357 19256
rect 18315 19207 18357 19216
rect 18316 18341 18356 19207
rect 18508 18677 18548 19384
rect 18604 19256 18644 19265
rect 18604 18929 18644 19216
rect 18603 18920 18645 18929
rect 18603 18880 18604 18920
rect 18644 18880 18645 18920
rect 18603 18871 18645 18880
rect 18507 18668 18549 18677
rect 18507 18628 18508 18668
rect 18548 18628 18549 18668
rect 18507 18619 18549 18628
rect 18412 18584 18452 18593
rect 18315 18332 18357 18341
rect 18315 18292 18316 18332
rect 18356 18292 18357 18332
rect 18315 18283 18357 18292
rect 18412 18257 18452 18544
rect 18604 18584 18644 18593
rect 18508 18500 18548 18509
rect 18411 18248 18453 18257
rect 18411 18208 18412 18248
rect 18452 18208 18453 18248
rect 18411 18199 18453 18208
rect 18315 17240 18357 17249
rect 18315 17200 18316 17240
rect 18356 17200 18357 17240
rect 18315 17191 18357 17200
rect 18316 16493 18356 17191
rect 18315 16484 18357 16493
rect 18315 16444 18316 16484
rect 18356 16444 18357 16484
rect 18315 16435 18357 16444
rect 18028 16360 18164 16400
rect 18028 16241 18068 16360
rect 17932 16183 17972 16192
rect 18027 16232 18069 16241
rect 18027 16192 18028 16232
rect 18068 16192 18069 16232
rect 18027 16183 18069 16192
rect 18124 16232 18164 16241
rect 18316 16232 18356 16435
rect 18508 16400 18548 18460
rect 18604 18005 18644 18544
rect 18603 17996 18645 18005
rect 18603 17956 18604 17996
rect 18644 17956 18645 17996
rect 18603 17947 18645 17956
rect 18603 17828 18645 17837
rect 18603 17788 18604 17828
rect 18644 17788 18645 17828
rect 18603 17779 18645 17788
rect 18604 17072 18644 17779
rect 18700 17501 18740 20056
rect 18796 20021 18836 20140
rect 18987 20140 18988 20180
rect 19028 20140 19029 20180
rect 18987 20131 19029 20140
rect 18988 20096 19028 20131
rect 18988 20045 19028 20056
rect 18795 20012 18837 20021
rect 18795 19972 18796 20012
rect 18836 19972 18837 20012
rect 18795 19963 18837 19972
rect 19083 20012 19125 20021
rect 19083 19972 19084 20012
rect 19124 19972 19125 20012
rect 19083 19963 19125 19972
rect 19084 19878 19124 19963
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 18795 18920 18837 18929
rect 18795 18880 18796 18920
rect 18836 18880 18837 18920
rect 18795 18871 18837 18880
rect 18796 18584 18836 18871
rect 19276 18593 19316 22567
rect 19372 22457 19412 24667
rect 19564 24632 19604 24641
rect 19467 23456 19509 23465
rect 19467 23416 19468 23456
rect 19508 23416 19509 23456
rect 19467 23407 19509 23416
rect 19371 22448 19413 22457
rect 19371 22408 19372 22448
rect 19412 22408 19413 22448
rect 19371 22399 19413 22408
rect 19468 21608 19508 23407
rect 19564 22625 19604 24592
rect 19563 22616 19605 22625
rect 19563 22576 19564 22616
rect 19604 22576 19605 22616
rect 19563 22567 19605 22576
rect 19564 22280 19604 22567
rect 19564 22231 19604 22240
rect 19468 20180 19508 21568
rect 19756 20768 19796 25264
rect 19851 23792 19893 23801
rect 19851 23752 19852 23792
rect 19892 23752 19893 23792
rect 19851 23743 19893 23752
rect 19852 23120 19892 23743
rect 19948 23288 19988 26104
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20235 24716 20277 24725
rect 20235 24676 20236 24716
rect 20276 24676 20277 24716
rect 20235 24667 20277 24676
rect 20044 24618 20084 24627
rect 20236 24582 20276 24667
rect 20044 23969 20084 24578
rect 20043 23960 20085 23969
rect 20043 23920 20044 23960
rect 20084 23920 20085 23960
rect 20043 23911 20085 23920
rect 20236 23960 20276 23969
rect 20524 23960 20564 28279
rect 20276 23920 20564 23960
rect 20236 23911 20276 23920
rect 20044 23792 20084 23803
rect 20044 23717 20084 23752
rect 20043 23708 20085 23717
rect 20043 23668 20044 23708
rect 20084 23668 20085 23708
rect 20043 23659 20085 23668
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 20140 23288 20180 23297
rect 19948 23248 20140 23288
rect 20140 23239 20180 23248
rect 19948 23120 19988 23129
rect 19852 23080 19948 23120
rect 19948 23071 19988 23080
rect 20044 22285 20084 22294
rect 20044 22112 20084 22245
rect 20236 22196 20276 22205
rect 20620 22196 20660 39787
rect 20715 36224 20757 36233
rect 20715 36184 20716 36224
rect 20756 36184 20757 36224
rect 20715 36175 20757 36184
rect 20716 34553 20756 36175
rect 20811 35972 20853 35981
rect 20811 35932 20812 35972
rect 20852 35932 20853 35972
rect 20811 35923 20853 35932
rect 20715 34544 20757 34553
rect 20715 34504 20716 34544
rect 20756 34504 20757 34544
rect 20715 34495 20757 34504
rect 20812 33881 20852 35923
rect 20908 34301 20948 42895
rect 21004 42449 21044 63055
rect 21100 52949 21140 72463
rect 21195 63776 21237 63785
rect 21195 63736 21196 63776
rect 21236 63736 21237 63776
rect 21195 63727 21237 63736
rect 21099 52940 21141 52949
rect 21099 52900 21100 52940
rect 21140 52900 21141 52940
rect 21099 52891 21141 52900
rect 21003 42440 21045 42449
rect 21003 42400 21004 42440
rect 21044 42400 21045 42440
rect 21003 42391 21045 42400
rect 21003 42272 21045 42281
rect 21003 42232 21004 42272
rect 21044 42232 21045 42272
rect 21003 42223 21045 42232
rect 21004 39929 21044 42223
rect 21099 42188 21141 42197
rect 21099 42148 21100 42188
rect 21140 42148 21141 42188
rect 21099 42139 21141 42148
rect 21100 41609 21140 42139
rect 21196 41861 21236 63727
rect 21292 62525 21332 74563
rect 21291 62516 21333 62525
rect 21291 62476 21292 62516
rect 21332 62476 21333 62516
rect 21291 62467 21333 62476
rect 21291 54200 21333 54209
rect 21291 54160 21292 54200
rect 21332 54160 21333 54200
rect 21291 54151 21333 54160
rect 21292 49001 21332 54151
rect 21387 49832 21429 49841
rect 21387 49792 21388 49832
rect 21428 49792 21429 49832
rect 21387 49783 21429 49792
rect 21388 49337 21428 49783
rect 21387 49328 21429 49337
rect 21387 49288 21388 49328
rect 21428 49288 21429 49328
rect 21387 49279 21429 49288
rect 21291 48992 21333 49001
rect 21291 48952 21292 48992
rect 21332 48952 21333 48992
rect 21291 48943 21333 48952
rect 21291 47396 21333 47405
rect 21291 47356 21292 47396
rect 21332 47356 21333 47396
rect 21291 47347 21333 47356
rect 21195 41852 21237 41861
rect 21195 41812 21196 41852
rect 21236 41812 21237 41852
rect 21195 41803 21237 41812
rect 21099 41600 21141 41609
rect 21099 41560 21100 41600
rect 21140 41560 21141 41600
rect 21099 41551 21141 41560
rect 21195 41264 21237 41273
rect 21195 41224 21196 41264
rect 21236 41224 21237 41264
rect 21195 41215 21237 41224
rect 21003 39920 21045 39929
rect 21003 39880 21004 39920
rect 21044 39880 21045 39920
rect 21003 39871 21045 39880
rect 21099 36644 21141 36653
rect 21099 36604 21100 36644
rect 21140 36604 21141 36644
rect 21099 36595 21141 36604
rect 21003 36392 21045 36401
rect 21003 36352 21004 36392
rect 21044 36352 21045 36392
rect 21003 36343 21045 36352
rect 20907 34292 20949 34301
rect 20907 34252 20908 34292
rect 20948 34252 20949 34292
rect 20907 34243 20949 34252
rect 20811 33872 20853 33881
rect 20811 33832 20812 33872
rect 20852 33832 20853 33872
rect 20811 33823 20853 33832
rect 20811 31856 20853 31865
rect 20811 31816 20812 31856
rect 20852 31816 20853 31856
rect 20811 31807 20853 31816
rect 20715 31184 20757 31193
rect 20715 31144 20716 31184
rect 20756 31144 20757 31184
rect 20715 31135 20757 31144
rect 20716 29513 20756 31135
rect 20715 29504 20757 29513
rect 20715 29464 20716 29504
rect 20756 29464 20757 29504
rect 20715 29455 20757 29464
rect 20715 29168 20757 29177
rect 20715 29128 20716 29168
rect 20756 29128 20757 29168
rect 20715 29119 20757 29128
rect 20716 24725 20756 29119
rect 20715 24716 20757 24725
rect 20715 24676 20716 24716
rect 20756 24676 20757 24716
rect 20715 24667 20757 24676
rect 20812 23960 20852 31807
rect 20907 28748 20949 28757
rect 20907 28708 20908 28748
rect 20948 28708 20949 28748
rect 20907 28699 20949 28708
rect 20908 27497 20948 28699
rect 20907 27488 20949 27497
rect 20907 27448 20908 27488
rect 20948 27448 20949 27488
rect 20907 27439 20949 27448
rect 20276 22156 20660 22196
rect 20716 23920 20852 23960
rect 20236 22147 20276 22156
rect 19948 22072 20084 22112
rect 19948 21692 19988 22072
rect 20716 22028 20756 23920
rect 21004 23129 21044 36343
rect 21100 32873 21140 36595
rect 21099 32864 21141 32873
rect 21099 32824 21100 32864
rect 21140 32824 21141 32864
rect 21099 32815 21141 32824
rect 21196 30689 21236 41215
rect 21292 33545 21332 47347
rect 21291 33536 21333 33545
rect 21291 33496 21292 33536
rect 21332 33496 21333 33536
rect 21291 33487 21333 33496
rect 21195 30680 21237 30689
rect 21195 30640 21196 30680
rect 21236 30640 21237 30680
rect 21195 30631 21237 30640
rect 21099 28580 21141 28589
rect 21099 28540 21100 28580
rect 21140 28540 21141 28580
rect 21099 28531 21141 28540
rect 21100 27161 21140 28531
rect 21099 27152 21141 27161
rect 21099 27112 21100 27152
rect 21140 27112 21141 27152
rect 21099 27103 21141 27112
rect 21003 23120 21045 23129
rect 21003 23080 21004 23120
rect 21044 23080 21045 23120
rect 21003 23071 21045 23080
rect 20524 21988 20756 22028
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20140 21776 20180 21785
rect 20524 21776 20564 21988
rect 20180 21736 20564 21776
rect 20140 21727 20180 21736
rect 19948 21652 20084 21692
rect 19948 21594 19988 21603
rect 19948 20768 19988 21554
rect 19372 20140 19604 20180
rect 18796 18509 18836 18544
rect 19275 18584 19317 18593
rect 19275 18544 19276 18584
rect 19316 18544 19317 18584
rect 19275 18535 19317 18544
rect 18795 18500 18837 18509
rect 18795 18460 18796 18500
rect 18836 18460 18837 18500
rect 18795 18451 18837 18460
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 19372 17996 19412 20140
rect 19564 20096 19604 20140
rect 19564 20047 19604 20056
rect 19467 20012 19509 20021
rect 19467 19972 19468 20012
rect 19508 19972 19509 20012
rect 19467 19963 19509 19972
rect 19084 17956 19412 17996
rect 19084 17576 19124 17956
rect 19179 17828 19221 17837
rect 19179 17788 19180 17828
rect 19220 17788 19221 17828
rect 19179 17779 19221 17788
rect 19180 17744 19220 17779
rect 19180 17693 19220 17704
rect 19372 17660 19412 17669
rect 19276 17620 19372 17660
rect 19084 17536 19220 17576
rect 18699 17492 18741 17501
rect 18699 17452 18700 17492
rect 18740 17452 18741 17492
rect 18699 17443 18741 17452
rect 18795 17240 18837 17249
rect 18795 17200 18796 17240
rect 18836 17200 18837 17240
rect 18795 17191 18837 17200
rect 19083 17240 19125 17249
rect 19083 17200 19084 17240
rect 19124 17200 19125 17240
rect 19083 17191 19125 17200
rect 18796 17106 18836 17191
rect 18604 16484 18644 17032
rect 19084 17072 19124 17191
rect 19084 17023 19124 17032
rect 19180 16988 19220 17536
rect 19276 17165 19316 17620
rect 19372 17611 19412 17620
rect 19371 17492 19413 17501
rect 19371 17452 19372 17492
rect 19412 17452 19413 17492
rect 19371 17443 19413 17452
rect 19275 17156 19317 17165
rect 19275 17116 19276 17156
rect 19316 17116 19317 17156
rect 19275 17107 19317 17116
rect 19372 17072 19412 17443
rect 19468 17156 19508 19963
rect 19756 19601 19796 20728
rect 19852 20728 19988 20768
rect 19852 20180 19892 20728
rect 19948 20600 19988 20609
rect 20044 20600 20084 21652
rect 19988 20560 20084 20600
rect 19948 20551 19988 20560
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 20235 20180 20277 20189
rect 19852 20140 19988 20180
rect 19755 19592 19797 19601
rect 19755 19552 19756 19592
rect 19796 19552 19797 19592
rect 19755 19543 19797 19552
rect 19659 18668 19701 18677
rect 19659 18628 19660 18668
rect 19700 18628 19701 18668
rect 19756 18668 19796 19543
rect 19948 19508 19988 20140
rect 20235 20140 20236 20180
rect 20276 20140 20277 20180
rect 20235 20131 20277 20140
rect 20044 20082 20084 20091
rect 20236 20046 20276 20131
rect 20044 19685 20084 20042
rect 20043 19676 20085 19685
rect 20043 19636 20044 19676
rect 20084 19636 20085 19676
rect 20043 19627 20085 19636
rect 20523 19676 20565 19685
rect 20523 19636 20524 19676
rect 20564 19636 20565 19676
rect 20523 19627 20565 19636
rect 20044 19508 20084 19517
rect 19948 19468 20044 19508
rect 20044 19459 20084 19468
rect 19851 19256 19893 19265
rect 19851 19216 19852 19256
rect 19892 19216 19893 19256
rect 19851 19207 19893 19216
rect 19852 19122 19892 19207
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 20236 18752 20276 18761
rect 20524 18752 20564 19627
rect 20276 18712 20564 18752
rect 20236 18703 20276 18712
rect 19756 18628 20084 18668
rect 19659 18619 19701 18628
rect 19563 17996 19605 18005
rect 19563 17956 19564 17996
rect 19604 17956 19605 17996
rect 19563 17947 19605 17956
rect 19564 17744 19604 17947
rect 19564 17695 19604 17704
rect 19660 17744 19700 18619
rect 20044 18584 20084 18628
rect 20044 18535 20084 18544
rect 19660 17695 19700 17704
rect 19756 17744 19796 17753
rect 20044 17744 20084 17753
rect 19796 17704 20044 17744
rect 19756 17695 19796 17704
rect 20044 17695 20084 17704
rect 20140 17744 20180 17753
rect 20180 17704 20564 17744
rect 20140 17695 20180 17704
rect 19851 17576 19893 17585
rect 19851 17536 19852 17576
rect 19892 17536 19893 17576
rect 19851 17527 19893 17536
rect 19852 17442 19892 17527
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 20043 17240 20085 17249
rect 20043 17200 20044 17240
rect 20084 17200 20085 17240
rect 20043 17191 20085 17200
rect 20236 17240 20276 17249
rect 20524 17240 20564 17704
rect 20276 17200 20564 17240
rect 20236 17191 20276 17200
rect 19468 17107 19508 17116
rect 19372 17023 19412 17032
rect 19947 17072 19989 17081
rect 19947 17032 19948 17072
rect 19988 17032 19989 17072
rect 19947 17023 19989 17032
rect 20044 17072 20084 17191
rect 20139 17156 20181 17165
rect 20139 17116 20140 17156
rect 20180 17116 20181 17156
rect 20139 17107 20181 17116
rect 20044 17023 20084 17032
rect 20140 17030 20180 17107
rect 19180 16948 19316 16988
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 18891 16484 18933 16493
rect 19276 16484 19316 16948
rect 19948 16938 19988 17023
rect 19756 16820 19796 16829
rect 19660 16780 19756 16820
rect 18604 16444 18836 16484
rect 18508 16360 18740 16400
rect 18164 16192 18260 16232
rect 18124 16183 18164 16192
rect 18028 16064 18068 16073
rect 18068 16024 18164 16064
rect 18028 16015 18068 16024
rect 18027 15896 18069 15905
rect 18027 15856 18028 15896
rect 18068 15856 18069 15896
rect 18027 15847 18069 15856
rect 17835 15392 17877 15401
rect 17835 15352 17836 15392
rect 17876 15352 17877 15392
rect 17835 15343 17877 15352
rect 18028 15149 18068 15847
rect 18124 15728 18164 16024
rect 18220 15812 18260 16192
rect 18316 16183 18356 16192
rect 18412 16232 18452 16241
rect 18412 16073 18452 16192
rect 18508 16232 18548 16243
rect 18508 16157 18548 16192
rect 18603 16232 18645 16241
rect 18603 16192 18604 16232
rect 18644 16192 18645 16232
rect 18603 16183 18645 16192
rect 18507 16148 18549 16157
rect 18507 16108 18508 16148
rect 18548 16108 18549 16148
rect 18507 16099 18549 16108
rect 18604 16098 18644 16183
rect 18700 16157 18740 16360
rect 18699 16148 18741 16157
rect 18699 16108 18700 16148
rect 18740 16108 18741 16148
rect 18699 16099 18741 16108
rect 18411 16064 18453 16073
rect 18411 16024 18412 16064
rect 18452 16024 18453 16064
rect 18796 16064 18836 16444
rect 18891 16444 18892 16484
rect 18932 16444 18933 16484
rect 18891 16435 18933 16444
rect 19084 16444 19316 16484
rect 19371 16484 19413 16493
rect 19371 16444 19372 16484
rect 19412 16444 19413 16484
rect 18892 16232 18932 16435
rect 18892 16183 18932 16192
rect 19084 16073 19124 16444
rect 19371 16435 19413 16444
rect 19372 16316 19412 16435
rect 19564 16400 19604 16409
rect 19180 16276 19412 16316
rect 19468 16360 19564 16400
rect 19180 16232 19220 16276
rect 19180 16183 19220 16192
rect 19276 16148 19316 16157
rect 19083 16064 19125 16073
rect 18796 16024 18932 16064
rect 18411 16015 18453 16024
rect 18220 15772 18356 15812
rect 18124 15688 18260 15728
rect 18124 15560 18164 15569
rect 18124 15317 18164 15520
rect 18123 15308 18165 15317
rect 18123 15268 18124 15308
rect 18164 15268 18165 15308
rect 18123 15259 18165 15268
rect 18027 15140 18069 15149
rect 18027 15100 18028 15140
rect 18068 15100 18069 15140
rect 18027 15091 18069 15100
rect 17452 13336 17684 13376
rect 17452 12545 17492 13336
rect 18124 13301 18164 13386
rect 17739 13292 17781 13301
rect 17739 13252 17740 13292
rect 17780 13252 17781 13292
rect 17739 13243 17781 13252
rect 18123 13292 18165 13301
rect 18123 13252 18124 13292
rect 18164 13252 18165 13292
rect 18123 13243 18165 13252
rect 17596 13217 17636 13226
rect 17636 13177 17684 13208
rect 17596 13168 17684 13177
rect 17547 12704 17589 12713
rect 17547 12664 17548 12704
rect 17588 12664 17589 12704
rect 17547 12655 17589 12664
rect 17451 12536 17493 12545
rect 17451 12496 17452 12536
rect 17492 12496 17493 12536
rect 17451 12487 17493 12496
rect 17548 12536 17588 12655
rect 17644 12620 17684 13168
rect 17740 13124 17780 13243
rect 17740 13075 17780 13084
rect 18123 13124 18165 13133
rect 18123 13084 18124 13124
rect 18164 13084 18165 13124
rect 18123 13075 18165 13084
rect 17931 13040 17973 13049
rect 17931 13000 17932 13040
rect 17972 13000 17973 13040
rect 17931 12991 17973 13000
rect 17932 12906 17972 12991
rect 18027 12956 18069 12965
rect 18027 12916 18028 12956
rect 18068 12916 18069 12956
rect 18027 12907 18069 12916
rect 17740 12620 17780 12629
rect 17644 12580 17740 12620
rect 17740 12571 17780 12580
rect 17452 11108 17492 11117
rect 17356 11068 17452 11108
rect 17260 11010 17300 11019
rect 17260 10445 17300 10970
rect 17259 10436 17301 10445
rect 17259 10396 17260 10436
rect 17300 10396 17301 10436
rect 17259 10387 17301 10396
rect 17163 10352 17205 10361
rect 17163 10312 17164 10352
rect 17204 10312 17205 10352
rect 17163 10303 17205 10312
rect 17164 10109 17204 10303
rect 17163 10100 17205 10109
rect 17163 10060 17164 10100
rect 17204 10060 17205 10100
rect 17163 10051 17205 10060
rect 17356 8849 17396 11068
rect 17452 11059 17492 11068
rect 17451 10520 17493 10529
rect 17451 10480 17452 10520
rect 17492 10480 17493 10520
rect 17451 10471 17493 10480
rect 17355 8840 17397 8849
rect 17355 8800 17356 8840
rect 17396 8800 17397 8840
rect 17355 8791 17397 8800
rect 17067 8000 17109 8009
rect 17067 7960 17068 8000
rect 17108 7960 17109 8000
rect 17067 7951 17109 7960
rect 17164 8000 17204 8009
rect 16779 6320 16821 6329
rect 16779 6280 16780 6320
rect 16820 6280 16821 6320
rect 16779 6271 16821 6280
rect 16780 5648 16820 5657
rect 16683 5564 16725 5573
rect 16683 5524 16684 5564
rect 16724 5524 16725 5564
rect 16683 5515 16725 5524
rect 16780 5405 16820 5608
rect 16876 5648 16916 5657
rect 16916 5608 17012 5648
rect 16876 5599 16916 5608
rect 16779 5396 16821 5405
rect 16779 5356 16780 5396
rect 16820 5356 16821 5396
rect 16779 5347 16821 5356
rect 16588 5020 16916 5060
rect 16587 4136 16629 4145
rect 16587 4096 16588 4136
rect 16628 4096 16629 4136
rect 16587 4087 16629 4096
rect 16588 4002 16628 4087
rect 16780 3968 16820 3977
rect 16684 3928 16780 3968
rect 16587 3380 16629 3389
rect 16587 3340 16588 3380
rect 16628 3340 16629 3380
rect 16587 3331 16629 3340
rect 16588 3246 16628 3331
rect 16587 3128 16629 3137
rect 16587 3088 16588 3128
rect 16628 3088 16629 3128
rect 16587 3079 16629 3088
rect 16396 2500 16532 2540
rect 16299 1112 16341 1121
rect 16299 1072 16300 1112
rect 16340 1072 16341 1112
rect 16299 1063 16341 1072
rect 16396 80 16436 2500
rect 16491 2204 16533 2213
rect 16491 2164 16492 2204
rect 16532 2164 16533 2204
rect 16491 2155 16533 2164
rect 16492 1952 16532 2155
rect 16492 1903 16532 1912
rect 16588 80 16628 3079
rect 16684 2638 16724 3928
rect 16780 3919 16820 3928
rect 16780 3212 16820 3221
rect 16780 2885 16820 3172
rect 16779 2876 16821 2885
rect 16779 2836 16780 2876
rect 16820 2836 16821 2876
rect 16779 2827 16821 2836
rect 16684 2589 16724 2598
rect 16876 2540 16916 5020
rect 16972 4565 17012 5608
rect 16971 4556 17013 4565
rect 16971 4516 16972 4556
rect 17012 4516 17013 4556
rect 16971 4507 17013 4516
rect 16971 3380 17013 3389
rect 16971 3340 16972 3380
rect 17012 3340 17013 3380
rect 16971 3331 17013 3340
rect 16972 3246 17012 3331
rect 17068 2969 17108 7951
rect 17164 7589 17204 7960
rect 17163 7580 17205 7589
rect 17163 7540 17164 7580
rect 17204 7540 17205 7580
rect 17163 7531 17205 7540
rect 17259 5900 17301 5909
rect 17259 5860 17260 5900
rect 17300 5860 17301 5900
rect 17259 5851 17301 5860
rect 17260 5732 17300 5851
rect 17355 5816 17397 5825
rect 17355 5776 17356 5816
rect 17396 5776 17397 5816
rect 17355 5767 17397 5776
rect 17260 5683 17300 5692
rect 17356 5732 17396 5767
rect 17356 5681 17396 5692
rect 17259 5564 17301 5573
rect 17259 5524 17260 5564
rect 17300 5524 17301 5564
rect 17259 5515 17301 5524
rect 17163 4976 17205 4985
rect 17163 4936 17164 4976
rect 17204 4936 17205 4976
rect 17260 4976 17300 5515
rect 17355 5396 17397 5405
rect 17355 5356 17356 5396
rect 17396 5356 17397 5396
rect 17355 5347 17397 5356
rect 17356 5144 17396 5347
rect 17356 5095 17396 5104
rect 17260 4936 17396 4976
rect 17163 4927 17205 4936
rect 17164 4842 17204 4927
rect 17356 3380 17396 4936
rect 17356 3331 17396 3340
rect 17164 3212 17204 3221
rect 17067 2960 17109 2969
rect 17067 2920 17068 2960
rect 17108 2920 17109 2960
rect 17067 2911 17109 2920
rect 17068 2624 17108 2911
rect 17068 2575 17108 2584
rect 16876 2491 16916 2500
rect 16683 1952 16725 1961
rect 16683 1912 16684 1952
rect 16724 1912 16725 1952
rect 16683 1903 16725 1912
rect 16684 197 16724 1903
rect 17164 1541 17204 3172
rect 17163 1532 17205 1541
rect 17163 1492 17164 1532
rect 17204 1492 17205 1532
rect 17163 1483 17205 1492
rect 16779 1364 16821 1373
rect 16779 1324 16780 1364
rect 16820 1324 16821 1364
rect 16779 1315 16821 1324
rect 16780 1112 16820 1315
rect 17163 1196 17205 1205
rect 17163 1156 17164 1196
rect 17204 1156 17205 1196
rect 17163 1147 17205 1156
rect 16780 1063 16820 1072
rect 17164 1062 17204 1147
rect 16972 944 17012 953
rect 16779 776 16821 785
rect 16779 736 16780 776
rect 16820 736 16821 776
rect 16779 727 16821 736
rect 16683 188 16725 197
rect 16683 148 16684 188
rect 16724 148 16725 188
rect 16683 139 16725 148
rect 16780 80 16820 727
rect 16972 281 17012 904
rect 17355 944 17397 953
rect 17355 904 17356 944
rect 17396 904 17397 944
rect 17355 895 17397 904
rect 17356 810 17396 895
rect 17452 692 17492 10471
rect 17548 3137 17588 12496
rect 17931 11696 17973 11705
rect 17931 11656 17932 11696
rect 17972 11656 17973 11696
rect 17931 11647 17973 11656
rect 17835 10436 17877 10445
rect 17835 10396 17836 10436
rect 17876 10396 17877 10436
rect 17835 10387 17877 10396
rect 17836 10302 17876 10387
rect 17644 10228 17780 10268
rect 17644 10184 17684 10228
rect 17740 10184 17780 10228
rect 17740 10144 17876 10184
rect 17644 10135 17684 10144
rect 17836 10100 17876 10144
rect 17836 10060 17879 10100
rect 17839 10016 17879 10060
rect 17836 9976 17879 10016
rect 17739 9932 17781 9941
rect 17739 9892 17740 9932
rect 17780 9892 17781 9932
rect 17739 9883 17781 9892
rect 17740 9512 17780 9883
rect 17836 9521 17876 9976
rect 17932 9941 17972 11647
rect 18028 10361 18068 12907
rect 18027 10352 18069 10361
rect 18027 10312 18028 10352
rect 18068 10312 18069 10352
rect 18027 10303 18069 10312
rect 17931 9932 17973 9941
rect 17931 9892 17932 9932
rect 17972 9892 17973 9932
rect 17931 9883 17973 9892
rect 17931 9680 17973 9689
rect 17931 9640 17932 9680
rect 17972 9640 17973 9680
rect 17931 9631 17973 9640
rect 17932 9546 17972 9631
rect 17740 9463 17780 9472
rect 17835 9512 17877 9521
rect 17835 9472 17836 9512
rect 17876 9472 17877 9512
rect 17835 9463 17877 9472
rect 17836 9344 17876 9463
rect 17740 9304 17876 9344
rect 17740 6488 17780 9304
rect 18027 9176 18069 9185
rect 18027 9136 18028 9176
rect 18068 9136 18069 9176
rect 18027 9127 18069 9136
rect 17932 8000 17972 8009
rect 17932 7328 17972 7960
rect 18028 8000 18068 9127
rect 18124 8840 18164 13075
rect 18220 10445 18260 15688
rect 18316 14981 18356 15772
rect 18315 14972 18357 14981
rect 18315 14932 18316 14972
rect 18356 14932 18357 14972
rect 18315 14923 18357 14932
rect 18412 14804 18452 16015
rect 18892 15569 18932 16024
rect 19083 16024 19084 16064
rect 19124 16024 19125 16064
rect 19083 16015 19125 16024
rect 19179 15980 19221 15989
rect 19179 15940 19180 15980
rect 19220 15940 19221 15980
rect 19179 15931 19221 15940
rect 18891 15560 18933 15569
rect 18891 15520 18892 15560
rect 18932 15520 18933 15560
rect 18891 15511 18933 15520
rect 19180 15317 19220 15931
rect 19276 15905 19316 16108
rect 19371 16064 19413 16073
rect 19371 16024 19372 16064
rect 19412 16024 19413 16064
rect 19371 16015 19413 16024
rect 19275 15896 19317 15905
rect 19275 15856 19276 15896
rect 19316 15856 19317 15896
rect 19275 15847 19317 15856
rect 19372 15728 19412 16015
rect 19276 15688 19412 15728
rect 19179 15308 19221 15317
rect 19179 15268 19180 15308
rect 19220 15268 19221 15308
rect 19179 15259 19221 15268
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 19179 14972 19221 14981
rect 19179 14932 19180 14972
rect 19220 14932 19221 14972
rect 19179 14923 19221 14932
rect 18795 14888 18837 14897
rect 18795 14848 18796 14888
rect 18836 14848 18837 14888
rect 18795 14839 18837 14848
rect 18316 14764 18452 14804
rect 18316 13133 18356 14764
rect 18796 14720 18836 14839
rect 19180 14838 19220 14923
rect 18411 14552 18453 14561
rect 18411 14512 18412 14552
rect 18452 14512 18453 14552
rect 18411 14503 18453 14512
rect 18412 14048 18452 14503
rect 18412 13999 18452 14008
rect 18508 14048 18548 14057
rect 18411 13712 18453 13721
rect 18411 13672 18412 13712
rect 18452 13672 18453 13712
rect 18411 13663 18453 13672
rect 18315 13124 18357 13133
rect 18315 13084 18316 13124
rect 18356 13084 18357 13124
rect 18315 13075 18357 13084
rect 18412 12965 18452 13663
rect 18411 12956 18453 12965
rect 18411 12916 18412 12956
rect 18452 12916 18453 12956
rect 18411 12907 18453 12916
rect 18316 12536 18356 12545
rect 18316 12041 18356 12496
rect 18412 12536 18452 12545
rect 18508 12536 18548 14008
rect 18699 14048 18741 14057
rect 18699 14008 18700 14048
rect 18740 14008 18741 14048
rect 18699 13999 18741 14008
rect 18603 13964 18645 13973
rect 18603 13924 18604 13964
rect 18644 13924 18645 13964
rect 18603 13915 18645 13924
rect 18452 12496 18548 12536
rect 18315 12032 18357 12041
rect 18315 11992 18316 12032
rect 18356 11992 18357 12032
rect 18315 11983 18357 11992
rect 18412 11696 18452 12496
rect 18604 12452 18644 13915
rect 18700 13460 18740 13999
rect 18796 13973 18836 14680
rect 19180 14720 19220 14729
rect 19276 14720 19316 15688
rect 19371 15560 19413 15569
rect 19371 15520 19372 15560
rect 19412 15520 19413 15560
rect 19371 15511 19413 15520
rect 19372 15426 19412 15511
rect 19220 14680 19316 14720
rect 19371 14720 19413 14729
rect 19371 14680 19372 14720
rect 19412 14680 19413 14720
rect 19180 14671 19220 14680
rect 19371 14671 19413 14680
rect 19468 14720 19508 16360
rect 19564 16351 19604 16360
rect 19563 15644 19605 15653
rect 19563 15604 19564 15644
rect 19604 15604 19605 15644
rect 19563 15595 19605 15604
rect 19564 15510 19604 15595
rect 19660 15560 19700 16780
rect 19756 16771 19796 16780
rect 20140 16652 20180 16990
rect 20044 16612 20180 16652
rect 20044 16325 20084 16612
rect 20043 16316 20085 16325
rect 20043 16276 20044 16316
rect 20084 16276 20085 16316
rect 20043 16267 20085 16276
rect 19756 16232 19796 16243
rect 19756 16157 19796 16192
rect 19851 16232 19893 16241
rect 19851 16192 19852 16232
rect 19892 16192 19893 16232
rect 19851 16183 19893 16192
rect 19948 16232 19988 16241
rect 19755 16148 19797 16157
rect 19755 16108 19756 16148
rect 19796 16108 19797 16148
rect 19755 16099 19797 16108
rect 19852 16098 19892 16183
rect 19948 15644 19988 16192
rect 20044 16073 20084 16158
rect 20043 16064 20085 16073
rect 20043 16024 20044 16064
rect 20084 16024 20085 16064
rect 20043 16015 20085 16024
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 20043 15644 20085 15653
rect 19948 15604 20044 15644
rect 20084 15604 20085 15644
rect 20043 15595 20085 15604
rect 19756 15560 19796 15569
rect 19660 15520 19756 15560
rect 19756 15511 19796 15520
rect 19852 15560 19892 15569
rect 19563 15308 19605 15317
rect 19563 15268 19564 15308
rect 19604 15268 19605 15308
rect 19563 15259 19605 15268
rect 19468 14671 19508 14680
rect 19372 14586 19412 14671
rect 18987 14552 19029 14561
rect 18987 14512 18988 14552
rect 19028 14512 19029 14552
rect 18987 14503 19029 14512
rect 18988 14418 19028 14503
rect 18987 14048 19029 14057
rect 18987 14008 18988 14048
rect 19028 14008 19029 14048
rect 18987 13999 19029 14008
rect 19468 14048 19508 14057
rect 18795 13964 18837 13973
rect 18795 13924 18796 13964
rect 18836 13924 18837 13964
rect 18795 13915 18837 13924
rect 18892 13964 18932 13975
rect 18892 13889 18932 13924
rect 18988 13914 19028 13999
rect 18891 13880 18933 13889
rect 18891 13840 18892 13880
rect 18932 13840 18933 13880
rect 18891 13831 18933 13840
rect 19275 13880 19317 13889
rect 19275 13840 19276 13880
rect 19316 13840 19317 13880
rect 19275 13831 19317 13840
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 18700 13420 18932 13460
rect 18796 13208 18836 13217
rect 18796 12881 18836 13168
rect 18795 12872 18837 12881
rect 18795 12832 18796 12872
rect 18836 12832 18837 12872
rect 18795 12823 18837 12832
rect 18795 12620 18837 12629
rect 18795 12580 18796 12620
rect 18836 12580 18837 12620
rect 18795 12571 18837 12580
rect 18796 12536 18836 12571
rect 18796 12485 18836 12496
rect 18892 12536 18932 13420
rect 19276 12629 19316 13831
rect 19275 12620 19317 12629
rect 19275 12580 19276 12620
rect 19316 12580 19317 12620
rect 19275 12571 19317 12580
rect 18508 12412 18644 12452
rect 18508 11705 18548 12412
rect 18892 12368 18932 12496
rect 18604 12328 18932 12368
rect 19372 12536 19412 12545
rect 19468 12536 19508 14008
rect 19412 12496 19508 12536
rect 18316 11656 18452 11696
rect 18507 11696 18549 11705
rect 18507 11656 18508 11696
rect 18548 11656 18549 11696
rect 18219 10436 18261 10445
rect 18219 10396 18220 10436
rect 18260 10396 18261 10436
rect 18219 10387 18261 10396
rect 18316 10193 18356 11656
rect 18507 11647 18549 11656
rect 18508 11562 18548 11647
rect 18604 11201 18644 12328
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18699 12032 18741 12041
rect 18699 11992 18700 12032
rect 18740 11992 18741 12032
rect 18699 11983 18741 11992
rect 18700 11948 18740 11983
rect 18700 11897 18740 11908
rect 19372 11360 19412 12496
rect 19564 11957 19604 15259
rect 19660 14972 19700 14981
rect 19852 14972 19892 15520
rect 20044 15560 20084 15595
rect 20044 15509 20084 15520
rect 19947 15476 19989 15485
rect 19947 15436 19948 15476
rect 19988 15436 19989 15476
rect 19947 15427 19989 15436
rect 19700 14932 19892 14972
rect 19660 14729 19700 14932
rect 19948 14888 19988 15427
rect 20043 15392 20085 15401
rect 20043 15352 20044 15392
rect 20084 15352 20085 15392
rect 20043 15343 20085 15352
rect 20044 15258 20084 15343
rect 19756 14848 19988 14888
rect 19659 14720 19701 14729
rect 19659 14680 19660 14720
rect 19700 14680 19701 14720
rect 19659 14671 19701 14680
rect 19756 14720 19796 14848
rect 19756 14671 19796 14680
rect 19851 14720 19893 14729
rect 19851 14680 19852 14720
rect 19892 14680 19893 14720
rect 19851 14671 19893 14680
rect 19659 14300 19701 14309
rect 19659 14260 19660 14300
rect 19700 14260 19701 14300
rect 19659 14251 19701 14260
rect 19563 11948 19605 11957
rect 19563 11908 19564 11948
rect 19604 11908 19605 11948
rect 19563 11899 19605 11908
rect 19467 11696 19509 11705
rect 19467 11656 19468 11696
rect 19508 11656 19509 11696
rect 19467 11647 19509 11656
rect 19276 11320 19412 11360
rect 18603 11192 18645 11201
rect 18603 11152 18604 11192
rect 18644 11152 18645 11192
rect 18603 11143 18645 11152
rect 18604 10529 18644 11143
rect 19276 11033 19316 11320
rect 18700 11024 18740 11033
rect 18700 10613 18740 10984
rect 19275 11024 19317 11033
rect 19275 10984 19276 11024
rect 19316 10984 19317 11024
rect 19275 10975 19317 10984
rect 18699 10604 18741 10613
rect 18699 10564 18700 10604
rect 18740 10564 18741 10604
rect 18699 10555 18741 10564
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18603 10520 18645 10529
rect 18603 10480 18604 10520
rect 18644 10480 18645 10520
rect 18603 10471 18645 10480
rect 18411 10436 18453 10445
rect 18411 10396 18412 10436
rect 18452 10396 18453 10436
rect 18411 10387 18453 10396
rect 18795 10436 18837 10445
rect 18795 10396 18796 10436
rect 18836 10396 18837 10436
rect 18795 10387 18837 10396
rect 18220 10184 18260 10193
rect 18220 9689 18260 10144
rect 18315 10184 18357 10193
rect 18315 10144 18316 10184
rect 18356 10144 18357 10184
rect 18315 10135 18357 10144
rect 18219 9680 18261 9689
rect 18219 9640 18220 9680
rect 18260 9640 18261 9680
rect 18219 9631 18261 9640
rect 18220 9512 18260 9521
rect 18220 8924 18260 9472
rect 18316 9512 18356 10135
rect 18316 9463 18356 9472
rect 18316 8924 18356 8933
rect 18220 8884 18316 8924
rect 18316 8875 18356 8884
rect 18412 8849 18452 10387
rect 18603 10352 18645 10361
rect 18603 10312 18604 10352
rect 18644 10312 18645 10352
rect 18603 10303 18645 10312
rect 18604 9512 18644 10303
rect 18699 10268 18741 10277
rect 18699 10228 18700 10268
rect 18740 10228 18741 10268
rect 18699 10219 18741 10228
rect 18796 10268 18836 10387
rect 18700 10134 18740 10219
rect 18700 9512 18740 9521
rect 18604 9472 18700 9512
rect 18700 9463 18740 9472
rect 18796 9512 18836 10228
rect 19276 10184 19316 10975
rect 19276 10135 19316 10144
rect 19371 9764 19413 9773
rect 19371 9724 19372 9764
rect 19412 9724 19413 9764
rect 19371 9715 19413 9724
rect 18796 9463 18836 9472
rect 19275 9512 19317 9521
rect 19275 9472 19276 9512
rect 19316 9472 19317 9512
rect 19275 9463 19317 9472
rect 19276 9269 19316 9463
rect 19275 9260 19317 9269
rect 19275 9220 19276 9260
rect 19316 9220 19317 9260
rect 19275 9211 19317 9220
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 18507 8924 18549 8933
rect 18507 8884 18508 8924
rect 18548 8884 18549 8924
rect 18507 8875 18549 8884
rect 18411 8840 18453 8849
rect 18124 8800 18260 8840
rect 18124 8672 18164 8681
rect 18124 8009 18164 8632
rect 18028 7673 18068 7960
rect 18123 8000 18165 8009
rect 18123 7960 18124 8000
rect 18164 7960 18165 8000
rect 18123 7951 18165 7960
rect 18027 7664 18069 7673
rect 18027 7624 18028 7664
rect 18068 7624 18069 7664
rect 18027 7615 18069 7624
rect 18028 7328 18068 7337
rect 17932 7288 18028 7328
rect 18028 7279 18068 7288
rect 17835 7160 17877 7169
rect 17835 7120 17836 7160
rect 17876 7120 17877 7160
rect 17835 7111 17877 7120
rect 17644 6448 17740 6488
rect 17644 4985 17684 6448
rect 17740 6439 17780 6448
rect 17836 5816 17876 7111
rect 18220 6413 18260 8800
rect 18411 8800 18412 8840
rect 18452 8800 18453 8840
rect 18411 8791 18453 8800
rect 18411 8504 18453 8513
rect 18411 8464 18412 8504
rect 18452 8464 18453 8504
rect 18411 8455 18453 8464
rect 18412 8000 18452 8455
rect 18219 6404 18261 6413
rect 18219 6364 18220 6404
rect 18260 6364 18261 6404
rect 18219 6355 18261 6364
rect 17932 6236 17972 6245
rect 17932 5825 17972 6196
rect 18412 5909 18452 7960
rect 18508 8000 18548 8875
rect 18603 8840 18645 8849
rect 18603 8800 18604 8840
rect 18644 8800 18645 8840
rect 18603 8791 18645 8800
rect 18508 7951 18548 7960
rect 18507 7580 18549 7589
rect 18604 7580 18644 8791
rect 18700 8672 18740 8681
rect 18700 8093 18740 8632
rect 18699 8084 18741 8093
rect 18699 8044 18700 8084
rect 18740 8044 18741 8084
rect 18699 8035 18741 8044
rect 18988 8000 19028 8009
rect 18988 7841 19028 7960
rect 18987 7832 19029 7841
rect 18987 7792 18988 7832
rect 19028 7792 19029 7832
rect 18987 7783 19029 7792
rect 19372 7757 19412 9715
rect 19468 8681 19508 11647
rect 19660 11360 19700 14251
rect 19852 13040 19892 14671
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 20043 14216 20085 14225
rect 20140 14216 20180 14225
rect 20043 14176 20044 14216
rect 20084 14176 20140 14216
rect 20043 14167 20085 14176
rect 20140 14167 20180 14176
rect 19996 14038 20036 14047
rect 20036 13998 20276 14034
rect 19996 13994 20276 13998
rect 19996 13989 20036 13994
rect 20043 13880 20085 13889
rect 20043 13840 20044 13880
rect 20084 13840 20085 13880
rect 20043 13831 20085 13840
rect 20044 13208 20084 13831
rect 20236 13460 20276 13994
rect 20236 13411 20276 13420
rect 20044 13159 20084 13168
rect 19564 11320 19700 11360
rect 19756 13000 19892 13040
rect 19467 8672 19509 8681
rect 19467 8632 19468 8672
rect 19508 8632 19509 8672
rect 19467 8623 19509 8632
rect 19468 7986 19508 7995
rect 19371 7748 19413 7757
rect 19371 7708 19372 7748
rect 19412 7708 19413 7748
rect 19371 7699 19413 7708
rect 18507 7540 18508 7580
rect 18548 7540 18644 7580
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18507 7531 18549 7540
rect 18808 7531 19176 7540
rect 18508 6992 18548 7531
rect 19371 7496 19413 7505
rect 19371 7456 19372 7496
rect 19412 7456 19413 7496
rect 19371 7447 19413 7456
rect 18603 7328 18645 7337
rect 18603 7288 18604 7328
rect 18644 7288 18645 7328
rect 18603 7279 18645 7288
rect 18604 7160 18644 7279
rect 18604 7111 18644 7120
rect 18508 6952 18644 6992
rect 18507 6572 18549 6581
rect 18507 6532 18508 6572
rect 18548 6532 18549 6572
rect 18507 6523 18549 6532
rect 18508 6488 18548 6523
rect 18508 6437 18548 6448
rect 18507 6320 18549 6329
rect 18507 6280 18508 6320
rect 18548 6280 18549 6320
rect 18507 6271 18549 6280
rect 18219 5900 18261 5909
rect 18219 5860 18220 5900
rect 18260 5860 18261 5900
rect 18219 5851 18261 5860
rect 18411 5900 18453 5909
rect 18411 5860 18412 5900
rect 18452 5860 18453 5900
rect 18411 5851 18453 5860
rect 17740 5776 17876 5816
rect 17931 5816 17973 5825
rect 17931 5776 17932 5816
rect 17972 5776 17973 5816
rect 17643 4976 17685 4985
rect 17643 4936 17644 4976
rect 17684 4936 17685 4976
rect 17643 4927 17685 4936
rect 17547 3128 17589 3137
rect 17547 3088 17548 3128
rect 17588 3088 17589 3128
rect 17547 3079 17589 3088
rect 17740 2633 17780 5776
rect 17931 5767 17973 5776
rect 17835 5648 17877 5657
rect 17835 5608 17836 5648
rect 17876 5608 17877 5648
rect 17835 5599 17877 5608
rect 17836 5514 17876 5599
rect 18220 4962 18260 5851
rect 18315 5816 18357 5825
rect 18315 5776 18316 5816
rect 18356 5776 18357 5816
rect 18315 5767 18357 5776
rect 18316 5662 18356 5767
rect 18508 5741 18548 6271
rect 18507 5732 18549 5741
rect 18507 5692 18508 5732
rect 18548 5692 18549 5732
rect 18507 5683 18549 5692
rect 18316 5613 18356 5622
rect 18508 5564 18548 5683
rect 18508 5515 18548 5524
rect 18315 5228 18357 5237
rect 18315 5188 18316 5228
rect 18356 5188 18357 5228
rect 18315 5179 18357 5188
rect 18316 5060 18356 5179
rect 18316 5011 18356 5020
rect 18411 5060 18453 5069
rect 18411 5020 18412 5060
rect 18452 5020 18453 5060
rect 18411 5011 18453 5020
rect 18220 4922 18356 4962
rect 18219 4724 18261 4733
rect 18219 4684 18220 4724
rect 18260 4684 18261 4724
rect 18219 4675 18261 4684
rect 17836 4136 17876 4145
rect 17836 2885 17876 4096
rect 17931 4136 17973 4145
rect 17931 4096 17932 4136
rect 17972 4096 18068 4136
rect 17931 4087 17973 4096
rect 17932 4002 17972 4087
rect 17932 3464 17972 3473
rect 17835 2876 17877 2885
rect 17835 2836 17836 2876
rect 17876 2836 17877 2876
rect 17835 2827 17877 2836
rect 17739 2624 17781 2633
rect 17739 2584 17740 2624
rect 17780 2584 17781 2624
rect 17739 2575 17781 2584
rect 17740 1952 17780 2575
rect 17932 2120 17972 3424
rect 18028 3464 18068 4096
rect 18028 3415 18068 3424
rect 18027 3044 18069 3053
rect 18027 3004 18028 3044
rect 18068 3004 18069 3044
rect 18027 2995 18069 3004
rect 17932 2071 17972 2080
rect 17644 1912 17740 1952
rect 17547 1196 17589 1205
rect 17547 1156 17548 1196
rect 17588 1156 17589 1196
rect 17547 1147 17589 1156
rect 17548 1062 17588 1147
rect 17644 1121 17684 1912
rect 17740 1903 17780 1912
rect 18028 1532 18068 2995
rect 17932 1492 18068 1532
rect 17739 1280 17781 1289
rect 17739 1240 17740 1280
rect 17780 1240 17781 1280
rect 17739 1231 17781 1240
rect 17643 1112 17685 1121
rect 17643 1072 17644 1112
rect 17684 1072 17685 1112
rect 17643 1063 17685 1072
rect 17547 944 17589 953
rect 17547 904 17548 944
rect 17588 904 17589 944
rect 17547 895 17589 904
rect 17356 652 17492 692
rect 17163 440 17205 449
rect 17163 400 17164 440
rect 17204 400 17205 440
rect 17163 391 17205 400
rect 16971 272 17013 281
rect 16971 232 16972 272
rect 17012 232 17013 272
rect 16971 223 17013 232
rect 16971 104 17013 113
rect 16971 80 16972 104
rect 7988 64 8008 80
rect 7928 0 8008 64
rect 8120 0 8200 80
rect 8312 0 8392 80
rect 8504 0 8584 80
rect 8696 0 8776 80
rect 8888 0 8968 80
rect 9080 0 9160 80
rect 9272 0 9352 80
rect 9464 0 9544 80
rect 9656 0 9736 80
rect 9848 0 9928 80
rect 10040 0 10120 80
rect 10232 0 10312 80
rect 10424 0 10504 80
rect 10616 0 10696 80
rect 10808 0 10888 80
rect 11000 0 11080 80
rect 11192 0 11272 80
rect 11384 0 11464 80
rect 11576 0 11656 80
rect 11768 0 11848 80
rect 11960 0 12040 80
rect 12152 0 12232 80
rect 12344 0 12424 80
rect 12536 0 12616 80
rect 12728 0 12808 80
rect 12920 0 13000 80
rect 13112 0 13192 80
rect 13304 0 13384 80
rect 13496 0 13576 80
rect 13688 0 13768 80
rect 13880 0 13960 80
rect 14072 0 14152 80
rect 14264 0 14344 80
rect 14456 0 14536 80
rect 14648 0 14728 80
rect 14840 0 14920 80
rect 15032 0 15112 80
rect 15224 0 15304 80
rect 15416 0 15496 80
rect 15608 0 15688 80
rect 15800 0 15880 80
rect 15992 0 16072 80
rect 16184 0 16264 80
rect 16376 0 16456 80
rect 16568 0 16648 80
rect 16760 0 16840 80
rect 16952 64 16972 80
rect 17012 80 17013 104
rect 17164 80 17204 391
rect 17356 80 17396 652
rect 17548 80 17588 895
rect 17644 869 17684 1063
rect 17643 860 17685 869
rect 17643 820 17644 860
rect 17684 820 17685 860
rect 17643 811 17685 820
rect 17740 80 17780 1231
rect 17932 80 17972 1492
rect 18123 1280 18165 1289
rect 18123 1240 18124 1280
rect 18164 1240 18165 1280
rect 18123 1231 18165 1240
rect 18028 944 18068 953
rect 18028 533 18068 904
rect 18027 524 18069 533
rect 18027 484 18028 524
rect 18068 484 18069 524
rect 18027 475 18069 484
rect 18124 80 18164 1231
rect 18220 1196 18260 4675
rect 18316 4220 18356 4922
rect 18316 3380 18356 4180
rect 18412 4220 18452 5011
rect 18412 3548 18452 4180
rect 18508 4962 18548 4971
rect 18508 3725 18548 4922
rect 18507 3716 18549 3725
rect 18507 3676 18508 3716
rect 18548 3676 18549 3716
rect 18507 3667 18549 3676
rect 18412 3508 18548 3548
rect 18508 3464 18548 3508
rect 18508 3415 18548 3424
rect 18412 3380 18452 3389
rect 18316 3340 18412 3380
rect 18412 3331 18452 3340
rect 18507 2876 18549 2885
rect 18507 2836 18508 2876
rect 18548 2836 18549 2876
rect 18507 2827 18549 2836
rect 18508 2742 18548 2827
rect 18316 2633 18356 2718
rect 18315 2624 18357 2633
rect 18315 2584 18316 2624
rect 18356 2584 18357 2624
rect 18315 2575 18357 2584
rect 18604 2540 18644 6952
rect 19275 6236 19317 6245
rect 19275 6196 19276 6236
rect 19316 6196 19317 6236
rect 19275 6187 19317 6196
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 18700 5648 18740 5657
rect 18700 5321 18740 5608
rect 18795 5648 18837 5657
rect 18795 5608 18796 5648
rect 18836 5608 18837 5648
rect 18795 5599 18837 5608
rect 18699 5312 18741 5321
rect 18699 5272 18700 5312
rect 18740 5272 18741 5312
rect 18699 5263 18741 5272
rect 18796 5144 18836 5599
rect 18700 5104 18836 5144
rect 18700 4388 18740 5104
rect 18987 4976 19029 4985
rect 18987 4936 18988 4976
rect 19028 4936 19029 4976
rect 18987 4927 19029 4936
rect 18988 4842 19028 4927
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 18700 4348 18932 4388
rect 18892 4136 18932 4348
rect 18892 3464 18932 4096
rect 19276 3968 19316 6187
rect 19372 4985 19412 7447
rect 19468 6665 19508 7946
rect 19467 6656 19509 6665
rect 19467 6616 19468 6656
rect 19508 6616 19509 6656
rect 19467 6607 19509 6616
rect 19467 5060 19509 5069
rect 19467 5020 19468 5060
rect 19508 5020 19509 5060
rect 19467 5011 19509 5020
rect 19371 4976 19413 4985
rect 19371 4936 19372 4976
rect 19412 4936 19413 4976
rect 19371 4927 19413 4936
rect 19468 4976 19508 5011
rect 19468 4925 19508 4936
rect 19564 4976 19604 11320
rect 19756 10352 19796 13000
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 20044 12620 20084 12631
rect 20044 12545 20084 12580
rect 20043 12536 20085 12545
rect 19900 12494 19940 12503
rect 20043 12496 20044 12536
rect 20084 12496 20085 12536
rect 20043 12487 20085 12496
rect 19900 12452 19940 12454
rect 19900 12412 19988 12452
rect 19851 11696 19893 11705
rect 19851 11656 19852 11696
rect 19892 11656 19893 11696
rect 19851 11647 19893 11656
rect 19852 11024 19892 11647
rect 19948 11192 19988 12412
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20140 11192 20180 11201
rect 19948 11152 20140 11192
rect 20140 11143 20180 11152
rect 19948 11024 19988 11033
rect 19852 10984 19948 11024
rect 19948 10975 19988 10984
rect 19660 10312 19796 10352
rect 19660 9521 19700 10312
rect 19804 10193 19844 10202
rect 19844 10153 19892 10184
rect 19804 10144 19892 10153
rect 19852 9596 19892 10144
rect 19947 10100 19989 10109
rect 19947 10060 19948 10100
rect 19988 10060 19989 10100
rect 19947 10051 19989 10060
rect 19948 9966 19988 10051
rect 20048 9848 20416 9857
rect 19948 9773 19988 9817
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 19947 9764 19989 9773
rect 19947 9724 19948 9764
rect 19988 9724 19989 9764
rect 19947 9722 19989 9724
rect 19947 9715 19948 9722
rect 19988 9715 19989 9722
rect 19948 9673 19988 9682
rect 19852 9556 20084 9596
rect 19659 9512 19701 9521
rect 19659 9472 19660 9512
rect 19700 9472 19701 9512
rect 19659 9463 19701 9472
rect 19804 9470 19844 9479
rect 19804 9428 19844 9430
rect 19804 9388 19892 9428
rect 19755 8672 19797 8681
rect 19755 8632 19756 8672
rect 19796 8632 19797 8672
rect 19755 8623 19797 8632
rect 19659 8168 19701 8177
rect 19659 8128 19660 8168
rect 19700 8128 19701 8168
rect 19659 8119 19701 8128
rect 19660 8034 19700 8119
rect 19756 7169 19796 8623
rect 19852 8168 19892 9388
rect 20044 8924 20084 9556
rect 20140 8924 20180 8933
rect 20044 8884 20140 8924
rect 20140 8875 20180 8884
rect 19947 8672 19989 8681
rect 19947 8632 19948 8672
rect 19988 8632 19989 8672
rect 19947 8623 19989 8632
rect 19948 8538 19988 8623
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19852 8128 20084 8168
rect 19851 8000 19893 8009
rect 19851 7960 19852 8000
rect 19892 7960 19893 8000
rect 19851 7951 19893 7960
rect 19755 7160 19797 7169
rect 19755 7120 19756 7160
rect 19796 7120 19797 7160
rect 19755 7111 19797 7120
rect 19852 7160 19892 7951
rect 20044 7412 20084 8128
rect 20044 7363 20084 7372
rect 19756 6488 19796 7111
rect 19756 6439 19796 6448
rect 19564 4927 19604 4936
rect 19852 5648 19892 7120
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19947 6656 19989 6665
rect 19947 6616 19948 6656
rect 19988 6616 19989 6656
rect 19947 6607 19989 6616
rect 19948 6522 19988 6607
rect 19948 5648 19988 5657
rect 19852 5608 19948 5648
rect 19852 4220 19892 5608
rect 19948 5599 19988 5608
rect 20140 5480 20180 5489
rect 19948 5440 20140 5480
rect 19948 5144 19988 5440
rect 20140 5431 20180 5440
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 19948 5104 20084 5144
rect 19948 4976 19988 4987
rect 19948 4901 19988 4936
rect 20044 4976 20084 5104
rect 20044 4927 20084 4936
rect 19947 4892 19989 4901
rect 19947 4852 19948 4892
rect 19988 4852 19989 4892
rect 19947 4843 19989 4852
rect 19852 4180 19988 4220
rect 19420 4145 19460 4154
rect 19460 4105 19892 4136
rect 19420 4096 19892 4105
rect 19564 3968 19604 3977
rect 19276 3928 19564 3968
rect 19564 3919 19604 3928
rect 19659 3632 19701 3641
rect 19659 3592 19660 3632
rect 19700 3592 19701 3632
rect 19659 3583 19701 3592
rect 19660 3498 19700 3583
rect 18988 3464 19028 3473
rect 18892 3424 18988 3464
rect 18988 3415 19028 3424
rect 19516 3422 19556 3431
rect 19516 3380 19556 3382
rect 19516 3340 19796 3380
rect 18699 3296 18741 3305
rect 18699 3256 18700 3296
rect 18740 3256 18741 3296
rect 18699 3247 18741 3256
rect 18700 2624 18740 3247
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 18796 2624 18836 2633
rect 18700 2584 18796 2624
rect 18796 2575 18836 2584
rect 19563 2624 19605 2633
rect 19563 2584 19564 2624
rect 19604 2584 19605 2624
rect 19563 2575 19605 2584
rect 18604 2500 18740 2540
rect 18412 1952 18452 1961
rect 18700 1952 18740 2500
rect 18452 1912 18740 1952
rect 18412 1903 18452 1912
rect 18411 1784 18453 1793
rect 18411 1744 18412 1784
rect 18452 1744 18453 1784
rect 18411 1735 18453 1744
rect 18220 1147 18260 1156
rect 18315 1196 18357 1205
rect 18315 1156 18316 1196
rect 18356 1156 18357 1196
rect 18315 1147 18357 1156
rect 18316 80 18356 1147
rect 18412 1112 18452 1735
rect 18508 1373 18548 1912
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18507 1364 18549 1373
rect 18507 1324 18508 1364
rect 18548 1324 18549 1364
rect 18507 1315 18549 1324
rect 18699 1280 18741 1289
rect 18699 1240 18700 1280
rect 18740 1240 18741 1280
rect 18699 1231 18741 1240
rect 18412 1063 18452 1072
rect 18507 860 18549 869
rect 18507 820 18508 860
rect 18548 820 18549 860
rect 18507 811 18549 820
rect 18508 80 18548 811
rect 18700 80 18740 1231
rect 19083 1028 19125 1037
rect 19083 988 19084 1028
rect 19124 988 19125 1028
rect 19083 979 19125 988
rect 18891 692 18933 701
rect 18891 652 18892 692
rect 18932 652 18933 692
rect 18891 643 18933 652
rect 18892 80 18932 643
rect 19084 80 19124 979
rect 19564 449 19604 2575
rect 19660 1952 19700 1961
rect 19660 1121 19700 1912
rect 19756 1280 19796 3340
rect 19852 2120 19892 4096
rect 19948 2633 19988 4180
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 20235 3548 20277 3557
rect 20235 3508 20236 3548
rect 20276 3508 20277 3548
rect 20235 3499 20277 3508
rect 20236 2876 20276 3499
rect 20236 2827 20276 2836
rect 19947 2624 19989 2633
rect 20044 2624 20084 2633
rect 19947 2584 19948 2624
rect 19988 2584 20044 2624
rect 19947 2575 19989 2584
rect 20044 2575 20084 2584
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 19852 2071 19892 2080
rect 20235 1868 20277 1877
rect 20235 1828 20236 1868
rect 20276 1828 20277 1868
rect 20235 1819 20277 1828
rect 20236 1734 20276 1819
rect 20044 1700 20084 1709
rect 19948 1660 20044 1700
rect 19852 1280 19892 1289
rect 19756 1240 19852 1280
rect 19852 1231 19892 1240
rect 19659 1112 19701 1121
rect 19659 1072 19660 1112
rect 19700 1072 19701 1112
rect 19659 1063 19701 1072
rect 19660 978 19700 1063
rect 19563 440 19605 449
rect 19563 400 19564 440
rect 19604 400 19605 440
rect 19563 391 19605 400
rect 19948 365 19988 1660
rect 20044 1651 20084 1660
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 19947 356 19989 365
rect 19947 316 19948 356
rect 19988 316 19989 356
rect 19947 307 19989 316
rect 19275 272 19317 281
rect 19275 232 19276 272
rect 19316 232 19317 272
rect 19275 223 19317 232
rect 19276 80 19316 223
rect 19467 188 19509 197
rect 19467 148 19468 188
rect 19508 148 19509 188
rect 19467 139 19509 148
rect 19468 80 19508 139
rect 17012 64 17032 80
rect 16952 0 17032 64
rect 17144 0 17224 80
rect 17336 0 17416 80
rect 17528 0 17608 80
rect 17720 0 17800 80
rect 17912 0 17992 80
rect 18104 0 18184 80
rect 18296 0 18376 80
rect 18488 0 18568 80
rect 18680 0 18760 80
rect 18872 0 18952 80
rect 19064 0 19144 80
rect 19256 0 19336 80
rect 19448 0 19528 80
<< via2 >>
rect 1516 84568 1556 84608
rect 1324 84316 1364 84356
rect 1708 84316 1748 84356
rect 1516 83812 1556 83852
rect 1324 83476 1364 83516
rect 1324 82216 1364 82256
rect 1900 84904 1940 84944
rect 1804 81880 1844 81920
rect 1516 81460 1556 81500
rect 1324 80536 1364 80576
rect 1036 79948 1076 79988
rect 748 79360 788 79400
rect 172 75580 212 75620
rect 76 67768 116 67808
rect 76 67264 116 67304
rect 76 66256 116 66296
rect 460 74908 500 74948
rect 268 71884 308 71924
rect 172 61888 212 61928
rect 364 69700 404 69740
rect 268 60544 308 60584
rect 748 73732 788 73772
rect 1228 79024 1268 79064
rect 1132 78688 1172 78728
rect 1612 80284 1652 80324
rect 1516 79864 1556 79904
rect 1420 79780 1460 79820
rect 1612 79696 1652 79736
rect 1516 79612 1556 79652
rect 1420 79528 1460 79568
rect 1420 78100 1460 78140
rect 1228 77512 1268 77552
rect 1228 75916 1268 75956
rect 1132 74824 1172 74864
rect 1036 73648 1076 73688
rect 1228 73144 1268 73184
rect 1516 76756 1556 76796
rect 2092 85744 2132 85784
rect 2092 83980 2132 84020
rect 2092 81460 2132 81500
rect 1996 80116 2036 80156
rect 1900 79948 1940 79988
rect 1804 79864 1844 79904
rect 2092 79864 2132 79904
rect 1900 79528 1940 79568
rect 1900 78436 1940 78476
rect 1804 77176 1844 77216
rect 1708 76756 1748 76796
rect 1420 76168 1460 76208
rect 1420 75244 1460 75284
rect 1612 76336 1652 76376
rect 1612 75748 1652 75788
rect 1612 75412 1652 75452
rect 1516 74404 1556 74444
rect 1420 72808 1460 72848
rect 1324 71800 1364 71840
rect 1420 71632 1460 71672
rect 1324 71548 1364 71588
rect 1036 70624 1076 70664
rect 1228 70624 1268 70664
rect 940 70288 980 70328
rect 940 66508 980 66548
rect 2092 79696 2132 79736
rect 2380 84988 2420 85028
rect 2284 84316 2324 84356
rect 2668 84484 2708 84524
rect 2572 83896 2612 83936
rect 2860 85324 2900 85364
rect 2860 84316 2900 84356
rect 3052 85156 3092 85196
rect 3052 84400 3092 84440
rect 3340 85324 3380 85364
rect 3244 84988 3284 85028
rect 3244 84736 3284 84776
rect 3916 84988 3956 85028
rect 3724 84904 3764 84944
rect 3532 84652 3572 84692
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 3436 84400 3476 84440
rect 2764 83812 2804 83852
rect 2764 83476 2804 83516
rect 2764 82888 2804 82928
rect 2668 82552 2708 82592
rect 2764 82384 2804 82424
rect 2956 83224 2996 83264
rect 3340 83812 3380 83852
rect 3340 83476 3380 83516
rect 3148 82972 3188 83012
rect 2860 82300 2900 82340
rect 2572 82216 2612 82256
rect 3052 82804 3092 82844
rect 2860 82132 2900 82172
rect 2764 81460 2804 81500
rect 3052 81460 3092 81500
rect 3244 82552 3284 82592
rect 3244 82300 3284 82340
rect 2380 80788 2420 80828
rect 2284 80368 2324 80408
rect 2284 80116 2324 80156
rect 2188 76840 2228 76880
rect 2188 76588 2228 76628
rect 1900 76504 1940 76544
rect 1804 75496 1844 75536
rect 1900 74824 1940 74864
rect 2860 81208 2900 81248
rect 3148 81208 3188 81248
rect 2572 79696 2612 79736
rect 3148 81040 3188 81080
rect 3052 80452 3092 80492
rect 2860 80200 2900 80240
rect 2476 78184 2516 78224
rect 2476 77512 2516 77552
rect 2380 76588 2420 76628
rect 2380 75580 2420 75620
rect 2476 75328 2516 75368
rect 2284 74656 2324 74696
rect 2188 73984 2228 74024
rect 1804 71800 1844 71840
rect 1420 71128 1460 71168
rect 1324 69952 1364 69992
rect 1228 69112 1268 69152
rect 1228 68356 1268 68396
rect 1132 66760 1172 66800
rect 1036 66424 1076 66464
rect 748 65164 788 65204
rect 460 64240 500 64280
rect 652 61300 692 61340
rect 364 60208 404 60248
rect 940 62980 980 63020
rect 844 60964 884 61004
rect 748 59200 788 59240
rect 1036 61720 1076 61760
rect 940 58864 980 58904
rect 652 55336 692 55376
rect 556 55252 596 55292
rect 172 51724 212 51764
rect 556 50884 596 50924
rect 748 51640 788 51680
rect 652 47104 692 47144
rect 940 55168 980 55208
rect 844 50884 884 50924
rect 556 39712 596 39752
rect 556 34000 596 34040
rect 748 33496 788 33536
rect 652 33160 692 33200
rect 172 32992 212 33032
rect 76 32152 116 32192
rect 556 32404 596 32444
rect 364 30976 404 31016
rect 748 28876 788 28916
rect 1420 69532 1460 69572
rect 1804 71380 1844 71420
rect 2092 71632 2132 71672
rect 2092 70624 2132 70664
rect 1900 69532 1940 69572
rect 1900 69364 1940 69404
rect 1516 68356 1556 68396
rect 1420 66256 1460 66296
rect 1516 65584 1556 65624
rect 1420 63988 1460 64028
rect 1420 63736 1460 63776
rect 1324 63652 1364 63692
rect 1708 68440 1748 68480
rect 1804 68356 1844 68396
rect 1612 63736 1652 63776
rect 1516 63232 1556 63272
rect 1516 62812 1556 62852
rect 1420 62728 1460 62768
rect 1228 62224 1268 62264
rect 1516 61216 1556 61256
rect 1708 63148 1748 63188
rect 2092 68188 2132 68228
rect 1996 66172 2036 66212
rect 2380 73900 2420 73940
rect 2668 78100 2708 78140
rect 2668 77260 2708 77300
rect 3052 79528 3092 79568
rect 2956 79360 2996 79400
rect 2860 78940 2900 78980
rect 3724 84232 3764 84272
rect 4300 84400 4340 84440
rect 4396 84064 4436 84104
rect 4108 83896 4148 83936
rect 4300 83560 4340 83600
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 4204 83140 4244 83180
rect 3532 82972 3572 83012
rect 4012 82972 4052 83012
rect 3436 81964 3476 82004
rect 3820 81964 3860 82004
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 4012 81460 4052 81500
rect 3532 81208 3572 81248
rect 3340 81040 3380 81080
rect 3916 81208 3956 81248
rect 3436 80872 3476 80912
rect 3340 80032 3380 80072
rect 4204 81964 4244 82004
rect 4588 84400 4628 84440
rect 5164 84652 5204 84692
rect 5068 84568 5108 84608
rect 5260 84484 5300 84524
rect 4972 84400 5012 84440
rect 4876 84064 4916 84104
rect 5068 84064 5108 84104
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 4780 83308 4820 83348
rect 4972 83560 5012 83600
rect 4684 83140 4724 83180
rect 4876 83140 4916 83180
rect 4588 82720 4628 82760
rect 4876 82888 4916 82928
rect 5356 83224 5396 83264
rect 5836 85240 5876 85280
rect 5644 84904 5684 84944
rect 5644 84484 5684 84524
rect 5548 84232 5588 84272
rect 5548 83812 5588 83852
rect 5548 83224 5588 83264
rect 5452 82972 5492 83012
rect 5164 82888 5204 82928
rect 5452 82804 5492 82844
rect 4972 82720 5012 82760
rect 4492 81964 4532 82004
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 4684 82132 4724 82172
rect 4492 81712 4532 81752
rect 4300 81460 4340 81500
rect 4204 81376 4244 81416
rect 4204 80956 4244 80996
rect 4108 80872 4148 80912
rect 3724 80788 3764 80828
rect 3532 80452 3572 80492
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 4012 79696 4052 79736
rect 3532 79528 3572 79568
rect 3244 78520 3284 78560
rect 2956 77680 2996 77720
rect 2860 77512 2900 77552
rect 2764 76588 2804 76628
rect 2956 77260 2996 77300
rect 2764 75160 2804 75200
rect 2572 74992 2612 75032
rect 2860 74740 2900 74780
rect 3148 78184 3188 78224
rect 4492 80788 4532 80828
rect 4396 80368 4436 80408
rect 4588 80704 4628 80744
rect 4492 80200 4532 80240
rect 4588 79864 4628 79904
rect 3820 78772 3860 78812
rect 3532 78688 3572 78728
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 3532 78352 3572 78392
rect 3436 78184 3476 78224
rect 4780 81880 4820 81920
rect 5164 82132 5204 82172
rect 5164 81460 5204 81500
rect 5356 81880 5396 81920
rect 6124 85240 6164 85280
rect 6028 84400 6068 84440
rect 5932 84148 5972 84188
rect 5740 82300 5780 82340
rect 6220 84988 6260 85028
rect 6988 85660 7028 85700
rect 6796 85576 6836 85616
rect 6796 85408 6836 85448
rect 6796 84568 6836 84608
rect 6412 84400 6452 84440
rect 6604 84400 6644 84440
rect 6988 84316 7028 84356
rect 6220 84064 6260 84104
rect 6700 83896 6740 83936
rect 6220 83560 6260 83600
rect 6220 82804 6260 82844
rect 6412 83140 6452 83180
rect 5932 82132 5972 82172
rect 6700 83308 6740 83348
rect 6892 82972 6932 83012
rect 6796 82720 6836 82760
rect 6796 82384 6836 82424
rect 6604 82132 6644 82172
rect 6700 81964 6740 82004
rect 5548 81292 5588 81332
rect 4780 80872 4820 80912
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 5452 81040 5492 81080
rect 4780 80704 4820 80744
rect 4972 80536 5012 80576
rect 4876 80452 4916 80492
rect 4780 80284 4820 80324
rect 5164 80200 5204 80240
rect 5740 81208 5780 81248
rect 5644 80620 5684 80660
rect 5740 80452 5780 80492
rect 5644 80200 5684 80240
rect 5356 80032 5396 80072
rect 5356 79612 5396 79652
rect 4972 79528 5012 79568
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 4780 79276 4820 79316
rect 5548 79780 5588 79820
rect 5452 79528 5492 79568
rect 4972 79192 5012 79232
rect 3436 77932 3476 77972
rect 3340 77176 3380 77216
rect 3244 76840 3284 76880
rect 3148 76756 3188 76796
rect 3244 76672 3284 76712
rect 3052 76588 3092 76628
rect 3724 77680 3764 77720
rect 3724 77260 3764 77300
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 4492 79024 4532 79064
rect 4492 78772 4532 78812
rect 4204 77512 4244 77552
rect 4684 78100 4724 78140
rect 5068 78940 5108 78980
rect 4876 78436 4916 78476
rect 4972 78184 5012 78224
rect 5068 78100 5108 78140
rect 5260 78520 5300 78560
rect 5836 80032 5876 80072
rect 5740 79864 5780 79904
rect 5740 79612 5780 79652
rect 5644 79108 5684 79148
rect 5644 78688 5684 78728
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 4876 77512 4916 77552
rect 3724 76672 3764 76712
rect 4108 76672 4148 76712
rect 2956 74404 2996 74444
rect 2860 74152 2900 74192
rect 2668 73564 2708 73604
rect 2476 72388 2516 72428
rect 2572 71716 2612 71756
rect 2572 71548 2612 71588
rect 2476 70792 2516 70832
rect 2380 70624 2420 70664
rect 2380 70456 2420 70496
rect 2668 70456 2708 70496
rect 2284 67684 2324 67724
rect 2956 72388 2996 72428
rect 2860 72304 2900 72344
rect 2956 71716 2996 71756
rect 2476 69196 2516 69236
rect 2668 69112 2708 69152
rect 2572 68440 2612 68480
rect 3244 75160 3284 75200
rect 3148 74908 3188 74948
rect 3148 74740 3188 74780
rect 4108 76000 4148 76040
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 4588 77176 4628 77216
rect 4780 77008 4820 77048
rect 4396 76924 4436 76964
rect 4588 76840 4628 76880
rect 4780 76756 4820 76796
rect 5164 77428 5204 77468
rect 4588 76504 4628 76544
rect 4396 76252 4436 76292
rect 4108 75244 4148 75284
rect 3628 75160 3668 75200
rect 3436 74992 3476 75032
rect 3148 74404 3188 74444
rect 3340 74236 3380 74276
rect 3724 75076 3764 75116
rect 4588 75748 4628 75788
rect 4588 75244 4628 75284
rect 4492 75160 4532 75200
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 4972 76084 5012 76124
rect 4876 76000 4916 76040
rect 4972 75832 5012 75872
rect 4876 75244 4916 75284
rect 5644 78184 5684 78224
rect 5548 78100 5588 78140
rect 5452 75076 5492 75116
rect 4876 74992 4916 75032
rect 4492 74824 4532 74864
rect 4300 74404 4340 74444
rect 3628 74236 3668 74276
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 3148 73816 3188 73856
rect 3532 73816 3572 73856
rect 3532 73648 3572 73688
rect 3340 73396 3380 73436
rect 3340 73228 3380 73268
rect 3244 71800 3284 71840
rect 3628 72976 3668 73016
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 3436 72304 3476 72344
rect 4012 72304 4052 72344
rect 3340 71716 3380 71756
rect 3340 71548 3380 71588
rect 3052 70624 3092 70664
rect 3148 70540 3188 70580
rect 3052 69196 3092 69236
rect 2956 68860 2996 68900
rect 2764 68440 2804 68480
rect 2668 68188 2708 68228
rect 2956 67180 2996 67220
rect 2380 66508 2420 66548
rect 2188 64912 2228 64952
rect 1996 63988 2036 64028
rect 1900 63232 1940 63272
rect 1612 60880 1652 60920
rect 1324 60796 1364 60836
rect 1708 60544 1748 60584
rect 1420 58780 1460 58820
rect 1324 58528 1364 58568
rect 1516 57772 1556 57812
rect 1420 57520 1460 57560
rect 1708 57268 1748 57308
rect 1228 57184 1268 57224
rect 1708 57100 1748 57140
rect 1324 56008 1364 56048
rect 1324 55000 1364 55040
rect 1708 56764 1748 56804
rect 1516 55420 1556 55460
rect 1612 55168 1652 55208
rect 1900 60880 1940 60920
rect 1900 56848 1940 56888
rect 2284 62980 2324 63020
rect 2188 62812 2228 62852
rect 2092 60376 2132 60416
rect 3532 71716 3572 71756
rect 4012 71212 4052 71252
rect 3532 71128 3572 71168
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 3532 70624 3572 70664
rect 4300 72304 4340 72344
rect 4300 72136 4340 72176
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 5356 74404 5396 74444
rect 4780 73816 4820 73856
rect 5356 73732 5396 73772
rect 4396 71716 4436 71756
rect 4300 71464 4340 71504
rect 4300 71212 4340 71252
rect 4396 70876 4436 70916
rect 4588 71716 4628 71756
rect 4492 70792 4532 70832
rect 4396 70708 4436 70748
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 4876 72976 4916 73016
rect 4780 72808 4820 72848
rect 5740 77512 5780 77552
rect 5932 79780 5972 79820
rect 5644 74068 5684 74108
rect 5644 73816 5684 73856
rect 5260 72724 5300 72764
rect 4876 72052 4916 72092
rect 5644 73228 5684 73268
rect 5452 72136 5492 72176
rect 5644 73060 5684 73100
rect 5260 71968 5300 72008
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 5356 71716 5396 71756
rect 4684 71464 4724 71504
rect 4876 71296 4916 71336
rect 5356 71296 5396 71336
rect 4780 70792 4820 70832
rect 4300 70540 4340 70580
rect 4204 70456 4244 70496
rect 3436 68524 3476 68564
rect 3340 68440 3380 68480
rect 2572 65416 2612 65456
rect 2860 65584 2900 65624
rect 2956 65416 2996 65456
rect 2668 64660 2708 64700
rect 2668 63988 2708 64028
rect 2572 63904 2612 63944
rect 2572 63148 2612 63188
rect 2860 63232 2900 63272
rect 2668 62980 2708 63020
rect 2476 62560 2516 62600
rect 2572 62308 2612 62348
rect 2764 62140 2804 62180
rect 2956 62644 2996 62684
rect 3148 65248 3188 65288
rect 4012 69868 4052 69908
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 4108 69364 4148 69404
rect 4108 69196 4148 69236
rect 4108 68944 4148 68984
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 3340 66088 3380 66128
rect 4876 70624 4916 70664
rect 4492 70036 4532 70076
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 4396 69364 4436 69404
rect 4300 68944 4340 68984
rect 4204 68860 4244 68900
rect 4204 67096 4244 67136
rect 3532 66760 3572 66800
rect 4108 66760 4148 66800
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 3436 65416 3476 65456
rect 3340 65332 3380 65372
rect 4204 66088 4244 66128
rect 3532 65332 3572 65372
rect 3244 64912 3284 64952
rect 3148 64744 3188 64784
rect 3148 62980 3188 63020
rect 3052 62476 3092 62516
rect 3052 62308 3092 62348
rect 3148 61132 3188 61172
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 3532 64912 3572 64952
rect 3340 64660 3380 64700
rect 3628 64660 3668 64700
rect 3820 64492 3860 64532
rect 3820 64156 3860 64196
rect 3820 63652 3860 63692
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 4492 69196 4532 69236
rect 4684 69112 4724 69152
rect 5164 70120 5204 70160
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 4492 67768 4532 67808
rect 4684 67768 4724 67808
rect 4780 67600 4820 67640
rect 5164 67768 5204 67808
rect 5260 67600 5300 67640
rect 4588 66340 4628 66380
rect 4492 65920 4532 65960
rect 4492 64576 4532 64616
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 5164 67096 5204 67136
rect 5068 66172 5108 66212
rect 4780 65920 4820 65960
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 4684 65080 4724 65120
rect 5260 64492 5300 64532
rect 4588 64324 4628 64364
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 5068 63988 5108 64028
rect 4588 63736 4628 63776
rect 4492 63568 4532 63608
rect 4204 63064 4244 63104
rect 4300 62980 4340 63020
rect 4396 62644 4436 62684
rect 3340 62476 3380 62516
rect 4012 62476 4052 62516
rect 3820 62308 3860 62348
rect 3916 62224 3956 62264
rect 4108 62224 4148 62264
rect 3436 62056 3476 62096
rect 3340 61384 3380 61424
rect 3244 61048 3284 61088
rect 3052 60628 3092 60668
rect 2956 60292 2996 60332
rect 2764 60208 2804 60248
rect 2092 57520 2132 57560
rect 1996 56008 2036 56048
rect 2668 59116 2708 59156
rect 2668 57940 2708 57980
rect 3340 60460 3380 60500
rect 3244 60208 3284 60248
rect 3340 58780 3380 58820
rect 3052 58528 3092 58568
rect 3532 61972 3572 62012
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 4492 62140 4532 62180
rect 4204 61888 4244 61928
rect 4396 61888 4436 61928
rect 4300 61720 4340 61760
rect 3628 61552 3668 61592
rect 3628 61384 3668 61424
rect 3532 60880 3572 60920
rect 4300 60628 4340 60668
rect 3532 60460 3572 60500
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 4108 60124 4148 60164
rect 3628 59956 3668 59996
rect 3820 60040 3860 60080
rect 4300 59956 4340 59996
rect 3724 59284 3764 59324
rect 4204 59284 4244 59324
rect 4204 59116 4244 59156
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 3628 58780 3668 58820
rect 3436 58528 3476 58568
rect 2764 56932 2804 56972
rect 2476 56596 2516 56636
rect 2092 55084 2132 55124
rect 2188 54916 2228 54956
rect 1804 54664 1844 54704
rect 1420 53992 1460 54032
rect 1516 53404 1556 53444
rect 1516 52648 1556 52688
rect 1900 54580 1940 54620
rect 1324 51136 1364 51176
rect 1612 52480 1652 52520
rect 1612 52312 1652 52352
rect 1516 51724 1556 51764
rect 1516 51556 1556 51596
rect 1900 53236 1940 53276
rect 2092 53908 2132 53948
rect 1804 52816 1844 52856
rect 1996 52816 2036 52856
rect 1708 51808 1748 51848
rect 2092 51724 2132 51764
rect 1996 51472 2036 51512
rect 1804 50464 1844 50504
rect 1708 50212 1748 50252
rect 1612 49876 1652 49916
rect 1516 49792 1556 49832
rect 1420 49540 1460 49580
rect 1708 49288 1748 49328
rect 1324 49120 1364 49160
rect 1612 48784 1652 48824
rect 2668 55336 2708 55376
rect 2476 54916 2516 54956
rect 2380 54580 2420 54620
rect 2572 54328 2612 54368
rect 2668 54160 2708 54200
rect 2572 53320 2612 53360
rect 2956 57940 2996 57980
rect 4108 58276 4148 58316
rect 3628 58024 3668 58064
rect 4012 57856 4052 57896
rect 3532 57688 3572 57728
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 3628 57184 3668 57224
rect 3820 57184 3860 57224
rect 3052 56428 3092 56468
rect 2956 56344 2996 56384
rect 3436 56344 3476 56384
rect 3052 55756 3092 55796
rect 3340 56092 3380 56132
rect 3244 55672 3284 55712
rect 3148 55504 3188 55544
rect 3628 56428 3668 56468
rect 4780 63652 4820 63692
rect 4684 63232 4724 63272
rect 4588 62056 4628 62096
rect 5260 63652 5300 63692
rect 5068 63064 5108 63104
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 5068 62560 5108 62600
rect 4588 61384 4628 61424
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 4780 61132 4820 61172
rect 5164 60880 5204 60920
rect 4588 59368 4628 59408
rect 4972 60628 5012 60668
rect 4780 60292 4820 60332
rect 4396 59284 4436 59324
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 5548 69112 5588 69152
rect 5548 68776 5588 68816
rect 6220 80536 6260 80576
rect 6124 79444 6164 79484
rect 6220 79024 6260 79064
rect 6028 78604 6068 78644
rect 7660 85156 7700 85196
rect 7564 84484 7604 84524
rect 7948 85240 7988 85280
rect 7756 84652 7796 84692
rect 7660 84316 7700 84356
rect 7276 83896 7316 83936
rect 7180 83812 7220 83852
rect 7084 83560 7124 83600
rect 7180 83392 7220 83432
rect 7276 82720 7316 82760
rect 7564 83308 7604 83348
rect 7372 82468 7412 82508
rect 7084 82384 7124 82424
rect 7372 82132 7412 82172
rect 7084 82048 7124 82088
rect 7852 84400 7892 84440
rect 8044 84736 8084 84776
rect 7948 83140 7988 83180
rect 7756 82720 7796 82760
rect 7660 82468 7700 82508
rect 6892 80704 6932 80744
rect 7372 81208 7412 81248
rect 6700 79192 6740 79232
rect 6508 79024 6548 79064
rect 6028 78184 6068 78224
rect 6124 77512 6164 77552
rect 6316 76756 6356 76796
rect 6220 76588 6260 76628
rect 5932 75412 5972 75452
rect 6700 78184 6740 78224
rect 6508 78100 6548 78140
rect 6508 77512 6548 77552
rect 6988 80452 7028 80492
rect 7180 80452 7220 80492
rect 7660 80956 7700 80996
rect 7564 80704 7604 80744
rect 7276 80284 7316 80324
rect 6892 79360 6932 79400
rect 6988 79192 7028 79232
rect 7180 79192 7220 79232
rect 6892 79024 6932 79064
rect 7660 80536 7700 80576
rect 7564 80452 7604 80492
rect 7468 80284 7508 80324
rect 7468 79780 7508 79820
rect 7564 79528 7604 79568
rect 7564 79360 7604 79400
rect 6988 78268 7028 78308
rect 6892 78184 6932 78224
rect 7084 77596 7124 77636
rect 7180 77512 7220 77552
rect 7372 78856 7412 78896
rect 7372 78100 7412 78140
rect 7276 77428 7316 77468
rect 6796 77344 6836 77384
rect 7084 76672 7124 76712
rect 6412 75916 6452 75956
rect 6700 76168 6740 76208
rect 6892 76168 6932 76208
rect 6796 76084 6836 76124
rect 6316 75580 6356 75620
rect 6220 75244 6260 75284
rect 5836 74236 5876 74276
rect 5740 72472 5780 72512
rect 5932 74068 5972 74108
rect 5932 73144 5972 73184
rect 5836 72388 5876 72428
rect 5932 72136 5972 72176
rect 5932 71884 5972 71924
rect 6124 72472 6164 72512
rect 6028 71800 6068 71840
rect 6028 71464 6068 71504
rect 6028 69280 6068 69320
rect 6028 69112 6068 69152
rect 6604 75580 6644 75620
rect 6796 75580 6836 75620
rect 6508 75160 6548 75200
rect 6508 74908 6548 74948
rect 6604 74488 6644 74528
rect 7180 76000 7220 76040
rect 7084 75832 7124 75872
rect 6604 73648 6644 73688
rect 6700 73312 6740 73352
rect 6220 71296 6260 71336
rect 6316 70288 6356 70328
rect 6316 69700 6356 69740
rect 5932 68776 5972 68816
rect 6796 72892 6836 72932
rect 6700 72724 6740 72764
rect 6604 72136 6644 72176
rect 6604 70120 6644 70160
rect 7084 75076 7124 75116
rect 7948 81208 7988 81248
rect 7852 80704 7892 80744
rect 7948 80452 7988 80492
rect 7852 79612 7892 79652
rect 8524 84400 8564 84440
rect 8332 83728 8372 83768
rect 8236 83644 8276 83684
rect 8332 83308 8372 83348
rect 8236 83140 8276 83180
rect 8524 84064 8564 84104
rect 8428 83056 8468 83096
rect 8428 82804 8468 82844
rect 8332 82552 8372 82592
rect 8332 82048 8372 82088
rect 8236 80956 8276 80996
rect 8332 80620 8372 80660
rect 8236 79696 8276 79736
rect 8140 79612 8180 79652
rect 8044 79528 8084 79568
rect 7756 79360 7796 79400
rect 7948 79360 7988 79400
rect 8620 83644 8660 83684
rect 8620 83140 8660 83180
rect 8908 84484 8948 84524
rect 9292 85324 9332 85364
rect 9292 84232 9332 84272
rect 9004 83728 9044 83768
rect 8812 83308 8852 83348
rect 8716 83056 8756 83096
rect 8908 82216 8948 82256
rect 8812 81964 8852 82004
rect 8620 80620 8660 80660
rect 7948 79024 7988 79064
rect 7852 78772 7892 78812
rect 7660 78184 7700 78224
rect 8236 78856 8276 78896
rect 8236 78352 8276 78392
rect 7660 77596 7700 77636
rect 8428 79192 8468 79232
rect 8428 78940 8468 78980
rect 8428 78352 8468 78392
rect 9004 81796 9044 81836
rect 9004 81544 9044 81584
rect 8716 79696 8756 79736
rect 9196 82804 9236 82844
rect 8812 79612 8852 79652
rect 8812 79360 8852 79400
rect 8620 79024 8660 79064
rect 8140 77428 8180 77468
rect 8044 77344 8084 77384
rect 7468 76252 7508 76292
rect 8812 78184 8852 78224
rect 8524 77596 8564 77636
rect 9292 81376 9332 81416
rect 9292 81040 9332 81080
rect 9100 79612 9140 79652
rect 9004 78688 9044 78728
rect 9100 78268 9140 78308
rect 9004 77764 9044 77804
rect 8524 76588 8564 76628
rect 7372 76168 7412 76208
rect 7948 76168 7988 76208
rect 7852 76084 7892 76124
rect 8044 76000 8084 76040
rect 7948 75832 7988 75872
rect 7564 74908 7604 74948
rect 7276 74824 7316 74864
rect 7756 74572 7796 74612
rect 8140 75328 8180 75368
rect 8044 74488 8084 74528
rect 7852 74236 7892 74276
rect 7276 73984 7316 74024
rect 7084 73648 7124 73688
rect 7468 73648 7508 73688
rect 6988 73480 7028 73520
rect 7372 73480 7412 73520
rect 7084 73312 7124 73352
rect 6892 71296 6932 71336
rect 6892 70708 6932 70748
rect 6892 70120 6932 70160
rect 6700 69280 6740 69320
rect 5740 67936 5780 67976
rect 5644 67768 5684 67808
rect 5740 66424 5780 66464
rect 5932 66088 5972 66128
rect 5836 65920 5876 65960
rect 5644 65332 5684 65372
rect 5452 64660 5492 64700
rect 5452 64408 5492 64448
rect 5452 63652 5492 63692
rect 5836 65248 5876 65288
rect 5740 64996 5780 65036
rect 5932 64660 5972 64700
rect 5740 64408 5780 64448
rect 5836 63904 5876 63944
rect 6124 67768 6164 67808
rect 6508 68440 6548 68480
rect 6508 66928 6548 66968
rect 6508 66760 6548 66800
rect 6604 66508 6644 66548
rect 6508 66424 6548 66464
rect 6412 66172 6452 66212
rect 6316 65584 6356 65624
rect 6892 69028 6932 69068
rect 7660 73648 7700 73688
rect 8140 73648 8180 73688
rect 8428 76336 8468 76376
rect 8332 76252 8372 76292
rect 8332 75328 8372 75368
rect 7660 73480 7700 73520
rect 7852 73480 7892 73520
rect 8236 73480 8276 73520
rect 7564 73144 7604 73184
rect 7756 72976 7796 73016
rect 8140 73396 8180 73436
rect 7948 73144 7988 73184
rect 7852 72892 7892 72932
rect 7180 72304 7220 72344
rect 7756 71968 7796 72008
rect 7660 71884 7700 71924
rect 7564 71800 7604 71840
rect 7468 71548 7508 71588
rect 7372 71464 7412 71504
rect 7276 69952 7316 69992
rect 7276 69364 7316 69404
rect 7276 68440 7316 68480
rect 7084 67432 7124 67472
rect 6844 66931 6879 66968
rect 6879 66931 6884 66968
rect 6844 66928 6884 66931
rect 7660 71044 7700 71084
rect 7564 69952 7604 69992
rect 7948 71884 7988 71924
rect 7756 70120 7796 70160
rect 7468 69280 7508 69320
rect 7365 67600 7372 67640
rect 7372 67600 7405 67640
rect 7468 67600 7508 67640
rect 7372 67432 7412 67472
rect 7372 67180 7412 67220
rect 7084 66508 7124 66548
rect 6700 66340 6740 66380
rect 7084 66172 7124 66212
rect 6508 65920 6548 65960
rect 6988 65920 7028 65960
rect 6796 65836 6836 65876
rect 6508 65332 6548 65372
rect 6220 64996 6260 65036
rect 6412 64996 6452 65036
rect 6124 64912 6164 64952
rect 6412 64744 6452 64784
rect 6316 64576 6356 64616
rect 6220 64324 6260 64364
rect 6412 64324 6452 64364
rect 6028 63904 6068 63944
rect 5932 63736 5972 63776
rect 5452 62728 5492 62768
rect 4780 59284 4820 59324
rect 5164 59284 5204 59324
rect 5356 59284 5396 59324
rect 4972 59200 5012 59240
rect 4300 58444 4340 58484
rect 4300 57940 4340 57980
rect 4492 57940 4532 57980
rect 4684 58528 4724 58568
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 5068 57940 5108 57980
rect 4300 57688 4340 57728
rect 4204 56260 4244 56300
rect 3724 56092 3764 56132
rect 4108 56092 4148 56132
rect 4492 56092 4532 56132
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 2956 54664 2996 54704
rect 2860 54244 2900 54284
rect 2572 52732 2612 52772
rect 2380 52144 2420 52184
rect 2380 51892 2420 51932
rect 2476 50464 2516 50504
rect 1996 49876 2036 49916
rect 1900 49456 1940 49496
rect 1708 48028 1748 48068
rect 1804 47860 1844 47900
rect 1420 47776 1460 47816
rect 1420 46348 1460 46388
rect 1324 46264 1364 46304
rect 1516 46096 1556 46136
rect 1708 47188 1748 47228
rect 1900 47440 1940 47480
rect 1900 47272 1940 47312
rect 2092 47692 2132 47732
rect 2476 49960 2516 50000
rect 3532 55168 3572 55208
rect 3628 54916 3668 54956
rect 4204 55336 4244 55376
rect 3340 54664 3380 54704
rect 3532 54664 3572 54704
rect 3340 53992 3380 54032
rect 3244 52732 3284 52772
rect 3340 52480 3380 52520
rect 3724 54580 3764 54620
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 3820 54244 3860 54284
rect 4012 54160 4052 54200
rect 3532 53404 3572 53444
rect 4012 53404 4052 53444
rect 2764 51724 2804 51764
rect 2956 51640 2996 51680
rect 2668 50296 2708 50336
rect 2860 50128 2900 50168
rect 2572 48784 2612 48824
rect 2476 48616 2516 48656
rect 2188 47440 2228 47480
rect 2284 46768 2324 46808
rect 2476 46600 2516 46640
rect 2860 46936 2900 46976
rect 1996 45592 2036 45632
rect 1612 45340 1652 45380
rect 1516 45088 1556 45128
rect 1804 45004 1844 45044
rect 1228 44416 1268 44456
rect 1228 41224 1268 41264
rect 1324 38452 1364 38492
rect 1324 38284 1364 38324
rect 1228 37360 1268 37400
rect 1324 37108 1364 37148
rect 1420 36856 1460 36896
rect 1420 36688 1460 36728
rect 1324 36352 1364 36392
rect 1324 34588 1364 34628
rect 1420 33916 1460 33956
rect 1132 33580 1172 33620
rect 1036 33496 1076 33536
rect 1132 33160 1172 33200
rect 940 30892 980 30932
rect 844 27028 884 27068
rect 940 25684 980 25724
rect 556 25264 596 25304
rect 364 23668 404 23708
rect 172 23164 212 23204
rect 76 19216 116 19256
rect 1324 32908 1364 32948
rect 1420 29968 1460 30008
rect 1324 29716 1364 29756
rect 1228 29632 1268 29672
rect 1228 27700 1268 27740
rect 1324 26524 1364 26564
rect 1228 26104 1268 26144
rect 1228 25264 1268 25304
rect 940 18880 980 18920
rect 76 16024 116 16064
rect 1228 22828 1268 22868
rect 1420 25012 1460 25052
rect 1132 21988 1172 22028
rect 1036 13672 1076 13712
rect 844 13168 884 13208
rect 172 10648 212 10688
rect 76 4432 116 4472
rect 1420 21568 1460 21608
rect 1324 21400 1364 21440
rect 1324 19384 1364 19424
rect 1324 19132 1364 19172
rect 1228 18964 1268 19004
rect 1420 18628 1460 18668
rect 1228 16024 1268 16064
rect 1228 15688 1268 15728
rect 1612 44752 1652 44792
rect 2380 45340 2420 45380
rect 2092 44836 2132 44876
rect 2668 45508 2708 45548
rect 2860 45844 2900 45884
rect 3052 51052 3092 51092
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 3820 52732 3860 52772
rect 3532 51724 3572 51764
rect 4204 52480 4244 52520
rect 3820 51808 3860 51848
rect 4108 51640 4148 51680
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 3244 50968 3284 51008
rect 3532 50968 3572 51008
rect 4300 52396 4340 52436
rect 5356 57772 5396 57812
rect 5260 56932 5300 56972
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 5164 56428 5204 56468
rect 4684 56344 4724 56384
rect 5452 55420 5492 55460
rect 5452 55252 5492 55292
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 4684 54832 4724 54872
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 5740 62728 5780 62768
rect 5644 57604 5684 57644
rect 5836 62644 5876 62684
rect 6124 61384 6164 61424
rect 6028 61216 6068 61256
rect 5836 59704 5876 59744
rect 5932 58444 5972 58484
rect 5932 58192 5972 58232
rect 5836 56428 5876 56468
rect 5836 56260 5876 56300
rect 5740 55420 5780 55460
rect 5644 53992 5684 54032
rect 6412 63232 6452 63272
rect 6508 63148 6548 63188
rect 6604 62980 6644 63020
rect 6316 62728 6356 62768
rect 6508 62140 6548 62180
rect 6508 61552 6548 61592
rect 6412 61048 6452 61088
rect 6316 60628 6356 60668
rect 6220 60040 6260 60080
rect 6220 59368 6260 59408
rect 6700 60208 6740 60248
rect 6700 60040 6740 60080
rect 7084 65416 7124 65456
rect 7084 64576 7124 64616
rect 6988 63400 7028 63440
rect 6892 63232 6932 63272
rect 6892 61552 6932 61592
rect 6892 60796 6932 60836
rect 7084 62308 7124 62348
rect 7276 65752 7316 65792
rect 8044 70540 8084 70580
rect 8236 73312 8276 73352
rect 8428 73648 8468 73688
rect 8620 73396 8660 73436
rect 8236 71044 8276 71084
rect 9292 78184 9332 78224
rect 9484 83392 9524 83432
rect 9484 82552 9524 82592
rect 9484 81544 9524 81584
rect 9676 84400 9716 84440
rect 9868 84400 9908 84440
rect 10060 84232 10100 84272
rect 9772 84148 9812 84188
rect 9676 83644 9716 83684
rect 9676 83392 9716 83432
rect 9868 83644 9908 83684
rect 9580 80704 9620 80744
rect 9484 80032 9524 80072
rect 8908 76504 8948 76544
rect 9004 76084 9044 76124
rect 9196 76672 9236 76712
rect 9100 72640 9140 72680
rect 9772 82804 9812 82844
rect 10156 83560 10196 83600
rect 10348 83560 10388 83600
rect 9868 82552 9908 82592
rect 9772 82468 9812 82508
rect 9964 81964 10004 82004
rect 9772 81796 9812 81836
rect 9964 81376 10004 81416
rect 9772 81208 9812 81248
rect 9868 80284 9908 80324
rect 10156 82636 10196 82676
rect 10156 82384 10196 82424
rect 10060 80788 10100 80828
rect 9772 79948 9812 79988
rect 9964 79948 10004 79988
rect 10060 79612 10100 79652
rect 9964 78688 10004 78728
rect 9580 77764 9620 77804
rect 9388 77008 9428 77048
rect 9388 75160 9428 75200
rect 9292 74068 9332 74108
rect 10732 84232 10772 84272
rect 10636 83896 10676 83936
rect 10540 83644 10580 83684
rect 10540 83476 10580 83516
rect 10636 83392 10676 83432
rect 10540 83140 10580 83180
rect 10252 82048 10292 82088
rect 10444 81964 10484 82004
rect 10348 81292 10388 81332
rect 10636 82216 10676 82256
rect 10924 83896 10964 83936
rect 10828 83476 10868 83516
rect 10924 83224 10964 83264
rect 11500 85492 11540 85532
rect 11212 84400 11252 84440
rect 11116 83560 11156 83600
rect 11020 83140 11060 83180
rect 10924 83056 10964 83096
rect 10828 82216 10868 82256
rect 10828 81964 10868 82004
rect 11500 84232 11540 84272
rect 12172 85492 12212 85532
rect 11980 84484 12020 84524
rect 11884 84400 11924 84440
rect 11788 84316 11828 84356
rect 11404 82720 11444 82760
rect 11596 82972 11636 83012
rect 11596 82552 11636 82592
rect 11308 82384 11348 82424
rect 11788 82972 11828 83012
rect 11884 82468 11924 82508
rect 11500 82384 11540 82424
rect 11020 82216 11060 82256
rect 10732 81628 10772 81668
rect 10636 80872 10676 80912
rect 10540 80368 10580 80408
rect 10828 80368 10868 80408
rect 10732 80200 10772 80240
rect 10732 79612 10772 79652
rect 10252 79108 10292 79148
rect 10444 79360 10484 79400
rect 10636 79360 10676 79400
rect 10636 79192 10676 79232
rect 10348 78856 10388 78896
rect 10252 78688 10292 78728
rect 10348 78436 10388 78476
rect 10540 78184 10580 78224
rect 10828 78352 10868 78392
rect 11212 81964 11252 82004
rect 11116 81460 11156 81500
rect 12268 85156 12308 85196
rect 12364 84736 12404 84776
rect 12460 84064 12500 84104
rect 12172 83644 12212 83684
rect 12268 83560 12308 83600
rect 12076 82720 12116 82760
rect 12172 82552 12212 82592
rect 12652 84652 12692 84692
rect 12556 83644 12596 83684
rect 12364 83308 12404 83348
rect 13132 85408 13172 85448
rect 13132 85072 13172 85112
rect 13036 84988 13076 85028
rect 12748 84400 12788 84440
rect 12748 84064 12788 84104
rect 12748 83140 12788 83180
rect 12652 82888 12692 82928
rect 12364 82720 12404 82760
rect 11980 82048 12020 82088
rect 11788 81796 11828 81836
rect 11500 81460 11540 81500
rect 11692 81460 11732 81500
rect 11500 81292 11540 81332
rect 11404 81208 11444 81248
rect 11788 81208 11828 81248
rect 11500 81040 11540 81080
rect 11308 80788 11348 80828
rect 11500 80620 11540 80660
rect 11212 80452 11252 80492
rect 11308 80368 11348 80408
rect 11500 80368 11540 80408
rect 11692 81040 11732 81080
rect 12460 82216 12500 82256
rect 12172 81376 12212 81416
rect 12172 81208 12212 81248
rect 12364 82048 12404 82088
rect 12465 82048 12500 82088
rect 12500 82048 12505 82088
rect 12364 81376 12404 81416
rect 12268 80620 12308 80660
rect 11212 80200 11252 80240
rect 11116 79696 11156 79736
rect 10924 78184 10964 78224
rect 10924 78016 10964 78056
rect 10348 77176 10388 77216
rect 10156 76672 10196 76712
rect 9676 76084 9716 76124
rect 10156 76336 10196 76376
rect 10060 75916 10100 75956
rect 9868 75664 9908 75704
rect 9772 75496 9812 75536
rect 9484 74572 9524 74612
rect 9772 74656 9812 74696
rect 9580 74488 9620 74528
rect 9484 74152 9524 74192
rect 9388 73228 9428 73268
rect 9388 72388 9428 72428
rect 9868 74152 9908 74192
rect 10060 74572 10100 74612
rect 10252 74488 10292 74528
rect 10636 77428 10676 77468
rect 10540 76756 10580 76796
rect 9964 73816 10004 73856
rect 10156 73816 10196 73856
rect 9868 73564 9908 73604
rect 9772 73312 9812 73352
rect 9676 73228 9716 73268
rect 10156 73480 10196 73520
rect 9196 72220 9236 72260
rect 8524 71464 8564 71504
rect 8812 71632 8852 71672
rect 9292 71800 9332 71840
rect 9100 71548 9140 71588
rect 8908 71464 8948 71504
rect 8812 71128 8852 71168
rect 8428 71044 8468 71084
rect 8332 70624 8372 70664
rect 7948 70372 7988 70412
rect 7948 70036 7988 70076
rect 7852 69196 7892 69236
rect 7756 68188 7796 68228
rect 7948 68020 7988 68060
rect 7660 67768 7700 67808
rect 7564 66844 7604 66884
rect 7468 66088 7508 66128
rect 7276 64744 7316 64784
rect 7756 65920 7796 65960
rect 7756 65668 7796 65708
rect 7564 65416 7604 65456
rect 7276 64240 7316 64280
rect 7276 63652 7316 63692
rect 7276 62308 7316 62348
rect 7084 62056 7124 62096
rect 7468 64324 7508 64364
rect 7660 64492 7700 64532
rect 7564 64240 7604 64280
rect 7468 63484 7508 63524
rect 7276 62140 7316 62180
rect 7180 60880 7220 60920
rect 7180 60712 7220 60752
rect 7084 60124 7124 60164
rect 6988 59956 7028 59996
rect 6412 59368 6452 59408
rect 6412 59116 6452 59156
rect 6124 58948 6164 58988
rect 6220 58696 6260 58736
rect 6316 58612 6356 58652
rect 8428 70372 8468 70412
rect 8140 66760 8180 66800
rect 8044 65248 8084 65288
rect 7948 65080 7988 65120
rect 7852 64576 7892 64616
rect 7852 64408 7892 64448
rect 7756 63736 7796 63776
rect 7660 63064 7700 63104
rect 7564 62560 7604 62600
rect 7468 61552 7508 61592
rect 7468 60796 7508 60836
rect 7372 59620 7412 59660
rect 6796 59200 6836 59240
rect 7180 59200 7220 59240
rect 6508 58948 6548 58988
rect 6412 56596 6452 56636
rect 6412 56260 6452 56300
rect 6988 58864 7028 58904
rect 6796 58444 6836 58484
rect 6796 57352 6836 57392
rect 6700 56176 6740 56216
rect 6604 54916 6644 54956
rect 6124 54496 6164 54536
rect 6316 54412 6356 54452
rect 4588 52984 4628 53024
rect 4492 52732 4532 52772
rect 5068 52900 5108 52940
rect 5356 52900 5396 52940
rect 4972 52816 5012 52856
rect 4684 52648 4724 52688
rect 4492 52396 4532 52436
rect 3148 50296 3188 50336
rect 4204 50884 4244 50924
rect 3916 50296 3956 50336
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 5068 51976 5108 52016
rect 4396 51724 4436 51764
rect 4396 51136 4436 51176
rect 4588 51136 4628 51176
rect 4492 50968 4532 51008
rect 4396 50884 4436 50924
rect 4300 50212 4340 50252
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 4108 49708 4148 49748
rect 3820 49204 3860 49244
rect 3340 48784 3380 48824
rect 4012 48532 4052 48572
rect 3244 47944 3284 47984
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 4204 48700 4244 48740
rect 4300 48532 4340 48572
rect 3820 47776 3860 47816
rect 4108 47776 4148 47816
rect 3340 47356 3380 47396
rect 3820 47356 3860 47396
rect 3916 47272 3956 47312
rect 4300 47272 4340 47312
rect 4780 51136 4820 51176
rect 4684 49708 4724 49748
rect 4588 49456 4628 49496
rect 5068 50884 5108 50924
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 4876 50212 4916 50252
rect 4492 49288 4532 49328
rect 4492 47860 4532 47900
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 3148 46684 3188 46724
rect 3052 46516 3092 46556
rect 3436 46516 3476 46556
rect 3244 46432 3284 46472
rect 3340 46180 3380 46220
rect 2764 45172 2804 45212
rect 3244 44920 3284 44960
rect 2476 44332 2516 44372
rect 4108 45760 4148 45800
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 3916 45172 3956 45212
rect 3436 44248 3476 44288
rect 1804 44164 1844 44204
rect 3820 44752 3860 44792
rect 3820 44248 3860 44288
rect 4396 46768 4436 46808
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 5740 53656 5780 53696
rect 5836 53404 5876 53444
rect 5740 53236 5780 53276
rect 5452 52732 5492 52772
rect 5836 51472 5876 51512
rect 5836 51304 5876 51344
rect 5548 50716 5588 50756
rect 5452 50464 5492 50504
rect 5740 50464 5780 50504
rect 5644 49708 5684 49748
rect 5644 49204 5684 49244
rect 5356 48784 5396 48824
rect 4780 48700 4820 48740
rect 4780 48364 4820 48404
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 6124 53992 6164 54032
rect 6028 53404 6068 53444
rect 6220 52144 6260 52184
rect 6028 51724 6068 51764
rect 6124 51472 6164 51512
rect 5932 50968 5972 51008
rect 5932 50128 5972 50168
rect 5932 49708 5972 49748
rect 6124 50296 6164 50336
rect 6028 49456 6068 49496
rect 5836 49288 5876 49328
rect 6028 48196 6068 48236
rect 6028 47608 6068 47648
rect 4396 45760 4436 45800
rect 4300 44416 4340 44456
rect 5548 46516 5588 46556
rect 5356 46180 5396 46220
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 4780 45340 4820 45380
rect 6028 46180 6068 46220
rect 6988 56932 7028 56972
rect 6988 56764 7028 56804
rect 7084 56344 7124 56384
rect 7468 58948 7508 58988
rect 7756 62560 7796 62600
rect 7660 61552 7700 61592
rect 7660 61132 7700 61172
rect 7756 61048 7796 61088
rect 7660 60208 7700 60248
rect 7660 59872 7700 59912
rect 8716 70876 8756 70916
rect 8812 70624 8852 70664
rect 9004 70876 9044 70916
rect 9100 70792 9140 70832
rect 8627 69952 8667 69992
rect 8428 69112 8468 69152
rect 8332 69028 8372 69068
rect 8044 63904 8084 63944
rect 7948 62140 7988 62180
rect 7852 60544 7892 60584
rect 8236 64072 8276 64112
rect 8620 68356 8660 68396
rect 8428 67684 8468 67724
rect 8428 67516 8468 67556
rect 8428 67012 8468 67052
rect 8620 67096 8660 67136
rect 8620 66760 8660 66800
rect 8524 66592 8564 66632
rect 8620 66424 8660 66464
rect 8908 69196 8948 69236
rect 8908 68020 8948 68060
rect 9100 68020 9140 68060
rect 8812 67768 8852 67808
rect 9388 70876 9428 70916
rect 9484 70624 9524 70664
rect 9388 68860 9428 68900
rect 10444 73816 10484 73856
rect 10348 73648 10388 73688
rect 10828 77176 10868 77216
rect 10828 76840 10868 76880
rect 11404 79948 11444 79988
rect 11692 79864 11732 79904
rect 11404 79696 11444 79736
rect 11500 79024 11540 79064
rect 11308 78016 11348 78056
rect 11116 77092 11156 77132
rect 11020 75160 11060 75200
rect 10828 74656 10868 74696
rect 10732 74404 10772 74444
rect 11020 74236 11060 74276
rect 10636 73648 10676 73688
rect 10540 73312 10580 73352
rect 10444 73228 10484 73268
rect 10252 73144 10292 73184
rect 10252 72976 10292 73016
rect 10540 72808 10580 72848
rect 9772 72220 9812 72260
rect 9676 72052 9716 72092
rect 9676 71380 9716 71420
rect 10252 72136 10292 72176
rect 10060 71632 10100 71672
rect 10060 70540 10100 70580
rect 10156 70372 10196 70412
rect 9772 69280 9812 69320
rect 9964 68860 10004 68900
rect 9388 68188 9428 68228
rect 9292 67936 9332 67976
rect 9484 67768 9524 67808
rect 9004 67684 9044 67724
rect 9580 67516 9620 67556
rect 9868 68356 9908 68396
rect 9772 68188 9812 68228
rect 8812 67096 8852 67136
rect 8812 66760 8852 66800
rect 8524 64576 8564 64616
rect 8428 64240 8468 64280
rect 8332 63904 8372 63944
rect 9004 66256 9044 66296
rect 9196 67432 9236 67472
rect 9676 67348 9716 67388
rect 9964 68020 10004 68060
rect 9868 67600 9908 67640
rect 10156 68440 10196 68480
rect 10156 67600 10196 67640
rect 10444 71968 10484 72008
rect 10348 71548 10388 71588
rect 10636 72052 10676 72092
rect 11020 73984 11060 74024
rect 10828 73648 10868 73688
rect 11308 76840 11348 76880
rect 11308 75916 11348 75956
rect 11692 76672 11732 76712
rect 11404 75580 11444 75620
rect 11212 75412 11252 75452
rect 11404 75412 11444 75452
rect 11308 75244 11348 75284
rect 11212 74992 11252 75032
rect 11788 75244 11828 75284
rect 11788 74992 11828 75032
rect 11404 74404 11444 74444
rect 11212 74068 11252 74108
rect 11404 74068 11444 74108
rect 10828 72136 10868 72176
rect 10828 71968 10868 72008
rect 10732 71548 10772 71588
rect 11404 72388 11444 72428
rect 11116 72052 11156 72092
rect 10540 71296 10580 71336
rect 10636 71212 10676 71252
rect 10540 70540 10580 70580
rect 10348 69112 10388 69152
rect 10348 67600 10388 67640
rect 9292 67012 9332 67052
rect 9484 66928 9524 66968
rect 9196 66844 9236 66884
rect 9292 66760 9332 66800
rect 9580 66760 9620 66800
rect 9484 66256 9524 66296
rect 9100 65500 9140 65540
rect 9004 64996 9044 65036
rect 8908 64660 8948 64700
rect 8428 63820 8468 63860
rect 8524 63568 8564 63608
rect 8428 62980 8468 63020
rect 8236 62140 8276 62180
rect 8140 61048 8180 61088
rect 8140 60880 8180 60920
rect 8332 60460 8372 60500
rect 8716 63904 8756 63944
rect 8812 62980 8852 63020
rect 8716 62812 8756 62852
rect 8620 62476 8660 62516
rect 8524 60880 8564 60920
rect 8524 60460 8564 60500
rect 7372 58444 7412 58484
rect 7564 58444 7604 58484
rect 7468 58192 7508 58232
rect 7276 57016 7316 57056
rect 7276 56764 7316 56804
rect 7660 57436 7700 57476
rect 7660 56764 7700 56804
rect 7084 55504 7124 55544
rect 6796 54916 6836 54956
rect 6892 54496 6932 54536
rect 6604 52480 6644 52520
rect 6604 52312 6644 52352
rect 6508 52144 6548 52184
rect 6412 50968 6452 51008
rect 6508 48784 6548 48824
rect 6316 48364 6356 48404
rect 6316 48196 6356 48236
rect 6412 47944 6452 47984
rect 6316 47860 6356 47900
rect 6700 49624 6740 49664
rect 6796 48784 6836 48824
rect 6604 48196 6644 48236
rect 6604 47104 6644 47144
rect 6412 46432 6452 46472
rect 6124 45844 6164 45884
rect 5644 44920 5684 44960
rect 5452 44836 5492 44876
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 5836 44920 5876 44960
rect 6412 45676 6452 45716
rect 4876 44416 4916 44456
rect 5548 44332 5588 44372
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 1612 43744 1652 43784
rect 2476 43408 2516 43448
rect 3436 43408 3476 43448
rect 2188 43324 2228 43364
rect 2092 43156 2132 43196
rect 1804 42316 1844 42356
rect 1612 41224 1652 41264
rect 1708 40048 1748 40088
rect 1612 34336 1652 34376
rect 1996 41140 2036 41180
rect 1900 41056 1940 41096
rect 1804 38284 1844 38324
rect 3532 42988 3572 43028
rect 3148 42820 3188 42860
rect 2764 42736 2804 42776
rect 2764 41980 2804 42020
rect 2284 41392 2324 41432
rect 2572 41308 2612 41348
rect 2092 39964 2132 40004
rect 2284 40384 2324 40424
rect 2668 41224 2708 41264
rect 2572 40384 2612 40424
rect 2668 40216 2708 40256
rect 3436 42736 3476 42776
rect 3724 43072 3764 43112
rect 3724 42904 3764 42944
rect 4012 43240 4052 43280
rect 3916 43156 3956 43196
rect 3628 42736 3668 42776
rect 3052 42484 3092 42524
rect 2956 41980 2996 42020
rect 3052 41896 3092 41936
rect 3244 42484 3284 42524
rect 2956 41812 2996 41852
rect 2860 41224 2900 41264
rect 3916 42736 3956 42776
rect 4108 42736 4148 42776
rect 4204 42568 4244 42608
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 3436 41308 3476 41348
rect 3340 41224 3380 41264
rect 3628 41896 3668 41936
rect 4012 41812 4052 41852
rect 4012 41476 4052 41516
rect 4492 42736 4532 42776
rect 4396 42568 4436 42608
rect 4684 42820 4724 42860
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 5356 43072 5396 43112
rect 4396 42148 4436 42188
rect 4588 41896 4628 41936
rect 3820 41392 3860 41432
rect 3724 41140 3764 41180
rect 4204 41308 4244 41348
rect 3916 41140 3956 41180
rect 3820 41056 3860 41096
rect 4108 41056 4148 41096
rect 3148 40972 3188 41012
rect 2956 40636 2996 40676
rect 2860 40552 2900 40592
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 4396 41224 4436 41264
rect 2860 40384 2900 40424
rect 2476 39880 2516 39920
rect 2956 40132 2996 40172
rect 3148 40048 3188 40088
rect 3340 39880 3380 39920
rect 2476 39544 2516 39584
rect 2380 39376 2420 39416
rect 2188 39124 2228 39164
rect 1900 38200 1940 38240
rect 1804 36856 1844 36896
rect 1804 34924 1844 34964
rect 1804 34000 1844 34040
rect 1708 32908 1748 32948
rect 1612 31396 1652 31436
rect 1708 31144 1748 31184
rect 1996 35176 2036 35216
rect 1996 34840 2036 34880
rect 1996 33664 2036 33704
rect 2764 38872 2804 38912
rect 2668 38788 2708 38828
rect 3148 38956 3188 38996
rect 3052 38872 3092 38912
rect 2956 38032 2996 38072
rect 2860 37612 2900 37652
rect 3148 37612 3188 37652
rect 2572 37528 2612 37568
rect 2860 37192 2900 37232
rect 3340 37528 3380 37568
rect 3148 37024 3188 37064
rect 2668 36520 2708 36560
rect 2476 33916 2516 33956
rect 1804 26776 1844 26816
rect 1708 25348 1748 25388
rect 1708 22492 1748 22532
rect 1612 22408 1652 22448
rect 1708 19888 1748 19928
rect 2092 32152 2132 32192
rect 2476 33748 2516 33788
rect 2284 31564 2324 31604
rect 2668 35176 2708 35216
rect 2956 35176 2996 35216
rect 2860 35008 2900 35048
rect 2860 34168 2900 34208
rect 2572 32068 2612 32108
rect 2476 31648 2516 31688
rect 2668 31564 2708 31604
rect 2572 31480 2612 31520
rect 2380 31228 2420 31268
rect 2476 30472 2516 30512
rect 2668 30556 2708 30596
rect 2572 30304 2612 30344
rect 1996 26272 2036 26312
rect 1996 23836 2036 23876
rect 2380 27868 2420 27908
rect 2572 29380 2612 29420
rect 2572 29128 2612 29168
rect 2668 28288 2708 28328
rect 2860 31480 2900 31520
rect 3052 33748 3092 33788
rect 3244 34672 3284 34712
rect 3148 33412 3188 33452
rect 3052 32152 3092 32192
rect 3340 32824 3380 32864
rect 3628 40468 3668 40508
rect 3532 40216 3572 40256
rect 3916 40552 3956 40592
rect 4108 40468 4148 40508
rect 4300 40552 4340 40592
rect 4204 40384 4244 40424
rect 4492 40804 4532 40844
rect 5548 42988 5588 43028
rect 4876 42652 4916 42692
rect 5260 42400 5300 42440
rect 5452 42400 5492 42440
rect 5260 42232 5300 42272
rect 4876 42148 4916 42188
rect 5260 41980 5300 42020
rect 5356 41728 5396 41768
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 4684 41392 4724 41432
rect 4876 41392 4916 41432
rect 4780 41224 4820 41264
rect 4684 41056 4724 41096
rect 4780 40636 4820 40676
rect 4396 40468 4436 40508
rect 4684 40552 4724 40592
rect 4588 40384 4628 40424
rect 5260 40552 5300 40592
rect 5356 40468 5396 40508
rect 4972 40300 5012 40340
rect 5356 40300 5396 40340
rect 3820 39796 3860 39836
rect 4492 39712 4532 39752
rect 4780 40048 4820 40088
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 4972 39796 5012 39836
rect 4876 39712 4916 39752
rect 4012 39460 4052 39500
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 4108 38956 4148 38996
rect 4396 38956 4436 38996
rect 3628 38872 3668 38912
rect 4204 38704 4244 38744
rect 3532 38620 3572 38660
rect 3916 38200 3956 38240
rect 3916 38032 3956 38072
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3532 37360 3572 37400
rect 4012 37360 4052 37400
rect 4108 37276 4148 37316
rect 4012 36772 4052 36812
rect 4108 36688 4148 36728
rect 4396 37360 4436 37400
rect 4492 37276 4532 37316
rect 4300 36856 4340 36896
rect 4492 36772 4532 36812
rect 4204 36352 4244 36392
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 4588 36520 4628 36560
rect 4492 35680 4532 35720
rect 4012 35428 4052 35468
rect 3724 35260 3764 35300
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 3532 34672 3572 34712
rect 4492 34588 4532 34628
rect 4012 34420 4052 34460
rect 4204 34336 4244 34376
rect 4012 34084 4052 34124
rect 4012 33832 4052 33872
rect 3820 33412 3860 33452
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 4300 33664 4340 33704
rect 4588 33328 4628 33368
rect 4492 32740 4532 32780
rect 3724 32236 3764 32276
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 2956 31312 2996 31352
rect 2860 31228 2900 31268
rect 2956 31060 2996 31100
rect 3148 31060 3188 31100
rect 3052 30724 3092 30764
rect 2860 30472 2900 30512
rect 2956 29884 2996 29924
rect 2860 29716 2900 29756
rect 2860 29044 2900 29084
rect 2956 27952 2996 27992
rect 2764 27196 2804 27236
rect 2956 27616 2996 27656
rect 2956 27280 2996 27320
rect 2476 26776 2516 26816
rect 2860 26776 2900 26816
rect 2476 26440 2516 26480
rect 2380 25516 2420 25556
rect 2476 25432 2516 25472
rect 2476 25180 2516 25220
rect 2188 24592 2228 24632
rect 2188 23920 2228 23960
rect 2092 23248 2132 23288
rect 1900 23080 1940 23120
rect 2188 22576 2228 22616
rect 2380 22492 2420 22532
rect 3436 31312 3476 31352
rect 3340 30724 3380 30764
rect 3340 30556 3380 30596
rect 3532 30556 3572 30596
rect 3148 29968 3188 30008
rect 3148 29296 3188 29336
rect 3148 29044 3188 29084
rect 3916 31312 3956 31352
rect 4396 31312 4436 31352
rect 3820 30976 3860 31016
rect 3820 30556 3860 30596
rect 3436 29548 3476 29588
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 3628 29968 3668 30008
rect 3532 29296 3572 29336
rect 3436 29044 3476 29084
rect 4108 29632 4148 29672
rect 4300 29800 4340 29840
rect 3148 28456 3188 28496
rect 3148 28288 3188 28328
rect 3340 27700 3380 27740
rect 3244 27616 3284 27656
rect 3148 26440 3188 26480
rect 2668 26272 2708 26312
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 3340 27112 3380 27152
rect 4012 28456 4052 28496
rect 3916 28204 3956 28244
rect 4108 28288 4148 28328
rect 4492 30472 4532 30512
rect 4492 28456 4532 28496
rect 3916 27448 3956 27488
rect 3628 27364 3668 27404
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3436 27028 3476 27068
rect 3628 27028 3668 27068
rect 3340 26944 3380 26984
rect 3244 26188 3284 26228
rect 3052 26104 3092 26144
rect 2956 26020 2996 26060
rect 2860 25516 2900 25556
rect 3244 25684 3284 25724
rect 3052 25432 3092 25472
rect 2956 25180 2996 25220
rect 2764 24592 2804 24632
rect 3244 24592 3284 24632
rect 3052 24508 3092 24548
rect 2956 24340 2996 24380
rect 2764 23920 2804 23960
rect 2860 23668 2900 23708
rect 2668 23248 2708 23288
rect 1804 19552 1844 19592
rect 1612 17872 1652 17912
rect 1612 15436 1652 15476
rect 1516 15352 1556 15392
rect 2860 22156 2900 22196
rect 2284 21484 2324 21524
rect 1996 20140 2036 20180
rect 1996 19720 2036 19760
rect 2092 19552 2132 19592
rect 1996 15688 2036 15728
rect 1900 15268 1940 15308
rect 2476 18628 2516 18668
rect 3436 26776 3476 26816
rect 4204 26776 4244 26816
rect 4108 26608 4148 26648
rect 5260 39628 5300 39668
rect 5356 39040 5396 39080
rect 4876 38956 4916 38996
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 4780 38284 4820 38324
rect 5164 38200 5204 38240
rect 5644 42820 5684 42860
rect 5548 41980 5588 42020
rect 5548 41308 5588 41348
rect 5548 38368 5588 38408
rect 5548 38116 5588 38156
rect 7084 53740 7124 53780
rect 7180 52480 7220 52520
rect 6988 47776 7028 47816
rect 6988 47356 7028 47396
rect 7180 50296 7220 50336
rect 7756 56596 7796 56636
rect 7756 55504 7796 55544
rect 7756 54916 7796 54956
rect 7660 54496 7700 54536
rect 7564 53992 7604 54032
rect 7564 52900 7604 52940
rect 7180 49036 7220 49076
rect 7180 48112 7220 48152
rect 7180 47944 7220 47984
rect 7276 47356 7316 47396
rect 7276 45424 7316 45464
rect 7084 45340 7124 45380
rect 6892 45088 6932 45128
rect 8044 58024 8084 58064
rect 8044 57856 8084 57896
rect 7948 57100 7988 57140
rect 7948 55420 7988 55460
rect 8140 57016 8180 57056
rect 8140 56680 8180 56720
rect 8044 55084 8084 55124
rect 8524 59620 8564 59660
rect 8428 59536 8468 59576
rect 8332 59368 8372 59408
rect 8428 57856 8468 57896
rect 9196 65080 9236 65120
rect 9100 64492 9140 64532
rect 9100 64324 9140 64364
rect 9004 62476 9044 62516
rect 8812 61552 8852 61592
rect 8908 61468 8948 61508
rect 8908 60880 8948 60920
rect 8620 59536 8660 59576
rect 8620 59368 8660 59408
rect 8716 58024 8756 58064
rect 8428 57436 8468 57476
rect 8332 57016 8372 57056
rect 8428 56764 8468 56804
rect 8236 56008 8276 56048
rect 8332 55504 8372 55544
rect 8236 55336 8276 55376
rect 8332 55252 8372 55292
rect 8140 54496 8180 54536
rect 8140 54328 8180 54368
rect 7852 53656 7892 53696
rect 8524 56680 8564 56720
rect 8908 58864 8948 58904
rect 8908 58192 8948 58232
rect 8908 57856 8948 57896
rect 9004 57772 9044 57812
rect 8812 57436 8852 57476
rect 8716 55672 8756 55712
rect 8524 55168 8564 55208
rect 7852 52816 7892 52856
rect 7756 51640 7796 51680
rect 8524 53992 8564 54032
rect 8716 53992 8756 54032
rect 8620 53824 8660 53864
rect 8716 53740 8756 53780
rect 8524 53656 8564 53696
rect 8428 52312 8468 52352
rect 8236 51892 8276 51932
rect 7948 51556 7988 51596
rect 7660 51136 7700 51176
rect 7660 50968 7700 51008
rect 7852 51220 7892 51260
rect 8716 53488 8756 53528
rect 8620 53068 8660 53108
rect 8716 52396 8756 52436
rect 8236 51640 8276 51680
rect 7756 50716 7796 50756
rect 7948 50296 7988 50336
rect 7564 49036 7604 49076
rect 7660 48280 7700 48320
rect 7660 47608 7700 47648
rect 8140 49792 8180 49832
rect 8620 51556 8660 51596
rect 8524 51220 8564 51260
rect 8428 50800 8468 50840
rect 8716 51220 8756 51260
rect 8620 50716 8660 50756
rect 8332 49960 8372 50000
rect 7948 49036 7988 49076
rect 8044 48784 8084 48824
rect 7948 48028 7988 48068
rect 7564 47188 7604 47228
rect 7660 46600 7700 46640
rect 8236 48952 8276 48992
rect 8236 47944 8276 47984
rect 8428 49792 8468 49832
rect 8524 49708 8564 49748
rect 8428 48700 8468 48740
rect 8908 52312 8948 52352
rect 9388 65416 9428 65456
rect 9292 64576 9332 64616
rect 9772 67180 9812 67220
rect 9868 67096 9908 67136
rect 9676 65248 9716 65288
rect 9580 65080 9620 65120
rect 9580 64660 9620 64700
rect 9388 64156 9428 64196
rect 9388 63904 9428 63944
rect 9292 63064 9332 63104
rect 9292 62476 9332 62516
rect 9868 64576 9908 64616
rect 10023 64576 10063 64616
rect 10060 64240 10100 64280
rect 9772 64072 9812 64112
rect 9964 63652 10004 63692
rect 9484 63232 9524 63272
rect 9868 63148 9908 63188
rect 9772 63064 9812 63104
rect 9484 62644 9524 62684
rect 9388 61468 9428 61508
rect 9676 61972 9716 62012
rect 9580 61636 9620 61676
rect 9484 59200 9524 59240
rect 9580 58864 9620 58904
rect 9292 58444 9332 58484
rect 9292 57856 9332 57896
rect 9772 61048 9812 61088
rect 9964 62476 10004 62516
rect 10636 70372 10676 70412
rect 10636 68860 10676 68900
rect 10540 66844 10580 66884
rect 10636 66760 10676 66800
rect 10540 66592 10580 66632
rect 10252 65248 10292 65288
rect 10444 65248 10484 65288
rect 10636 66508 10676 66548
rect 10636 65080 10676 65120
rect 10348 64576 10388 64616
rect 10252 64324 10292 64364
rect 10540 64912 10580 64952
rect 10156 63904 10196 63944
rect 10444 63904 10484 63944
rect 10348 63316 10388 63356
rect 10252 63232 10292 63272
rect 10348 63148 10388 63188
rect 10156 63064 10196 63104
rect 10252 62980 10292 63020
rect 10252 62308 10292 62348
rect 10444 62308 10484 62348
rect 10156 61636 10196 61676
rect 10156 61300 10196 61340
rect 9868 60796 9908 60836
rect 9772 60544 9812 60584
rect 10060 60880 10100 60920
rect 10252 60964 10292 61004
rect 10924 70876 10964 70916
rect 10924 70624 10964 70664
rect 11308 71968 11348 72008
rect 11980 79360 12020 79400
rect 12268 80200 12308 80240
rect 12268 79948 12308 79988
rect 12652 82636 12692 82676
rect 12652 82216 12692 82256
rect 12652 81880 12692 81920
rect 12556 81292 12596 81332
rect 12460 80200 12500 80240
rect 12364 79864 12404 79904
rect 12268 79780 12308 79820
rect 12172 79276 12212 79316
rect 12076 79192 12116 79232
rect 12556 79024 12596 79064
rect 12364 78772 12404 78812
rect 12076 78604 12116 78644
rect 12076 78189 12116 78224
rect 12076 78184 12116 78189
rect 12172 78100 12212 78140
rect 12364 78100 12404 78140
rect 11980 75580 12020 75620
rect 11980 75412 12020 75452
rect 11980 75244 12020 75284
rect 12364 77596 12404 77636
rect 12268 77260 12308 77300
rect 12268 76924 12308 76964
rect 12172 76336 12212 76376
rect 12364 76672 12404 76712
rect 12364 76336 12404 76376
rect 12172 75580 12212 75620
rect 11980 74656 12020 74696
rect 11692 72388 11732 72428
rect 11884 72220 11924 72260
rect 11692 72136 11732 72176
rect 11788 71800 11828 71840
rect 11308 71212 11348 71252
rect 11116 70540 11156 70580
rect 11308 70372 11348 70412
rect 11212 70120 11252 70160
rect 11596 71212 11636 71252
rect 11500 70624 11540 70664
rect 11692 70876 11732 70916
rect 12076 74152 12116 74192
rect 12076 73564 12116 73604
rect 12076 71212 12116 71252
rect 12076 70960 12116 71000
rect 11788 70624 11828 70664
rect 11308 69700 11348 69740
rect 10828 69112 10868 69152
rect 11212 69280 11252 69320
rect 10828 68860 10868 68900
rect 11212 68692 11252 68732
rect 11692 69952 11732 69992
rect 11596 69868 11636 69908
rect 11692 69700 11732 69740
rect 11404 68692 11444 68732
rect 11692 66844 11732 66884
rect 11116 66592 11156 66632
rect 11020 66508 11060 66548
rect 10828 66004 10868 66044
rect 11212 66004 11252 66044
rect 10924 65080 10964 65120
rect 10828 64576 10868 64616
rect 10924 64492 10964 64532
rect 10828 63652 10868 63692
rect 10732 63148 10772 63188
rect 10636 63064 10676 63104
rect 10828 62560 10868 62600
rect 10732 61888 10772 61928
rect 10636 61384 10676 61424
rect 10444 61132 10484 61172
rect 9964 59620 10004 59660
rect 10252 59620 10292 59660
rect 10156 59200 10196 59240
rect 9388 57772 9428 57812
rect 9388 57436 9428 57476
rect 9388 57184 9428 57224
rect 9676 58360 9716 58400
rect 10540 60964 10580 61004
rect 10732 60208 10772 60248
rect 10636 59788 10676 59828
rect 10444 59704 10484 59744
rect 10540 59368 10580 59408
rect 10060 58360 10100 58400
rect 9964 57520 10004 57560
rect 9100 52900 9140 52940
rect 9580 56344 9620 56384
rect 9580 56092 9620 56132
rect 9484 55756 9524 55796
rect 9772 57016 9812 57056
rect 9772 56596 9812 56636
rect 10156 57016 10196 57056
rect 10060 56512 10100 56552
rect 9772 56092 9812 56132
rect 9676 54916 9716 54956
rect 10444 58444 10484 58484
rect 10348 56428 10388 56468
rect 10252 56008 10292 56048
rect 10252 55756 10292 55796
rect 10156 55000 10196 55040
rect 9868 54076 9908 54116
rect 9868 53236 9908 53276
rect 9484 52816 9524 52856
rect 9772 52816 9812 52856
rect 9388 52480 9428 52520
rect 9292 51976 9332 52016
rect 9292 51556 9332 51596
rect 10060 53908 10100 53948
rect 10060 51640 10100 51680
rect 9004 50296 9044 50336
rect 9196 50296 9236 50336
rect 8908 49876 8948 49916
rect 9004 49540 9044 49580
rect 9004 49204 9044 49244
rect 8716 48028 8756 48068
rect 8620 47944 8660 47984
rect 8812 47944 8852 47984
rect 9484 49792 9524 49832
rect 9484 49456 9524 49496
rect 9484 49120 9524 49160
rect 9388 48784 9428 48824
rect 8428 46768 8468 46808
rect 7756 45844 7796 45884
rect 8140 45844 8180 45884
rect 7660 45424 7700 45464
rect 7372 45340 7412 45380
rect 7948 44920 7988 44960
rect 6412 43660 6452 43700
rect 7084 43660 7124 43700
rect 6316 43408 6356 43448
rect 6124 41644 6164 41684
rect 5836 41392 5876 41432
rect 5740 40384 5780 40424
rect 5932 40804 5972 40844
rect 5740 40216 5780 40256
rect 6316 41896 6356 41936
rect 6604 43408 6644 43448
rect 6796 43408 6836 43448
rect 6508 42316 6548 42356
rect 6508 41896 6548 41936
rect 6700 42484 6740 42524
rect 6700 41896 6740 41936
rect 6604 41560 6644 41600
rect 6412 41392 6452 41432
rect 7180 43324 7220 43364
rect 6892 43156 6932 43196
rect 6988 42904 7028 42944
rect 6988 42484 7028 42524
rect 6988 42148 7028 42188
rect 6892 41980 6932 42020
rect 6988 41728 7028 41768
rect 7372 43324 7412 43364
rect 7372 42904 7412 42944
rect 7276 42736 7316 42776
rect 7180 42568 7220 42608
rect 7180 42400 7220 42440
rect 7372 42400 7412 42440
rect 7276 41896 7316 41936
rect 7180 41812 7220 41852
rect 7276 41644 7316 41684
rect 8236 44920 8276 44960
rect 8332 44836 8372 44876
rect 8236 43408 8276 43448
rect 7948 43156 7988 43196
rect 7660 42316 7700 42356
rect 8428 43324 8468 43364
rect 8716 46768 8756 46808
rect 9004 46264 9044 46304
rect 8716 45760 8756 45800
rect 8908 45256 8948 45296
rect 9196 45256 9236 45296
rect 10060 50548 10100 50588
rect 9868 50296 9908 50336
rect 9772 50212 9812 50252
rect 10252 51556 10292 51596
rect 10156 50380 10196 50420
rect 10060 50044 10100 50084
rect 10060 49792 10100 49832
rect 9868 49456 9908 49496
rect 9772 49120 9812 49160
rect 9676 49036 9716 49076
rect 10732 59200 10772 59240
rect 10828 58444 10868 58484
rect 11308 65248 11348 65288
rect 11020 64156 11060 64196
rect 11020 63736 11060 63776
rect 11404 64492 11444 64532
rect 11116 62560 11156 62600
rect 11116 61720 11156 61760
rect 11020 61552 11060 61592
rect 11116 61468 11156 61508
rect 11020 61384 11060 61424
rect 11308 63069 11348 63104
rect 11308 63064 11348 63069
rect 11308 61720 11348 61760
rect 11020 60628 11060 60668
rect 11212 60208 11252 60248
rect 11020 60124 11060 60164
rect 11127 60124 11156 60164
rect 11156 60124 11167 60164
rect 11116 59872 11156 59912
rect 11020 59368 11060 59408
rect 11212 59620 11252 59660
rect 11596 65416 11636 65456
rect 12076 70792 12116 70832
rect 12076 70624 12116 70664
rect 12076 70372 12116 70412
rect 11980 70036 12020 70076
rect 12076 69952 12116 69992
rect 12268 72976 12308 73016
rect 12748 81040 12788 81080
rect 12652 75664 12692 75704
rect 13324 84736 13364 84776
rect 13516 84652 13556 84692
rect 13804 85240 13844 85280
rect 13036 84400 13076 84440
rect 13708 84400 13748 84440
rect 13132 84316 13172 84356
rect 13516 84316 13556 84356
rect 12940 84064 12980 84104
rect 12940 82552 12980 82592
rect 13420 84232 13460 84272
rect 13324 84064 13364 84104
rect 13324 83644 13364 83684
rect 13900 84400 13940 84440
rect 14092 84232 14132 84272
rect 13516 84064 13556 84104
rect 13516 83644 13556 83684
rect 13708 84064 13748 84104
rect 13324 83224 13364 83264
rect 13612 83308 13652 83348
rect 13516 82972 13556 83012
rect 13804 83476 13844 83516
rect 14380 85324 14420 85364
rect 14284 83476 14324 83516
rect 14764 85408 14804 85448
rect 14668 85156 14708 85196
rect 14668 84652 14708 84692
rect 14476 84316 14516 84356
rect 14572 83980 14612 84020
rect 13996 83056 14036 83096
rect 14380 83056 14420 83096
rect 13420 82552 13460 82592
rect 14380 82720 14420 82760
rect 14572 82552 14612 82592
rect 14380 81964 14420 82004
rect 14284 81880 14324 81920
rect 13420 80872 13460 80912
rect 13324 80536 13364 80576
rect 13324 79780 13364 79820
rect 13516 80620 13556 80660
rect 13900 81208 13940 81248
rect 13900 80872 13940 80912
rect 13804 80620 13844 80660
rect 13420 78520 13460 78560
rect 13228 78268 13268 78308
rect 13324 78184 13364 78224
rect 13036 77848 13076 77888
rect 13420 76672 13460 76712
rect 13324 76588 13364 76628
rect 12844 75580 12884 75620
rect 13036 75244 13076 75284
rect 12556 75160 12596 75200
rect 12460 74824 12500 74864
rect 12556 74488 12596 74528
rect 12460 73144 12500 73184
rect 12364 71800 12404 71840
rect 12364 71548 12404 71588
rect 12268 71464 12308 71504
rect 12364 70960 12404 71000
rect 12268 70876 12308 70916
rect 12460 70792 12500 70832
rect 13516 76420 13556 76460
rect 13420 76000 13460 76040
rect 13516 75916 13556 75956
rect 13516 75328 13556 75368
rect 13612 75244 13652 75284
rect 12844 74488 12884 74528
rect 13132 74488 13172 74528
rect 13420 73900 13460 73940
rect 12940 73564 12980 73604
rect 12652 72892 12692 72932
rect 12844 72640 12884 72680
rect 13132 73648 13172 73688
rect 13612 74488 13652 74528
rect 13516 73648 13556 73688
rect 14284 80452 14324 80492
rect 14380 79444 14420 79484
rect 13900 79360 13940 79400
rect 14572 81712 14612 81752
rect 14476 79276 14516 79316
rect 13804 79024 13844 79064
rect 14380 79024 14420 79064
rect 14092 78940 14132 78980
rect 13900 78688 13940 78728
rect 13804 78352 13844 78392
rect 13996 78184 14036 78224
rect 13900 78100 13940 78140
rect 13900 75664 13940 75704
rect 13804 75076 13844 75116
rect 13708 74068 13748 74108
rect 13708 73732 13748 73772
rect 13516 73060 13556 73100
rect 13132 72892 13172 72932
rect 13612 72976 13652 73016
rect 13516 72808 13556 72848
rect 13420 72136 13460 72176
rect 13996 75580 14036 75620
rect 13996 74908 14036 74948
rect 13900 74656 13940 74696
rect 13996 74320 14036 74360
rect 13900 73900 13940 73940
rect 13804 73144 13844 73184
rect 13996 73480 14036 73520
rect 13900 73060 13940 73100
rect 13804 72976 13844 73016
rect 13036 71884 13076 71924
rect 12652 71548 12692 71588
rect 12748 70792 12788 70832
rect 12844 70624 12884 70664
rect 12652 70456 12692 70496
rect 11980 69700 12020 69740
rect 11980 67684 12020 67724
rect 12172 69700 12212 69740
rect 12076 66844 12116 66884
rect 12460 69112 12500 69152
rect 12364 68188 12404 68228
rect 12364 67936 12404 67976
rect 12364 67684 12404 67724
rect 12268 66928 12308 66968
rect 12556 68692 12596 68732
rect 12556 67936 12596 67976
rect 12844 69196 12884 69236
rect 12556 66928 12596 66968
rect 12460 66508 12500 66548
rect 12364 66340 12404 66380
rect 12364 65668 12404 65708
rect 12172 65416 12212 65456
rect 11788 64324 11828 64364
rect 11500 64240 11540 64280
rect 11500 64072 11540 64112
rect 11596 63904 11636 63944
rect 12460 64240 12500 64280
rect 12076 64072 12116 64112
rect 12364 64072 12404 64112
rect 11596 63484 11636 63524
rect 11884 63316 11924 63356
rect 11884 63064 11924 63104
rect 11500 62728 11540 62768
rect 11404 61216 11444 61256
rect 11596 60208 11636 60248
rect 11596 59956 11636 59996
rect 11020 59200 11060 59240
rect 11020 58780 11060 58820
rect 11020 57184 11060 57224
rect 11020 57016 11060 57056
rect 10540 55672 10580 55712
rect 10540 51976 10580 52016
rect 10636 51808 10676 51848
rect 10444 51724 10484 51764
rect 10348 50884 10388 50924
rect 10348 50296 10388 50336
rect 10636 50548 10676 50588
rect 10444 49624 10484 49664
rect 10156 49372 10196 49412
rect 9868 47692 9908 47732
rect 9772 46852 9812 46892
rect 9676 46684 9716 46724
rect 10540 49464 10580 49496
rect 10540 49456 10580 49464
rect 10636 49036 10676 49076
rect 10348 48784 10388 48824
rect 10636 48784 10676 48824
rect 10252 48280 10292 48320
rect 11308 58864 11348 58904
rect 11212 58528 11252 58568
rect 11404 58780 11444 58820
rect 11404 57940 11444 57980
rect 11308 57436 11348 57476
rect 11500 56764 11540 56804
rect 11308 56680 11348 56720
rect 11596 56680 11636 56720
rect 11404 56596 11444 56636
rect 11308 56512 11348 56552
rect 11212 56428 11252 56468
rect 11308 56176 11348 56216
rect 11500 56176 11540 56216
rect 10828 51640 10868 51680
rect 10828 50296 10868 50336
rect 11884 62812 11924 62852
rect 12076 62812 12116 62852
rect 11788 61384 11828 61424
rect 11788 61132 11828 61172
rect 11788 59956 11828 59996
rect 11788 59452 11828 59492
rect 12364 63232 12404 63272
rect 12172 62728 12212 62768
rect 12172 62140 12212 62180
rect 11980 61720 12020 61760
rect 12460 62980 12500 63020
rect 12748 67012 12788 67052
rect 12652 66592 12692 66632
rect 13228 71800 13268 71840
rect 13420 71968 13460 72008
rect 13420 71800 13460 71840
rect 13132 71464 13172 71504
rect 13036 70792 13076 70832
rect 13036 68188 13076 68228
rect 13420 71632 13460 71672
rect 13324 71464 13364 71504
rect 13324 70960 13364 71000
rect 13228 69952 13268 69992
rect 13228 69280 13268 69320
rect 13228 68524 13268 68564
rect 13420 69952 13460 69992
rect 13804 71968 13844 72008
rect 13420 69028 13460 69068
rect 13324 68272 13364 68312
rect 13228 67432 13268 67472
rect 12940 67096 12980 67136
rect 13036 66592 13076 66632
rect 12844 65668 12884 65708
rect 12748 64324 12788 64364
rect 13036 64996 13076 65036
rect 12652 64240 12692 64280
rect 12844 64240 12884 64280
rect 12364 62308 12404 62348
rect 12268 61552 12308 61592
rect 12172 61216 12212 61256
rect 12556 62140 12596 62180
rect 12460 61216 12500 61256
rect 12268 60376 12308 60416
rect 11980 59536 12020 59576
rect 11980 59200 12020 59240
rect 12076 56932 12116 56972
rect 11980 56764 12020 56804
rect 11788 56512 11828 56552
rect 11692 56176 11732 56216
rect 11884 56344 11924 56384
rect 12364 59704 12404 59744
rect 12844 63988 12884 64028
rect 12748 63736 12788 63776
rect 12940 62056 12980 62096
rect 13036 61804 13076 61844
rect 12844 61132 12884 61172
rect 12748 61048 12788 61088
rect 13036 60796 13076 60836
rect 12652 60292 12692 60332
rect 12652 60124 12692 60164
rect 12556 60040 12596 60080
rect 12652 59872 12692 59912
rect 13036 60628 13076 60668
rect 12844 59536 12884 59576
rect 13036 59536 13076 59576
rect 12364 58528 12404 58568
rect 12364 57772 12404 57812
rect 12268 57184 12308 57224
rect 12268 56932 12308 56972
rect 12268 56680 12308 56720
rect 11116 55924 11156 55964
rect 11020 55672 11060 55712
rect 11308 54916 11348 54956
rect 11308 54160 11348 54200
rect 11116 53908 11156 53948
rect 11116 53656 11156 53696
rect 11596 55504 11636 55544
rect 11596 54076 11636 54116
rect 11404 53908 11444 53948
rect 11404 53740 11444 53780
rect 11308 53656 11348 53696
rect 11212 53488 11252 53528
rect 11788 55924 11828 55964
rect 11788 55504 11828 55544
rect 12172 55588 12212 55628
rect 11212 53236 11252 53276
rect 11020 52900 11060 52940
rect 11116 52648 11156 52688
rect 11020 52480 11060 52520
rect 11116 51892 11156 51932
rect 11020 51808 11060 51848
rect 11308 53152 11348 53192
rect 11212 50884 11252 50924
rect 11212 50380 11252 50420
rect 11116 50296 11156 50336
rect 11020 49456 11060 49496
rect 10828 49372 10868 49412
rect 10156 47272 10196 47312
rect 10060 47104 10100 47144
rect 9964 46852 10004 46892
rect 9964 46684 10004 46724
rect 9964 45256 10004 45296
rect 8620 44836 8660 44876
rect 8524 43156 8564 43196
rect 8428 43072 8468 43112
rect 8236 42400 8276 42440
rect 8428 42736 8468 42776
rect 7852 42232 7892 42272
rect 7564 41896 7604 41936
rect 7468 41644 7508 41684
rect 7756 41896 7796 41936
rect 7660 41728 7700 41768
rect 7852 41728 7892 41768
rect 7756 41560 7796 41600
rect 8428 42232 8468 42272
rect 8236 42148 8276 42188
rect 8044 41896 8084 41936
rect 8236 41812 8276 41852
rect 8140 41728 8180 41768
rect 7372 41392 7412 41432
rect 7564 41392 7604 41432
rect 6700 41056 6740 41096
rect 6508 40804 6548 40844
rect 6316 40720 6356 40760
rect 6028 40300 6068 40340
rect 6892 40804 6932 40844
rect 6988 40636 7028 40676
rect 7372 41056 7412 41096
rect 7468 40636 7508 40676
rect 7372 40552 7412 40592
rect 7276 40468 7316 40508
rect 6796 40384 6836 40424
rect 7276 40300 7316 40340
rect 6700 39880 6740 39920
rect 7276 39880 7316 39920
rect 8044 41392 8084 41432
rect 7948 41308 7988 41348
rect 7660 40468 7700 40508
rect 7468 40384 7508 40424
rect 7852 40552 7892 40592
rect 7948 40384 7988 40424
rect 8236 41560 8276 41600
rect 8332 41476 8372 41516
rect 8428 41392 8468 41432
rect 8716 42736 8756 42776
rect 8716 41728 8756 41768
rect 8716 41560 8756 41600
rect 8620 41392 8660 41432
rect 8332 41308 8372 41348
rect 9580 45004 9620 45044
rect 9388 44248 9428 44288
rect 9388 43492 9428 43532
rect 9964 44248 10004 44288
rect 9100 42736 9140 42776
rect 9196 42568 9236 42608
rect 9100 42484 9140 42524
rect 9388 42568 9428 42608
rect 9100 41728 9140 41768
rect 9004 41560 9044 41600
rect 8908 41476 8948 41516
rect 9484 41728 9524 41768
rect 9292 41644 9332 41684
rect 9868 41812 9908 41852
rect 9676 41560 9716 41600
rect 9292 41392 9332 41432
rect 8716 41224 8756 41264
rect 8428 40888 8468 40928
rect 8620 40888 8660 40928
rect 8332 40636 8372 40676
rect 8236 40216 8276 40256
rect 7852 40132 7892 40172
rect 7756 39964 7796 40004
rect 6508 39712 6548 39752
rect 6892 39712 6932 39752
rect 6508 39292 6548 39332
rect 6988 39544 7028 39584
rect 6892 39040 6932 39080
rect 6028 38536 6068 38576
rect 6220 38116 6260 38156
rect 6220 37780 6260 37820
rect 5452 37696 5492 37736
rect 5836 37612 5876 37652
rect 5740 37528 5780 37568
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 5260 36688 5300 36728
rect 5260 35680 5300 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 6412 38872 6452 38912
rect 7372 39712 7412 39752
rect 7660 39880 7700 39920
rect 8044 40048 8084 40088
rect 7948 39880 7988 39920
rect 7564 39292 7604 39332
rect 6988 38788 7028 38828
rect 6796 38200 6836 38240
rect 7468 38620 7508 38660
rect 5452 36856 5492 36896
rect 6028 37360 6068 37400
rect 5740 36688 5780 36728
rect 5644 36604 5684 36644
rect 5452 36520 5492 36560
rect 5452 36100 5492 36140
rect 6412 37360 6452 37400
rect 6220 37192 6260 37232
rect 6412 37024 6452 37064
rect 6796 37528 6836 37568
rect 7084 37192 7124 37232
rect 6700 37024 6740 37064
rect 6220 36772 6260 36812
rect 6316 36688 6356 36728
rect 6316 36436 6356 36476
rect 6028 36268 6068 36308
rect 5836 36100 5876 36140
rect 5644 35680 5684 35720
rect 5452 35344 5492 35384
rect 4972 34924 5012 34964
rect 4972 34336 5012 34376
rect 5260 35176 5300 35216
rect 5260 34840 5300 34880
rect 5452 35176 5492 35216
rect 5932 35848 5972 35888
rect 6412 36100 6452 36140
rect 5932 35344 5972 35384
rect 5644 34840 5684 34880
rect 6028 35260 6068 35300
rect 6124 35176 6164 35216
rect 5836 35092 5876 35132
rect 5548 34672 5588 34712
rect 5836 34672 5876 34712
rect 5452 34504 5492 34544
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 6412 35176 6452 35216
rect 6316 35092 6356 35132
rect 6220 35008 6260 35048
rect 6220 34756 6260 34796
rect 5836 34336 5876 34376
rect 5740 33748 5780 33788
rect 6316 34504 6356 34544
rect 6028 34168 6068 34208
rect 6220 34084 6260 34124
rect 6124 33832 6164 33872
rect 6028 33664 6068 33704
rect 5932 32908 5972 32948
rect 5836 32824 5876 32864
rect 5932 32656 5972 32696
rect 5740 31816 5780 31856
rect 5644 31648 5684 31688
rect 5548 31564 5588 31604
rect 5452 31480 5492 31520
rect 4684 31396 4724 31436
rect 5068 31228 5108 31268
rect 4684 30976 4724 31016
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4780 30808 4820 30848
rect 5260 30808 5300 30848
rect 5644 31396 5684 31436
rect 5548 30640 5588 30680
rect 5836 30976 5876 31016
rect 5740 30640 5780 30680
rect 5068 30472 5108 30512
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 4684 28624 4724 28664
rect 4684 28036 4724 28076
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4588 27700 4628 27740
rect 4492 26440 4532 26480
rect 3820 26104 3860 26144
rect 3532 25768 3572 25808
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 3532 25012 3572 25052
rect 3436 24928 3476 24968
rect 3916 24760 3956 24800
rect 3532 24592 3572 24632
rect 4300 26104 4340 26144
rect 4300 25432 4340 25472
rect 4492 25264 4532 25304
rect 4300 24424 4340 24464
rect 3724 24340 3764 24380
rect 4204 24340 4244 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3532 24004 3572 24044
rect 3340 23584 3380 23624
rect 3244 21568 3284 21608
rect 3148 20728 3188 20768
rect 2668 20056 2708 20096
rect 2764 19216 2804 19256
rect 2668 18124 2708 18164
rect 2476 17704 2516 17744
rect 2092 15604 2132 15644
rect 1708 14428 1748 14468
rect 1420 13168 1460 13208
rect 1420 13000 1460 13040
rect 1804 14176 1844 14216
rect 2092 13588 2132 13628
rect 1612 13252 1652 13292
rect 1996 13084 2036 13124
rect 1708 12412 1748 12452
rect 1804 12244 1844 12284
rect 1708 11068 1748 11108
rect 1516 10144 1556 10184
rect 1516 9976 1556 10016
rect 1324 9892 1364 9932
rect 1132 8716 1172 8756
rect 1420 9808 1460 9848
rect 1420 8464 1460 8504
rect 1228 7960 1268 8000
rect 1324 7876 1364 7916
rect 1132 7792 1172 7832
rect 1036 7120 1076 7160
rect 844 6784 884 6824
rect 172 1744 212 1784
rect 1228 6448 1268 6488
rect 1612 9388 1652 9428
rect 1612 7456 1652 7496
rect 1420 5188 1460 5228
rect 1420 3676 1460 3716
rect 1132 2164 1172 2204
rect 1324 3508 1364 3548
rect 1900 11824 1940 11864
rect 1900 11152 1940 11192
rect 2092 12412 2132 12452
rect 2092 12076 2132 12116
rect 2284 14512 2324 14552
rect 2668 17620 2708 17660
rect 2668 16780 2708 16820
rect 3532 23584 3572 23624
rect 4012 23584 4052 23624
rect 3724 23164 3764 23204
rect 3724 22996 3764 23036
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 4012 22492 4052 22532
rect 4300 22072 4340 22112
rect 4012 21652 4052 21692
rect 3628 21484 3668 21524
rect 3436 19468 3476 19508
rect 2860 16612 2900 16652
rect 2476 15352 2516 15392
rect 2476 14596 2516 14636
rect 2380 13588 2420 13628
rect 2476 12580 2516 12620
rect 2188 11992 2228 12032
rect 2188 11152 2228 11192
rect 1996 10396 2036 10436
rect 1804 9388 1844 9428
rect 1996 9388 2036 9428
rect 1900 9136 1940 9176
rect 1804 8128 1844 8168
rect 1708 6196 1748 6236
rect 1708 4432 1748 4472
rect 1996 8044 2036 8084
rect 2188 10480 2228 10520
rect 2284 9640 2324 9680
rect 2476 11992 2516 12032
rect 2476 11824 2516 11864
rect 2764 15940 2804 15980
rect 2860 15520 2900 15560
rect 3244 19216 3284 19256
rect 3148 18796 3188 18836
rect 3148 17368 3188 17408
rect 3340 18460 3380 18500
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 4012 20812 4052 20852
rect 3724 19972 3764 20012
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3628 19468 3668 19508
rect 3532 19048 3572 19088
rect 4012 19216 4052 19256
rect 4012 18796 4052 18836
rect 4204 21568 4244 21608
rect 4684 26104 4724 26144
rect 5356 27700 5396 27740
rect 4876 27616 4916 27656
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 5164 24592 5204 24632
rect 5260 24508 5300 24548
rect 5164 23752 5204 23792
rect 5260 23668 5300 23708
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 5548 30220 5588 30260
rect 5740 29632 5780 29672
rect 5740 28960 5780 29000
rect 5740 28540 5780 28580
rect 6124 31228 6164 31268
rect 6028 30976 6068 31016
rect 5836 28372 5876 28412
rect 5644 28288 5684 28328
rect 5548 28204 5588 28244
rect 5548 27700 5588 27740
rect 5548 27364 5588 27404
rect 5452 25348 5492 25388
rect 5836 28120 5876 28160
rect 5740 27280 5780 27320
rect 5740 26524 5780 26564
rect 6124 30640 6164 30680
rect 6796 36856 6836 36896
rect 6604 36772 6644 36812
rect 6604 36436 6644 36476
rect 6700 36268 6740 36308
rect 6988 36100 7028 36140
rect 6604 36016 6644 36056
rect 7468 37276 7508 37316
rect 7468 37108 7508 37148
rect 7276 36688 7316 36728
rect 7660 39124 7700 39164
rect 7756 38956 7796 38996
rect 7852 38872 7892 38912
rect 7660 38032 7700 38072
rect 7660 36940 7700 36980
rect 7564 36856 7604 36896
rect 7948 37528 7988 37568
rect 6700 35764 6740 35804
rect 6604 35680 6644 35720
rect 6988 35596 7028 35636
rect 6604 34840 6644 34880
rect 7756 36604 7796 36644
rect 7372 35596 7412 35636
rect 7180 35344 7220 35384
rect 7564 35848 7604 35888
rect 7756 35848 7796 35888
rect 7468 35260 7508 35300
rect 7084 35176 7124 35216
rect 6700 34672 6740 34712
rect 6508 34588 6548 34628
rect 7180 34504 7220 34544
rect 6700 34252 6740 34292
rect 6796 34168 6836 34208
rect 6508 34000 6548 34040
rect 6508 33748 6548 33788
rect 6604 33496 6644 33536
rect 6604 33244 6644 33284
rect 6508 32824 6548 32864
rect 7084 34336 7124 34376
rect 7660 34840 7700 34880
rect 7180 34084 7220 34124
rect 7564 34336 7604 34376
rect 7660 34252 7700 34292
rect 7564 34000 7604 34040
rect 7468 33832 7508 33872
rect 7276 33664 7316 33704
rect 6988 33076 7028 33116
rect 6604 31480 6644 31520
rect 6412 31396 6452 31436
rect 6508 31312 6548 31352
rect 6220 30556 6260 30596
rect 6124 30472 6164 30512
rect 6604 30976 6644 31016
rect 6604 30304 6644 30344
rect 6508 30220 6548 30260
rect 6028 29128 6068 29168
rect 7180 32908 7220 32948
rect 7660 33748 7700 33788
rect 7372 32824 7412 32864
rect 7852 33664 7892 33704
rect 7852 33412 7892 33452
rect 7084 32740 7124 32780
rect 6892 31984 6932 32024
rect 6796 31816 6836 31856
rect 6796 31480 6836 31520
rect 6796 30220 6836 30260
rect 6700 30136 6740 30176
rect 6604 29464 6644 29504
rect 6700 29296 6740 29336
rect 6412 29044 6452 29084
rect 6988 31900 7028 31940
rect 7468 32656 7508 32696
rect 6988 31564 7028 31604
rect 6892 29464 6932 29504
rect 8140 39376 8180 39416
rect 8524 40468 8564 40508
rect 9004 41224 9044 41264
rect 9196 41224 9236 41264
rect 8908 40636 8948 40676
rect 8908 40468 8948 40508
rect 8812 40384 8852 40424
rect 9100 40552 9140 40592
rect 9292 41140 9332 41180
rect 9004 40216 9044 40256
rect 8428 40048 8468 40088
rect 8332 39880 8372 39920
rect 8524 39880 8564 39920
rect 8428 39796 8468 39836
rect 8908 40048 8948 40088
rect 8524 39628 8564 39668
rect 8332 38872 8372 38912
rect 8140 37192 8180 37232
rect 8140 36856 8180 36896
rect 8044 33160 8084 33200
rect 7948 33076 7988 33116
rect 8332 37444 8372 37484
rect 8332 37192 8372 37232
rect 8428 36100 8468 36140
rect 8428 35680 8468 35720
rect 8620 38872 8660 38912
rect 9292 40384 9332 40424
rect 9292 40216 9332 40256
rect 9580 40972 9620 41012
rect 10444 46936 10484 46976
rect 10252 46348 10292 46388
rect 10252 45844 10292 45884
rect 10348 45592 10388 45632
rect 10444 45088 10484 45128
rect 11020 49120 11060 49160
rect 10924 47944 10964 47984
rect 11212 49204 11252 49244
rect 11212 48868 11252 48908
rect 11212 48700 11252 48740
rect 11212 47860 11252 47900
rect 11020 47608 11060 47648
rect 10924 47272 10964 47312
rect 10828 47188 10868 47228
rect 10924 46432 10964 46472
rect 10924 45592 10964 45632
rect 10636 44920 10676 44960
rect 10060 41644 10100 41684
rect 10252 41560 10292 41600
rect 9772 41308 9812 41348
rect 9964 41308 10004 41348
rect 9868 41224 9908 41264
rect 9772 40972 9812 41012
rect 9484 40384 9524 40424
rect 9676 40636 9716 40676
rect 10252 41224 10292 41264
rect 10060 40720 10100 40760
rect 9964 40636 10004 40676
rect 9868 40552 9908 40592
rect 10060 40552 10100 40592
rect 9580 40216 9620 40256
rect 9484 40048 9524 40088
rect 9196 39628 9236 39668
rect 9772 39628 9812 39668
rect 9580 39544 9620 39584
rect 9676 39292 9716 39332
rect 9292 38452 9332 38492
rect 8716 37612 8756 37652
rect 8716 37360 8756 37400
rect 8620 35260 8660 35300
rect 8524 34336 8564 34376
rect 8908 36604 8948 36644
rect 9580 37528 9620 37568
rect 10924 43492 10964 43532
rect 11116 42148 11156 42188
rect 11116 41896 11156 41936
rect 11692 52060 11732 52100
rect 11980 54244 12020 54284
rect 11884 52984 11924 53024
rect 11500 51304 11540 51344
rect 11788 51220 11828 51260
rect 11404 51052 11444 51092
rect 11404 50548 11444 50588
rect 11404 49120 11444 49160
rect 11788 51052 11828 51092
rect 11692 50632 11732 50672
rect 11596 48784 11636 48824
rect 11596 48196 11636 48236
rect 11404 47356 11444 47396
rect 12364 56176 12404 56216
rect 12364 55588 12404 55628
rect 12364 55420 12404 55460
rect 12268 54244 12308 54284
rect 12076 53488 12116 53528
rect 12172 53236 12212 53276
rect 11980 52228 12020 52268
rect 12076 51640 12116 51680
rect 12268 51556 12308 51596
rect 12172 51052 12212 51092
rect 12076 50968 12116 51008
rect 11980 50548 12020 50588
rect 11884 50044 11924 50084
rect 12268 50716 12308 50756
rect 12364 50548 12404 50588
rect 12652 59368 12692 59408
rect 12748 58360 12788 58400
rect 12652 58024 12692 58064
rect 12556 57352 12596 57392
rect 12556 56428 12596 56468
rect 12556 56176 12596 56216
rect 12556 55924 12596 55964
rect 12748 57940 12788 57980
rect 12652 53656 12692 53696
rect 12652 53152 12692 53192
rect 13228 66676 13268 66716
rect 13228 66340 13268 66380
rect 13612 67684 13652 67724
rect 13516 63904 13556 63944
rect 13324 63652 13364 63692
rect 13516 62140 13556 62180
rect 13324 61888 13364 61928
rect 13228 60544 13268 60584
rect 13228 60040 13268 60080
rect 13132 58024 13172 58064
rect 13420 61216 13460 61256
rect 13324 57940 13364 57980
rect 13132 57856 13172 57896
rect 13804 68944 13844 68984
rect 13804 68272 13844 68312
rect 13708 63988 13748 64028
rect 13708 63652 13748 63692
rect 13708 62056 13748 62096
rect 13612 60712 13652 60752
rect 13516 59032 13556 59072
rect 13996 72052 14036 72092
rect 13996 71548 14036 71588
rect 14188 78772 14228 78812
rect 14284 78604 14324 78644
rect 14188 78100 14228 78140
rect 14476 76672 14516 76712
rect 14860 84064 14900 84104
rect 14956 83560 14996 83600
rect 15244 84736 15284 84776
rect 15340 84232 15380 84272
rect 15148 83812 15188 83852
rect 15052 83476 15092 83516
rect 14764 83056 14804 83096
rect 14956 82720 14996 82760
rect 14764 81964 14804 82004
rect 15052 81964 15092 82004
rect 14956 81880 14996 81920
rect 15052 81628 15092 81668
rect 15052 81208 15092 81248
rect 14860 80704 14900 80744
rect 14764 80200 14804 80240
rect 14668 78940 14708 78980
rect 14668 77680 14708 77720
rect 15244 83560 15284 83600
rect 15436 83896 15476 83936
rect 16012 84820 16052 84860
rect 15820 84568 15860 84608
rect 15628 83308 15668 83348
rect 15532 82720 15572 82760
rect 15628 82468 15668 82508
rect 15244 81628 15284 81668
rect 15436 81040 15476 81080
rect 14956 79780 14996 79820
rect 15148 79612 15188 79652
rect 14860 78772 14900 78812
rect 14956 78352 14996 78392
rect 16204 84736 16244 84776
rect 16108 83812 16148 83852
rect 15820 83476 15860 83516
rect 15916 83392 15956 83432
rect 15820 82972 15860 83012
rect 16012 83308 16052 83348
rect 16300 83308 16340 83348
rect 16012 83140 16052 83180
rect 16108 82468 16148 82508
rect 16204 82300 16244 82340
rect 16204 82048 16244 82088
rect 15628 80704 15668 80744
rect 15628 80536 15668 80576
rect 15532 80284 15572 80324
rect 15532 79696 15572 79736
rect 15436 79276 15476 79316
rect 15340 79108 15380 79148
rect 15244 78268 15284 78308
rect 14956 78184 14996 78224
rect 15340 78184 15380 78224
rect 15628 79192 15668 79232
rect 15532 79024 15572 79064
rect 14668 77008 14708 77048
rect 14764 76756 14804 76796
rect 14380 76504 14420 76544
rect 14380 75664 14420 75704
rect 14476 74488 14516 74528
rect 14284 73480 14324 73520
rect 14284 72976 14324 73016
rect 14188 71884 14228 71924
rect 14188 71716 14228 71756
rect 14188 70456 14228 70496
rect 14092 69280 14132 69320
rect 14668 76672 14708 76712
rect 14668 74740 14708 74780
rect 14764 73732 14804 73772
rect 15436 78100 15476 78140
rect 15628 78604 15668 78644
rect 15052 77260 15092 77300
rect 15244 76840 15284 76880
rect 15052 75916 15092 75956
rect 15820 80536 15860 80576
rect 16108 81040 16148 81080
rect 15820 80284 15860 80324
rect 15916 80116 15956 80156
rect 15820 79612 15860 79652
rect 15820 79444 15860 79484
rect 15916 79360 15956 79400
rect 15916 79024 15956 79064
rect 15820 78520 15860 78560
rect 16012 78688 16052 78728
rect 15916 78184 15956 78224
rect 15916 77680 15956 77720
rect 15436 76252 15476 76292
rect 15436 76084 15476 76124
rect 15340 75496 15380 75536
rect 15916 76840 15956 76880
rect 16588 83560 16628 83600
rect 16492 83224 16532 83264
rect 16492 81796 16532 81836
rect 16396 81040 16436 81080
rect 16588 81460 16628 81500
rect 16972 84400 17012 84440
rect 16780 84232 16820 84272
rect 17068 84064 17108 84104
rect 16972 83644 17012 83684
rect 16780 83140 16820 83180
rect 16780 82384 16820 82424
rect 16972 80872 17012 80912
rect 16300 80620 16340 80660
rect 16396 80284 16436 80324
rect 16300 80200 16340 80240
rect 16300 80032 16340 80072
rect 16396 79948 16436 79988
rect 16492 79864 16532 79904
rect 16300 79612 16340 79652
rect 16204 79024 16244 79064
rect 16492 79192 16532 79232
rect 16396 78520 16436 78560
rect 16396 78352 16436 78392
rect 16300 77680 16340 77720
rect 15628 76000 15668 76040
rect 15916 76084 15956 76124
rect 15340 75160 15380 75200
rect 15052 74740 15092 74780
rect 14668 72136 14708 72176
rect 14572 72052 14612 72092
rect 14380 71548 14420 71588
rect 14572 71464 14612 71504
rect 14380 70876 14420 70916
rect 14572 70876 14612 70916
rect 14284 69952 14324 69992
rect 14188 69112 14228 69152
rect 14188 68440 14228 68480
rect 14476 69112 14516 69152
rect 14284 68356 14324 68396
rect 14668 70036 14708 70076
rect 15148 74572 15188 74612
rect 15052 72136 15092 72176
rect 15532 74992 15572 75032
rect 15916 75160 15956 75200
rect 16108 76084 16148 76124
rect 15820 74992 15860 75032
rect 16012 74236 16052 74276
rect 15340 73816 15380 73856
rect 15244 73144 15284 73184
rect 15436 72808 15476 72848
rect 16204 74320 16244 74360
rect 16108 73732 16148 73772
rect 15724 72808 15764 72848
rect 15340 72388 15380 72428
rect 15244 72304 15284 72344
rect 15244 72136 15284 72176
rect 15148 71380 15188 71420
rect 15052 70876 15092 70916
rect 14956 70708 14996 70748
rect 15244 70876 15284 70916
rect 15148 70708 15188 70748
rect 15244 70624 15284 70664
rect 15148 70540 15188 70580
rect 14764 69364 14804 69404
rect 14956 70036 14996 70076
rect 15436 71968 15476 72008
rect 15916 72892 15956 72932
rect 15628 71464 15668 71504
rect 15820 71464 15860 71504
rect 15724 71380 15764 71420
rect 15436 71296 15476 71336
rect 15820 70876 15860 70916
rect 15532 70540 15572 70580
rect 14668 68944 14708 68984
rect 15436 70120 15476 70160
rect 14572 68524 14612 68564
rect 14092 66088 14132 66128
rect 14572 65836 14612 65876
rect 14188 65080 14228 65120
rect 13900 64576 13940 64616
rect 14092 63064 14132 63104
rect 13996 62980 14036 63020
rect 13900 61804 13940 61844
rect 13804 60460 13844 60500
rect 13996 61468 14036 61508
rect 13900 60376 13940 60416
rect 13900 60040 13940 60080
rect 13708 58864 13748 58904
rect 13708 58696 13748 58736
rect 13708 57940 13748 57980
rect 13420 57016 13460 57056
rect 13420 56680 13460 56720
rect 13612 56764 13652 56804
rect 12940 55840 12980 55880
rect 12940 55420 12980 55460
rect 13516 55336 13556 55376
rect 13420 55252 13460 55292
rect 12844 54160 12884 54200
rect 13228 53908 13268 53948
rect 12844 53656 12884 53696
rect 13228 53320 13268 53360
rect 13324 53236 13364 53276
rect 12940 52480 12980 52520
rect 13324 52480 13364 52520
rect 12844 51976 12884 52016
rect 12748 51136 12788 51176
rect 11980 49624 12020 49664
rect 11884 48784 11924 48824
rect 13036 52060 13076 52100
rect 12940 50296 12980 50336
rect 13708 53320 13748 53360
rect 13612 52984 13652 53024
rect 13516 52396 13556 52436
rect 13516 51724 13556 51764
rect 13036 50212 13076 50252
rect 13804 52900 13844 52940
rect 13804 51976 13844 52016
rect 13804 51640 13844 51680
rect 14092 60964 14132 61004
rect 14092 60712 14132 60752
rect 14092 60460 14132 60500
rect 14092 59368 14132 59408
rect 14092 57772 14132 57812
rect 13996 57352 14036 57392
rect 14092 57184 14132 57224
rect 13996 56596 14036 56636
rect 13708 51136 13748 51176
rect 13228 50212 13268 50252
rect 13516 50212 13556 50252
rect 13420 50128 13460 50168
rect 12652 49876 12692 49916
rect 13036 49876 13076 49916
rect 11980 48700 12020 48740
rect 11788 48364 11828 48404
rect 11692 47104 11732 47144
rect 11404 46096 11444 46136
rect 11308 42652 11348 42692
rect 11308 42400 11348 42440
rect 11212 41812 11252 41852
rect 10540 41728 10580 41768
rect 10444 41224 10484 41264
rect 11308 41644 11348 41684
rect 10636 41560 10676 41600
rect 11020 41392 11060 41432
rect 10732 41308 10772 41348
rect 10924 41224 10964 41264
rect 11212 41224 11252 41264
rect 11020 41140 11060 41180
rect 10828 40804 10868 40844
rect 10444 40636 10484 40676
rect 10348 40552 10388 40592
rect 10252 40468 10292 40508
rect 10156 40384 10196 40424
rect 10348 40384 10388 40424
rect 10252 40216 10292 40256
rect 9868 39544 9908 39584
rect 10924 40636 10964 40676
rect 10636 40132 10676 40172
rect 10732 39964 10772 40004
rect 10540 39796 10580 39836
rect 10348 39712 10388 39752
rect 9772 38872 9812 38912
rect 9964 38788 10004 38828
rect 9964 38368 10004 38408
rect 9292 36268 9332 36308
rect 9292 35932 9332 35972
rect 9196 35680 9236 35720
rect 9004 35176 9044 35216
rect 8908 34672 8948 34712
rect 8812 34336 8852 34376
rect 9004 34336 9044 34376
rect 8716 34000 8756 34040
rect 9004 34000 9044 34040
rect 8236 33832 8276 33872
rect 8428 33748 8468 33788
rect 8716 33748 8756 33788
rect 8236 33160 8276 33200
rect 7276 31312 7316 31352
rect 7276 30220 7316 30260
rect 7660 31144 7700 31184
rect 6988 29380 7028 29420
rect 7564 29884 7604 29924
rect 7276 29296 7316 29336
rect 6988 29044 7028 29084
rect 6508 28960 6548 29000
rect 6220 28708 6260 28748
rect 6124 28540 6164 28580
rect 6028 28456 6068 28496
rect 6028 28120 6068 28160
rect 5932 28036 5972 28076
rect 6028 27700 6068 27740
rect 6124 27616 6164 27656
rect 7084 28708 7124 28748
rect 7372 28456 7412 28496
rect 6604 28372 6644 28412
rect 6412 28288 6452 28328
rect 6412 28120 6452 28160
rect 6220 27028 6260 27068
rect 6316 26776 6356 26816
rect 6508 28036 6548 28076
rect 6700 28288 6740 28328
rect 6796 28120 6836 28160
rect 7564 28708 7604 28748
rect 6604 26944 6644 26984
rect 6028 26104 6068 26144
rect 5932 25852 5972 25892
rect 5836 25768 5876 25808
rect 6124 26020 6164 26060
rect 6124 25852 6164 25892
rect 5740 25264 5780 25304
rect 6124 25432 6164 25472
rect 6316 26524 6356 26564
rect 6700 26776 6740 26816
rect 6988 27616 7028 27656
rect 7276 27952 7316 27992
rect 7372 27700 7412 27740
rect 7180 27364 7220 27404
rect 6892 27028 6932 27068
rect 7276 26944 7316 26984
rect 6892 26860 6932 26900
rect 6796 26608 6836 26648
rect 6604 26524 6644 26564
rect 6508 26356 6548 26396
rect 6412 26104 6452 26144
rect 6316 25768 6356 25808
rect 5644 25180 5684 25220
rect 5548 24592 5588 24632
rect 5932 25012 5972 25052
rect 5740 24592 5780 24632
rect 5452 23752 5492 23792
rect 5356 23332 5396 23372
rect 4972 23248 5012 23288
rect 5452 23248 5492 23288
rect 4780 22576 4820 22616
rect 5356 23080 5396 23120
rect 5644 23836 5684 23876
rect 4972 22744 5012 22784
rect 5164 22576 5204 22616
rect 4876 22324 4916 22364
rect 4684 22156 4724 22196
rect 5260 22408 5300 22448
rect 5548 22828 5588 22868
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 5644 22744 5684 22784
rect 6124 24928 6164 24968
rect 6604 25852 6644 25892
rect 6508 25768 6548 25808
rect 6316 25096 6356 25136
rect 6220 24760 6260 24800
rect 6028 24508 6068 24548
rect 6316 24172 6356 24212
rect 6988 26776 7028 26816
rect 7180 26608 7220 26648
rect 7084 26524 7124 26564
rect 7468 27532 7508 27572
rect 7468 26944 7508 26984
rect 7468 26776 7508 26816
rect 7084 26104 7124 26144
rect 6892 25768 6932 25808
rect 7084 25432 7124 25472
rect 6700 25096 6740 25136
rect 6892 25096 6932 25136
rect 5932 23836 5972 23876
rect 5836 23752 5876 23792
rect 6124 23752 6164 23792
rect 5932 23248 5972 23288
rect 6124 23248 6164 23288
rect 6316 23080 6356 23120
rect 5836 22240 5876 22280
rect 5836 22072 5876 22112
rect 5740 21568 5780 21608
rect 5548 21400 5588 21440
rect 5740 21148 5780 21188
rect 5164 20560 5204 20600
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 6028 21568 6068 21608
rect 6028 21400 6068 21440
rect 4780 20308 4820 20348
rect 4492 19972 4532 20012
rect 4492 19804 4532 19844
rect 4396 19300 4436 19340
rect 4300 19216 4340 19256
rect 4684 18880 4724 18920
rect 3628 18460 3668 18500
rect 3436 17620 3476 17660
rect 3340 17368 3380 17408
rect 3244 17200 3284 17240
rect 3052 16444 3092 16484
rect 3148 16360 3188 16400
rect 3340 16948 3380 16988
rect 3436 16780 3476 16820
rect 3340 16612 3380 16652
rect 3244 15940 3284 15980
rect 3148 15268 3188 15308
rect 3052 15184 3092 15224
rect 3052 15016 3092 15056
rect 2668 14176 2708 14216
rect 2860 13924 2900 13964
rect 2764 13336 2804 13376
rect 2764 12832 2804 12872
rect 2764 12076 2804 12116
rect 2572 11572 2612 11612
rect 2476 11404 2516 11444
rect 2572 10984 2612 11024
rect 2668 10396 2708 10436
rect 2092 7960 2132 8000
rect 2380 8968 2420 9008
rect 2572 9808 2612 9848
rect 2956 12916 2996 12956
rect 3244 15100 3284 15140
rect 3244 14680 3284 14720
rect 3244 14092 3284 14132
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3820 17032 3860 17072
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3532 16444 3572 16484
rect 3724 16360 3764 16400
rect 3532 16276 3572 16316
rect 3724 15604 3764 15644
rect 3820 15352 3860 15392
rect 4396 16360 4436 16400
rect 4012 15268 4052 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3820 14764 3860 14804
rect 3532 14008 3572 14048
rect 4204 14848 4244 14888
rect 4108 14176 4148 14216
rect 4012 13924 4052 13964
rect 3628 13840 3668 13880
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3436 13336 3476 13376
rect 3244 12832 3284 12872
rect 3340 12244 3380 12284
rect 3148 12076 3188 12116
rect 3052 11740 3092 11780
rect 2860 11488 2900 11528
rect 2956 10984 2996 11024
rect 2860 10312 2900 10352
rect 2764 9808 2804 9848
rect 2764 9640 2804 9680
rect 2764 9304 2804 9344
rect 2668 9052 2708 9092
rect 2380 8548 2420 8588
rect 2188 7708 2228 7748
rect 2188 6952 2228 6992
rect 1996 5524 2036 5564
rect 1900 4516 1940 4556
rect 1804 3928 1844 3968
rect 1420 1408 1460 1448
rect 1036 904 1076 944
rect 1900 3760 1940 3800
rect 1900 148 1940 188
rect 2092 5356 2132 5396
rect 2284 6616 2324 6656
rect 2476 8296 2516 8336
rect 2476 7960 2516 8000
rect 2476 7708 2516 7748
rect 2860 8632 2900 8672
rect 3244 11656 3284 11696
rect 3052 10564 3092 10604
rect 3052 10228 3092 10268
rect 3148 9556 3188 9596
rect 3052 9472 3092 9512
rect 3244 8800 3284 8840
rect 3052 8632 3092 8672
rect 2860 8380 2900 8420
rect 3148 8380 3188 8420
rect 2668 7960 2708 8000
rect 2572 7120 2612 7160
rect 2476 5272 2516 5312
rect 2764 7120 2804 7160
rect 2668 6280 2708 6320
rect 2668 5692 2708 5732
rect 2764 5272 2804 5312
rect 4012 12832 4052 12872
rect 3820 12244 3860 12284
rect 4012 12244 4052 12284
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 4204 12916 4244 12956
rect 4684 17032 4724 17072
rect 4492 15940 4532 15980
rect 4396 15100 4436 15140
rect 5356 19888 5396 19928
rect 5164 19804 5204 19844
rect 5452 19720 5492 19760
rect 5356 19552 5396 19592
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 5356 18880 5396 18920
rect 5452 18796 5492 18836
rect 5452 17704 5492 17744
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 6220 21316 6260 21356
rect 6124 21148 6164 21188
rect 6316 20896 6356 20936
rect 6124 19720 6164 19760
rect 6028 18796 6068 18836
rect 6316 20644 6356 20684
rect 6316 19048 6356 19088
rect 6124 18376 6164 18416
rect 6028 18208 6068 18248
rect 5644 17704 5684 17744
rect 5356 17032 5396 17072
rect 5548 17032 5588 17072
rect 5836 16948 5876 16988
rect 6028 17704 6068 17744
rect 5932 16696 5972 16736
rect 5740 16528 5780 16568
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4972 15520 5012 15560
rect 5260 15436 5300 15476
rect 4780 15268 4820 15308
rect 4684 15016 4724 15056
rect 4684 14512 4724 14552
rect 4396 13672 4436 13712
rect 4684 12748 4724 12788
rect 4492 12244 4532 12284
rect 3628 11488 3668 11528
rect 4204 11824 4244 11864
rect 4108 11656 4148 11696
rect 4012 11152 4052 11192
rect 3820 10984 3860 11024
rect 4311 10984 4351 11024
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3532 10396 3572 10436
rect 3820 10396 3860 10436
rect 3436 10312 3476 10352
rect 3724 10144 3764 10184
rect 3532 10060 3572 10100
rect 3436 9976 3476 10016
rect 3724 9640 3764 9680
rect 3724 9472 3764 9512
rect 3532 9052 3572 9092
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3628 8884 3668 8924
rect 4204 10900 4244 10940
rect 4492 10900 4532 10940
rect 4492 10732 4532 10772
rect 4396 10564 4436 10604
rect 4300 9976 4340 10016
rect 4204 9507 4244 9512
rect 4204 9472 4244 9507
rect 4684 12076 4724 12116
rect 4684 10732 4724 10772
rect 4588 10480 4628 10520
rect 5356 15100 5396 15140
rect 5548 15100 5588 15140
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 5260 12580 5300 12620
rect 5452 14680 5492 14720
rect 5740 15940 5780 15980
rect 5740 12832 5780 12872
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 5260 10984 5300 11024
rect 4876 10900 4916 10940
rect 4972 10480 5012 10520
rect 4396 9472 4436 9512
rect 4108 8800 4148 8840
rect 3820 8716 3860 8756
rect 3628 8464 3668 8504
rect 3532 8128 3572 8168
rect 3436 8044 3476 8084
rect 3436 7876 3476 7916
rect 4108 8548 4148 8588
rect 4300 8800 4340 8840
rect 4204 8296 4244 8336
rect 4204 7960 4244 8000
rect 4012 7792 4052 7832
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3340 7456 3380 7496
rect 2956 7372 2996 7412
rect 3820 7372 3860 7412
rect 3724 7288 3764 7328
rect 3148 6784 3188 6824
rect 3052 6448 3092 6488
rect 3052 5692 3092 5732
rect 2188 4516 2228 4556
rect 2092 3592 2132 3632
rect 2284 3424 2324 3464
rect 2956 4852 2996 4892
rect 2860 4600 2900 4640
rect 2860 4264 2900 4304
rect 2572 3844 2612 3884
rect 2476 3592 2516 3632
rect 2764 3508 2804 3548
rect 2764 3004 2804 3044
rect 2668 2500 2708 2540
rect 2668 2080 2708 2120
rect 2860 2752 2900 2792
rect 2860 2164 2900 2204
rect 2572 1072 2612 1112
rect 3340 7120 3380 7160
rect 3628 7120 3668 7160
rect 3628 6784 3668 6824
rect 3436 6700 3476 6740
rect 3244 4852 3284 4892
rect 4012 7120 4052 7160
rect 4684 10060 4724 10100
rect 4588 8884 4628 8924
rect 4588 8716 4628 8756
rect 5164 10648 5204 10688
rect 5644 11152 5684 11192
rect 4780 9976 4820 10016
rect 5068 9976 5108 10016
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4588 8548 4628 8588
rect 4972 9220 5012 9260
rect 5164 8884 5204 8924
rect 4876 8716 4916 8756
rect 4876 8464 4916 8504
rect 5548 10984 5588 11024
rect 5452 8800 5492 8840
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4588 7708 4628 7748
rect 4300 7120 4340 7160
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3820 5860 3860 5900
rect 3628 5272 3668 5312
rect 4204 5608 4244 5648
rect 4204 5104 4244 5144
rect 4012 4684 4052 4724
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 3148 4180 3188 4220
rect 3148 3676 3188 3716
rect 3532 3592 3572 3632
rect 5260 8128 5300 8168
rect 5164 7456 5204 7496
rect 5260 7204 5300 7244
rect 4780 6784 4820 6824
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 5260 6616 5300 6656
rect 4396 5944 4436 5984
rect 4396 5104 4436 5144
rect 4204 4684 4244 4724
rect 4204 3928 4244 3968
rect 5164 6532 5204 6572
rect 5452 8128 5492 8168
rect 5452 7708 5492 7748
rect 5644 10480 5684 10520
rect 5644 9472 5684 9512
rect 5644 8716 5684 8756
rect 6220 18292 6260 18332
rect 6124 16948 6164 16988
rect 6028 16276 6068 16316
rect 6508 23836 6548 23876
rect 7084 24760 7124 24800
rect 6796 24172 6836 24212
rect 6796 23080 6836 23120
rect 6700 22240 6740 22280
rect 6508 22072 6548 22112
rect 7084 21316 7124 21356
rect 6796 20728 6836 20768
rect 7372 26188 7412 26228
rect 7276 26104 7316 26144
rect 7564 26608 7604 26648
rect 7852 29632 7892 29672
rect 7852 29464 7892 29504
rect 7852 29128 7892 29168
rect 7756 29044 7796 29084
rect 8140 32740 8180 32780
rect 8044 31648 8084 31688
rect 8044 29800 8084 29840
rect 8236 30640 8276 30680
rect 7756 28372 7796 28412
rect 7852 28288 7892 28328
rect 7756 27868 7796 27908
rect 8044 27616 8084 27656
rect 7660 26524 7700 26564
rect 7660 26104 7700 26144
rect 7468 26020 7508 26060
rect 7564 25684 7604 25724
rect 7372 24928 7412 24968
rect 8044 26524 8084 26564
rect 7852 26356 7892 26396
rect 7948 26188 7988 26228
rect 7852 26020 7892 26060
rect 7756 24760 7796 24800
rect 7372 23752 7412 23792
rect 7852 23836 7892 23876
rect 8044 23836 8084 23876
rect 7756 23752 7796 23792
rect 7564 23500 7604 23540
rect 7372 22492 7412 22532
rect 7948 23668 7988 23708
rect 8044 23332 8084 23372
rect 8044 23080 8084 23120
rect 7852 22660 7892 22700
rect 7660 21904 7700 21944
rect 7852 21904 7892 21944
rect 7276 20896 7316 20936
rect 7180 20644 7220 20684
rect 6988 20056 7028 20096
rect 6604 19720 6644 19760
rect 6988 19300 7028 19340
rect 6700 19132 6740 19172
rect 6604 18796 6644 18836
rect 7084 18880 7124 18920
rect 6700 18460 6740 18500
rect 6700 17368 6740 17408
rect 6316 17032 6356 17072
rect 6508 16780 6548 16820
rect 6412 16360 6452 16400
rect 6220 15856 6260 15896
rect 6412 15268 6452 15308
rect 6028 14932 6068 14972
rect 6316 14260 6356 14300
rect 5932 13336 5972 13376
rect 5932 12580 5972 12620
rect 5932 11656 5972 11696
rect 5932 11236 5972 11276
rect 6124 12832 6164 12872
rect 6412 14008 6452 14048
rect 6700 16612 6740 16652
rect 6700 16360 6740 16400
rect 7180 16780 7220 16820
rect 7372 17200 7412 17240
rect 6604 15520 6644 15560
rect 6988 14848 7028 14888
rect 7180 15268 7220 15308
rect 7372 16024 7412 16064
rect 7564 20308 7604 20348
rect 7564 20140 7604 20180
rect 7564 18208 7604 18248
rect 7468 15436 7508 15476
rect 7084 14764 7124 14804
rect 6988 14344 7028 14384
rect 6508 13840 6548 13880
rect 6508 13672 6548 13712
rect 6124 11656 6164 11696
rect 6316 11656 6356 11696
rect 6508 10648 6548 10688
rect 6220 10480 6260 10520
rect 6508 10396 6548 10436
rect 6316 10312 6356 10352
rect 6220 10144 6260 10184
rect 6124 10060 6164 10100
rect 6220 9976 6260 10016
rect 5932 9556 5972 9596
rect 6124 9472 6164 9512
rect 5932 8716 5972 8756
rect 5932 8548 5972 8588
rect 5740 7960 5780 8000
rect 5836 7372 5876 7412
rect 5740 6700 5780 6740
rect 4972 6280 5012 6320
rect 4876 5692 4916 5732
rect 5068 5608 5108 5648
rect 4780 5272 4820 5312
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5548 6532 5588 6572
rect 5740 6532 5780 6572
rect 5548 6112 5588 6152
rect 4588 4768 4628 4808
rect 4588 4348 4628 4388
rect 4108 3844 4148 3884
rect 4204 3508 4244 3548
rect 3052 3088 3092 3128
rect 3532 3004 3572 3044
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 3436 2836 3476 2876
rect 3244 2500 3284 2540
rect 3244 2248 3284 2288
rect 3148 1828 3188 1868
rect 2764 1072 2804 1112
rect 3148 988 3188 1028
rect 2956 904 2996 944
rect 2956 568 2996 608
rect 4492 3928 4532 3968
rect 4396 3172 4436 3212
rect 4204 2920 4244 2960
rect 3628 2752 3668 2792
rect 4012 2752 4052 2792
rect 3340 2080 3380 2120
rect 3340 1912 3380 1952
rect 3532 2164 3572 2204
rect 4396 2332 4436 2372
rect 4300 1744 4340 1784
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 3724 1240 3764 1280
rect 3340 484 3380 524
rect 3916 652 3956 692
rect 4972 4516 5012 4556
rect 5452 4936 5492 4976
rect 5356 4348 5396 4388
rect 5644 5608 5684 5648
rect 5164 3928 5204 3968
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4684 3172 4724 3212
rect 5452 3592 5492 3632
rect 5260 3424 5300 3464
rect 5164 3256 5204 3296
rect 4876 2584 4916 2624
rect 5356 3256 5396 3296
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 4684 1744 4724 1784
rect 4876 1576 4916 1616
rect 4684 1492 4724 1532
rect 4684 1324 4724 1364
rect 4876 1324 4916 1364
rect 4492 988 4532 1028
rect 5260 1912 5300 1952
rect 5260 1240 5300 1280
rect 4684 904 4724 944
rect 4492 820 4532 860
rect 5356 820 5396 860
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 5068 568 5108 608
rect 5740 5524 5780 5564
rect 5548 3340 5588 3380
rect 6220 9052 6260 9092
rect 6220 8800 6260 8840
rect 6124 8044 6164 8084
rect 6028 7540 6068 7580
rect 6220 7372 6260 7412
rect 6412 9976 6452 10016
rect 6412 8128 6452 8168
rect 6700 14176 6740 14216
rect 6796 14008 6836 14048
rect 7372 14764 7412 14804
rect 7276 14680 7316 14720
rect 7372 13840 7412 13880
rect 6796 13756 6836 13796
rect 6700 13336 6740 13376
rect 6892 11824 6932 11864
rect 6892 11404 6932 11444
rect 6892 9472 6932 9512
rect 6892 9304 6932 9344
rect 6796 9136 6836 9176
rect 6604 7708 6644 7748
rect 7468 13168 7508 13208
rect 7180 13084 7220 13124
rect 7276 12916 7316 12956
rect 7852 21568 7892 21608
rect 7852 20056 7892 20096
rect 7756 18208 7796 18248
rect 7756 18040 7796 18080
rect 7660 16192 7700 16232
rect 7852 16864 7892 16904
rect 7948 15184 7988 15224
rect 8428 33160 8468 33200
rect 8428 32320 8468 32360
rect 8620 33160 8660 33200
rect 8620 32992 8660 33032
rect 8524 32152 8564 32192
rect 8812 33496 8852 33536
rect 8812 33328 8852 33368
rect 8716 32740 8756 32780
rect 8332 26188 8372 26228
rect 8236 25684 8276 25724
rect 8620 31312 8660 31352
rect 8524 30640 8564 30680
rect 9004 32572 9044 32612
rect 9676 36520 9716 36560
rect 9484 36268 9524 36308
rect 9580 35932 9620 35972
rect 9292 34000 9332 34040
rect 9388 33328 9428 33368
rect 9388 33160 9428 33200
rect 9196 32992 9236 33032
rect 9100 32488 9140 32528
rect 9100 32320 9140 32360
rect 8908 31900 8948 31940
rect 8908 30640 8948 30680
rect 8812 30388 8852 30428
rect 8812 30220 8852 30260
rect 9388 32824 9428 32864
rect 9292 32656 9332 32696
rect 9388 32488 9428 32528
rect 9292 32152 9332 32192
rect 9676 35260 9716 35300
rect 10252 39208 10292 39248
rect 9868 36100 9908 36140
rect 9868 35932 9908 35972
rect 9580 32992 9620 33032
rect 9772 34336 9812 34376
rect 9772 33328 9812 33368
rect 9964 34336 10004 34376
rect 9868 33076 9908 33116
rect 9772 32740 9812 32780
rect 9676 32572 9716 32612
rect 9580 32320 9620 32360
rect 9676 32152 9716 32192
rect 9292 31312 9332 31352
rect 9292 31144 9332 31184
rect 9196 30220 9236 30260
rect 9004 29296 9044 29336
rect 9292 29296 9332 29336
rect 10156 33076 10196 33116
rect 10060 32740 10100 32780
rect 10156 32152 10196 32192
rect 10060 31732 10100 31772
rect 10156 31648 10196 31688
rect 9868 30724 9908 30764
rect 9484 30640 9524 30680
rect 9484 30388 9524 30428
rect 9484 30220 9524 30260
rect 9388 29128 9428 29168
rect 9292 28960 9332 29000
rect 8812 28204 8852 28244
rect 8716 27616 8756 27656
rect 8524 27532 8564 27572
rect 8524 26944 8564 26984
rect 8620 26608 8660 26648
rect 8524 26524 8564 26564
rect 8620 26188 8660 26228
rect 8524 26104 8564 26144
rect 8332 25264 8372 25304
rect 8428 25180 8468 25220
rect 8524 25012 8564 25052
rect 8428 24592 8468 24632
rect 8428 23920 8468 23960
rect 8332 23668 8372 23708
rect 8236 23500 8276 23540
rect 8332 22408 8372 22448
rect 8236 21232 8276 21272
rect 8812 26104 8852 26144
rect 8716 25768 8756 25808
rect 9004 26860 9044 26900
rect 9292 26440 9332 26480
rect 9292 26188 9332 26228
rect 9196 26020 9236 26060
rect 9004 25768 9044 25808
rect 8716 25180 8756 25220
rect 8908 24928 8948 24968
rect 9484 27616 9524 27656
rect 9484 26776 9524 26816
rect 9196 25264 9236 25304
rect 9388 25180 9428 25220
rect 9292 25012 9332 25052
rect 8812 23752 8852 23792
rect 8908 23668 8948 23708
rect 8812 23416 8852 23456
rect 8332 19888 8372 19928
rect 8332 19468 8372 19508
rect 9100 22492 9140 22532
rect 9100 21568 9140 21608
rect 9100 20812 9140 20852
rect 8716 20056 8756 20096
rect 8236 18964 8276 19004
rect 9868 29128 9908 29168
rect 10060 29464 10100 29504
rect 9772 27616 9812 27656
rect 9676 27532 9716 27572
rect 9868 27448 9908 27488
rect 10732 38872 10772 38912
rect 10540 38536 10580 38576
rect 10348 38200 10388 38240
rect 10828 38452 10868 38492
rect 10636 38032 10676 38072
rect 10540 37948 10580 37988
rect 10348 36268 10388 36308
rect 10348 35764 10388 35804
rect 10444 35176 10484 35216
rect 10348 35008 10388 35048
rect 10348 32740 10388 32780
rect 10348 31648 10388 31688
rect 10828 36100 10868 36140
rect 11884 48112 11924 48152
rect 12172 48196 12212 48236
rect 12076 47440 12116 47480
rect 13132 48784 13172 48824
rect 13612 49456 13652 49496
rect 13612 49204 13652 49244
rect 12268 47272 12308 47312
rect 11788 46012 11828 46052
rect 11596 45340 11636 45380
rect 11500 45256 11540 45296
rect 11692 45256 11732 45296
rect 11884 44500 11924 44540
rect 12940 47020 12980 47060
rect 12940 46852 12980 46892
rect 12172 46012 12212 46052
rect 12076 44248 12116 44288
rect 11692 42820 11732 42860
rect 12076 42736 12116 42776
rect 11500 42568 11540 42608
rect 11692 42316 11732 42356
rect 11500 41980 11540 42020
rect 11500 40468 11540 40508
rect 11308 39292 11348 39332
rect 11212 38620 11252 38660
rect 11404 38620 11444 38660
rect 11116 38536 11156 38576
rect 11212 38200 11252 38240
rect 11884 38956 11924 38996
rect 11788 38620 11828 38660
rect 11308 38032 11348 38072
rect 11212 35596 11252 35636
rect 10924 35176 10964 35216
rect 11020 34840 11060 34880
rect 11020 34588 11060 34628
rect 10636 34168 10676 34208
rect 11020 33748 11060 33788
rect 11020 33244 11060 33284
rect 10636 32908 10676 32948
rect 10732 32656 10772 32696
rect 10636 31564 10676 31604
rect 10540 30640 10580 30680
rect 10348 28288 10388 28328
rect 10732 30472 10772 30512
rect 10636 29884 10676 29924
rect 11020 32656 11060 32696
rect 11692 38200 11732 38240
rect 11596 37528 11636 37568
rect 11404 36268 11444 36308
rect 11404 36100 11444 36140
rect 11404 34756 11444 34796
rect 11500 33916 11540 33956
rect 11404 33832 11444 33872
rect 11500 33580 11540 33620
rect 11980 38872 12020 38912
rect 11884 38116 11924 38156
rect 12076 37528 12116 37568
rect 11788 36772 11828 36812
rect 11692 36436 11732 36476
rect 11596 32908 11636 32948
rect 11308 31312 11348 31352
rect 11500 30892 11540 30932
rect 11116 30640 11156 30680
rect 11404 30640 11444 30680
rect 11212 30472 11252 30512
rect 11116 30220 11156 30260
rect 11020 29884 11060 29924
rect 10924 29464 10964 29504
rect 10924 29044 10964 29084
rect 11116 28708 11156 28748
rect 11020 28456 11060 28496
rect 9676 27196 9716 27236
rect 9580 26104 9620 26144
rect 9772 26188 9812 26228
rect 9484 24928 9524 24968
rect 9580 24676 9620 24716
rect 9484 24424 9524 24464
rect 9292 23164 9332 23204
rect 9292 20812 9332 20852
rect 9196 19384 9236 19424
rect 9100 18460 9140 18500
rect 9004 18208 9044 18248
rect 9100 17788 9140 17828
rect 9964 26104 10004 26144
rect 9868 25684 9908 25724
rect 9772 25264 9812 25304
rect 9676 23416 9716 23456
rect 9484 23080 9524 23120
rect 10252 27364 10292 27404
rect 10252 26776 10292 26816
rect 10252 26608 10292 26648
rect 10156 26188 10196 26228
rect 10924 27700 10964 27740
rect 10348 26440 10388 26480
rect 10636 26440 10676 26480
rect 10444 26188 10484 26228
rect 10348 26104 10388 26144
rect 10636 26104 10676 26144
rect 10156 25684 10196 25724
rect 10156 25264 10196 25304
rect 10252 24592 10292 24632
rect 10732 24592 10772 24632
rect 9964 23920 10004 23960
rect 9868 23080 9908 23120
rect 9580 22492 9620 22532
rect 9484 22072 9524 22112
rect 9484 20980 9524 21020
rect 9388 20056 9428 20096
rect 8332 17200 8372 17240
rect 8140 16864 8180 16904
rect 8044 14176 8084 14216
rect 7756 13168 7796 13208
rect 7180 11068 7220 11108
rect 7564 11740 7604 11780
rect 7084 9640 7124 9680
rect 7084 9472 7124 9512
rect 7084 8800 7124 8840
rect 6988 8128 7028 8168
rect 6892 7876 6932 7916
rect 7084 7876 7124 7916
rect 7084 7708 7124 7748
rect 6796 7540 6836 7580
rect 6412 7120 6452 7160
rect 6316 6952 6356 6992
rect 6124 6784 6164 6824
rect 5932 5524 5972 5564
rect 6028 5188 6068 5228
rect 5932 4852 5972 4892
rect 5932 4600 5972 4640
rect 5548 904 5588 944
rect 6028 3172 6068 3212
rect 6412 6196 6452 6236
rect 6220 5944 6260 5984
rect 6796 6952 6836 6992
rect 6604 6700 6644 6740
rect 6988 6700 7028 6740
rect 6316 5272 6356 5312
rect 6412 4768 6452 4808
rect 6220 4600 6260 4640
rect 6316 4180 6356 4220
rect 6220 2584 6260 2624
rect 5932 568 5972 608
rect 6124 2080 6164 2120
rect 6412 3172 6452 3212
rect 6892 5608 6932 5648
rect 7276 9976 7316 10016
rect 7948 12748 7988 12788
rect 7852 11656 7892 11696
rect 7756 11572 7796 11612
rect 7468 10900 7508 10940
rect 7468 10060 7508 10100
rect 7372 9640 7412 9680
rect 7276 9304 7316 9344
rect 7276 8128 7316 8168
rect 7276 7120 7316 7160
rect 7276 6616 7316 6656
rect 7756 9304 7796 9344
rect 7564 8632 7604 8672
rect 7468 7708 7508 7748
rect 7468 7120 7508 7160
rect 7372 5860 7412 5900
rect 7276 5692 7316 5732
rect 7180 5104 7220 5144
rect 6796 4768 6836 4808
rect 6796 4348 6836 4388
rect 6796 2752 6836 2792
rect 6412 2500 6452 2540
rect 6316 2164 6356 2204
rect 6700 2080 6740 2120
rect 6412 1660 6452 1700
rect 6508 1492 6548 1532
rect 6412 1156 6452 1196
rect 6124 232 6164 272
rect 6220 148 6260 188
rect 7180 4936 7220 4976
rect 6988 4684 7028 4724
rect 7084 3088 7124 3128
rect 6988 2668 7028 2708
rect 7084 2584 7124 2624
rect 6892 2500 6932 2540
rect 7468 5272 7508 5312
rect 7468 5020 7508 5060
rect 8044 12580 8084 12620
rect 8620 17032 8660 17072
rect 9196 17116 9236 17156
rect 9580 20728 9620 20768
rect 9580 18628 9620 18668
rect 9484 17116 9524 17156
rect 8236 15436 8276 15476
rect 8428 14932 8468 14972
rect 8428 14680 8468 14720
rect 8428 14176 8468 14216
rect 8332 14008 8372 14048
rect 8236 13168 8276 13208
rect 8140 11824 8180 11864
rect 8140 11656 8180 11696
rect 8044 11404 8084 11444
rect 8044 10984 8084 11024
rect 8044 8128 8084 8168
rect 7660 7120 7700 7160
rect 7660 6700 7700 6740
rect 7660 6280 7700 6320
rect 7660 6028 7700 6068
rect 7372 4852 7412 4892
rect 7564 4768 7604 4808
rect 7276 4516 7316 4556
rect 6796 1072 6836 1112
rect 6508 736 6548 776
rect 6604 652 6644 692
rect 7084 2248 7124 2288
rect 6988 2164 7028 2204
rect 7180 1744 7220 1784
rect 6892 568 6932 608
rect 6988 316 7028 356
rect 7564 4096 7604 4136
rect 7468 3676 7508 3716
rect 7468 3424 7508 3464
rect 8044 7708 8084 7748
rect 7948 7288 7988 7328
rect 7948 7120 7988 7160
rect 7852 7036 7892 7076
rect 8044 7036 8084 7076
rect 7852 6700 7892 6740
rect 7948 6280 7988 6320
rect 7756 3928 7796 3968
rect 7660 3424 7700 3464
rect 7756 3340 7796 3380
rect 7564 2668 7604 2708
rect 7468 1324 7508 1364
rect 8716 16192 8756 16232
rect 8620 15352 8660 15392
rect 8620 14848 8660 14888
rect 9100 16192 9140 16232
rect 9388 16696 9428 16736
rect 9292 16612 9332 16652
rect 8908 15940 8948 15980
rect 8812 15352 8852 15392
rect 8524 14008 8564 14048
rect 8716 14008 8756 14048
rect 8620 13588 8660 13628
rect 9100 14092 9140 14132
rect 8908 13672 8948 13712
rect 8812 13588 8852 13628
rect 8716 12580 8756 12620
rect 8716 12244 8756 12284
rect 8716 11824 8756 11864
rect 8620 11656 8660 11696
rect 8524 10984 8564 11024
rect 8428 10648 8468 10688
rect 8524 10564 8564 10604
rect 8908 12328 8948 12368
rect 8812 9976 8852 10016
rect 9100 13336 9140 13376
rect 9484 16276 9524 16316
rect 9772 20728 9812 20768
rect 10060 23668 10100 23708
rect 10156 23584 10196 23624
rect 10060 23080 10100 23120
rect 10540 24172 10580 24212
rect 10828 24340 10868 24380
rect 11020 26440 11060 26480
rect 11020 25432 11060 25472
rect 10732 23920 10772 23960
rect 10636 23752 10676 23792
rect 10540 23080 10580 23120
rect 10636 22744 10676 22784
rect 10252 22492 10292 22532
rect 10924 23752 10964 23792
rect 10156 22240 10196 22280
rect 9964 20812 10004 20852
rect 10252 20644 10292 20684
rect 10252 20476 10292 20516
rect 10060 19384 10100 19424
rect 9964 18964 10004 19004
rect 9868 18460 9908 18500
rect 9964 16948 10004 16988
rect 9868 16612 9908 16652
rect 9964 16276 10004 16316
rect 9676 15940 9716 15980
rect 9676 15436 9716 15476
rect 9772 15352 9812 15392
rect 9772 15016 9812 15056
rect 10252 19221 10292 19256
rect 10252 19216 10292 19221
rect 10252 18964 10292 19004
rect 10252 18796 10292 18836
rect 10732 21568 10772 21608
rect 11116 24172 11156 24212
rect 11116 24004 11156 24044
rect 10732 21148 10772 21188
rect 10636 20476 10676 20516
rect 10828 19972 10868 20012
rect 10540 19216 10580 19256
rect 10444 18964 10484 19004
rect 10348 18712 10388 18752
rect 10828 19552 10868 19592
rect 10732 18880 10772 18920
rect 11500 30556 11540 30596
rect 11596 30388 11636 30428
rect 11308 29296 11348 29336
rect 11404 29128 11444 29168
rect 11500 28036 11540 28076
rect 11404 27868 11444 27908
rect 11308 23500 11348 23540
rect 11308 22744 11348 22784
rect 11212 21232 11252 21272
rect 11116 20812 11156 20852
rect 11020 20728 11060 20768
rect 11020 20224 11060 20264
rect 10156 17284 10196 17324
rect 10156 17032 10196 17072
rect 10444 17200 10484 17240
rect 10252 16360 10292 16400
rect 10156 15940 10196 15980
rect 10828 18712 10868 18752
rect 10732 17032 10772 17072
rect 10540 16108 10580 16148
rect 10540 15856 10580 15896
rect 10060 15520 10100 15560
rect 10348 15520 10388 15560
rect 10060 15352 10100 15392
rect 9964 14932 10004 14972
rect 10828 16276 10868 16316
rect 10732 16192 10772 16232
rect 11116 17536 11156 17576
rect 11116 17368 11156 17408
rect 10732 15856 10772 15896
rect 10636 14764 10676 14804
rect 10540 14680 10580 14720
rect 9484 13336 9524 13376
rect 9100 12832 9140 12872
rect 9580 12748 9620 12788
rect 9484 11908 9524 11948
rect 9196 11656 9236 11696
rect 10348 13252 10388 13292
rect 10732 13168 10772 13208
rect 10636 12916 10676 12956
rect 10444 12664 10484 12704
rect 10060 12580 10100 12620
rect 10732 12580 10772 12620
rect 9868 11404 9908 11444
rect 9100 9976 9140 10016
rect 8908 9892 8948 9932
rect 8524 9220 8564 9260
rect 8620 8800 8660 8840
rect 8332 8296 8372 8336
rect 8236 8212 8276 8252
rect 8332 7120 8372 7160
rect 9100 9136 9140 9176
rect 8812 9052 8852 9092
rect 8716 7456 8756 7496
rect 9100 8632 9140 8672
rect 8812 7204 8852 7244
rect 8140 6784 8180 6824
rect 8236 6280 8276 6320
rect 8044 5692 8084 5732
rect 8044 4852 8084 4892
rect 7948 4600 7988 4640
rect 7852 3172 7892 3212
rect 8332 5860 8372 5900
rect 8524 6952 8564 6992
rect 8140 4096 8180 4136
rect 8236 3844 8276 3884
rect 8140 3760 8180 3800
rect 8428 5608 8468 5648
rect 8908 6616 8948 6656
rect 8812 6532 8852 6572
rect 8716 6196 8756 6236
rect 9100 6196 9140 6236
rect 9004 6028 9044 6068
rect 8908 5692 8948 5732
rect 10540 12244 10580 12284
rect 10444 11908 10484 11948
rect 10156 9640 10196 9680
rect 9580 8632 9620 8672
rect 9580 8464 9620 8504
rect 9388 6952 9428 6992
rect 9292 6112 9332 6152
rect 9292 5860 9332 5900
rect 9196 5776 9236 5816
rect 8812 4936 8852 4976
rect 8620 4348 8660 4388
rect 9004 5104 9044 5144
rect 8620 3928 8660 3968
rect 8716 3508 8756 3548
rect 7756 3088 7796 3128
rect 7660 1156 7700 1196
rect 7564 988 7604 1028
rect 8044 2500 8084 2540
rect 8044 2164 8084 2204
rect 7948 1240 7988 1280
rect 7948 64 7988 104
rect 8332 3172 8372 3212
rect 8236 2500 8276 2540
rect 8236 2332 8276 2372
rect 8716 3088 8756 3128
rect 8524 2752 8564 2792
rect 8620 2500 8660 2540
rect 8524 2164 8564 2204
rect 8428 2080 8468 2120
rect 9868 9304 9908 9344
rect 10060 9220 10100 9260
rect 10060 7995 10100 8000
rect 10060 7960 10100 7995
rect 10060 7624 10100 7664
rect 9580 7372 9620 7412
rect 9484 6112 9524 6152
rect 9772 5860 9812 5900
rect 9388 5440 9428 5480
rect 9292 5020 9332 5060
rect 9196 4348 9236 4388
rect 9196 4180 9236 4220
rect 8908 2668 8948 2708
rect 8812 1996 8852 2036
rect 9292 3760 9332 3800
rect 9292 3424 9332 3464
rect 9196 3340 9236 3380
rect 9100 2584 9140 2624
rect 9100 1828 9140 1868
rect 8428 1492 8468 1532
rect 8908 1492 8948 1532
rect 8908 1240 8948 1280
rect 8620 1156 8660 1196
rect 8428 1072 8468 1112
rect 8716 1072 8756 1112
rect 8428 484 8468 524
rect 8524 232 8564 272
rect 8812 820 8852 860
rect 9292 1660 9332 1700
rect 9772 5272 9812 5312
rect 9676 5104 9716 5144
rect 9868 4180 9908 4220
rect 9676 3760 9716 3800
rect 9580 3340 9620 3380
rect 9484 2836 9524 2876
rect 9484 1828 9524 1868
rect 9676 2668 9716 2708
rect 10540 11656 10580 11696
rect 11116 15856 11156 15896
rect 11116 15520 11156 15560
rect 11020 15268 11060 15308
rect 10924 14008 10964 14048
rect 11308 20728 11348 20768
rect 11596 27616 11636 27656
rect 11980 36688 12020 36728
rect 12076 35092 12116 35132
rect 11788 29044 11828 29084
rect 12556 46180 12596 46220
rect 12652 44752 12692 44792
rect 12748 44248 12788 44288
rect 12460 44164 12500 44204
rect 12652 44164 12692 44204
rect 12460 42400 12500 42440
rect 12268 39376 12308 39416
rect 12268 39040 12308 39080
rect 12556 40804 12596 40844
rect 12748 42736 12788 42776
rect 13132 46432 13172 46472
rect 13612 47944 13652 47984
rect 13516 47356 13556 47396
rect 14092 56512 14132 56552
rect 14092 56176 14132 56216
rect 14092 54748 14132 54788
rect 14380 65248 14420 65288
rect 14476 64492 14516 64532
rect 14956 68356 14996 68396
rect 14764 67852 14804 67892
rect 14860 67684 14900 67724
rect 14860 66760 14900 66800
rect 14860 65836 14900 65876
rect 14764 65332 14804 65372
rect 14764 65164 14804 65204
rect 14668 63904 14708 63944
rect 14476 63736 14516 63776
rect 14476 61804 14516 61844
rect 14956 65080 14996 65120
rect 14860 63316 14900 63356
rect 14476 61468 14516 61508
rect 14860 61636 14900 61676
rect 15340 69952 15380 69992
rect 15532 69868 15572 69908
rect 15436 69784 15476 69824
rect 15436 68608 15476 68648
rect 15244 65500 15284 65540
rect 15148 61468 15188 61508
rect 14860 61132 14900 61172
rect 15052 61132 15092 61172
rect 15436 66760 15476 66800
rect 15340 65416 15380 65456
rect 15532 65668 15572 65708
rect 15532 64408 15572 64448
rect 15532 63232 15572 63272
rect 15532 62476 15572 62516
rect 15340 62224 15380 62264
rect 15340 61216 15380 61256
rect 14956 61048 14996 61088
rect 14572 60880 14612 60920
rect 14476 60796 14516 60836
rect 14476 60376 14516 60416
rect 14380 59872 14420 59912
rect 14284 59704 14324 59744
rect 14284 56344 14324 56384
rect 14284 56092 14324 56132
rect 14188 54160 14228 54200
rect 14476 59704 14516 59744
rect 14476 59452 14516 59492
rect 14476 59284 14516 59324
rect 14764 60460 14804 60500
rect 15017 60544 15057 60584
rect 14956 60376 14996 60416
rect 14668 59536 14708 59576
rect 14860 60040 14900 60080
rect 14956 59788 14996 59828
rect 14668 59368 14708 59408
rect 14572 59200 14612 59240
rect 14572 57016 14612 57056
rect 14476 55504 14516 55544
rect 15436 61048 15476 61088
rect 15244 60544 15284 60584
rect 15532 60880 15572 60920
rect 15244 59536 15284 59576
rect 15148 57184 15188 57224
rect 15052 57025 15092 57056
rect 15052 57016 15092 57025
rect 15340 58948 15380 58988
rect 15340 58612 15380 58652
rect 15436 57688 15476 57728
rect 15148 56932 15188 56972
rect 14956 56680 14996 56720
rect 15052 56512 15092 56552
rect 14860 56428 14900 56468
rect 14764 55924 14804 55964
rect 14476 55336 14516 55376
rect 14380 55000 14420 55040
rect 14572 55084 14612 55124
rect 14476 54832 14516 54872
rect 14380 54244 14420 54284
rect 14476 53992 14516 54032
rect 14284 53236 14324 53276
rect 14188 53152 14228 53192
rect 14476 53404 14516 53444
rect 14188 52396 14228 52436
rect 14092 51808 14132 51848
rect 14092 51472 14132 51512
rect 13804 50128 13844 50168
rect 13804 49456 13844 49496
rect 13804 47944 13844 47984
rect 13228 46180 13268 46220
rect 13420 45256 13460 45296
rect 13708 45760 13748 45800
rect 13228 44248 13268 44288
rect 13036 44164 13076 44204
rect 13132 43576 13172 43616
rect 13132 42652 13172 42692
rect 12748 41560 12788 41600
rect 12652 40552 12692 40592
rect 12748 39712 12788 39752
rect 12556 39544 12596 39584
rect 12364 38872 12404 38912
rect 12460 38368 12500 38408
rect 12460 36436 12500 36476
rect 12364 35932 12404 35972
rect 12268 35680 12308 35720
rect 13132 42232 13172 42272
rect 13132 41896 13172 41936
rect 13420 43660 13460 43700
rect 13516 41812 13556 41852
rect 13612 41560 13652 41600
rect 13036 39964 13076 40004
rect 13996 50968 14036 51008
rect 13996 50548 14036 50588
rect 14188 50968 14228 51008
rect 14380 52648 14420 52688
rect 14668 54244 14708 54284
rect 14956 55000 14996 55040
rect 14860 54748 14900 54788
rect 14764 53824 14804 53864
rect 14668 53320 14708 53360
rect 14860 53740 14900 53780
rect 14572 51892 14612 51932
rect 14572 51640 14612 51680
rect 14476 51472 14516 51512
rect 14860 53152 14900 53192
rect 14860 52648 14900 52688
rect 14860 51808 14900 51848
rect 14860 51640 14900 51680
rect 15052 52816 15092 52856
rect 15244 56848 15284 56888
rect 15532 57604 15572 57644
rect 16012 71212 16052 71252
rect 16012 70960 16052 71000
rect 16396 77512 16436 77552
rect 16876 80452 16916 80492
rect 16684 79948 16724 79988
rect 16684 79612 16724 79652
rect 16684 79444 16724 79484
rect 16588 78436 16628 78476
rect 16876 79948 16916 79988
rect 16876 79444 16916 79484
rect 17068 79780 17108 79820
rect 17068 79612 17108 79652
rect 17260 83980 17300 84020
rect 17260 83224 17300 83264
rect 17356 83140 17396 83180
rect 17452 82720 17492 82760
rect 17740 84484 17780 84524
rect 18220 84988 18260 85028
rect 18124 84736 18164 84776
rect 17932 84400 17972 84440
rect 18028 84232 18068 84272
rect 17740 83644 17780 83684
rect 17740 82720 17780 82760
rect 17260 80620 17300 80660
rect 17164 78772 17204 78812
rect 17068 78688 17108 78728
rect 17068 78520 17108 78560
rect 16972 78100 17012 78140
rect 16780 77512 16820 77552
rect 16684 75832 16724 75872
rect 16588 75160 16628 75200
rect 18124 83308 18164 83348
rect 18412 84652 18452 84692
rect 18316 84064 18356 84104
rect 18316 83896 18356 83936
rect 18220 83140 18260 83180
rect 18124 83056 18164 83096
rect 17740 80368 17780 80408
rect 17740 79948 17780 79988
rect 17644 79780 17684 79820
rect 17548 79528 17588 79568
rect 17441 79276 17481 79316
rect 17548 79276 17588 79316
rect 17740 79612 17780 79652
rect 17932 81880 17972 81920
rect 18220 81964 18260 82004
rect 19276 85072 19316 85112
rect 19084 84988 19124 85028
rect 19468 84904 19508 84944
rect 18700 84652 18740 84692
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 18892 84484 18932 84524
rect 19276 84400 19316 84440
rect 18508 84232 18548 84272
rect 18700 84232 18740 84272
rect 19084 84148 19124 84188
rect 19564 84820 19604 84860
rect 19468 84316 19508 84356
rect 18508 83728 18548 83768
rect 18412 83140 18452 83180
rect 18508 82972 18548 83012
rect 18700 83476 18740 83516
rect 19084 83392 19124 83432
rect 18700 83140 18740 83180
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 18700 82720 18740 82760
rect 18220 81040 18260 81080
rect 18028 80620 18068 80660
rect 18124 80536 18164 80576
rect 17932 80368 17972 80408
rect 18124 79948 18164 79988
rect 17932 79864 17972 79904
rect 18124 79612 18164 79652
rect 17356 78772 17396 78812
rect 17932 79192 17972 79232
rect 17836 79024 17876 79064
rect 18028 79024 18068 79064
rect 19084 82972 19124 83012
rect 18892 82636 18932 82676
rect 19756 84736 19796 84776
rect 19660 84064 19700 84104
rect 20044 84568 20084 84608
rect 19852 84316 19892 84356
rect 19948 84232 19988 84272
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 19756 83476 19796 83516
rect 20121 83224 20161 83264
rect 19372 82972 19412 83012
rect 19372 82552 19412 82592
rect 19468 82468 19508 82508
rect 19276 81880 19316 81920
rect 18796 81796 18836 81836
rect 19276 81712 19316 81752
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 18604 81376 18644 81416
rect 18796 81208 18836 81248
rect 18604 81040 18644 81080
rect 18508 80956 18548 80996
rect 18508 80368 18548 80408
rect 18412 79612 18452 79652
rect 18508 79108 18548 79148
rect 18220 78940 18260 78980
rect 18508 78940 18548 78980
rect 17644 78436 17684 78476
rect 18124 78604 18164 78644
rect 17260 78184 17300 78224
rect 17260 78016 17300 78056
rect 17356 77680 17396 77720
rect 17164 77428 17204 77468
rect 16972 75832 17012 75872
rect 16876 75412 16916 75452
rect 16492 74488 16532 74528
rect 16396 73564 16436 73604
rect 16396 72892 16436 72932
rect 16396 71968 16436 72008
rect 16204 71380 16244 71420
rect 15916 69112 15956 69152
rect 15916 67180 15956 67220
rect 16108 68944 16148 68984
rect 16108 67180 16148 67220
rect 16108 67012 16148 67052
rect 16012 66760 16052 66800
rect 15724 66088 15764 66128
rect 16012 65500 16052 65540
rect 15724 64576 15764 64616
rect 15916 64408 15956 64448
rect 16108 64324 16148 64364
rect 15820 64240 15860 64280
rect 15724 63232 15764 63272
rect 15724 63064 15764 63104
rect 16300 69868 16340 69908
rect 16492 71212 16532 71252
rect 18028 78268 18068 78308
rect 17548 78184 17588 78224
rect 17740 77512 17780 77552
rect 17452 76000 17492 76040
rect 17356 75580 17396 75620
rect 17260 75328 17300 75368
rect 17164 75244 17204 75284
rect 16972 74488 17012 74528
rect 16876 72892 16916 72932
rect 16780 71884 16820 71924
rect 16684 70288 16724 70328
rect 16396 69616 16436 69656
rect 16300 69112 16340 69152
rect 16300 64072 16340 64112
rect 16300 63820 16340 63860
rect 16204 63064 16244 63104
rect 15916 62980 15956 63020
rect 16108 62560 16148 62600
rect 16204 61804 16244 61844
rect 16108 61720 16148 61760
rect 15916 61384 15956 61424
rect 16300 61636 16340 61676
rect 16300 61300 16340 61340
rect 16204 60628 16244 60668
rect 16108 59872 16148 59912
rect 15916 59536 15956 59576
rect 15724 57856 15764 57896
rect 15724 57604 15764 57644
rect 15436 56932 15476 56972
rect 15340 56596 15380 56636
rect 15340 56344 15380 56384
rect 15244 56176 15284 56216
rect 15724 57016 15764 57056
rect 15916 57436 15956 57476
rect 16012 57100 16052 57140
rect 15724 56596 15764 56636
rect 15628 56176 15668 56216
rect 15532 55504 15572 55544
rect 15340 54916 15380 54956
rect 15244 52648 15284 52688
rect 15052 52396 15092 52436
rect 15244 52480 15284 52520
rect 15148 52312 15188 52352
rect 15052 51724 15092 51764
rect 15148 51640 15188 51680
rect 14764 51136 14804 51176
rect 13996 49456 14036 49496
rect 13996 49120 14036 49160
rect 13996 48028 14036 48068
rect 14188 50128 14228 50168
rect 14380 50296 14420 50336
rect 14284 50044 14324 50084
rect 14284 49456 14324 49496
rect 14572 50044 14612 50084
rect 14572 49792 14612 49832
rect 15052 51136 15092 51176
rect 14956 50968 14996 51008
rect 15436 54748 15476 54788
rect 15436 53404 15476 53444
rect 15628 53320 15668 53360
rect 15820 56260 15860 56300
rect 15820 55756 15860 55796
rect 15820 55336 15860 55376
rect 15724 53236 15764 53276
rect 15532 52816 15572 52856
rect 15340 51304 15380 51344
rect 15436 51220 15476 51260
rect 15532 50968 15572 51008
rect 15724 52480 15764 52520
rect 16012 56260 16052 56300
rect 16012 55420 16052 55460
rect 16204 57184 16244 57224
rect 16204 56680 16244 56720
rect 16492 64576 16532 64616
rect 16492 62980 16532 63020
rect 16396 59704 16436 59744
rect 16396 59536 16436 59576
rect 16876 69616 16916 69656
rect 16876 69448 16916 69488
rect 16684 66928 16724 66968
rect 16684 65920 16724 65960
rect 16684 65248 16724 65288
rect 17260 73011 17300 73016
rect 17260 72976 17300 73011
rect 17644 75580 17684 75620
rect 17932 78100 17972 78140
rect 18124 78100 18164 78140
rect 18892 80620 18932 80660
rect 18604 78520 18644 78560
rect 18508 78436 18548 78476
rect 18604 78352 18644 78392
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 19180 79948 19220 79988
rect 18988 79696 19028 79736
rect 18796 79360 18836 79400
rect 19756 82636 19796 82676
rect 19660 81796 19700 81836
rect 19564 81460 19604 81500
rect 19468 79780 19508 79820
rect 19180 79276 19220 79316
rect 19468 79444 19508 79484
rect 19564 79360 19604 79400
rect 19372 79024 19412 79064
rect 18892 78940 18932 78980
rect 18988 78856 19028 78896
rect 19276 78856 19316 78896
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 18220 77848 18260 77888
rect 18220 77680 18260 77720
rect 17932 76840 17972 76880
rect 18124 76756 18164 76796
rect 18028 76672 18068 76712
rect 17836 76000 17876 76040
rect 18028 76000 18068 76040
rect 17548 73144 17588 73184
rect 17740 75160 17780 75200
rect 17740 74992 17780 75032
rect 17644 73060 17684 73100
rect 17452 72892 17492 72932
rect 17548 72808 17588 72848
rect 17452 71968 17492 72008
rect 17164 71464 17204 71504
rect 17452 71464 17492 71504
rect 17260 70960 17300 71000
rect 17548 70960 17588 71000
rect 17164 68440 17204 68480
rect 17452 70288 17492 70328
rect 17644 70540 17684 70580
rect 18412 78268 18452 78308
rect 18316 77344 18356 77384
rect 18316 77092 18356 77132
rect 18220 75664 18260 75704
rect 18220 75328 18260 75368
rect 18028 74488 18068 74528
rect 17932 74404 17972 74444
rect 17836 73480 17876 73520
rect 17932 70624 17972 70664
rect 17068 66844 17108 66884
rect 17164 66088 17204 66128
rect 17836 70288 17876 70328
rect 18124 73648 18164 73688
rect 18508 78100 18548 78140
rect 18508 77848 18548 77888
rect 18604 77428 18644 77468
rect 18508 76840 18548 76880
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 18700 76840 18740 76880
rect 18892 76840 18932 76880
rect 18412 74992 18452 75032
rect 19372 76756 19412 76796
rect 19276 75748 19316 75788
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 20044 81796 20084 81836
rect 20524 81376 20564 81416
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 19948 80620 19988 80660
rect 20140 80368 20180 80408
rect 19852 80284 19892 80324
rect 19756 79864 19796 79904
rect 19948 79780 19988 79820
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 19948 79192 19988 79232
rect 20620 80452 20660 80492
rect 19948 79059 19988 79064
rect 19948 79024 19988 79059
rect 19756 77848 19796 77888
rect 19564 77260 19604 77300
rect 18124 73144 18164 73184
rect 18508 73480 18548 73520
rect 18412 73396 18452 73436
rect 18124 72808 18164 72848
rect 18124 70456 18164 70496
rect 18028 69616 18068 69656
rect 17932 69196 17972 69236
rect 17644 68440 17684 68480
rect 17452 67600 17492 67640
rect 19084 74236 19124 74276
rect 19276 74236 19316 74276
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 18700 73396 18740 73436
rect 18604 71296 18644 71336
rect 18316 71212 18356 71252
rect 18508 70456 18548 70496
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 19660 76252 19700 76292
rect 19660 75664 19700 75704
rect 18988 72052 19028 72092
rect 19372 72052 19412 72092
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 19372 70456 19412 70496
rect 18700 70288 18740 70328
rect 18316 69616 18356 69656
rect 18796 69952 18836 69992
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 19660 74320 19700 74360
rect 20140 78016 20180 78056
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 20044 77260 20084 77300
rect 20044 77092 20084 77132
rect 19852 76000 19892 76040
rect 20140 76504 20180 76544
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 20044 76168 20084 76208
rect 20044 74992 20084 75032
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 20236 74572 20276 74612
rect 19756 73648 19796 73688
rect 19852 73144 19892 73184
rect 19852 72724 19892 72764
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 20044 73144 20084 73184
rect 20716 77092 20756 77132
rect 21292 74572 21332 74612
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 19660 71464 19700 71504
rect 19564 70960 19604 71000
rect 19756 71044 19796 71084
rect 19660 70708 19700 70748
rect 19468 69784 19508 69824
rect 18028 67600 18068 67640
rect 18124 67096 18164 67136
rect 19180 69112 19220 69152
rect 18412 68188 18452 68228
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 18604 67264 18644 67304
rect 17644 66256 17684 66296
rect 17932 66256 17972 66296
rect 17548 65332 17588 65372
rect 18220 66172 18260 66212
rect 18124 65500 18164 65540
rect 17932 65080 17972 65120
rect 16876 63232 16916 63272
rect 16876 62560 16916 62600
rect 16780 61972 16820 62012
rect 16684 61552 16724 61592
rect 16972 60964 17012 61004
rect 16876 60460 16916 60500
rect 16588 59452 16628 59492
rect 16780 60040 16820 60080
rect 16780 59704 16820 59744
rect 16684 59200 16724 59240
rect 16492 57940 16532 57980
rect 16684 58108 16724 58148
rect 16588 57688 16628 57728
rect 17740 63400 17780 63440
rect 17932 63400 17972 63440
rect 18028 63148 18068 63188
rect 17548 61552 17588 61592
rect 17452 61384 17492 61424
rect 17356 60880 17396 60920
rect 17164 60712 17204 60752
rect 17356 60124 17396 60164
rect 17164 59200 17204 59240
rect 17260 58612 17300 58652
rect 17548 60880 17588 60920
rect 17548 60376 17588 60416
rect 18316 65920 18356 65960
rect 18988 66844 19028 66884
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 18988 66172 19028 66212
rect 18412 64996 18452 65036
rect 18316 64492 18356 64532
rect 18316 63484 18356 63524
rect 18412 63232 18452 63272
rect 18220 63148 18260 63188
rect 18220 61468 18260 61508
rect 17548 59116 17588 59156
rect 17452 58360 17492 58400
rect 19180 65164 19220 65204
rect 18604 64996 18644 65036
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 19372 69112 19412 69152
rect 19468 69028 19508 69068
rect 19372 68608 19412 68648
rect 19948 70456 19988 70496
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 20524 70204 20564 70244
rect 19948 70036 19988 70076
rect 19852 69784 19892 69824
rect 20524 69112 20564 69152
rect 20044 68944 20084 68984
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 19660 68608 19700 68648
rect 19660 67180 19700 67220
rect 19660 67012 19700 67052
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 19852 67180 19892 67220
rect 19756 66172 19796 66212
rect 19468 66088 19508 66128
rect 19372 65500 19412 65540
rect 19276 64408 19316 64448
rect 18604 63568 18644 63608
rect 18508 60796 18548 60836
rect 18412 60208 18452 60248
rect 18220 59368 18260 59408
rect 17644 58528 17684 58568
rect 17356 58024 17396 58064
rect 17068 57856 17108 57896
rect 16972 57688 17012 57728
rect 16780 57184 16820 57224
rect 17356 57604 17396 57644
rect 17548 57940 17588 57980
rect 18124 58528 18164 58568
rect 17836 57772 17876 57812
rect 17836 57604 17876 57644
rect 16876 57100 16916 57140
rect 16108 55084 16148 55124
rect 15916 55000 15956 55040
rect 16108 54916 16148 54956
rect 16012 54412 16052 54452
rect 15916 54244 15956 54284
rect 15916 52480 15956 52520
rect 16108 53992 16148 54032
rect 16492 57016 16532 57056
rect 16972 57016 17012 57056
rect 17260 57016 17300 57056
rect 16780 56680 16820 56720
rect 16588 56344 16628 56384
rect 16972 56596 17012 56636
rect 17644 56596 17684 56636
rect 17932 57520 17972 57560
rect 17836 56344 17876 56384
rect 17740 56260 17780 56300
rect 17356 56176 17396 56216
rect 17644 56092 17684 56132
rect 17164 55924 17204 55964
rect 16972 55588 17012 55628
rect 16492 55000 16532 55040
rect 16300 54412 16340 54452
rect 16492 54412 16532 54452
rect 16300 54244 16340 54284
rect 16204 53572 16244 53612
rect 16108 53236 16148 53276
rect 16108 52228 16148 52268
rect 16012 52060 16052 52100
rect 15724 51892 15764 51932
rect 15820 51724 15860 51764
rect 15724 50968 15764 51008
rect 15724 50716 15764 50756
rect 15052 50548 15092 50588
rect 14380 48784 14420 48824
rect 14764 49204 14804 49244
rect 14668 48952 14708 48992
rect 14284 48532 14324 48572
rect 14380 48028 14420 48068
rect 14572 48532 14612 48572
rect 14188 47272 14228 47312
rect 14476 47272 14516 47312
rect 14092 42736 14132 42776
rect 14380 42736 14420 42776
rect 13996 41560 14036 41600
rect 13708 41392 13748 41432
rect 13420 40972 13460 41012
rect 13132 39880 13172 39920
rect 13132 39712 13172 39752
rect 12940 39628 12980 39668
rect 12652 38284 12692 38324
rect 12844 38872 12884 38912
rect 13036 39460 13076 39500
rect 13708 40888 13748 40928
rect 13324 40636 13364 40676
rect 13516 40552 13556 40592
rect 13324 39712 13364 39752
rect 13228 38956 13268 38996
rect 13708 40216 13748 40256
rect 13612 40132 13652 40172
rect 13516 39964 13556 40004
rect 13420 39544 13460 39584
rect 13228 38788 13268 38828
rect 13132 38704 13172 38744
rect 13132 38536 13172 38576
rect 13132 38116 13172 38156
rect 12844 37276 12884 37316
rect 12748 36688 12788 36728
rect 12844 36604 12884 36644
rect 12268 34840 12308 34880
rect 12556 34840 12596 34880
rect 11980 32152 12020 32192
rect 11980 31312 12020 31352
rect 11980 30556 12020 30596
rect 12556 34672 12596 34712
rect 12364 34336 12404 34376
rect 12268 33160 12308 33200
rect 12268 32908 12308 32948
rect 12172 32236 12212 32276
rect 12460 32236 12500 32276
rect 12844 35680 12884 35720
rect 12748 35092 12788 35132
rect 12844 35008 12884 35048
rect 12748 34672 12788 34712
rect 12652 34000 12692 34040
rect 13036 36520 13076 36560
rect 12652 33832 12692 33872
rect 12556 32068 12596 32108
rect 12652 31312 12692 31352
rect 12652 30556 12692 30596
rect 12268 30388 12308 30428
rect 12652 30220 12692 30260
rect 13228 37444 13268 37484
rect 13324 37360 13364 37400
rect 13228 37276 13268 37316
rect 13132 35428 13172 35468
rect 13324 36604 13364 36644
rect 13420 35428 13460 35468
rect 13132 35008 13172 35048
rect 12940 31984 12980 32024
rect 13132 31984 13172 32024
rect 13804 39460 13844 39500
rect 13708 39292 13748 39332
rect 14284 41728 14324 41768
rect 14188 41476 14228 41516
rect 14092 40300 14132 40340
rect 14188 39880 14228 39920
rect 14380 41308 14420 41348
rect 16588 53404 16628 53444
rect 16492 51892 16532 51932
rect 16684 52060 16724 52100
rect 16108 51724 16148 51764
rect 16108 51556 16148 51596
rect 15628 49708 15668 49748
rect 15052 48784 15092 48824
rect 15532 48784 15572 48824
rect 15916 50296 15956 50336
rect 16300 51724 16340 51764
rect 16204 51220 16244 51260
rect 16300 51052 16340 51092
rect 16300 50884 16340 50924
rect 16588 50380 16628 50420
rect 16204 50296 16244 50336
rect 16108 50128 16148 50168
rect 15916 48784 15956 48824
rect 16396 50128 16436 50168
rect 16300 49540 16340 49580
rect 16588 49456 16628 49496
rect 16396 49120 16436 49160
rect 16492 49036 16532 49076
rect 15724 48700 15764 48740
rect 16012 48616 16052 48656
rect 15436 47776 15476 47816
rect 14956 47440 14996 47480
rect 15916 47944 15956 47984
rect 16108 47776 16148 47816
rect 16588 48784 16628 48824
rect 16492 48364 16532 48404
rect 16588 48028 16628 48068
rect 16492 47944 16532 47984
rect 16300 47776 16340 47816
rect 14956 46432 14996 46472
rect 16300 47356 16340 47396
rect 15724 46348 15764 46388
rect 16204 45340 16244 45380
rect 15052 44248 15092 44288
rect 15148 44164 15188 44204
rect 16012 45004 16052 45044
rect 16204 44248 16244 44288
rect 15436 44164 15476 44204
rect 14956 44080 14996 44120
rect 15244 43408 15284 43448
rect 16204 43408 16244 43448
rect 15148 42568 15188 42608
rect 15148 42148 15188 42188
rect 14956 41560 14996 41600
rect 14860 41476 14900 41516
rect 14668 41308 14708 41348
rect 14668 40972 14708 41012
rect 14380 40804 14420 40844
rect 14476 39880 14516 39920
rect 14284 39796 14324 39836
rect 14188 39712 14228 39752
rect 14860 40888 14900 40928
rect 14764 39880 14804 39920
rect 14380 39628 14420 39668
rect 14476 39544 14516 39584
rect 14668 39544 14708 39584
rect 14380 39460 14420 39500
rect 13996 39292 14036 39332
rect 13804 38620 13844 38660
rect 13996 38284 14036 38324
rect 13900 38200 13940 38240
rect 13804 38032 13844 38072
rect 14092 38032 14132 38072
rect 14284 39292 14324 39332
rect 14572 38872 14612 38912
rect 14860 39124 14900 39164
rect 14476 37612 14516 37652
rect 14668 38200 14708 38240
rect 14284 36772 14324 36812
rect 14572 36772 14612 36812
rect 13612 36688 13652 36728
rect 13612 34504 13652 34544
rect 14092 36604 14132 36644
rect 13804 34420 13844 34460
rect 13708 34252 13748 34292
rect 13612 34000 13652 34040
rect 13516 33832 13556 33872
rect 13324 33664 13364 33704
rect 13228 31312 13268 31352
rect 13420 33580 13460 33620
rect 13420 32908 13460 32948
rect 13036 30976 13076 31016
rect 13324 30976 13364 31016
rect 13228 30808 13268 30848
rect 13132 30640 13172 30680
rect 13516 30808 13556 30848
rect 12940 29884 12980 29924
rect 12364 29128 12404 29168
rect 13036 29800 13076 29840
rect 12940 29548 12980 29588
rect 13132 29548 13172 29588
rect 12652 29212 12692 29252
rect 12460 29044 12500 29084
rect 13132 29128 13172 29168
rect 12652 28960 12692 29000
rect 12844 28708 12884 28748
rect 12748 28288 12788 28328
rect 13612 30556 13652 30596
rect 13996 33664 14036 33704
rect 13900 32572 13940 32612
rect 14476 35680 14516 35720
rect 14476 34756 14516 34796
rect 14188 34336 14228 34376
rect 14188 34000 14228 34040
rect 14092 32404 14132 32444
rect 13900 32152 13940 32192
rect 13996 31564 14036 31604
rect 13900 30640 13940 30680
rect 13516 29884 13556 29924
rect 13708 29968 13748 30008
rect 13420 29716 13460 29756
rect 13420 29044 13460 29084
rect 13036 28876 13076 28916
rect 12652 28120 12692 28160
rect 12076 27868 12116 27908
rect 12268 27868 12308 27908
rect 12556 27868 12596 27908
rect 12940 27784 12980 27824
rect 11980 27616 12020 27656
rect 11500 27448 11540 27488
rect 11822 27448 11862 27488
rect 11500 26020 11540 26060
rect 11500 24592 11540 24632
rect 11500 23920 11540 23960
rect 11884 27280 11924 27320
rect 11692 27028 11732 27068
rect 11692 25012 11732 25052
rect 11692 24592 11732 24632
rect 11980 26860 12020 26900
rect 11884 26608 11924 26648
rect 12268 27616 12308 27656
rect 12172 27448 12212 27488
rect 12364 27364 12404 27404
rect 12844 27616 12884 27656
rect 12652 27448 12692 27488
rect 12556 27364 12596 27404
rect 12076 26776 12116 26816
rect 12268 26776 12308 26816
rect 12556 26776 12596 26816
rect 12172 26104 12212 26144
rect 11884 24928 11924 24968
rect 12844 26524 12884 26564
rect 12652 25264 12692 25304
rect 12268 24928 12308 24968
rect 12364 24592 12404 24632
rect 11596 23752 11636 23792
rect 11692 23416 11732 23456
rect 11596 21652 11636 21692
rect 11308 19888 11348 19928
rect 11404 19552 11444 19592
rect 11308 19300 11348 19340
rect 11308 17368 11348 17408
rect 11308 17032 11348 17072
rect 11308 16108 11348 16148
rect 11308 14428 11348 14468
rect 11212 14008 11252 14048
rect 11308 13756 11348 13796
rect 10540 10900 10580 10940
rect 10540 10312 10580 10352
rect 10348 9220 10388 9260
rect 10348 8884 10388 8924
rect 10252 7456 10292 7496
rect 10156 5944 10196 5984
rect 10252 5692 10292 5732
rect 9868 2752 9908 2792
rect 9868 2416 9908 2456
rect 9772 2332 9812 2372
rect 9388 988 9428 1028
rect 9292 484 9332 524
rect 9580 1492 9620 1532
rect 10252 4768 10292 4808
rect 11116 12916 11156 12956
rect 11116 12496 11156 12536
rect 11020 11740 11060 11780
rect 11212 11740 11252 11780
rect 10828 10900 10868 10940
rect 11596 20140 11636 20180
rect 11596 19132 11636 19172
rect 11596 17032 11636 17072
rect 11500 15352 11540 15392
rect 11500 12496 11540 12536
rect 11884 23752 11924 23792
rect 11884 23416 11924 23456
rect 11884 23080 11924 23120
rect 12172 24340 12212 24380
rect 12364 24172 12404 24212
rect 12748 24424 12788 24464
rect 14764 36100 14804 36140
rect 14956 38872 14996 38912
rect 15532 41392 15572 41432
rect 15820 41896 15860 41936
rect 15916 41476 15956 41516
rect 15244 41140 15284 41180
rect 15436 41140 15476 41180
rect 15436 40636 15476 40676
rect 15340 40552 15380 40592
rect 15148 39964 15188 40004
rect 15244 39880 15284 39920
rect 15148 39544 15188 39584
rect 15436 39712 15476 39752
rect 15340 39040 15380 39080
rect 16492 47272 16532 47312
rect 16588 46768 16628 46808
rect 17068 55504 17108 55544
rect 17068 55000 17108 55040
rect 17452 55672 17492 55712
rect 17260 55168 17300 55208
rect 17836 55168 17876 55208
rect 18124 56008 18164 56048
rect 18124 55672 18164 55712
rect 17164 54412 17204 54452
rect 17836 54328 17876 54368
rect 16972 53992 17012 54032
rect 16876 52984 16916 53024
rect 16780 51976 16820 52016
rect 16780 51640 16820 51680
rect 16972 50296 17012 50336
rect 17740 54160 17780 54200
rect 17644 54076 17684 54116
rect 17164 52396 17204 52436
rect 17164 51976 17204 52016
rect 17644 52900 17684 52940
rect 17548 52816 17588 52856
rect 17452 52396 17492 52436
rect 17548 50968 17588 51008
rect 17356 50716 17396 50756
rect 17548 50716 17588 50756
rect 17164 50380 17204 50420
rect 18028 53656 18068 53696
rect 17740 50464 17780 50504
rect 17644 50380 17684 50420
rect 18028 50464 18068 50504
rect 17932 50296 17972 50336
rect 17068 49036 17108 49076
rect 16972 48364 17012 48404
rect 17260 48280 17300 48320
rect 17260 47944 17300 47984
rect 16972 47776 17012 47816
rect 17164 46768 17204 46808
rect 16972 46432 17012 46472
rect 17356 46432 17396 46472
rect 17452 46012 17492 46052
rect 17356 45760 17396 45800
rect 17356 45592 17396 45632
rect 16972 45340 17012 45380
rect 16108 40888 16148 40928
rect 15532 39544 15572 39584
rect 15244 38788 15284 38828
rect 15244 38368 15284 38408
rect 15148 37528 15188 37568
rect 16108 40636 16148 40676
rect 16396 41728 16436 41768
rect 15724 40552 15764 40592
rect 15820 40468 15860 40508
rect 15724 39964 15764 40004
rect 15724 38368 15764 38408
rect 15436 37864 15476 37904
rect 16108 40300 16148 40340
rect 15244 37360 15284 37400
rect 15052 36856 15092 36896
rect 14956 36100 14996 36140
rect 14860 35680 14900 35720
rect 14668 34336 14708 34376
rect 14668 33664 14708 33704
rect 14476 33160 14516 33200
rect 14380 32992 14420 33032
rect 14572 32656 14612 32696
rect 14284 32068 14324 32108
rect 13132 27952 13172 27992
rect 13516 28624 13556 28664
rect 13516 27952 13556 27992
rect 13708 29464 13748 29504
rect 13804 29296 13844 29336
rect 13804 29044 13844 29084
rect 13900 28960 13940 29000
rect 13804 28876 13844 28916
rect 13708 28624 13748 28664
rect 13708 28372 13748 28412
rect 13708 28120 13748 28160
rect 13324 27784 13364 27824
rect 13228 27700 13268 27740
rect 13324 27616 13364 27656
rect 13228 27448 13268 27488
rect 13132 26104 13172 26144
rect 12460 23920 12500 23960
rect 12844 23920 12884 23960
rect 12844 23752 12884 23792
rect 12748 23500 12788 23540
rect 12268 23080 12308 23120
rect 12556 22996 12596 23036
rect 12652 22660 12692 22700
rect 11884 22576 11924 22616
rect 12556 22576 12596 22616
rect 11788 21484 11828 21524
rect 12364 22408 12404 22448
rect 12364 21904 12404 21944
rect 11980 21652 12020 21692
rect 12268 21400 12308 21440
rect 11980 19720 12020 19760
rect 12076 19636 12116 19676
rect 11980 18880 12020 18920
rect 12076 18796 12116 18836
rect 11884 17032 11924 17072
rect 11692 15604 11732 15644
rect 11692 15436 11732 15476
rect 11788 15352 11828 15392
rect 12844 23416 12884 23456
rect 12748 22408 12788 22448
rect 13036 25348 13076 25388
rect 13132 25264 13172 25304
rect 13324 27112 13364 27152
rect 12748 22240 12788 22280
rect 12844 21316 12884 21356
rect 12844 19972 12884 20012
rect 12364 18880 12404 18920
rect 12268 18796 12308 18836
rect 12268 18544 12308 18584
rect 11884 14092 11924 14132
rect 11692 13840 11732 13880
rect 12172 16024 12212 16064
rect 12460 17788 12500 17828
rect 12460 17620 12500 17660
rect 12556 17200 12596 17240
rect 12268 15184 12308 15224
rect 12076 13756 12116 13796
rect 11596 12328 11636 12368
rect 11596 12160 11636 12200
rect 11596 10060 11636 10100
rect 11404 9976 11444 10016
rect 11788 12328 11828 12368
rect 11788 11404 11828 11444
rect 11980 11152 12020 11192
rect 12172 13504 12212 13544
rect 13228 23920 13268 23960
rect 13132 23752 13172 23792
rect 13324 23332 13364 23372
rect 13228 22996 13268 23036
rect 13132 22744 13172 22784
rect 13228 22492 13268 22532
rect 13132 22240 13172 22280
rect 13324 22240 13364 22280
rect 13228 20476 13268 20516
rect 13516 27364 13556 27404
rect 13708 27280 13748 27320
rect 13612 26104 13652 26144
rect 14188 29968 14228 30008
rect 14188 29716 14228 29756
rect 14092 29380 14132 29420
rect 14380 30052 14420 30092
rect 14572 30052 14612 30092
rect 14476 29884 14516 29924
rect 14284 29464 14324 29504
rect 14284 29296 14324 29336
rect 14476 29044 14516 29084
rect 14572 28708 14612 28748
rect 14375 28624 14415 28664
rect 14476 28624 14516 28664
rect 14092 28372 14132 28412
rect 14380 28120 14420 28160
rect 14284 27616 14324 27656
rect 14188 27196 14228 27236
rect 13900 25264 13940 25304
rect 13516 22240 13556 22280
rect 13516 21484 13556 21524
rect 14764 32992 14804 33032
rect 14764 31144 14804 31184
rect 14860 30640 14900 30680
rect 14860 30136 14900 30176
rect 14764 29548 14804 29588
rect 15436 36940 15476 36980
rect 15628 36940 15668 36980
rect 15532 36520 15572 36560
rect 15724 36688 15764 36728
rect 16300 40300 16340 40340
rect 16300 39040 16340 39080
rect 16012 37444 16052 37484
rect 15916 37360 15956 37400
rect 15820 36604 15860 36644
rect 16108 36604 16148 36644
rect 16300 37780 16340 37820
rect 15628 35680 15668 35720
rect 15820 34336 15860 34376
rect 15244 32992 15284 33032
rect 15052 32320 15092 32360
rect 15052 32152 15092 32192
rect 15340 31648 15380 31688
rect 15148 31144 15188 31184
rect 15244 30640 15284 30680
rect 15244 29800 15284 29840
rect 14860 29296 14900 29336
rect 14956 29212 14996 29252
rect 14956 28960 14996 29000
rect 14860 28708 14900 28748
rect 14668 28372 14708 28412
rect 15244 28876 15284 28916
rect 15820 34000 15860 34040
rect 15724 33832 15764 33872
rect 15724 31564 15764 31604
rect 16012 32824 16052 32864
rect 15628 30556 15668 30596
rect 15628 29800 15668 29840
rect 15436 29464 15476 29504
rect 15532 29380 15572 29420
rect 15148 28624 15188 28664
rect 15052 28288 15092 28328
rect 14956 28120 14996 28160
rect 14860 27616 14900 27656
rect 14956 27280 14996 27320
rect 14764 27028 14804 27068
rect 14572 26944 14612 26984
rect 14956 27028 14996 27068
rect 15148 27112 15188 27152
rect 14572 26608 14612 26648
rect 14476 26440 14516 26480
rect 14284 24928 14324 24968
rect 13996 24508 14036 24548
rect 14092 23920 14132 23960
rect 13996 23248 14036 23288
rect 13996 23080 14036 23120
rect 14380 23836 14420 23876
rect 14380 23668 14420 23708
rect 14188 23080 14228 23120
rect 14092 22660 14132 22700
rect 14284 22660 14324 22700
rect 13900 21820 13940 21860
rect 13708 21568 13748 21608
rect 13900 21568 13940 21608
rect 13996 21064 14036 21104
rect 13420 18964 13460 19004
rect 13612 19216 13652 19256
rect 13516 18628 13556 18668
rect 13420 17536 13460 17576
rect 13324 17032 13364 17072
rect 13132 15604 13172 15644
rect 12940 15268 12980 15308
rect 13228 15520 13268 15560
rect 13996 20728 14036 20768
rect 13900 19384 13940 19424
rect 13804 19216 13844 19256
rect 13804 16192 13844 16232
rect 13324 15436 13364 15476
rect 13228 15268 13268 15308
rect 12844 14428 12884 14468
rect 12652 13252 12692 13292
rect 12364 13168 12404 13208
rect 12748 13168 12788 13208
rect 13036 14176 13076 14216
rect 12940 14092 12980 14132
rect 13228 14176 13268 14216
rect 13324 14008 13364 14048
rect 13228 13756 13268 13796
rect 12844 12496 12884 12536
rect 12748 12328 12788 12368
rect 12652 11572 12692 11612
rect 12364 11152 12404 11192
rect 12556 10396 12596 10436
rect 11788 9976 11828 10016
rect 11980 9976 12020 10016
rect 11020 9640 11060 9680
rect 10924 8716 10964 8756
rect 10444 7960 10484 8000
rect 10732 7960 10772 8000
rect 10540 7456 10580 7496
rect 10828 7288 10868 7328
rect 10540 7120 10580 7160
rect 10732 7120 10772 7160
rect 10732 6616 10772 6656
rect 11116 6952 11156 6992
rect 10924 6280 10964 6320
rect 11500 9556 11540 9596
rect 11500 9220 11540 9260
rect 11692 8380 11732 8420
rect 11500 7120 11540 7160
rect 11404 6280 11444 6320
rect 10732 5608 10772 5648
rect 10444 4936 10484 4976
rect 10828 4516 10868 4556
rect 10636 4432 10676 4472
rect 10156 3592 10196 3632
rect 10348 3928 10388 3968
rect 10828 4180 10868 4220
rect 10252 3508 10292 3548
rect 10060 3340 10100 3380
rect 10156 2584 10196 2624
rect 10060 2164 10100 2204
rect 9772 1408 9812 1448
rect 9676 1240 9716 1280
rect 10540 3340 10580 3380
rect 10540 3172 10580 3212
rect 10348 1996 10388 2036
rect 10060 568 10100 608
rect 10444 904 10484 944
rect 11116 6028 11156 6068
rect 11212 4432 11252 4472
rect 11212 4180 11252 4220
rect 11404 5020 11444 5060
rect 11692 7372 11732 7412
rect 11596 6616 11636 6656
rect 11884 9556 11924 9596
rect 11884 8632 11924 8672
rect 12748 10396 12788 10436
rect 12652 9976 12692 10016
rect 12556 9808 12596 9848
rect 12076 9472 12116 9512
rect 12268 9472 12308 9512
rect 12460 8548 12500 8588
rect 11788 5944 11828 5984
rect 11596 5860 11636 5900
rect 11692 5776 11732 5816
rect 11596 5608 11636 5648
rect 11980 5272 12020 5312
rect 13324 13336 13364 13376
rect 13612 14932 13652 14972
rect 13804 14176 13844 14216
rect 13804 13756 13844 13796
rect 14092 19636 14132 19676
rect 14380 22408 14420 22448
rect 14668 24172 14708 24212
rect 14860 26608 14900 26648
rect 15244 26776 15284 26816
rect 15052 26440 15092 26480
rect 14860 26104 14900 26144
rect 15916 30052 15956 30092
rect 15820 29128 15860 29168
rect 15724 28708 15764 28748
rect 15916 28708 15956 28748
rect 15436 28036 15476 28076
rect 15916 27952 15956 27992
rect 15820 27700 15860 27740
rect 15436 27616 15476 27656
rect 15724 26944 15764 26984
rect 15340 26020 15380 26060
rect 15436 25936 15476 25976
rect 15820 26440 15860 26480
rect 16300 36520 16340 36560
rect 16300 35428 16340 35468
rect 16204 33832 16244 33872
rect 16588 41476 16628 41516
rect 16588 40132 16628 40172
rect 16492 38704 16532 38744
rect 16780 42568 16820 42608
rect 16780 41896 16820 41936
rect 16876 41560 16916 41600
rect 16972 41140 17012 41180
rect 16780 40132 16820 40172
rect 17356 44080 17396 44120
rect 17548 43912 17588 43952
rect 17548 43492 17588 43532
rect 17452 43408 17492 43448
rect 17164 42652 17204 42692
rect 17356 42652 17396 42692
rect 17260 42400 17300 42440
rect 17740 49120 17780 49160
rect 18124 49372 18164 49412
rect 18124 49120 18164 49160
rect 18124 48364 18164 48404
rect 17836 47944 17876 47984
rect 17932 47272 17972 47312
rect 18412 54832 18452 54872
rect 18316 53656 18356 53696
rect 18700 63484 18740 63524
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 18604 58696 18644 58736
rect 18988 63064 19028 63104
rect 19372 63820 19412 63860
rect 19756 65668 19796 65708
rect 19660 64408 19700 64448
rect 20620 68104 20660 68144
rect 20524 66760 20564 66800
rect 20524 66088 20564 66128
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 21100 72472 21140 72512
rect 20716 67096 20756 67136
rect 20620 64996 20660 65036
rect 20524 64912 20564 64952
rect 19852 64828 19892 64868
rect 19852 64576 19892 64616
rect 20044 64408 20084 64448
rect 20620 64408 20660 64448
rect 19756 63316 19796 63356
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 19948 63652 19988 63692
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 19660 62644 19700 62684
rect 19564 61552 19604 61592
rect 19372 61468 19412 61508
rect 19852 62308 19892 62348
rect 19756 61636 19796 61676
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 20524 62728 20564 62768
rect 19276 60880 19316 60920
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 18892 60292 18932 60332
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 19564 59872 19604 59912
rect 19756 61048 19796 61088
rect 19756 59620 19796 59660
rect 19564 59452 19604 59492
rect 19756 59284 19796 59324
rect 19756 59116 19796 59156
rect 19660 58612 19700 58652
rect 19276 57940 19316 57980
rect 19084 57856 19124 57896
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 18700 56176 18740 56216
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 18604 55756 18644 55796
rect 18700 55588 18740 55628
rect 19372 56344 19412 56384
rect 19372 56176 19412 56216
rect 19372 55420 19412 55460
rect 18892 55084 18932 55124
rect 19276 55084 19316 55124
rect 19276 54916 19316 54956
rect 18892 54664 18932 54704
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 19084 53992 19124 54032
rect 18892 53824 18932 53864
rect 20524 61888 20564 61928
rect 20044 61468 20084 61508
rect 19948 61384 19988 61424
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 20044 60796 20084 60836
rect 20236 60628 20276 60668
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 19948 59116 19988 59156
rect 19852 58696 19892 58736
rect 19564 56848 19604 56888
rect 19756 57268 19796 57308
rect 19756 56932 19796 56972
rect 20044 58612 20084 58652
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 19948 57016 19988 57056
rect 19852 56764 19892 56804
rect 19756 56428 19796 56468
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 19756 56092 19796 56132
rect 19948 56092 19988 56132
rect 19660 56008 19700 56048
rect 19756 55756 19796 55796
rect 20524 55672 20564 55712
rect 19564 55504 19604 55544
rect 20044 55504 20084 55544
rect 19564 54916 19604 54956
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 19756 54748 19796 54788
rect 19948 54748 19988 54788
rect 19564 54160 19604 54200
rect 19276 53992 19316 54032
rect 19660 54076 19700 54116
rect 19180 53488 19220 53528
rect 19084 53320 19124 53360
rect 18892 53068 18932 53108
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 18412 51808 18452 51848
rect 18988 52648 19028 52688
rect 19180 52312 19220 52352
rect 19084 51892 19124 51932
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 18316 50800 18356 50840
rect 19180 50296 19220 50336
rect 19564 53320 19604 53360
rect 19756 53740 19796 53780
rect 19660 52900 19700 52940
rect 20236 53992 20276 54032
rect 20044 53824 20084 53864
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 19948 53404 19988 53444
rect 19948 53236 19988 53276
rect 19852 52984 19892 53024
rect 19468 52648 19508 52688
rect 19756 52564 19796 52604
rect 19372 52144 19412 52184
rect 19564 51976 19604 52016
rect 19756 51724 19796 51764
rect 19564 51640 19604 51680
rect 19564 50968 19604 51008
rect 19564 50296 19604 50336
rect 18604 50044 18644 50084
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 18508 49372 18548 49412
rect 18412 49120 18452 49160
rect 18316 48952 18356 48992
rect 18316 47524 18356 47564
rect 18316 47272 18356 47312
rect 19084 49456 19124 49496
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 19276 48196 19316 48236
rect 18892 47440 18932 47480
rect 18508 47272 18548 47312
rect 18796 47272 18836 47312
rect 18892 47020 18932 47060
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 17836 46012 17876 46052
rect 17932 44668 17972 44708
rect 17740 43660 17780 43700
rect 17644 42400 17684 42440
rect 18988 46684 19028 46724
rect 18412 45928 18452 45968
rect 18796 45928 18836 45968
rect 18700 45760 18740 45800
rect 18700 45424 18740 45464
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 18316 45172 18356 45212
rect 18508 44920 18548 44960
rect 18316 44500 18356 44540
rect 18124 44416 18164 44456
rect 18124 42904 18164 42944
rect 17932 42736 17972 42776
rect 17932 42568 17972 42608
rect 17836 42148 17876 42188
rect 17836 41560 17876 41600
rect 17740 41476 17780 41516
rect 17644 41308 17684 41348
rect 17164 41140 17204 41180
rect 17068 40132 17108 40172
rect 16972 38872 17012 38912
rect 16684 37528 16724 37568
rect 16684 36772 16724 36812
rect 16492 35680 16532 35720
rect 16588 33664 16628 33704
rect 16684 33412 16724 33452
rect 16588 33328 16628 33368
rect 16300 32068 16340 32108
rect 16300 30976 16340 31016
rect 16684 30976 16724 31016
rect 16492 30808 16532 30848
rect 16492 30640 16532 30680
rect 16396 30472 16436 30512
rect 17452 40636 17492 40676
rect 17452 40132 17492 40172
rect 17740 40972 17780 41012
rect 18220 42316 18260 42356
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 20140 52648 20180 52688
rect 19948 52312 19988 52352
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 20140 51640 20180 51680
rect 20140 50968 20180 51008
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 19948 50548 19988 50588
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 19372 47944 19412 47984
rect 19372 47524 19412 47564
rect 19564 47272 19604 47312
rect 19372 46096 19412 46136
rect 19468 45844 19508 45884
rect 18796 43660 18836 43700
rect 18604 43324 18644 43364
rect 18796 42652 18836 42692
rect 19180 43240 19220 43280
rect 18988 42820 19028 42860
rect 18604 42400 18644 42440
rect 18124 42064 18164 42104
rect 17932 41140 17972 41180
rect 17836 40720 17876 40760
rect 17740 39796 17780 39836
rect 17548 39124 17588 39164
rect 17836 39040 17876 39080
rect 17644 38788 17684 38828
rect 16876 37696 16916 37736
rect 17068 36856 17108 36896
rect 16972 36268 17012 36308
rect 16876 35596 16916 35636
rect 16876 35428 16916 35468
rect 16876 35008 16916 35048
rect 16780 30136 16820 30176
rect 17068 35176 17108 35216
rect 17356 36604 17396 36644
rect 17452 36520 17492 36560
rect 17836 38452 17876 38492
rect 17836 38200 17876 38240
rect 17548 36268 17588 36308
rect 17260 35428 17300 35468
rect 17452 35428 17492 35468
rect 17356 35176 17396 35216
rect 17260 35092 17300 35132
rect 17068 34756 17108 34796
rect 16972 30472 17012 30512
rect 16876 29044 16916 29084
rect 16396 28120 16436 28160
rect 16204 27784 16244 27824
rect 16588 28120 16628 28160
rect 16588 27616 16628 27656
rect 16396 26776 16436 26816
rect 16108 26440 16148 26480
rect 15628 25684 15668 25724
rect 15148 25264 15188 25304
rect 14764 23836 14804 23876
rect 14572 23584 14612 23624
rect 14860 23584 14900 23624
rect 14764 23248 14804 23288
rect 15244 25180 15284 25220
rect 15532 25180 15572 25220
rect 15340 24592 15380 24632
rect 15244 24508 15284 24548
rect 15148 23752 15188 23792
rect 15052 23248 15092 23288
rect 14764 23080 14804 23120
rect 15148 23080 15188 23120
rect 15436 23836 15476 23876
rect 15532 23668 15572 23708
rect 14572 22744 14612 22784
rect 15052 22744 15092 22784
rect 14471 21988 14511 22028
rect 14476 21820 14516 21860
rect 14284 20056 14324 20096
rect 14188 19384 14228 19424
rect 14092 19048 14132 19088
rect 13996 17200 14036 17240
rect 14284 18964 14324 19004
rect 14476 18964 14516 19004
rect 14764 21568 14804 21608
rect 14764 21400 14804 21440
rect 14956 21736 14996 21776
rect 16204 26104 16244 26144
rect 16780 28288 16820 28328
rect 16780 27532 16820 27572
rect 17068 27532 17108 27572
rect 16972 26944 17012 26984
rect 16780 26776 16820 26816
rect 16588 26440 16628 26480
rect 16492 26272 16532 26312
rect 16204 25936 16244 25976
rect 16396 25936 16436 25976
rect 16108 25516 16148 25556
rect 16108 25348 16148 25388
rect 16012 25264 16052 25304
rect 16300 25264 16340 25304
rect 16492 25264 16532 25304
rect 16204 24928 16244 24968
rect 15916 24508 15956 24548
rect 16108 24508 16148 24548
rect 15724 24340 15764 24380
rect 16108 24340 16148 24380
rect 16396 24844 16436 24884
rect 16300 24592 16340 24632
rect 16684 25684 16724 25724
rect 16972 26608 17012 26648
rect 16876 26104 16916 26144
rect 16780 25432 16820 25472
rect 16588 25180 16628 25220
rect 16492 24088 16532 24128
rect 15724 23836 15764 23876
rect 15724 23500 15764 23540
rect 15628 23332 15668 23372
rect 15532 22912 15572 22952
rect 16300 23836 16340 23876
rect 16204 23164 16244 23204
rect 15820 23080 15860 23120
rect 15724 22744 15764 22784
rect 15724 22240 15764 22280
rect 15340 21736 15380 21776
rect 15916 21988 15956 22028
rect 15820 21736 15860 21776
rect 15532 21568 15572 21608
rect 15244 21484 15284 21524
rect 14956 21400 14996 21440
rect 15148 21400 15188 21440
rect 14956 20728 14996 20768
rect 15340 21400 15380 21440
rect 15436 20728 15476 20768
rect 15340 20560 15380 20600
rect 15724 21484 15764 21524
rect 16017 21400 16057 21440
rect 15724 20980 15764 21020
rect 16108 20728 16148 20768
rect 15244 20224 15284 20264
rect 15052 19804 15092 19844
rect 14860 19552 14900 19592
rect 14668 19132 14708 19172
rect 14860 19132 14900 19172
rect 14764 19048 14804 19088
rect 14668 18880 14708 18920
rect 14188 18712 14228 18752
rect 14572 18712 14612 18752
rect 14764 18712 14804 18752
rect 14092 16024 14132 16064
rect 13996 13420 14036 13460
rect 14476 18628 14516 18668
rect 14668 18544 14708 18584
rect 14476 18208 14516 18248
rect 14284 17956 14324 17996
rect 14284 16780 14324 16820
rect 15436 19720 15476 19760
rect 15148 18964 15188 19004
rect 15052 18544 15092 18584
rect 14860 17956 14900 17996
rect 14572 17200 14612 17240
rect 14572 16948 14612 16988
rect 14476 16024 14516 16064
rect 14764 16780 14804 16820
rect 14668 15520 14708 15560
rect 14380 14764 14420 14804
rect 14764 14764 14804 14804
rect 14188 14344 14228 14384
rect 14956 15100 14996 15140
rect 14092 12748 14132 12788
rect 14956 14428 14996 14468
rect 14380 13168 14420 13208
rect 14284 12832 14324 12872
rect 15724 19384 15764 19424
rect 15628 19216 15668 19256
rect 15532 18964 15572 19004
rect 15628 18880 15668 18920
rect 15436 18544 15476 18584
rect 15436 17788 15476 17828
rect 15244 17620 15284 17660
rect 15148 17032 15188 17072
rect 15244 16948 15284 16988
rect 15916 20056 15956 20096
rect 15820 19132 15860 19172
rect 16108 19720 16148 19760
rect 16012 19552 16052 19592
rect 15724 17200 15764 17240
rect 15724 17032 15764 17072
rect 15532 16024 15572 16064
rect 15724 16192 15764 16232
rect 15724 16024 15764 16064
rect 15724 15688 15764 15728
rect 15436 15520 15476 15560
rect 15340 15436 15380 15476
rect 15244 15016 15284 15056
rect 15244 14764 15284 14804
rect 15628 15520 15668 15560
rect 15532 15100 15572 15140
rect 16108 19132 16148 19172
rect 16108 18628 16148 18668
rect 15916 16108 15956 16148
rect 16684 24004 16724 24044
rect 16684 23752 16724 23792
rect 16492 22996 16532 23036
rect 16396 22576 16436 22616
rect 16972 25264 17012 25304
rect 17068 24172 17108 24212
rect 16972 24088 17012 24128
rect 17356 33412 17396 33452
rect 17260 31396 17300 31436
rect 17260 30640 17300 30680
rect 17740 35176 17780 35216
rect 18316 41392 18356 41432
rect 18220 40636 18260 40676
rect 18124 39964 18164 40004
rect 18114 39796 18154 39836
rect 18508 41308 18548 41348
rect 18412 39880 18452 39920
rect 18124 38620 18164 38660
rect 18124 36856 18164 36896
rect 17932 36520 17972 36560
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 18988 42148 19028 42188
rect 19180 41980 19220 42020
rect 18796 41140 18836 41180
rect 19180 40972 19220 41012
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 19372 43156 19412 43196
rect 19372 42484 19412 42524
rect 19372 42148 19412 42188
rect 19372 40972 19412 41012
rect 19276 40636 19316 40676
rect 19756 45844 19796 45884
rect 19564 45508 19604 45548
rect 19564 44080 19604 44120
rect 19564 42736 19604 42776
rect 19564 41728 19604 41768
rect 19756 45676 19796 45716
rect 19756 45424 19796 45464
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 20044 47356 20084 47396
rect 19948 46936 19988 46976
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 19948 45508 19988 45548
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 19852 44248 19892 44288
rect 20524 44248 20564 44288
rect 20908 67768 20948 67808
rect 20812 66004 20852 66044
rect 20812 65752 20852 65792
rect 20812 64156 20852 64196
rect 21004 66760 21044 66800
rect 21004 64660 21044 64700
rect 20908 63820 20948 63860
rect 20716 63736 20756 63776
rect 20812 63652 20852 63692
rect 20716 60628 20756 60668
rect 21004 63064 21044 63104
rect 20908 59872 20948 59912
rect 20812 59704 20852 59744
rect 20716 57016 20756 57056
rect 20812 56848 20852 56888
rect 20716 52816 20756 52856
rect 20908 47272 20948 47312
rect 20812 45928 20852 45968
rect 20716 44584 20756 44624
rect 20620 44080 20660 44120
rect 19756 43996 19796 44036
rect 19756 43744 19796 43784
rect 19948 43660 19988 43700
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 20908 42904 20948 42944
rect 19948 42484 19988 42524
rect 20140 42148 20180 42188
rect 19756 42064 19796 42104
rect 19756 41728 19796 41768
rect 19948 41560 19988 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 20236 41392 20276 41432
rect 19564 41224 19604 41264
rect 19660 40972 19700 41012
rect 19180 40132 19220 40172
rect 18508 39040 18548 39080
rect 18412 38872 18452 38912
rect 18604 38788 18644 38828
rect 18316 38620 18356 38660
rect 18508 38620 18548 38660
rect 19180 39460 19220 39500
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 19084 39124 19124 39164
rect 18796 38872 18836 38912
rect 18700 38536 18740 38576
rect 18316 38200 18356 38240
rect 18316 37192 18356 37232
rect 18988 38872 19028 38912
rect 18892 38788 18932 38828
rect 18604 38200 18644 38240
rect 20044 41140 20084 41180
rect 19948 40384 19988 40424
rect 19468 40300 19508 40340
rect 20524 40216 20564 40256
rect 19468 39124 19508 39164
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 19852 39880 19892 39920
rect 20140 39544 20180 39584
rect 19468 38956 19508 38996
rect 19372 37948 19412 37988
rect 19276 37864 19316 37904
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18220 35764 18260 35804
rect 18124 35680 18164 35720
rect 18124 35428 18164 35468
rect 17932 35260 17972 35300
rect 17836 35092 17876 35132
rect 18700 37360 18740 37400
rect 18892 37192 18932 37232
rect 19372 36688 19412 36728
rect 18508 36520 18548 36560
rect 18796 36520 18836 36560
rect 19564 38368 19604 38408
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 19468 36268 19508 36308
rect 18508 35764 18548 35804
rect 18508 35176 18548 35216
rect 17740 34336 17780 34376
rect 17644 34000 17684 34040
rect 17644 33748 17684 33788
rect 17932 34000 17972 34040
rect 17932 33076 17972 33116
rect 17932 32824 17972 32864
rect 18412 34000 18452 34040
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18700 34000 18740 34040
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 19756 38116 19796 38156
rect 19948 38032 19988 38072
rect 19756 37360 19796 37400
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 19756 35764 19796 35804
rect 19852 35260 19892 35300
rect 19756 35176 19796 35216
rect 18892 33748 18932 33788
rect 18316 32068 18356 32108
rect 17452 31396 17492 31436
rect 17932 31312 17972 31352
rect 18124 31312 18164 31352
rect 17452 30724 17492 30764
rect 19084 33496 19124 33536
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 19180 33076 19220 33116
rect 19660 34336 19700 34376
rect 19564 34252 19604 34292
rect 19468 33748 19508 33788
rect 18796 32740 18836 32780
rect 19564 33580 19604 33620
rect 19468 32740 19508 32780
rect 18604 32068 18644 32108
rect 18508 31228 18548 31268
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18988 31396 19028 31436
rect 17836 29632 17876 29672
rect 17644 29212 17684 29252
rect 17548 29044 17588 29084
rect 17260 28876 17300 28916
rect 17356 27448 17396 27488
rect 17260 26944 17300 26984
rect 17356 26104 17396 26144
rect 17164 23920 17204 23960
rect 17260 23752 17300 23792
rect 16876 23164 16916 23204
rect 16972 23080 17012 23120
rect 16684 22828 16724 22868
rect 16780 22660 16820 22700
rect 16588 22492 16628 22532
rect 16300 21316 16340 21356
rect 16396 20728 16436 20768
rect 17548 24088 17588 24128
rect 17740 29044 17780 29084
rect 17932 29128 17972 29168
rect 18124 29632 18164 29672
rect 18220 29380 18260 29420
rect 18028 28876 18068 28916
rect 17932 28624 17972 28664
rect 17836 28288 17876 28328
rect 17932 28036 17972 28076
rect 17836 27868 17876 27908
rect 17932 27700 17972 27740
rect 17740 26860 17780 26900
rect 18028 27616 18068 27656
rect 17740 26356 17780 26396
rect 17740 25936 17780 25976
rect 17740 24508 17780 24548
rect 17356 23668 17396 23708
rect 17260 23416 17300 23456
rect 17452 23332 17492 23372
rect 17356 23248 17396 23288
rect 17452 23080 17492 23120
rect 17068 21484 17108 21524
rect 16684 20644 16724 20684
rect 16588 20392 16628 20432
rect 16492 19384 16532 19424
rect 16396 19300 16436 19340
rect 16300 19132 16340 19172
rect 16300 18544 16340 18584
rect 16300 17956 16340 17996
rect 16204 17788 16244 17828
rect 16876 20728 16916 20768
rect 16972 20560 17012 20600
rect 17260 20560 17300 20600
rect 16876 20308 16916 20348
rect 17068 20308 17108 20348
rect 16972 20140 17012 20180
rect 17356 20308 17396 20348
rect 16972 19888 17012 19928
rect 17260 19888 17300 19928
rect 17164 19300 17204 19340
rect 16684 19132 16724 19172
rect 16588 18544 16628 18584
rect 17164 19048 17204 19088
rect 16780 18796 16820 18836
rect 17644 23836 17684 23876
rect 17644 23584 17684 23624
rect 17644 20728 17684 20768
rect 17548 20560 17588 20600
rect 17452 20224 17492 20264
rect 17452 19804 17492 19844
rect 16684 17956 16724 17996
rect 16684 17788 16724 17828
rect 16876 18544 16916 18584
rect 17740 19888 17780 19928
rect 17644 18544 17684 18584
rect 17452 18376 17492 18416
rect 16780 17620 16820 17660
rect 16396 17032 16436 17072
rect 16012 16024 16052 16064
rect 16300 16024 16340 16064
rect 16204 15940 16244 15980
rect 16108 15772 16148 15812
rect 16012 15688 16052 15728
rect 15724 15100 15764 15140
rect 14668 13840 14708 13880
rect 14572 12496 14612 12536
rect 13708 11404 13748 11444
rect 13036 10648 13076 10688
rect 13228 10648 13268 10688
rect 12844 9472 12884 9512
rect 12652 8800 12692 8840
rect 12172 5608 12212 5648
rect 12460 7456 12500 7496
rect 12364 6364 12404 6404
rect 12076 5104 12116 5144
rect 12076 4936 12116 4976
rect 11596 4768 11636 4808
rect 12268 5020 12308 5060
rect 12172 4684 12212 4724
rect 11884 4264 11924 4304
rect 11308 4096 11348 4136
rect 11404 3928 11444 3968
rect 11980 3928 12020 3968
rect 11020 3256 11060 3296
rect 10828 2836 10868 2876
rect 11116 2836 11156 2876
rect 10732 2584 10772 2624
rect 10636 1996 10676 2036
rect 11116 2332 11156 2372
rect 11116 2164 11156 2204
rect 10636 1408 10676 1448
rect 11308 2332 11348 2372
rect 11308 2080 11348 2120
rect 10348 568 10388 608
rect 11212 988 11252 1028
rect 11020 232 11060 272
rect 11884 3508 11924 3548
rect 11500 3340 11540 3380
rect 11692 2584 11732 2624
rect 11596 2164 11636 2204
rect 11500 1744 11540 1784
rect 11500 1324 11540 1364
rect 11788 2080 11828 2120
rect 11980 1912 12020 1952
rect 11980 1660 12020 1700
rect 11884 1156 11924 1196
rect 11884 820 11924 860
rect 12556 7036 12596 7076
rect 12556 6448 12596 6488
rect 12940 8716 12980 8756
rect 12844 8632 12884 8672
rect 12940 8380 12980 8420
rect 13036 8212 13076 8252
rect 12844 7792 12884 7832
rect 12844 6868 12884 6908
rect 12652 6112 12692 6152
rect 12556 4768 12596 4808
rect 12556 3844 12596 3884
rect 12172 2836 12212 2876
rect 12268 2752 12308 2792
rect 12268 2332 12308 2372
rect 12268 1912 12308 1952
rect 12364 1240 12404 1280
rect 12748 4348 12788 4388
rect 12844 3088 12884 3128
rect 12940 2584 12980 2624
rect 13132 6868 13172 6908
rect 13420 10228 13460 10268
rect 13324 9472 13364 9512
rect 13228 6448 13268 6488
rect 13132 6280 13172 6320
rect 13516 10060 13556 10100
rect 13420 8632 13460 8672
rect 13900 10228 13940 10268
rect 13708 8548 13748 8588
rect 13708 7960 13748 8000
rect 13612 7456 13652 7496
rect 13324 6112 13364 6152
rect 13228 4852 13268 4892
rect 13132 4348 13172 4388
rect 13132 3592 13172 3632
rect 13132 3256 13172 3296
rect 13132 2836 13172 2876
rect 13036 2332 13076 2372
rect 12748 1912 12788 1952
rect 13516 6448 13556 6488
rect 13804 7876 13844 7916
rect 14092 8548 14132 8588
rect 14572 11992 14612 12032
rect 14764 12832 14804 12872
rect 14764 12076 14804 12116
rect 14284 11488 14324 11528
rect 14284 10228 14324 10268
rect 14284 10060 14324 10100
rect 14476 11488 14516 11528
rect 14476 11152 14516 11192
rect 14476 10816 14516 10856
rect 14668 11152 14708 11192
rect 14764 10228 14804 10268
rect 14188 8212 14228 8252
rect 14380 9640 14420 9680
rect 15340 14008 15380 14048
rect 15148 13504 15188 13544
rect 15052 11824 15092 11864
rect 15628 14596 15668 14636
rect 15244 13168 15284 13208
rect 15244 11740 15284 11780
rect 14956 9976 14996 10016
rect 14860 9136 14900 9176
rect 14764 8632 14804 8672
rect 14284 8128 14324 8168
rect 14092 7960 14132 8000
rect 14188 7540 14228 7580
rect 13516 4936 13556 4976
rect 13804 4936 13844 4976
rect 13516 4348 13556 4388
rect 13516 4180 13556 4220
rect 13708 4096 13748 4136
rect 14092 6448 14132 6488
rect 14092 5608 14132 5648
rect 14668 7456 14708 7496
rect 14860 7540 14900 7580
rect 14764 7372 14804 7412
rect 15052 8128 15092 8168
rect 15244 8548 15284 8588
rect 15532 13420 15572 13460
rect 15724 13420 15764 13460
rect 15724 13252 15764 13292
rect 15628 11740 15668 11780
rect 15820 13168 15860 13208
rect 15820 12664 15860 12704
rect 15820 10984 15860 11024
rect 16300 15520 16340 15560
rect 16204 15352 16244 15392
rect 16012 15268 16052 15308
rect 16300 15268 16340 15308
rect 16204 14932 16244 14972
rect 16012 14008 16052 14048
rect 16204 13420 16244 13460
rect 16108 13168 16148 13208
rect 16300 12496 16340 12536
rect 15916 10480 15956 10520
rect 16300 12328 16340 12368
rect 16588 16192 16628 16232
rect 16492 16024 16532 16064
rect 16588 15688 16628 15728
rect 16492 15604 16532 15644
rect 16492 15352 16532 15392
rect 16684 15268 16724 15308
rect 16588 14764 16628 14804
rect 16588 14008 16628 14048
rect 16492 13840 16532 13880
rect 16588 13420 16628 13460
rect 16492 13252 16532 13292
rect 16300 11152 16340 11192
rect 16204 10900 16244 10940
rect 15628 9472 15668 9512
rect 15436 8716 15476 8756
rect 15532 8548 15572 8588
rect 15340 8296 15380 8336
rect 15244 8212 15284 8252
rect 15532 8212 15572 8252
rect 15244 7624 15284 7664
rect 14284 7036 14324 7076
rect 14572 7036 14612 7076
rect 14380 6364 14420 6404
rect 14188 5356 14228 5396
rect 14476 5776 14516 5816
rect 14572 5692 14612 5732
rect 14284 4264 14324 4304
rect 14092 3508 14132 3548
rect 13708 3340 13748 3380
rect 13612 2920 13652 2960
rect 13324 2416 13364 2456
rect 12748 1240 12788 1280
rect 13324 1240 13364 1280
rect 12652 1156 12692 1196
rect 12556 904 12596 944
rect 13132 1156 13172 1196
rect 12940 904 12980 944
rect 13900 1324 13940 1364
rect 13900 1156 13940 1196
rect 13996 1072 14036 1112
rect 13900 904 13940 944
rect 13516 820 13556 860
rect 13708 736 13748 776
rect 14284 2836 14324 2876
rect 14188 2668 14228 2708
rect 14188 2416 14228 2456
rect 14380 2416 14420 2456
rect 15340 7540 15380 7580
rect 14860 7036 14900 7076
rect 15052 7036 15092 7076
rect 14860 6532 14900 6572
rect 14764 5776 14804 5816
rect 15052 5608 15092 5648
rect 14956 4852 14996 4892
rect 14956 4096 14996 4136
rect 14572 2668 14612 2708
rect 15052 3424 15092 3464
rect 15052 3172 15092 3212
rect 14668 2584 14708 2624
rect 14380 1912 14420 1952
rect 14764 1912 14804 1952
rect 14284 904 14324 944
rect 14188 484 14228 524
rect 14860 484 14900 524
rect 14668 316 14708 356
rect 16396 10144 16436 10184
rect 16012 9976 16052 10016
rect 16204 9976 16244 10016
rect 16108 8716 16148 8756
rect 15820 8296 15860 8336
rect 15724 8128 15764 8168
rect 15628 6280 15668 6320
rect 15436 6196 15476 6236
rect 16012 8128 16052 8168
rect 15916 7876 15956 7916
rect 16492 9640 16532 9680
rect 16492 9052 16532 9092
rect 16396 8968 16436 9008
rect 16204 7876 16244 7916
rect 16300 6952 16340 6992
rect 17548 18292 17588 18332
rect 17356 17032 17396 17072
rect 17260 16276 17300 16316
rect 17164 16024 17204 16064
rect 16972 15772 17012 15812
rect 16876 15604 16916 15644
rect 16972 15268 17012 15308
rect 16876 14764 16916 14804
rect 17068 14512 17108 14552
rect 16588 8212 16628 8252
rect 16492 7456 16532 7496
rect 16588 7288 16628 7328
rect 16588 6868 16628 6908
rect 16108 6448 16148 6488
rect 16492 6448 16532 6488
rect 16204 6280 16244 6320
rect 16492 6280 16532 6320
rect 15532 4936 15572 4976
rect 15724 4936 15764 4976
rect 15532 4096 15572 4136
rect 15916 4852 15956 4892
rect 15820 4012 15860 4052
rect 15340 3844 15380 3884
rect 15244 3424 15284 3464
rect 15820 3844 15860 3884
rect 15628 3676 15668 3716
rect 15724 3508 15764 3548
rect 15628 2752 15668 2792
rect 15244 2584 15284 2624
rect 15148 2080 15188 2120
rect 16204 5020 16244 5060
rect 16300 4936 16340 4976
rect 16108 3676 16148 3716
rect 16204 3592 16244 3632
rect 16012 3508 16052 3548
rect 16204 3088 16244 3128
rect 15244 1912 15284 1952
rect 15820 1912 15860 1952
rect 16012 1912 16052 1952
rect 16204 1660 16244 1700
rect 15340 1576 15380 1616
rect 15244 1324 15284 1364
rect 15436 1492 15476 1532
rect 15244 232 15284 272
rect 15532 1072 15572 1112
rect 15820 1072 15860 1112
rect 15628 736 15668 776
rect 16012 820 16052 860
rect 16396 3172 16436 3212
rect 16780 10984 16820 11024
rect 16972 14008 17012 14048
rect 17068 13084 17108 13124
rect 16972 12496 17012 12536
rect 16972 10144 17012 10184
rect 16876 8632 16916 8672
rect 17452 15856 17492 15896
rect 17452 15604 17492 15644
rect 17260 14764 17300 14804
rect 17644 17956 17684 17996
rect 17932 26272 17972 26312
rect 19276 30724 19316 30764
rect 18796 30640 18836 30680
rect 18604 29716 18644 29756
rect 18412 29044 18452 29084
rect 18508 28624 18548 28664
rect 19468 32236 19508 32276
rect 19660 30640 19700 30680
rect 19372 30556 19412 30596
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 19468 30472 19508 30512
rect 19372 29800 19412 29840
rect 19276 29380 19316 29420
rect 18796 29212 18836 29252
rect 18988 29212 19028 29252
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18604 28288 18644 28328
rect 18988 28288 19028 28328
rect 19084 27952 19124 27992
rect 19276 27784 19316 27824
rect 18796 27700 18836 27740
rect 18124 27448 18164 27488
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18316 26608 18356 26648
rect 18508 26356 18548 26396
rect 19276 26440 19316 26480
rect 19564 28204 19604 28244
rect 18700 26272 18740 26312
rect 18316 26104 18356 26144
rect 18508 26104 18548 26144
rect 18796 26104 18836 26144
rect 18700 25852 18740 25892
rect 19276 25852 19316 25892
rect 18604 25600 18644 25640
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18700 25348 18740 25388
rect 18316 25264 18356 25304
rect 18124 25180 18164 25220
rect 18604 24256 18644 24296
rect 18124 23836 18164 23876
rect 18028 23752 18068 23792
rect 17932 23248 17972 23288
rect 18028 23164 18068 23204
rect 17932 22660 17972 22700
rect 17932 21316 17972 21356
rect 17932 20392 17972 20432
rect 18412 23752 18452 23792
rect 18220 23080 18260 23120
rect 18316 22744 18356 22784
rect 18220 22408 18260 22448
rect 18412 22660 18452 22700
rect 18604 23920 18644 23960
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 19948 34672 19988 34712
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 20620 39796 20660 39836
rect 20044 33244 20084 33284
rect 20524 33244 20564 33284
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20140 31144 20180 31184
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20044 30556 20084 30596
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20236 28792 20276 28832
rect 20044 28293 20084 28328
rect 20044 28288 20084 28293
rect 20524 28288 20564 28328
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 20044 27616 20084 27656
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 18988 24676 19028 24716
rect 19372 24676 19412 24716
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 18700 23080 18740 23120
rect 18796 22996 18836 23036
rect 18508 22408 18548 22448
rect 18604 22240 18644 22280
rect 18124 21652 18164 21692
rect 18412 21652 18452 21692
rect 18028 20140 18068 20180
rect 18028 19216 18068 19256
rect 17740 17200 17780 17240
rect 17932 17536 17972 17576
rect 17644 16276 17684 16316
rect 17548 15268 17588 15308
rect 17548 14680 17588 14720
rect 17260 11656 17300 11696
rect 17164 11404 17204 11444
rect 17164 11236 17204 11276
rect 17740 15520 17780 15560
rect 18316 21316 18356 21356
rect 18508 21316 18548 21356
rect 18220 20140 18260 20180
rect 18220 19552 18260 19592
rect 19276 22912 19316 22952
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 19276 22576 19316 22616
rect 19084 22492 19124 22532
rect 18988 22408 19028 22448
rect 18892 22240 18932 22280
rect 18988 21568 19028 21608
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18604 19888 18644 19928
rect 18316 19216 18356 19256
rect 18604 18880 18644 18920
rect 18508 18628 18548 18668
rect 18316 18292 18356 18332
rect 18412 18208 18452 18248
rect 18316 17200 18356 17240
rect 18316 16444 18356 16484
rect 18028 16192 18068 16232
rect 18604 17956 18644 17996
rect 18604 17788 18644 17828
rect 18988 20140 19028 20180
rect 18796 19972 18836 20012
rect 19084 19972 19124 20012
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 18796 18880 18836 18920
rect 19468 23416 19508 23456
rect 19372 22408 19412 22448
rect 19564 22576 19604 22616
rect 19852 23752 19892 23792
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20236 24676 20276 24716
rect 20044 23920 20084 23960
rect 20044 23668 20084 23708
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 20716 36184 20756 36224
rect 20812 35932 20852 35972
rect 20716 34504 20756 34544
rect 21196 63736 21236 63776
rect 21100 52900 21140 52940
rect 21004 42400 21044 42440
rect 21004 42232 21044 42272
rect 21100 42148 21140 42188
rect 21292 62476 21332 62516
rect 21292 54160 21332 54200
rect 21388 49792 21428 49832
rect 21388 49288 21428 49328
rect 21292 48952 21332 48992
rect 21292 47356 21332 47396
rect 21196 41812 21236 41852
rect 21100 41560 21140 41600
rect 21196 41224 21236 41264
rect 21004 39880 21044 39920
rect 21100 36604 21140 36644
rect 21004 36352 21044 36392
rect 20908 34252 20948 34292
rect 20812 33832 20852 33872
rect 20812 31816 20852 31856
rect 20716 31144 20756 31184
rect 20716 29464 20756 29504
rect 20716 29128 20756 29168
rect 20716 24676 20756 24716
rect 20908 28708 20948 28748
rect 20908 27448 20948 27488
rect 21100 32824 21140 32864
rect 21292 33496 21332 33536
rect 21196 30640 21236 30680
rect 21100 28540 21140 28580
rect 21100 27112 21140 27152
rect 21004 23080 21044 23120
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 19276 18544 19316 18584
rect 18796 18460 18836 18500
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 19468 19972 19508 20012
rect 19180 17788 19220 17828
rect 18700 17452 18740 17492
rect 18796 17200 18836 17240
rect 19084 17200 19124 17240
rect 19372 17452 19412 17492
rect 19276 17116 19316 17156
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 19756 19552 19796 19592
rect 19660 18628 19700 18668
rect 20236 20140 20276 20180
rect 20044 19636 20084 19676
rect 20524 19636 20564 19676
rect 19852 19216 19892 19256
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 19564 17956 19604 17996
rect 19852 17536 19892 17576
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20044 17200 20084 17240
rect 19948 17032 19988 17072
rect 20140 17116 20180 17156
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18028 15856 18068 15896
rect 17836 15352 17876 15392
rect 18604 16192 18644 16232
rect 18508 16108 18548 16148
rect 18700 16108 18740 16148
rect 18412 16024 18452 16064
rect 18892 16444 18932 16484
rect 19372 16444 19412 16484
rect 18124 15268 18164 15308
rect 18028 15100 18068 15140
rect 17740 13252 17780 13292
rect 18124 13252 18164 13292
rect 17548 12664 17588 12704
rect 17452 12496 17492 12536
rect 18124 13084 18164 13124
rect 17932 13000 17972 13040
rect 18028 12916 18068 12956
rect 17260 10396 17300 10436
rect 17164 10312 17204 10352
rect 17164 10060 17204 10100
rect 17452 10480 17492 10520
rect 17356 8800 17396 8840
rect 17068 7960 17108 8000
rect 16780 6280 16820 6320
rect 16684 5524 16724 5564
rect 16780 5356 16820 5396
rect 16588 4096 16628 4136
rect 16588 3340 16628 3380
rect 16588 3088 16628 3128
rect 16300 1072 16340 1112
rect 16492 2164 16532 2204
rect 16780 2836 16820 2876
rect 16972 4516 17012 4556
rect 16972 3340 17012 3380
rect 17164 7540 17204 7580
rect 17260 5860 17300 5900
rect 17356 5776 17396 5816
rect 17260 5524 17300 5564
rect 17164 4936 17204 4976
rect 17356 5356 17396 5396
rect 17068 2920 17108 2960
rect 16684 1912 16724 1952
rect 17164 1492 17204 1532
rect 16780 1324 16820 1364
rect 17164 1156 17204 1196
rect 16780 736 16820 776
rect 16684 148 16724 188
rect 17356 904 17396 944
rect 17932 11656 17972 11696
rect 17836 10396 17876 10436
rect 17740 9892 17780 9932
rect 18028 10312 18068 10352
rect 17932 9892 17972 9932
rect 17932 9640 17972 9680
rect 17836 9472 17876 9512
rect 18028 9136 18068 9176
rect 18316 14932 18356 14972
rect 19084 16024 19124 16064
rect 19180 15940 19220 15980
rect 18892 15520 18932 15560
rect 19372 16024 19412 16064
rect 19276 15856 19316 15896
rect 19180 15268 19220 15308
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 19180 14932 19220 14972
rect 18796 14848 18836 14888
rect 18412 14512 18452 14552
rect 18412 13672 18452 13712
rect 18316 13084 18356 13124
rect 18412 12916 18452 12956
rect 18700 14008 18740 14048
rect 18604 13924 18644 13964
rect 18316 11992 18356 12032
rect 19372 15520 19412 15560
rect 19372 14680 19412 14720
rect 19564 15604 19604 15644
rect 20044 16276 20084 16316
rect 19852 16192 19892 16232
rect 19756 16108 19796 16148
rect 20044 16024 20084 16064
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20044 15604 20084 15644
rect 19564 15268 19604 15308
rect 18988 14512 19028 14552
rect 18988 14008 19028 14048
rect 18796 13924 18836 13964
rect 18892 13840 18932 13880
rect 19276 13840 19316 13880
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 18796 12832 18836 12872
rect 18796 12580 18836 12620
rect 19276 12580 19316 12620
rect 18508 11656 18548 11696
rect 18220 10396 18260 10436
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18700 11992 18740 12032
rect 19948 15436 19988 15476
rect 20044 15352 20084 15392
rect 19660 14680 19700 14720
rect 19852 14680 19892 14720
rect 19660 14260 19700 14300
rect 19564 11908 19604 11948
rect 19468 11656 19508 11696
rect 18604 11152 18644 11192
rect 19276 10984 19316 11024
rect 18700 10564 18740 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18604 10480 18644 10520
rect 18412 10396 18452 10436
rect 18796 10396 18836 10436
rect 18316 10144 18356 10184
rect 18220 9640 18260 9680
rect 18604 10312 18644 10352
rect 18700 10228 18740 10268
rect 19372 9724 19412 9764
rect 19276 9472 19316 9512
rect 19276 9220 19316 9260
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 18508 8884 18548 8924
rect 18124 7960 18164 8000
rect 18028 7624 18068 7664
rect 17836 7120 17876 7160
rect 18412 8800 18452 8840
rect 18412 8464 18452 8504
rect 18220 6364 18260 6404
rect 18604 8800 18644 8840
rect 18700 8044 18740 8084
rect 18988 7792 19028 7832
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20044 14176 20084 14216
rect 20044 13840 20084 13880
rect 19468 8632 19508 8672
rect 19372 7708 19412 7748
rect 18508 7540 18548 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 19372 7456 19412 7496
rect 18604 7288 18644 7328
rect 18508 6532 18548 6572
rect 18508 6280 18548 6320
rect 18220 5860 18260 5900
rect 18412 5860 18452 5900
rect 17932 5776 17972 5816
rect 17644 4936 17684 4976
rect 17548 3088 17588 3128
rect 17836 5608 17876 5648
rect 18316 5776 18356 5816
rect 18508 5692 18548 5732
rect 18316 5188 18356 5228
rect 18412 5020 18452 5060
rect 18220 4684 18260 4724
rect 17932 4096 17972 4136
rect 17836 2836 17876 2876
rect 17740 2584 17780 2624
rect 18028 3004 18068 3044
rect 17548 1156 17588 1196
rect 17740 1240 17780 1280
rect 17644 1072 17684 1112
rect 17548 904 17588 944
rect 17164 400 17204 440
rect 16972 232 17012 272
rect 16972 64 17012 104
rect 17644 820 17684 860
rect 18124 1240 18164 1280
rect 18028 484 18068 524
rect 18508 3676 18548 3716
rect 18508 2836 18548 2876
rect 18316 2584 18356 2624
rect 19276 6196 19316 6236
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 18796 5608 18836 5648
rect 18700 5272 18740 5312
rect 18988 4936 19028 4976
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 19468 6616 19508 6656
rect 19468 5020 19508 5060
rect 19372 4936 19412 4976
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 20044 12496 20084 12536
rect 19852 11656 19892 11696
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 19948 10060 19988 10100
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 19948 9724 19988 9764
rect 19660 9472 19700 9512
rect 19756 8632 19796 8672
rect 19660 8128 19700 8168
rect 19948 8632 19988 8672
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 19852 7960 19892 8000
rect 19756 7120 19796 7160
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 19948 6616 19988 6656
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 19948 4852 19988 4892
rect 19660 3592 19700 3632
rect 18700 3256 18740 3296
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 19564 2584 19604 2624
rect 18412 1744 18452 1784
rect 18316 1156 18356 1196
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 18508 1324 18548 1364
rect 18700 1240 18740 1280
rect 18508 820 18548 860
rect 19084 988 19124 1028
rect 18892 652 18932 692
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 20236 3508 20276 3548
rect 19948 2584 19988 2624
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 20236 1828 20276 1868
rect 19660 1072 19700 1112
rect 19564 400 19604 440
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 19948 316 19988 356
rect 19276 232 19316 272
rect 19468 148 19508 188
<< metal3 >>
rect 0 85784 80 85804
rect 0 85744 2092 85784
rect 2132 85744 2141 85784
rect 0 85724 80 85744
rect 7267 85700 7325 85701
rect 6979 85660 6988 85700
rect 7028 85660 7276 85700
rect 7316 85660 7325 85700
rect 7267 85659 7325 85660
rect 7747 85616 7805 85617
rect 6787 85576 6796 85616
rect 6836 85576 7756 85616
rect 7796 85576 7805 85616
rect 7747 85575 7805 85576
rect 11491 85492 11500 85532
rect 11540 85492 12172 85532
rect 12212 85492 12221 85532
rect 0 85448 80 85468
rect 0 85408 6796 85448
rect 6836 85408 6845 85448
rect 13123 85408 13132 85448
rect 13172 85408 14764 85448
rect 14804 85408 14813 85448
rect 0 85388 80 85408
rect 2851 85324 2860 85364
rect 2900 85324 3340 85364
rect 3380 85324 3389 85364
rect 9283 85324 9292 85364
rect 9332 85324 14380 85364
rect 14420 85324 14429 85364
rect 931 85280 989 85281
rect 931 85240 940 85280
rect 980 85240 5836 85280
rect 5876 85240 5885 85280
rect 6115 85240 6124 85280
rect 6164 85240 7948 85280
rect 7988 85240 7997 85280
rect 11320 85240 13804 85280
rect 13844 85240 13853 85280
rect 931 85239 989 85240
rect 3043 85156 3052 85196
rect 3092 85156 7660 85196
rect 7700 85156 7709 85196
rect 0 85112 80 85132
rect 11320 85112 11360 85240
rect 12259 85156 12268 85196
rect 12308 85156 14668 85196
rect 14708 85156 14717 85196
rect 0 85072 11360 85112
rect 13123 85072 13132 85112
rect 13172 85072 19276 85112
rect 19316 85072 19325 85112
rect 0 85052 80 85072
rect 8515 85028 8573 85029
rect 2371 84988 2380 85028
rect 2420 84988 3244 85028
rect 3284 84988 3293 85028
rect 3340 84988 3916 85028
rect 3956 84988 3965 85028
rect 6211 84988 6220 85028
rect 6260 84988 8524 85028
rect 8564 84988 8573 85028
rect 3340 84944 3380 84988
rect 8515 84987 8573 84988
rect 11320 84988 13036 85028
rect 13076 84988 13085 85028
rect 18211 84988 18220 85028
rect 18260 84988 19084 85028
rect 19124 84988 19133 85028
rect 1891 84904 1900 84944
rect 1940 84904 3380 84944
rect 3427 84944 3485 84945
rect 7651 84944 7709 84945
rect 3427 84904 3436 84944
rect 3476 84904 3724 84944
rect 3764 84904 3773 84944
rect 5635 84904 5644 84944
rect 5684 84904 7660 84944
rect 7700 84904 7709 84944
rect 3427 84903 3485 84904
rect 7651 84903 7709 84904
rect 11320 84860 11360 84988
rect 12355 84944 12413 84945
rect 12355 84904 12364 84944
rect 12404 84904 19468 84944
rect 19508 84904 19517 84944
rect 12355 84903 12413 84904
rect 2500 84820 11360 84860
rect 16003 84820 16012 84860
rect 16052 84820 19564 84860
rect 19604 84820 19613 84860
rect 0 84776 80 84796
rect 2500 84776 2540 84820
rect 12835 84776 12893 84777
rect 0 84736 2540 84776
rect 3235 84736 3244 84776
rect 3284 84736 8044 84776
rect 8084 84736 8093 84776
rect 8140 84736 12364 84776
rect 12404 84736 12413 84776
rect 12835 84736 12844 84776
rect 12884 84736 13324 84776
rect 13364 84736 13373 84776
rect 15235 84736 15244 84776
rect 15284 84736 16204 84776
rect 16244 84736 16253 84776
rect 18115 84736 18124 84776
rect 18164 84736 19756 84776
rect 19796 84736 19805 84776
rect 0 84716 80 84736
rect 2947 84692 3005 84693
rect 4771 84692 4829 84693
rect 8140 84692 8180 84736
rect 12835 84735 12893 84736
rect 2947 84652 2956 84692
rect 2996 84652 3532 84692
rect 3572 84652 3581 84692
rect 3679 84652 3688 84692
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 4056 84652 4065 84692
rect 4771 84652 4780 84692
rect 4820 84652 5164 84692
rect 5204 84652 5213 84692
rect 7747 84652 7756 84692
rect 7796 84652 8180 84692
rect 11320 84652 12652 84692
rect 12692 84652 12701 84692
rect 13507 84652 13516 84692
rect 13556 84652 14668 84692
rect 14708 84652 14717 84692
rect 18403 84652 18412 84692
rect 18452 84652 18700 84692
rect 18740 84652 18749 84692
rect 18799 84652 18808 84692
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 19176 84652 19185 84692
rect 2947 84651 3005 84652
rect 4771 84651 4829 84652
rect 11320 84608 11360 84652
rect 1507 84568 1516 84608
rect 1556 84568 5068 84608
rect 5108 84568 5117 84608
rect 6787 84568 6796 84608
rect 6836 84568 11360 84608
rect 15811 84568 15820 84608
rect 15860 84568 20044 84608
rect 20084 84568 20093 84608
rect 11011 84524 11069 84525
rect 11971 84524 12029 84525
rect 2659 84484 2668 84524
rect 2708 84484 5260 84524
rect 5300 84484 5309 84524
rect 5635 84484 5644 84524
rect 5684 84484 7564 84524
rect 7604 84484 7613 84524
rect 8899 84484 8908 84524
rect 8948 84484 11020 84524
rect 11060 84484 11069 84524
rect 11886 84484 11980 84524
rect 12020 84484 12029 84524
rect 17731 84484 17740 84524
rect 17780 84484 18892 84524
rect 18932 84484 18941 84524
rect 11011 84483 11069 84484
rect 11971 84483 12029 84484
rect 0 84440 80 84460
rect 6019 84440 6077 84441
rect 6403 84440 6461 84441
rect 6595 84440 6653 84441
rect 9667 84440 9725 84441
rect 9859 84440 9917 84441
rect 11203 84440 11261 84441
rect 12739 84440 12797 84441
rect 13891 84440 13949 84441
rect 0 84400 3052 84440
rect 3092 84400 3101 84440
rect 3427 84400 3436 84440
rect 3476 84400 4300 84440
rect 4340 84400 4349 84440
rect 4579 84400 4588 84440
rect 4628 84400 4972 84440
rect 5012 84400 5021 84440
rect 5934 84400 6028 84440
rect 6068 84400 6077 84440
rect 6318 84400 6412 84440
rect 6452 84400 6461 84440
rect 6510 84400 6604 84440
rect 6644 84400 6653 84440
rect 7843 84400 7852 84440
rect 7892 84400 8524 84440
rect 8564 84400 8573 84440
rect 9582 84400 9676 84440
rect 9716 84400 9725 84440
rect 9774 84400 9868 84440
rect 9908 84400 9917 84440
rect 11118 84400 11212 84440
rect 11252 84400 11261 84440
rect 11875 84400 11884 84440
rect 11924 84400 11933 84440
rect 12654 84400 12748 84440
rect 12788 84400 12797 84440
rect 13027 84400 13036 84440
rect 13076 84400 13085 84440
rect 13420 84400 13708 84440
rect 13748 84400 13757 84440
rect 13806 84400 13900 84440
rect 13940 84400 13949 84440
rect 0 84380 80 84400
rect 6019 84399 6077 84400
rect 6403 84399 6461 84400
rect 6595 84399 6653 84400
rect 9667 84399 9725 84400
rect 9859 84399 9917 84400
rect 11203 84399 11261 84400
rect 1315 84356 1373 84357
rect 1230 84316 1324 84356
rect 1364 84316 1373 84356
rect 1699 84316 1708 84356
rect 1748 84316 2284 84356
rect 2324 84316 2333 84356
rect 2851 84316 2860 84356
rect 2900 84316 6988 84356
rect 7028 84316 7037 84356
rect 7651 84316 7660 84356
rect 7700 84316 11788 84356
rect 11828 84316 11837 84356
rect 1315 84315 1373 84316
rect 3523 84272 3581 84273
rect 3523 84232 3532 84272
rect 3572 84232 3724 84272
rect 3764 84232 3773 84272
rect 5539 84232 5548 84272
rect 5588 84232 9292 84272
rect 9332 84232 9341 84272
rect 10051 84232 10060 84272
rect 10100 84232 10732 84272
rect 10772 84232 10781 84272
rect 11320 84232 11500 84272
rect 11540 84232 11549 84272
rect 3523 84231 3581 84232
rect 11320 84188 11360 84232
rect 2500 84148 5932 84188
rect 5972 84148 5981 84188
rect 9763 84148 9772 84188
rect 9812 84148 11360 84188
rect 0 84104 80 84124
rect 2500 84104 2540 84148
rect 11884 84104 11924 84400
rect 12739 84399 12797 84400
rect 13036 84188 13076 84400
rect 13420 84356 13460 84400
rect 13891 84399 13949 84400
rect 16867 84440 16925 84441
rect 16867 84400 16876 84440
rect 16916 84400 16972 84440
rect 17012 84400 17021 84440
rect 17923 84400 17932 84440
rect 17972 84400 19276 84440
rect 19316 84400 19325 84440
rect 16867 84399 16925 84400
rect 18019 84356 18077 84357
rect 19651 84356 19709 84357
rect 13123 84316 13132 84356
rect 13172 84316 13460 84356
rect 13507 84316 13516 84356
rect 13556 84316 14476 84356
rect 14516 84316 14525 84356
rect 18019 84316 18028 84356
rect 18068 84316 19468 84356
rect 19508 84316 19517 84356
rect 19651 84316 19660 84356
rect 19700 84316 19852 84356
rect 19892 84316 19901 84356
rect 18019 84315 18077 84316
rect 19651 84315 19709 84316
rect 16579 84272 16637 84273
rect 13411 84232 13420 84272
rect 13460 84232 14092 84272
rect 14132 84232 14141 84272
rect 14956 84232 15340 84272
rect 15380 84232 15389 84272
rect 16579 84232 16588 84272
rect 16628 84232 16780 84272
rect 16820 84232 16829 84272
rect 18019 84232 18028 84272
rect 18068 84232 18508 84272
rect 18548 84232 18557 84272
rect 18691 84232 18700 84272
rect 18740 84232 19948 84272
rect 19988 84232 19997 84272
rect 13036 84148 13556 84188
rect 12451 84104 12509 84105
rect 13219 84104 13277 84105
rect 13516 84104 13556 84148
rect 0 84064 2540 84104
rect 4387 84064 4396 84104
rect 4436 84064 4876 84104
rect 4916 84064 4925 84104
rect 5059 84064 5068 84104
rect 5108 84064 6220 84104
rect 6260 84064 6269 84104
rect 8515 84064 8524 84104
rect 8564 84064 11924 84104
rect 12366 84064 12460 84104
rect 12500 84064 12509 84104
rect 12739 84064 12748 84104
rect 12788 84064 12940 84104
rect 12980 84064 12989 84104
rect 13219 84064 13228 84104
rect 13268 84064 13324 84104
rect 13364 84064 13373 84104
rect 13507 84064 13516 84104
rect 13556 84064 13565 84104
rect 13699 84064 13708 84104
rect 13748 84064 14860 84104
rect 14900 84064 14909 84104
rect 0 84044 80 84064
rect 12451 84063 12509 84064
rect 13219 84063 13277 84064
rect 14956 84020 14996 84232
rect 16579 84231 16637 84232
rect 17740 84148 19084 84188
rect 19124 84148 19133 84188
rect 17740 84105 17780 84148
rect 17731 84104 17789 84105
rect 17059 84064 17068 84104
rect 17108 84064 17740 84104
rect 17780 84064 17789 84104
rect 18307 84064 18316 84104
rect 18356 84064 19660 84104
rect 19700 84064 19709 84104
rect 17731 84063 17789 84064
rect 2083 83980 2092 84020
rect 2132 83980 14572 84020
rect 14612 83980 14996 84020
rect 15340 83980 17260 84020
rect 17300 83980 17309 84020
rect 2563 83936 2621 83937
rect 4291 83936 4349 83937
rect 15340 83936 15380 83980
rect 2563 83896 2572 83936
rect 2612 83896 2706 83936
rect 4099 83896 4108 83936
rect 4148 83896 4300 83936
rect 4340 83896 4349 83936
rect 4919 83896 4928 83936
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 5296 83896 5305 83936
rect 6691 83896 6700 83936
rect 6740 83896 7276 83936
rect 7316 83896 10636 83936
rect 10676 83896 10685 83936
rect 10915 83896 10924 83936
rect 10964 83896 15380 83936
rect 15427 83896 15436 83936
rect 15476 83896 18316 83936
rect 18356 83896 18365 83936
rect 20039 83896 20048 83936
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20416 83896 20425 83936
rect 2563 83895 2621 83896
rect 4291 83895 4349 83896
rect 1507 83812 1516 83852
rect 1556 83812 2764 83852
rect 2804 83812 2813 83852
rect 3331 83812 3340 83852
rect 3380 83812 5548 83852
rect 5588 83812 5597 83852
rect 7171 83812 7180 83852
rect 7220 83812 9140 83852
rect 15139 83812 15148 83852
rect 15188 83812 16108 83852
rect 16148 83812 16157 83852
rect 0 83768 80 83788
rect 9100 83768 9140 83812
rect 0 83728 2540 83768
rect 8323 83728 8332 83768
rect 8372 83728 9004 83768
rect 9044 83728 9053 83768
rect 9100 83728 18508 83768
rect 18548 83728 18557 83768
rect 0 83708 80 83728
rect 2500 83684 2540 83728
rect 10435 83684 10493 83685
rect 2500 83644 8236 83684
rect 8276 83644 8285 83684
rect 8611 83644 8620 83684
rect 8660 83644 9676 83684
rect 9716 83644 9868 83684
rect 9908 83644 9917 83684
rect 10435 83644 10444 83684
rect 10484 83644 10540 83684
rect 10580 83644 10589 83684
rect 12163 83644 12172 83684
rect 12212 83644 12221 83684
rect 12547 83644 12556 83684
rect 12596 83644 12605 83684
rect 13315 83644 13324 83684
rect 13364 83644 13516 83684
rect 13556 83644 13565 83684
rect 14956 83644 16972 83684
rect 17012 83644 17740 83684
rect 17780 83644 17789 83684
rect 8620 83600 8660 83644
rect 10435 83643 10493 83644
rect 4291 83560 4300 83600
rect 4340 83560 4972 83600
rect 5012 83560 5021 83600
rect 6211 83560 6220 83600
rect 6260 83560 7084 83600
rect 7124 83560 8660 83600
rect 10051 83600 10109 83601
rect 12172 83600 12212 83644
rect 12556 83600 12596 83644
rect 14956 83600 14996 83644
rect 10051 83560 10060 83600
rect 10100 83560 10156 83600
rect 10196 83560 10205 83600
rect 10339 83560 10348 83600
rect 10388 83560 10964 83600
rect 11107 83560 11116 83600
rect 11156 83560 12212 83600
rect 12259 83560 12268 83600
rect 12308 83560 12596 83600
rect 13708 83560 14956 83600
rect 14996 83560 15005 83600
rect 15235 83560 15244 83600
rect 15284 83560 16588 83600
rect 16628 83560 19796 83600
rect 10051 83559 10109 83560
rect 1507 83516 1565 83517
rect 3331 83516 3389 83517
rect 10531 83516 10589 83517
rect 10924 83516 10964 83560
rect 13708 83516 13748 83560
rect 16963 83516 17021 83517
rect 19756 83516 19796 83560
rect 1315 83476 1324 83516
rect 1364 83476 1516 83516
rect 1556 83476 1565 83516
rect 2755 83476 2764 83516
rect 2804 83476 3340 83516
rect 3380 83476 3389 83516
rect 10446 83476 10540 83516
rect 10580 83476 10828 83516
rect 10868 83476 10877 83516
rect 10924 83476 13748 83516
rect 13795 83476 13804 83516
rect 13844 83476 14284 83516
rect 14324 83476 14333 83516
rect 15043 83476 15052 83516
rect 15092 83476 15820 83516
rect 15860 83476 15869 83516
rect 16963 83476 16972 83516
rect 17012 83476 18700 83516
rect 18740 83476 18749 83516
rect 19747 83476 19756 83516
rect 19796 83476 19805 83516
rect 1507 83475 1565 83476
rect 3331 83475 3389 83476
rect 10531 83475 10589 83476
rect 16963 83475 17021 83476
rect 0 83432 80 83452
rect 8899 83432 8957 83433
rect 0 83392 7124 83432
rect 7171 83392 7180 83432
rect 7220 83392 8908 83432
rect 8948 83392 8957 83432
rect 0 83372 80 83392
rect 7084 83348 7124 83392
rect 8899 83391 8957 83392
rect 9283 83432 9341 83433
rect 9283 83392 9292 83432
rect 9332 83392 9484 83432
rect 9524 83392 9676 83432
rect 9716 83392 10636 83432
rect 10676 83392 10685 83432
rect 15907 83392 15916 83432
rect 15956 83392 19084 83432
rect 19124 83392 19133 83432
rect 9283 83391 9341 83392
rect 12355 83348 12413 83349
rect 13603 83348 13661 83349
rect 4771 83308 4780 83348
rect 4820 83308 6700 83348
rect 6740 83308 6749 83348
rect 7084 83308 7564 83348
rect 7604 83308 7613 83348
rect 8323 83308 8332 83348
rect 8372 83308 8812 83348
rect 8852 83308 8861 83348
rect 12270 83308 12364 83348
rect 12404 83308 12413 83348
rect 13518 83308 13612 83348
rect 13652 83308 13661 83348
rect 12355 83307 12413 83308
rect 13603 83307 13661 83308
rect 14947 83348 15005 83349
rect 16003 83348 16061 83349
rect 14947 83308 14956 83348
rect 14996 83308 15628 83348
rect 15668 83308 15677 83348
rect 15918 83308 16012 83348
rect 16052 83308 16061 83348
rect 16291 83308 16300 83348
rect 16340 83308 18124 83348
rect 18164 83308 18173 83348
rect 14947 83307 15005 83308
rect 16003 83307 16061 83308
rect 6307 83264 6365 83265
rect 2947 83224 2956 83264
rect 2996 83224 4244 83264
rect 5347 83224 5356 83264
rect 5396 83224 5548 83264
rect 5588 83224 5597 83264
rect 6307 83224 6316 83264
rect 6356 83224 10924 83264
rect 10964 83224 10973 83264
rect 13315 83224 13324 83264
rect 13364 83224 16492 83264
rect 16532 83224 16541 83264
rect 17251 83224 17260 83264
rect 17300 83224 17876 83264
rect 4204 83180 4244 83224
rect 6307 83223 6365 83224
rect 13987 83180 14045 83181
rect 17443 83180 17501 83181
rect 2500 83140 3092 83180
rect 3679 83140 3688 83180
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 4056 83140 4065 83180
rect 4195 83140 4204 83180
rect 4244 83140 4684 83180
rect 4724 83140 4733 83180
rect 4867 83140 4876 83180
rect 4916 83140 6356 83180
rect 6403 83140 6412 83180
rect 6452 83140 7948 83180
rect 7988 83140 7997 83180
rect 8227 83140 8236 83180
rect 8276 83140 8620 83180
rect 8660 83140 8669 83180
rect 10531 83140 10540 83180
rect 10580 83140 11020 83180
rect 11060 83140 11069 83180
rect 12739 83140 12748 83180
rect 12788 83140 13996 83180
rect 14036 83140 14045 83180
rect 16003 83140 16012 83180
rect 16052 83140 16780 83180
rect 16820 83140 16829 83180
rect 17347 83140 17356 83180
rect 17396 83140 17452 83180
rect 17492 83140 17501 83180
rect 0 83096 80 83116
rect 2500 83096 2540 83140
rect 0 83056 2540 83096
rect 0 83036 80 83056
rect 2380 82972 2996 83012
rect 0 82760 80 82780
rect 2380 82760 2420 82972
rect 0 82720 2420 82760
rect 2476 82888 2764 82928
rect 2804 82888 2813 82928
rect 0 82700 80 82720
rect 2476 82592 2516 82888
rect 2956 82676 2996 82972
rect 3052 82928 3092 83140
rect 3331 83096 3389 83097
rect 6316 83096 6356 83140
rect 13987 83139 14045 83140
rect 17443 83139 17501 83140
rect 3331 83056 3340 83096
rect 3380 83056 5588 83096
rect 6316 83056 8428 83096
rect 8468 83056 8477 83096
rect 8707 83056 8716 83096
rect 8756 83056 10924 83096
rect 10964 83056 10973 83096
rect 11320 83056 13996 83096
rect 14036 83056 14045 83096
rect 14371 83056 14380 83096
rect 14420 83056 14764 83096
rect 14804 83056 14813 83096
rect 3331 83055 3389 83056
rect 5548 83012 5588 83056
rect 6307 83012 6365 83013
rect 10435 83012 10493 83013
rect 3139 82972 3148 83012
rect 3188 82972 3532 83012
rect 3572 82972 3581 83012
rect 4003 82972 4012 83012
rect 4052 82972 5452 83012
rect 5492 82972 5501 83012
rect 5548 82972 6316 83012
rect 6356 82972 6365 83012
rect 6883 82972 6892 83012
rect 6932 82972 10444 83012
rect 10484 82972 10493 83012
rect 6307 82971 6365 82972
rect 5347 82928 5405 82929
rect 6892 82928 6932 82972
rect 10435 82971 10493 82972
rect 11320 82928 11360 83056
rect 13795 83012 13853 83013
rect 17836 83012 17876 83224
rect 18220 83224 20121 83264
rect 20161 83224 20170 83264
rect 18220 83180 18260 83224
rect 18403 83180 18461 83181
rect 18211 83140 18220 83180
rect 18260 83140 18269 83180
rect 18318 83140 18412 83180
rect 18452 83140 18461 83180
rect 18691 83140 18700 83180
rect 18740 83140 18749 83180
rect 18799 83140 18808 83180
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 19176 83140 19185 83180
rect 18403 83139 18461 83140
rect 18700 83096 18740 83140
rect 18115 83056 18124 83096
rect 18164 83056 18740 83096
rect 11587 82972 11596 83012
rect 11636 82972 11788 83012
rect 11828 82972 11837 83012
rect 13507 82972 13516 83012
rect 13556 82972 13804 83012
rect 13844 82972 15820 83012
rect 15860 82972 15869 83012
rect 17836 82972 18508 83012
rect 18548 82972 18557 83012
rect 19075 82972 19084 83012
rect 19124 82972 19372 83012
rect 19412 82972 19421 83012
rect 13795 82971 13853 82972
rect 12643 82928 12701 82929
rect 3052 82888 4876 82928
rect 4916 82888 4925 82928
rect 5155 82888 5164 82928
rect 5204 82888 5356 82928
rect 5396 82888 6932 82928
rect 9196 82888 11360 82928
rect 12558 82888 12652 82928
rect 12692 82888 12701 82928
rect 5347 82887 5405 82888
rect 5443 82844 5501 82845
rect 7459 82844 7517 82845
rect 9196 82844 9236 82888
rect 12643 82887 12701 82888
rect 3043 82804 3052 82844
rect 3092 82804 5204 82844
rect 5358 82804 5452 82844
rect 5492 82804 5501 82844
rect 6211 82804 6220 82844
rect 6260 82804 7468 82844
rect 7508 82804 7517 82844
rect 8419 82804 8428 82844
rect 8468 82804 9196 82844
rect 9236 82804 9245 82844
rect 9763 82804 9772 82844
rect 9812 82804 17492 82844
rect 5164 82760 5204 82804
rect 5443 82803 5501 82804
rect 7459 82803 7517 82804
rect 5731 82760 5789 82761
rect 7363 82760 7421 82761
rect 14371 82760 14429 82761
rect 17452 82760 17492 82804
rect 4579 82720 4588 82760
rect 4628 82720 4972 82760
rect 5012 82720 5021 82760
rect 5164 82720 5740 82760
rect 5780 82720 6796 82760
rect 6836 82720 6845 82760
rect 7267 82720 7276 82760
rect 7316 82720 7372 82760
rect 7412 82720 7421 82760
rect 7747 82720 7756 82760
rect 7796 82720 11404 82760
rect 11444 82720 11453 82760
rect 12067 82720 12076 82760
rect 12116 82720 12364 82760
rect 12404 82720 12413 82760
rect 14286 82720 14380 82760
rect 14420 82720 14429 82760
rect 14947 82720 14956 82760
rect 14996 82720 15532 82760
rect 15572 82720 15581 82760
rect 17443 82720 17452 82760
rect 17492 82720 17501 82760
rect 17731 82720 17740 82760
rect 17780 82720 18700 82760
rect 18740 82720 18749 82760
rect 5731 82719 5789 82720
rect 7363 82719 7421 82720
rect 14371 82719 14429 82720
rect 2956 82636 8372 82676
rect 10147 82636 10156 82676
rect 10196 82636 12652 82676
rect 12692 82636 12701 82676
rect 18883 82636 18892 82676
rect 18932 82636 19756 82676
rect 19796 82636 19805 82676
rect 8332 82592 8372 82636
rect 12163 82592 12221 82593
rect 12931 82592 12989 82593
rect 748 82552 2516 82592
rect 2659 82552 2668 82592
rect 2708 82552 3244 82592
rect 3284 82552 3293 82592
rect 8323 82552 8332 82592
rect 8372 82552 8381 82592
rect 9475 82552 9484 82592
rect 9524 82552 9868 82592
rect 9908 82552 11596 82592
rect 11636 82552 11645 82592
rect 12078 82552 12172 82592
rect 12212 82552 12221 82592
rect 12846 82552 12940 82592
rect 12980 82552 12989 82592
rect 0 82424 80 82444
rect 748 82424 788 82552
rect 12163 82551 12221 82552
rect 12931 82551 12989 82552
rect 13123 82592 13181 82593
rect 14755 82592 14813 82593
rect 19555 82592 19613 82593
rect 13123 82552 13132 82592
rect 13172 82552 13420 82592
rect 13460 82552 13469 82592
rect 14563 82552 14572 82592
rect 14612 82552 14764 82592
rect 14804 82552 14813 82592
rect 19363 82552 19372 82592
rect 19412 82552 19564 82592
rect 19604 82552 19613 82592
rect 13123 82551 13181 82552
rect 14755 82551 14813 82552
rect 19555 82551 19613 82552
rect 0 82384 788 82424
rect 844 82468 7372 82508
rect 7412 82468 7421 82508
rect 7651 82468 7660 82508
rect 7700 82468 9772 82508
rect 9812 82468 9821 82508
rect 11875 82468 11884 82508
rect 11924 82468 15628 82508
rect 15668 82468 16108 82508
rect 16148 82468 19468 82508
rect 19508 82468 19517 82508
rect 0 82364 80 82384
rect 0 82088 80 82108
rect 844 82088 884 82468
rect 2755 82424 2813 82425
rect 11587 82424 11645 82425
rect 2670 82384 2764 82424
rect 2804 82384 2813 82424
rect 4919 82384 4928 82424
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 5296 82384 5305 82424
rect 6787 82384 6796 82424
rect 6836 82384 7084 82424
rect 7124 82384 7133 82424
rect 10147 82384 10156 82424
rect 10196 82384 11308 82424
rect 11348 82384 11357 82424
rect 11491 82384 11500 82424
rect 11540 82384 11596 82424
rect 11636 82384 11645 82424
rect 2755 82383 2813 82384
rect 11587 82383 11645 82384
rect 11875 82424 11933 82425
rect 11875 82384 11884 82424
rect 11924 82384 16780 82424
rect 16820 82384 16829 82424
rect 20039 82384 20048 82424
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20416 82384 20425 82424
rect 11875 82383 11933 82384
rect 11971 82340 12029 82341
rect 19555 82340 19613 82341
rect 2851 82300 2860 82340
rect 2900 82300 3244 82340
rect 3284 82300 3293 82340
rect 5731 82300 5740 82340
rect 5780 82300 11980 82340
rect 12020 82300 12029 82340
rect 16195 82300 16204 82340
rect 16244 82300 19564 82340
rect 19604 82300 19613 82340
rect 11971 82299 12029 82300
rect 19555 82299 19613 82300
rect 1315 82256 1373 82257
rect 1230 82216 1324 82256
rect 1364 82216 1373 82256
rect 2563 82216 2572 82256
rect 2612 82216 8908 82256
rect 8948 82216 8957 82256
rect 10627 82216 10636 82256
rect 10676 82216 10828 82256
rect 10868 82216 10877 82256
rect 11011 82216 11020 82256
rect 11060 82216 12460 82256
rect 12500 82216 12509 82256
rect 12643 82216 12652 82256
rect 12692 82216 12701 82256
rect 1315 82215 1373 82216
rect 4099 82172 4157 82173
rect 4771 82172 4829 82173
rect 5347 82172 5405 82173
rect 2851 82132 2860 82172
rect 2900 82132 4108 82172
rect 4148 82132 4157 82172
rect 4675 82132 4684 82172
rect 4724 82132 4780 82172
rect 4820 82132 4829 82172
rect 5155 82132 5164 82172
rect 5204 82132 5356 82172
rect 5396 82132 5405 82172
rect 4099 82131 4157 82132
rect 4771 82131 4829 82132
rect 5347 82131 5405 82132
rect 5827 82172 5885 82173
rect 6499 82172 6557 82173
rect 11779 82172 11837 82173
rect 5827 82132 5836 82172
rect 5876 82132 5932 82172
rect 5972 82132 5981 82172
rect 6499 82132 6508 82172
rect 6548 82132 6604 82172
rect 6644 82132 6653 82172
rect 7363 82132 7372 82172
rect 7412 82132 11788 82172
rect 11828 82132 11837 82172
rect 5827 82131 5885 82132
rect 6499 82131 6557 82132
rect 11779 82131 11837 82132
rect 0 82048 884 82088
rect 1027 82088 1085 82089
rect 10339 82088 10397 82089
rect 12652 82088 12692 82216
rect 1027 82048 1036 82088
rect 1076 82048 2540 82088
rect 0 82028 80 82048
rect 1027 82047 1085 82048
rect 2500 82004 2540 82048
rect 4204 82048 7084 82088
rect 7124 82048 7133 82088
rect 8323 82048 8332 82088
rect 8372 82048 10252 82088
rect 10292 82048 10348 82088
rect 10388 82048 10397 82088
rect 11971 82048 11980 82088
rect 12020 82048 12364 82088
rect 12404 82048 12413 82088
rect 12456 82048 12465 82088
rect 12505 82048 12692 82088
rect 16108 82048 16204 82088
rect 16244 82048 16253 82088
rect 3811 82004 3869 82005
rect 4204 82004 4244 82048
rect 10339 82047 10397 82048
rect 2500 81964 3436 82004
rect 3476 81964 3485 82004
rect 3726 81964 3820 82004
rect 3860 81964 3869 82004
rect 4195 81964 4204 82004
rect 4244 81964 4253 82004
rect 4483 81964 4492 82004
rect 4532 81964 5396 82004
rect 6691 81964 6700 82004
rect 6740 81964 8812 82004
rect 8852 81964 9964 82004
rect 10004 81964 10444 82004
rect 10484 81964 10493 82004
rect 10819 81964 10828 82004
rect 10868 81964 11212 82004
rect 11252 81964 11261 82004
rect 14371 81964 14380 82004
rect 14420 81964 14764 82004
rect 14804 81964 15052 82004
rect 15092 81964 15101 82004
rect 3811 81963 3869 81964
rect 1795 81920 1853 81921
rect 4771 81920 4829 81921
rect 5356 81920 5396 81964
rect 12643 81920 12701 81921
rect 14371 81920 14429 81921
rect 1710 81880 1804 81920
rect 1844 81880 1853 81920
rect 4686 81880 4780 81920
rect 4820 81880 4829 81920
rect 5316 81880 5356 81920
rect 5396 81880 5405 81920
rect 12558 81880 12652 81920
rect 12692 81880 12701 81920
rect 14275 81880 14284 81920
rect 14324 81880 14380 81920
rect 14420 81880 14956 81920
rect 14996 81880 15005 81920
rect 1795 81879 1853 81880
rect 4771 81879 4829 81880
rect 12643 81879 12701 81880
rect 14371 81879 14429 81880
rect 11971 81836 12029 81837
rect 16108 81836 16148 82048
rect 17932 81964 18220 82004
rect 18260 81964 18269 82004
rect 17932 81920 17972 81964
rect 19267 81920 19325 81921
rect 17892 81880 17932 81920
rect 17972 81880 17981 81920
rect 19182 81880 19276 81920
rect 19316 81880 19325 81920
rect 19267 81879 19325 81880
rect 8995 81796 9004 81836
rect 9044 81796 9772 81836
rect 9812 81796 9821 81836
rect 11779 81796 11788 81836
rect 11828 81796 11980 81836
rect 12020 81796 16148 81836
rect 16387 81836 16445 81837
rect 16387 81796 16396 81836
rect 16436 81796 16492 81836
rect 16532 81796 16541 81836
rect 18787 81796 18796 81836
rect 18836 81796 18845 81836
rect 19651 81796 19660 81836
rect 19700 81796 20044 81836
rect 20084 81796 20093 81836
rect 11971 81795 12029 81796
rect 16387 81795 16445 81796
rect 0 81752 80 81772
rect 3523 81752 3581 81753
rect 11587 81752 11645 81753
rect 14755 81752 14813 81753
rect 0 81712 3532 81752
rect 3572 81712 3581 81752
rect 4483 81712 4492 81752
rect 4532 81712 11596 81752
rect 11636 81712 11645 81752
rect 14563 81712 14572 81752
rect 14612 81712 14764 81752
rect 14804 81712 14813 81752
rect 18796 81752 18836 81796
rect 18796 81712 19276 81752
rect 19316 81712 19325 81752
rect 0 81692 80 81712
rect 3523 81711 3581 81712
rect 11587 81711 11645 81712
rect 14755 81711 14813 81712
rect 3679 81628 3688 81668
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 4056 81628 4065 81668
rect 4204 81628 10732 81668
rect 10772 81628 10781 81668
rect 15043 81628 15052 81668
rect 15092 81628 15244 81668
rect 15284 81628 15293 81668
rect 18799 81628 18808 81668
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 19176 81628 19185 81668
rect 1603 81500 1661 81501
rect 4204 81500 4244 81628
rect 8995 81544 9004 81584
rect 9044 81544 9484 81584
rect 9524 81544 9533 81584
rect 1507 81460 1516 81500
rect 1556 81460 1612 81500
rect 1652 81460 1661 81500
rect 2083 81460 2092 81500
rect 2132 81460 2764 81500
rect 2804 81460 2813 81500
rect 3043 81460 3052 81500
rect 3092 81460 4012 81500
rect 4052 81460 4244 81500
rect 4291 81460 4300 81500
rect 4340 81460 5164 81500
rect 5204 81460 11116 81500
rect 11156 81460 11165 81500
rect 11491 81460 11500 81500
rect 11540 81460 11692 81500
rect 11732 81460 11741 81500
rect 16579 81460 16588 81500
rect 16628 81460 19564 81500
rect 19604 81460 19613 81500
rect 1603 81459 1661 81460
rect 0 81416 80 81436
rect 0 81376 4204 81416
rect 4244 81376 4253 81416
rect 9283 81376 9292 81416
rect 9332 81376 9964 81416
rect 10004 81376 10013 81416
rect 12163 81376 12172 81416
rect 12212 81376 12364 81416
rect 12404 81376 12413 81416
rect 18595 81376 18604 81416
rect 18644 81376 20524 81416
rect 20564 81376 20573 81416
rect 0 81356 80 81376
rect 7843 81332 7901 81333
rect 2500 81292 5492 81332
rect 5539 81292 5548 81332
rect 5588 81292 7852 81332
rect 7892 81292 7901 81332
rect 0 81080 80 81100
rect 2500 81080 2540 81292
rect 3523 81248 3581 81249
rect 3907 81248 3965 81249
rect 2851 81208 2860 81248
rect 2900 81208 3148 81248
rect 3188 81208 3197 81248
rect 3438 81208 3532 81248
rect 3572 81208 3581 81248
rect 3822 81208 3916 81248
rect 3956 81208 3965 81248
rect 5452 81248 5492 81292
rect 7843 81291 7901 81292
rect 7948 81292 10348 81332
rect 10388 81292 10397 81332
rect 11491 81292 11500 81332
rect 11540 81292 12556 81332
rect 12596 81292 12605 81332
rect 7948 81248 7988 81292
rect 18691 81248 18749 81249
rect 5452 81208 5740 81248
rect 5780 81208 5789 81248
rect 7363 81208 7372 81248
rect 7412 81208 7948 81248
rect 7988 81208 7997 81248
rect 9763 81208 9772 81248
rect 9812 81208 11404 81248
rect 11444 81208 11788 81248
rect 11828 81208 11837 81248
rect 12163 81208 12172 81248
rect 12212 81208 12221 81248
rect 13891 81208 13900 81248
rect 13940 81208 15052 81248
rect 15092 81208 15101 81248
rect 18691 81208 18700 81248
rect 18740 81208 18796 81248
rect 18836 81208 18845 81248
rect 3523 81207 3581 81208
rect 3907 81207 3965 81208
rect 3619 81164 3677 81165
rect 10339 81164 10397 81165
rect 12172 81164 12212 81208
rect 18691 81207 18749 81208
rect 3619 81124 3628 81164
rect 3668 81124 9428 81164
rect 3619 81123 3677 81124
rect 9388 81080 9428 81124
rect 10339 81124 10348 81164
rect 10388 81124 12212 81164
rect 10339 81123 10397 81124
rect 16387 81080 16445 81081
rect 0 81040 2540 81080
rect 3139 81040 3148 81080
rect 3188 81040 3340 81080
rect 3380 81040 3389 81080
rect 5443 81040 5452 81080
rect 5492 81040 9292 81080
rect 9332 81040 9341 81080
rect 9388 81040 11500 81080
rect 11540 81040 11549 81080
rect 11683 81040 11692 81080
rect 11732 81040 12748 81080
rect 12788 81040 12797 81080
rect 15427 81040 15436 81080
rect 15476 81040 16108 81080
rect 16148 81040 16396 81080
rect 16436 81040 16445 81080
rect 18211 81040 18220 81080
rect 18260 81040 18604 81080
rect 18644 81040 18653 81080
rect 0 81020 80 81040
rect 16387 81039 16445 81040
rect 16003 80996 16061 80997
rect 4195 80956 4204 80996
rect 4244 80956 7604 80996
rect 7651 80956 7660 80996
rect 7700 80956 8236 80996
rect 8276 80956 8285 80996
rect 16003 80956 16012 80996
rect 16052 80956 18508 80996
rect 18548 80956 18557 80996
rect 7564 80912 7604 80956
rect 16003 80955 16061 80956
rect 17059 80912 17117 80913
rect 3427 80872 3436 80912
rect 3476 80872 4108 80912
rect 4148 80872 4157 80912
rect 4204 80872 4780 80912
rect 4820 80872 4829 80912
rect 4919 80872 4928 80912
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 5296 80872 5305 80912
rect 7564 80872 10636 80912
rect 10676 80872 10685 80912
rect 13411 80872 13420 80912
rect 13460 80872 13900 80912
rect 13940 80872 13949 80912
rect 16963 80872 16972 80912
rect 17012 80872 17068 80912
rect 17108 80872 17117 80912
rect 20039 80872 20048 80912
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20416 80872 20425 80912
rect 1315 80828 1373 80829
rect 1891 80828 1949 80829
rect 4204 80828 4244 80872
rect 1315 80788 1324 80828
rect 1364 80788 1900 80828
rect 1940 80788 1949 80828
rect 2371 80788 2380 80828
rect 2420 80788 3724 80828
rect 3764 80788 4244 80828
rect 4483 80788 4492 80828
rect 4532 80788 10060 80828
rect 10100 80788 10109 80828
rect 11299 80788 11308 80828
rect 11348 80788 11357 80828
rect 1315 80787 1373 80788
rect 1891 80787 1949 80788
rect 0 80744 80 80764
rect 0 80704 4588 80744
rect 4628 80704 4637 80744
rect 4771 80704 4780 80744
rect 4820 80704 6892 80744
rect 6932 80704 6941 80744
rect 7555 80704 7564 80744
rect 7604 80704 7852 80744
rect 7892 80704 7901 80744
rect 7948 80704 9580 80744
rect 9620 80704 9629 80744
rect 0 80684 80 80704
rect 7948 80660 7988 80704
rect 1324 80620 5644 80660
rect 5684 80620 5693 80660
rect 5740 80620 7988 80660
rect 8323 80620 8332 80660
rect 8372 80620 8620 80660
rect 8660 80620 8669 80660
rect 1324 80576 1364 80620
rect 5740 80576 5780 80620
rect 1315 80536 1324 80576
rect 1364 80536 1373 80576
rect 4963 80536 4972 80576
rect 5012 80536 5780 80576
rect 6211 80536 6220 80576
rect 6260 80536 7660 80576
rect 7700 80536 7709 80576
rect 4771 80492 4829 80493
rect 6979 80492 7037 80493
rect 7459 80492 7517 80493
rect 8035 80492 8093 80493
rect 11308 80492 11348 80788
rect 11491 80620 11500 80660
rect 11540 80620 12268 80660
rect 12308 80620 12317 80660
rect 13420 80576 13460 80872
rect 17059 80871 17117 80872
rect 14851 80704 14860 80744
rect 14900 80704 15628 80744
rect 15668 80704 15677 80744
rect 14851 80660 14909 80661
rect 13507 80620 13516 80660
rect 13556 80620 13804 80660
rect 13844 80620 13853 80660
rect 14851 80620 14860 80660
rect 14900 80620 16300 80660
rect 16340 80620 16349 80660
rect 17251 80620 17260 80660
rect 17300 80620 18028 80660
rect 18068 80620 18892 80660
rect 18932 80620 19948 80660
rect 19988 80620 19997 80660
rect 14851 80619 14909 80620
rect 17923 80576 17981 80577
rect 13315 80536 13324 80576
rect 13364 80536 13460 80576
rect 15619 80536 15628 80576
rect 15668 80536 15820 80576
rect 15860 80536 15869 80576
rect 17923 80536 17932 80576
rect 17972 80536 18124 80576
rect 18164 80536 18173 80576
rect 17923 80535 17981 80536
rect 14275 80492 14333 80493
rect 1228 80452 3052 80492
rect 3092 80452 3532 80492
rect 3572 80452 3581 80492
rect 4771 80452 4780 80492
rect 4820 80452 4876 80492
rect 4916 80452 5740 80492
rect 5780 80452 5789 80492
rect 6894 80452 6988 80492
rect 7028 80452 7037 80492
rect 7171 80452 7180 80492
rect 7220 80452 7468 80492
rect 7508 80452 7564 80492
rect 7604 80452 7613 80492
rect 7939 80452 7948 80492
rect 7988 80452 8044 80492
rect 8084 80452 8093 80492
rect 11203 80452 11212 80492
rect 11252 80452 11348 80492
rect 14190 80452 14284 80492
rect 14324 80452 14333 80492
rect 16867 80452 16876 80492
rect 16916 80452 20620 80492
rect 20660 80452 20669 80492
rect 0 80408 80 80428
rect 1228 80408 1268 80452
rect 4771 80451 4829 80452
rect 6979 80451 7037 80452
rect 7459 80451 7517 80452
rect 8035 80451 8093 80452
rect 14275 80451 14333 80452
rect 3139 80408 3197 80409
rect 18595 80408 18653 80409
rect 0 80368 1268 80408
rect 2275 80368 2284 80408
rect 2324 80368 3148 80408
rect 3188 80368 3197 80408
rect 4387 80368 4396 80408
rect 4436 80368 10540 80408
rect 10580 80368 10589 80408
rect 10819 80368 10828 80408
rect 10868 80368 11308 80408
rect 11348 80368 11357 80408
rect 11491 80368 11500 80408
rect 11540 80368 14228 80408
rect 0 80348 80 80368
rect 3139 80367 3197 80368
rect 14188 80324 14228 80368
rect 15532 80368 17740 80408
rect 17780 80368 17789 80408
rect 17923 80368 17932 80408
rect 17972 80368 18508 80408
rect 18548 80368 18604 80408
rect 18644 80368 18653 80408
rect 15532 80324 15572 80368
rect 18595 80367 18653 80368
rect 19939 80408 19997 80409
rect 19939 80368 19948 80408
rect 19988 80368 20140 80408
rect 20180 80368 20189 80408
rect 19939 80367 19997 80368
rect 15811 80324 15869 80325
rect 1420 80284 1612 80324
rect 1652 80284 4780 80324
rect 4820 80284 4829 80324
rect 7267 80284 7276 80324
rect 7316 80284 7468 80324
rect 7508 80284 7517 80324
rect 9859 80284 9868 80324
rect 9908 80284 12404 80324
rect 14188 80284 15532 80324
rect 15572 80284 15581 80324
rect 15726 80284 15820 80324
rect 15860 80284 15869 80324
rect 16387 80284 16396 80324
rect 16436 80284 19852 80324
rect 19892 80284 19901 80324
rect 0 80072 80 80092
rect 1420 80072 1460 80284
rect 2851 80200 2860 80240
rect 2900 80200 4492 80240
rect 4532 80200 4541 80240
rect 5155 80200 5164 80240
rect 5204 80200 5644 80240
rect 5684 80200 10732 80240
rect 10772 80200 10781 80240
rect 11203 80200 11212 80240
rect 11252 80200 12268 80240
rect 12308 80200 12317 80240
rect 7651 80156 7709 80157
rect 11395 80156 11453 80157
rect 1987 80116 1996 80156
rect 2036 80116 2284 80156
rect 2324 80116 2333 80156
rect 3679 80116 3688 80156
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 4056 80116 4065 80156
rect 7651 80116 7660 80156
rect 7700 80116 11404 80156
rect 11444 80116 11453 80156
rect 12364 80156 12404 80284
rect 15811 80283 15869 80284
rect 12451 80200 12460 80240
rect 12500 80200 14764 80240
rect 14804 80200 16300 80240
rect 16340 80200 16349 80240
rect 12364 80116 15916 80156
rect 15956 80116 15965 80156
rect 18799 80116 18808 80156
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 19176 80116 19185 80156
rect 7651 80115 7709 80116
rect 11395 80115 11453 80116
rect 4483 80072 4541 80073
rect 5539 80072 5597 80073
rect 18499 80072 18557 80073
rect 0 80032 1460 80072
rect 3331 80032 3340 80072
rect 3380 80032 4492 80072
rect 4532 80032 4541 80072
rect 5347 80032 5356 80072
rect 5396 80032 5548 80072
rect 5588 80032 5597 80072
rect 5827 80032 5836 80072
rect 5876 80032 9484 80072
rect 9524 80032 9533 80072
rect 11500 80032 16300 80072
rect 16340 80032 18508 80072
rect 18548 80032 18557 80072
rect 0 80012 80 80032
rect 4483 80031 4541 80032
rect 5539 80031 5597 80032
rect 1027 79948 1036 79988
rect 1076 79948 1900 79988
rect 1940 79948 6932 79988
rect 9763 79948 9772 79988
rect 9812 79948 9964 79988
rect 10004 79948 11404 79988
rect 11444 79948 11453 79988
rect 1411 79904 1469 79905
rect 6892 79904 6932 79948
rect 11500 79904 11540 80032
rect 18499 80031 18557 80032
rect 19267 79988 19325 79989
rect 12259 79948 12268 79988
rect 12308 79948 16396 79988
rect 16436 79948 16445 79988
rect 16675 79948 16684 79988
rect 16724 79948 16876 79988
rect 16916 79948 16925 79988
rect 17731 79948 17740 79988
rect 17780 79948 18124 79988
rect 18164 79948 18173 79988
rect 19171 79948 19180 79988
rect 19220 79948 19276 79988
rect 19316 79948 19325 79988
rect 19267 79947 19325 79948
rect 1411 79864 1420 79904
rect 1460 79864 1516 79904
rect 1556 79864 1565 79904
rect 1795 79864 1804 79904
rect 1844 79864 2092 79904
rect 2132 79864 2141 79904
rect 4579 79864 4588 79904
rect 4628 79864 5740 79904
rect 5780 79864 5789 79904
rect 6892 79864 11540 79904
rect 11683 79864 11692 79904
rect 11732 79864 12364 79904
rect 12404 79864 12413 79904
rect 16483 79864 16492 79904
rect 16532 79864 17932 79904
rect 17972 79864 19756 79904
rect 19796 79864 19805 79904
rect 1411 79863 1469 79864
rect 5827 79820 5885 79821
rect 8035 79820 8093 79821
rect 17155 79820 17213 79821
rect 1411 79780 1420 79820
rect 1460 79780 5548 79820
rect 5588 79780 5597 79820
rect 5827 79780 5836 79820
rect 5876 79780 5932 79820
rect 5972 79780 5981 79820
rect 7459 79780 7468 79820
rect 7508 79780 8044 79820
rect 8084 79780 8093 79820
rect 5827 79779 5885 79780
rect 8035 79779 8093 79780
rect 11212 79780 12268 79820
rect 12308 79780 13324 79820
rect 13364 79780 13373 79820
rect 14947 79780 14956 79820
rect 14996 79780 17068 79820
rect 17108 79780 17164 79820
rect 17204 79780 17213 79820
rect 17635 79780 17644 79820
rect 17684 79780 19468 79820
rect 19508 79780 19948 79820
rect 19988 79780 19997 79820
rect 0 79736 80 79756
rect 1315 79736 1373 79737
rect 1987 79736 2045 79737
rect 4675 79736 4733 79737
rect 6787 79736 6845 79737
rect 8611 79736 8669 79737
rect 0 79696 1324 79736
rect 1364 79696 1373 79736
rect 1603 79696 1612 79736
rect 1652 79696 1661 79736
rect 1987 79696 1996 79736
rect 2036 79696 2092 79736
rect 2132 79696 2141 79736
rect 2563 79696 2572 79736
rect 2612 79696 4012 79736
rect 4052 79696 4061 79736
rect 4675 79696 4684 79736
rect 4724 79696 6796 79736
rect 6836 79696 6845 79736
rect 0 79676 80 79696
rect 1315 79695 1373 79696
rect 1612 79652 1652 79696
rect 1987 79695 2045 79696
rect 4675 79695 4733 79696
rect 6787 79695 6845 79696
rect 7852 79696 8236 79736
rect 8276 79696 8285 79736
rect 8592 79696 8620 79736
rect 8660 79696 8716 79736
rect 8756 79696 11116 79736
rect 11156 79696 11165 79736
rect 7852 79652 7892 79696
rect 8611 79695 8669 79696
rect 11212 79652 11252 79780
rect 14956 79736 14996 79780
rect 17155 79779 17213 79780
rect 18499 79736 18557 79737
rect 11395 79696 11404 79736
rect 11444 79696 14996 79736
rect 15523 79696 15532 79736
rect 15572 79696 17780 79736
rect 17059 79652 17117 79653
rect 17740 79652 17780 79696
rect 18499 79696 18508 79736
rect 18548 79696 18988 79736
rect 19028 79696 19037 79736
rect 18499 79695 18557 79696
rect 18211 79652 18269 79653
rect 1507 79612 1516 79652
rect 1556 79612 1565 79652
rect 1612 79612 5356 79652
rect 5396 79612 5405 79652
rect 5731 79612 5740 79652
rect 5780 79612 7852 79652
rect 7892 79612 7901 79652
rect 8131 79612 8140 79652
rect 8180 79612 8189 79652
rect 8803 79612 8812 79652
rect 8852 79612 9100 79652
rect 9140 79612 10060 79652
rect 10100 79612 10732 79652
rect 10772 79612 11252 79652
rect 15139 79612 15148 79652
rect 15188 79612 15820 79652
rect 15860 79612 15869 79652
rect 16291 79612 16300 79652
rect 16340 79612 16684 79652
rect 16724 79612 16733 79652
rect 16974 79612 17068 79652
rect 17108 79612 17117 79652
rect 17731 79612 17740 79652
rect 17780 79612 17789 79652
rect 18115 79612 18124 79652
rect 18164 79612 18220 79652
rect 18260 79612 18412 79652
rect 18452 79612 18461 79652
rect 643 79568 701 79569
rect 1516 79568 1556 79612
rect 2755 79568 2813 79569
rect 6115 79568 6173 79569
rect 8140 79568 8180 79612
rect 17059 79611 17117 79612
rect 18211 79611 18269 79612
rect 643 79528 652 79568
rect 692 79528 1420 79568
rect 1460 79528 1469 79568
rect 1516 79528 1900 79568
rect 1940 79528 2764 79568
rect 2804 79528 2813 79568
rect 3043 79528 3052 79568
rect 3092 79528 3532 79568
rect 3572 79528 3581 79568
rect 4963 79528 4972 79568
rect 5012 79528 5021 79568
rect 5443 79528 5452 79568
rect 5492 79528 6124 79568
rect 6164 79528 6173 79568
rect 7555 79528 7564 79568
rect 7604 79528 8044 79568
rect 8084 79528 8093 79568
rect 8140 79528 17548 79568
rect 17588 79528 17597 79568
rect 643 79527 701 79528
rect 2755 79527 2813 79528
rect 1123 79484 1181 79485
rect 4972 79484 5012 79528
rect 6115 79527 6173 79528
rect 8227 79484 8285 79485
rect 1123 79444 1132 79484
rect 1172 79444 5012 79484
rect 6115 79444 6124 79484
rect 6164 79444 8236 79484
rect 8276 79444 8285 79484
rect 14371 79444 14380 79484
rect 14420 79444 15820 79484
rect 15860 79444 15869 79484
rect 16675 79444 16684 79484
rect 16724 79444 16876 79484
rect 16916 79444 16925 79484
rect 17548 79444 19468 79484
rect 19508 79444 19517 79484
rect 1123 79443 1181 79444
rect 8227 79443 8285 79444
rect 0 79400 80 79420
rect 2947 79400 3005 79401
rect 6883 79400 6941 79401
rect 10435 79400 10493 79401
rect 10627 79400 10685 79401
rect 11971 79400 12029 79401
rect 17548 79400 17588 79444
rect 0 79360 748 79400
rect 788 79360 797 79400
rect 2862 79360 2956 79400
rect 2996 79360 3005 79400
rect 4919 79360 4928 79400
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 5296 79360 5305 79400
rect 6798 79360 6892 79400
rect 6932 79360 6941 79400
rect 7555 79360 7564 79400
rect 7604 79360 7756 79400
rect 7796 79360 7805 79400
rect 7939 79360 7948 79400
rect 7988 79360 8812 79400
rect 8852 79360 8861 79400
rect 10350 79360 10444 79400
rect 10484 79360 10493 79400
rect 10542 79360 10636 79400
rect 10676 79360 10685 79400
rect 11886 79360 11980 79400
rect 12020 79360 12029 79400
rect 13891 79360 13900 79400
rect 13940 79360 13949 79400
rect 15907 79360 15916 79400
rect 15956 79360 17588 79400
rect 17635 79400 17693 79401
rect 19555 79400 19613 79401
rect 17635 79360 17644 79400
rect 17684 79360 18796 79400
rect 18836 79360 18845 79400
rect 19470 79360 19564 79400
rect 19604 79360 19613 79400
rect 20039 79360 20048 79400
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20416 79360 20425 79400
rect 0 79340 80 79360
rect 2947 79359 3005 79360
rect 6883 79359 6941 79360
rect 10435 79359 10493 79360
rect 10627 79359 10685 79360
rect 11971 79359 12029 79360
rect 2275 79316 2333 79317
rect 12547 79316 12605 79317
rect 2275 79276 2284 79316
rect 2324 79276 4724 79316
rect 4771 79276 4780 79316
rect 4820 79276 11360 79316
rect 12163 79276 12172 79316
rect 12212 79276 12556 79316
rect 12596 79276 12605 79316
rect 13900 79316 13940 79360
rect 13900 79276 14476 79316
rect 14516 79276 15436 79316
rect 15476 79276 15485 79316
rect 2275 79275 2333 79276
rect 1315 79148 1373 79149
rect 4684 79148 4724 79276
rect 4972 79232 5012 79276
rect 7171 79232 7229 79233
rect 7939 79232 7997 79233
rect 11320 79232 11360 79276
rect 12547 79275 12605 79276
rect 16492 79232 16532 79360
rect 17635 79359 17693 79360
rect 19555 79359 19613 79360
rect 17356 79276 17441 79316
rect 17481 79276 17490 79316
rect 17539 79276 17548 79316
rect 17588 79276 19180 79316
rect 19220 79276 19229 79316
rect 17356 79233 17396 79276
rect 17347 79232 17405 79233
rect 4963 79192 4972 79232
rect 5012 79192 5021 79232
rect 6220 79192 6700 79232
rect 6740 79192 6988 79232
rect 7028 79192 7037 79232
rect 7171 79192 7180 79232
rect 7220 79192 7314 79232
rect 7939 79192 7948 79232
rect 7988 79192 8428 79232
rect 8468 79192 8477 79232
rect 10252 79192 10636 79232
rect 10676 79192 10685 79232
rect 11320 79192 12076 79232
rect 12116 79192 12125 79232
rect 15244 79192 15628 79232
rect 15668 79192 15677 79232
rect 16483 79192 16492 79232
rect 16532 79192 16541 79232
rect 17347 79192 17356 79232
rect 17396 79192 17405 79232
rect 17923 79192 17932 79232
rect 17972 79192 19948 79232
rect 19988 79192 19997 79232
rect 1315 79108 1324 79148
rect 1364 79108 4148 79148
rect 4684 79108 5644 79148
rect 5684 79108 5693 79148
rect 1315 79107 1373 79108
rect 0 79064 80 79084
rect 1603 79064 1661 79065
rect 0 79024 212 79064
rect 1219 79024 1228 79064
rect 1268 79024 1612 79064
rect 1652 79024 1661 79064
rect 0 79004 80 79024
rect 172 78896 212 79024
rect 1603 79023 1661 79024
rect 2467 78980 2525 78981
rect 4108 78980 4148 79108
rect 6220 79064 6260 79192
rect 7171 79191 7229 79192
rect 7939 79191 7997 79192
rect 10252 79148 10292 79192
rect 15244 79148 15284 79192
rect 17347 79191 17405 79192
rect 18307 79148 18365 79149
rect 6316 79108 8840 79148
rect 10243 79108 10252 79148
rect 10292 79108 10301 79148
rect 11404 79108 15284 79148
rect 15331 79108 15340 79148
rect 15380 79108 18068 79148
rect 4483 79024 4492 79064
rect 4532 79024 6220 79064
rect 6260 79024 6269 79064
rect 6316 78980 6356 79108
rect 8800 79064 8840 79108
rect 11404 79064 11444 79108
rect 18028 79064 18068 79108
rect 18307 79108 18316 79148
rect 18356 79108 18508 79148
rect 18548 79108 18557 79148
rect 18307 79107 18365 79108
rect 6499 79024 6508 79064
rect 6548 79024 6892 79064
rect 6932 79024 6941 79064
rect 7939 79024 7948 79064
rect 7988 79024 8620 79064
rect 8660 79024 8669 79064
rect 8800 79024 11444 79064
rect 11491 79024 11500 79064
rect 11540 79024 12556 79064
rect 12596 79024 12605 79064
rect 13795 79024 13804 79064
rect 13844 79024 14380 79064
rect 14420 79024 14429 79064
rect 15523 79024 15532 79064
rect 15572 79024 15916 79064
rect 15956 79024 15965 79064
rect 16195 79024 16204 79064
rect 16244 79024 17836 79064
rect 17876 79024 17885 79064
rect 18019 79024 18028 79064
rect 18068 79024 18077 79064
rect 19363 79024 19372 79064
rect 19412 79024 19948 79064
rect 19988 79024 19997 79064
rect 2467 78940 2476 78980
rect 2516 78940 2860 78980
rect 2900 78940 2909 78980
rect 4108 78940 5068 78980
rect 5108 78940 6356 78980
rect 7171 78980 7229 78981
rect 19267 78980 19325 78981
rect 7171 78940 7180 78980
rect 7220 78940 8428 78980
rect 8468 78940 8477 78980
rect 14083 78940 14092 78980
rect 14132 78940 14668 78980
rect 14708 78940 14717 78980
rect 18211 78940 18220 78980
rect 18260 78940 18508 78980
rect 18548 78940 18557 78980
rect 18883 78940 18892 78980
rect 18932 78940 19276 78980
rect 19316 78940 19325 78980
rect 2467 78939 2525 78940
rect 7171 78939 7229 78940
rect 19267 78939 19325 78940
rect 3331 78896 3389 78897
rect 172 78856 3340 78896
rect 3380 78856 3389 78896
rect 3331 78855 3389 78856
rect 7075 78896 7133 78897
rect 8227 78896 8285 78897
rect 17251 78896 17309 78897
rect 7075 78856 7084 78896
rect 7124 78856 7372 78896
rect 7412 78856 7421 78896
rect 8142 78856 8236 78896
rect 8276 78856 8285 78896
rect 10339 78856 10348 78896
rect 10388 78856 17260 78896
rect 17300 78856 18988 78896
rect 19028 78856 19276 78896
rect 19316 78856 19325 78896
rect 7075 78855 7133 78856
rect 8227 78855 8285 78856
rect 17251 78855 17309 78856
rect 3811 78772 3820 78812
rect 3860 78772 4492 78812
rect 4532 78772 4541 78812
rect 7843 78772 7852 78812
rect 7892 78772 12364 78812
rect 12404 78772 12413 78812
rect 14179 78772 14188 78812
rect 14228 78772 14860 78812
rect 14900 78772 14909 78812
rect 17155 78772 17164 78812
rect 17204 78772 17356 78812
rect 17396 78772 17405 78812
rect 0 78728 80 78748
rect 17059 78728 17117 78729
rect 0 78688 1132 78728
rect 1172 78688 1181 78728
rect 3523 78688 3532 78728
rect 3572 78688 4148 78728
rect 5635 78688 5644 78728
rect 5684 78688 9004 78728
rect 9044 78688 9053 78728
rect 9955 78688 9964 78728
rect 10004 78688 10252 78728
rect 10292 78688 10301 78728
rect 10828 78688 13900 78728
rect 13940 78688 16012 78728
rect 16052 78688 16061 78728
rect 16974 78688 17068 78728
rect 17108 78688 17117 78728
rect 0 78668 80 78688
rect 4108 78644 4148 78688
rect 10828 78644 10868 78688
rect 17059 78687 17117 78688
rect 3679 78604 3688 78644
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 4056 78604 4065 78644
rect 4108 78604 6028 78644
rect 6068 78604 10868 78644
rect 12067 78604 12076 78644
rect 12116 78604 14284 78644
rect 14324 78604 14333 78644
rect 15619 78604 15628 78644
rect 15668 78604 18124 78644
rect 18164 78604 18173 78644
rect 18799 78604 18808 78644
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 19176 78604 19185 78644
rect 3235 78560 3293 78561
rect 13027 78560 13085 78561
rect 14275 78560 14333 78561
rect 3150 78520 3244 78560
rect 3284 78520 5260 78560
rect 5300 78520 10868 78560
rect 3235 78519 3293 78520
rect 10828 78476 10868 78520
rect 13027 78520 13036 78560
rect 13076 78520 13420 78560
rect 13460 78520 14284 78560
rect 14324 78520 15820 78560
rect 15860 78520 15869 78560
rect 16387 78520 16396 78560
rect 16436 78520 17068 78560
rect 17108 78520 17117 78560
rect 18595 78520 18604 78560
rect 18644 78520 18932 78560
rect 13027 78519 13085 78520
rect 14275 78519 14333 78520
rect 18307 78476 18365 78477
rect 1891 78436 1900 78476
rect 1940 78436 4876 78476
rect 4916 78436 4925 78476
rect 8140 78436 10348 78476
rect 10388 78436 10397 78476
rect 10828 78436 16532 78476
rect 16579 78436 16588 78476
rect 16628 78436 17644 78476
rect 17684 78436 17693 78476
rect 18307 78436 18316 78476
rect 18356 78436 18508 78476
rect 18548 78436 18557 78476
rect 0 78392 80 78412
rect 1219 78392 1277 78393
rect 8140 78392 8180 78436
rect 10819 78392 10877 78393
rect 16492 78392 16532 78436
rect 18307 78435 18365 78436
rect 18691 78392 18749 78393
rect 0 78352 1172 78392
rect 0 78332 80 78352
rect 1132 78308 1172 78352
rect 1219 78352 1228 78392
rect 1268 78352 3532 78392
rect 3572 78352 8180 78392
rect 8227 78352 8236 78392
rect 8276 78352 8428 78392
rect 8468 78352 8477 78392
rect 10734 78352 10828 78392
rect 10868 78352 10877 78392
rect 13795 78352 13804 78392
rect 13844 78352 14956 78392
rect 14996 78352 16396 78392
rect 16436 78352 16445 78392
rect 16492 78352 18604 78392
rect 18644 78352 18700 78392
rect 18740 78352 18768 78392
rect 1219 78351 1277 78352
rect 10819 78351 10877 78352
rect 18691 78351 18749 78352
rect 2275 78308 2333 78309
rect 11779 78308 11837 78309
rect 18019 78308 18077 78309
rect 18892 78308 18932 78520
rect 1132 78268 2284 78308
rect 2324 78268 2333 78308
rect 6979 78268 6988 78308
rect 7028 78268 9100 78308
rect 9140 78268 9149 78308
rect 11779 78268 11788 78308
rect 11828 78268 13228 78308
rect 13268 78268 13277 78308
rect 15235 78268 15244 78308
rect 15284 78268 16244 78308
rect 17934 78268 18028 78308
rect 18068 78268 18077 78308
rect 18403 78268 18412 78308
rect 18452 78268 18932 78308
rect 2275 78267 2333 78268
rect 11779 78267 11837 78268
rect 8419 78224 8477 78225
rect 15715 78224 15773 78225
rect 2467 78184 2476 78224
rect 2516 78184 3092 78224
rect 3139 78184 3148 78224
rect 3188 78184 3436 78224
rect 3476 78184 4972 78224
rect 5012 78184 5021 78224
rect 5635 78184 5644 78224
rect 5684 78184 6028 78224
rect 6068 78184 6077 78224
rect 6691 78184 6700 78224
rect 6740 78184 6892 78224
rect 6932 78184 6941 78224
rect 7651 78184 7660 78224
rect 7700 78184 7709 78224
rect 8419 78184 8428 78224
rect 8468 78184 8812 78224
rect 8852 78184 8861 78224
rect 9283 78184 9292 78224
rect 9332 78184 10540 78224
rect 10580 78184 10589 78224
rect 10915 78184 10924 78224
rect 10964 78184 12076 78224
rect 12116 78184 12125 78224
rect 13315 78184 13324 78224
rect 13364 78184 13996 78224
rect 14036 78184 14045 78224
rect 14947 78184 14956 78224
rect 14996 78184 15340 78224
rect 15380 78184 15389 78224
rect 15715 78184 15724 78224
rect 15764 78184 15916 78224
rect 15956 78184 15965 78224
rect 3052 78140 3092 78184
rect 4675 78140 4733 78141
rect 7660 78140 7700 78184
rect 8419 78183 8477 78184
rect 15715 78183 15773 78184
rect 15523 78140 15581 78141
rect 1411 78100 1420 78140
rect 1460 78100 2668 78140
rect 2708 78100 2717 78140
rect 3052 78100 3476 78140
rect 4590 78100 4684 78140
rect 4724 78100 4733 78140
rect 5059 78100 5068 78140
rect 5108 78100 5548 78140
rect 5588 78100 5597 78140
rect 6499 78100 6508 78140
rect 6548 78100 7372 78140
rect 7412 78100 7421 78140
rect 7660 78100 12172 78140
rect 12212 78100 12221 78140
rect 12355 78100 12364 78140
rect 12404 78100 13900 78140
rect 13940 78100 14188 78140
rect 14228 78100 14237 78140
rect 15427 78100 15436 78140
rect 15476 78100 15532 78140
rect 15572 78100 15581 78140
rect 16204 78140 16244 78268
rect 18019 78267 18077 78268
rect 17251 78184 17260 78224
rect 17300 78184 17548 78224
rect 17588 78184 17597 78224
rect 16204 78100 16916 78140
rect 16963 78100 16972 78140
rect 17012 78100 17932 78140
rect 17972 78100 17981 78140
rect 18115 78100 18124 78140
rect 18164 78100 18508 78140
rect 18548 78100 18557 78140
rect 0 78056 80 78076
rect 1987 78056 2045 78057
rect 0 78016 1996 78056
rect 2036 78016 2045 78056
rect 0 77996 80 78016
rect 1987 78015 2045 78016
rect 3436 77972 3476 78100
rect 4675 78099 4733 78100
rect 15523 78099 15581 78100
rect 16876 78056 16916 78100
rect 10915 78016 10924 78056
rect 10964 78016 11308 78056
rect 11348 78016 11357 78056
rect 16876 78016 17260 78056
rect 17300 78016 17309 78056
rect 19756 78016 20140 78056
rect 20180 78016 20189 78056
rect 10435 77972 10493 77973
rect 3427 77932 3436 77972
rect 3476 77932 3485 77972
rect 10435 77932 10444 77972
rect 10484 77932 13172 77972
rect 10435 77931 10493 77932
rect 9571 77888 9629 77889
rect 13132 77888 13172 77932
rect 19756 77888 19796 78016
rect 4919 77848 4928 77888
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 5296 77848 5305 77888
rect 9571 77848 9580 77888
rect 9620 77848 13036 77888
rect 13076 77848 13085 77888
rect 13132 77848 18220 77888
rect 18260 77848 18508 77888
rect 18548 77848 18557 77888
rect 19747 77848 19756 77888
rect 19796 77848 19805 77888
rect 20039 77848 20048 77888
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20416 77848 20425 77888
rect 9571 77847 9629 77848
rect 1987 77804 2045 77805
rect 1987 77764 1996 77804
rect 2036 77764 9004 77804
rect 9044 77764 9580 77804
rect 9620 77764 9629 77804
rect 1987 77763 2045 77764
rect 0 77720 80 77740
rect 1891 77720 1949 77721
rect 17347 77720 17405 77721
rect 18211 77720 18269 77721
rect 0 77680 1900 77720
rect 1940 77680 2956 77720
rect 2996 77680 3724 77720
rect 3764 77680 3773 77720
rect 14659 77680 14668 77720
rect 14708 77680 15916 77720
rect 15956 77680 16300 77720
rect 16340 77680 16349 77720
rect 17262 77680 17356 77720
rect 17396 77680 17405 77720
rect 18126 77680 18220 77720
rect 18260 77680 18269 77720
rect 0 77660 80 77680
rect 1891 77679 1949 77680
rect 17347 77679 17405 77680
rect 18211 77679 18269 77680
rect 13315 77636 13373 77637
rect 7075 77596 7084 77636
rect 7124 77596 7660 77636
rect 7700 77596 8524 77636
rect 8564 77596 8573 77636
rect 11320 77596 12364 77636
rect 12404 77596 13324 77636
rect 13364 77596 13373 77636
rect 1315 77552 1373 77553
rect 11320 77552 11360 77596
rect 13315 77595 13373 77596
rect 17059 77552 17117 77553
rect 1219 77512 1228 77552
rect 1268 77512 1324 77552
rect 1364 77512 1373 77552
rect 2467 77512 2476 77552
rect 2516 77512 2860 77552
rect 2900 77512 4204 77552
rect 4244 77512 4253 77552
rect 4867 77512 4876 77552
rect 4916 77512 5740 77552
rect 5780 77512 5789 77552
rect 6115 77512 6124 77552
rect 6164 77512 6508 77552
rect 6548 77512 6557 77552
rect 7171 77512 7180 77552
rect 7220 77512 11360 77552
rect 16387 77512 16396 77552
rect 16436 77512 16780 77552
rect 16820 77512 17068 77552
rect 17108 77512 17740 77552
rect 17780 77512 17789 77552
rect 1315 77511 1373 77512
rect 17059 77511 17117 77512
rect 3523 77468 3581 77469
rect 4195 77468 4253 77469
rect 10627 77468 10685 77469
rect 17155 77468 17213 77469
rect 3523 77428 3532 77468
rect 3572 77428 4204 77468
rect 4244 77428 5164 77468
rect 5204 77428 5213 77468
rect 7267 77428 7276 77468
rect 7316 77428 8140 77468
rect 8180 77428 8189 77468
rect 10542 77428 10636 77468
rect 10676 77428 10685 77468
rect 17070 77428 17164 77468
rect 17204 77428 17213 77468
rect 18595 77428 18604 77468
rect 18644 77428 18653 77468
rect 3523 77427 3581 77428
rect 4195 77427 4253 77428
rect 10627 77427 10685 77428
rect 17155 77427 17213 77428
rect 0 77384 80 77404
rect 1603 77384 1661 77385
rect 2371 77384 2429 77385
rect 18307 77384 18365 77385
rect 0 77344 1612 77384
rect 1652 77344 2380 77384
rect 2420 77344 2429 77384
rect 6787 77344 6796 77384
rect 6836 77344 8044 77384
rect 8084 77344 8093 77384
rect 18222 77344 18316 77384
rect 18356 77344 18365 77384
rect 0 77324 80 77344
rect 1603 77343 1661 77344
rect 2371 77343 2429 77344
rect 18307 77343 18365 77344
rect 15043 77300 15101 77301
rect 2659 77260 2668 77300
rect 2708 77260 2956 77300
rect 2996 77260 3005 77300
rect 3715 77260 3724 77300
rect 3764 77260 12268 77300
rect 12308 77260 12317 77300
rect 14958 77260 15052 77300
rect 15092 77260 15101 77300
rect 15043 77259 15101 77260
rect 2083 77216 2141 77217
rect 1795 77176 1804 77216
rect 1844 77176 2092 77216
rect 2132 77176 2141 77216
rect 3331 77176 3340 77216
rect 3380 77176 4588 77216
rect 4628 77176 4637 77216
rect 10339 77176 10348 77216
rect 10388 77176 10828 77216
rect 10868 77176 10877 77216
rect 2083 77175 2141 77176
rect 2851 77132 2909 77133
rect 3235 77132 3293 77133
rect 10819 77132 10877 77133
rect 18604 77132 18644 77428
rect 19555 77260 19564 77300
rect 19604 77260 20044 77300
rect 20084 77260 20093 77300
rect 556 77092 2860 77132
rect 2900 77092 3244 77132
rect 3284 77092 3293 77132
rect 3679 77092 3688 77132
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 4056 77092 4065 77132
rect 10819 77092 10828 77132
rect 10868 77092 11116 77132
rect 11156 77092 11165 77132
rect 18307 77092 18316 77132
rect 18356 77092 18644 77132
rect 18799 77092 18808 77132
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 19176 77092 19185 77132
rect 20035 77092 20044 77132
rect 20084 77092 20716 77132
rect 20756 77092 20765 77132
rect 0 77048 80 77068
rect 556 77048 596 77092
rect 2851 77091 2909 77092
rect 3235 77091 3293 77092
rect 10819 77091 10877 77092
rect 0 77008 596 77048
rect 3523 77048 3581 77049
rect 3523 77008 3532 77048
rect 3572 77008 4780 77048
rect 4820 77008 4829 77048
rect 9379 77008 9388 77048
rect 9428 77008 14668 77048
rect 14708 77008 14717 77048
rect 0 76988 80 77008
rect 3523 77007 3581 77008
rect 4099 76964 4157 76965
rect 17923 76964 17981 76965
rect 4099 76924 4108 76964
rect 4148 76924 4396 76964
rect 4436 76924 4445 76964
rect 12259 76924 12268 76964
rect 12308 76924 17932 76964
rect 17972 76924 17981 76964
rect 4099 76923 4157 76924
rect 17923 76923 17981 76924
rect 3427 76880 3485 76881
rect 8227 76880 8285 76881
rect 10435 76880 10493 76881
rect 17443 76880 17501 76881
rect 19267 76880 19325 76881
rect 1516 76840 2188 76880
rect 2228 76840 2237 76880
rect 2500 76840 3244 76880
rect 3284 76840 3293 76880
rect 3427 76840 3436 76880
rect 3476 76840 4588 76880
rect 4628 76840 4637 76880
rect 8227 76840 8236 76880
rect 8276 76840 10444 76880
rect 10484 76840 10493 76880
rect 10819 76840 10828 76880
rect 10868 76840 11308 76880
rect 11348 76840 11357 76880
rect 15235 76840 15244 76880
rect 15284 76840 15916 76880
rect 15956 76840 15965 76880
rect 17443 76840 17452 76880
rect 17492 76840 17932 76880
rect 17972 76840 17981 76880
rect 18499 76840 18508 76880
rect 18548 76840 18700 76880
rect 18740 76840 18749 76880
rect 18883 76840 18892 76880
rect 18932 76840 19276 76880
rect 19316 76840 19412 76880
rect 1516 76796 1556 76840
rect 2500 76796 2540 76840
rect 3427 76839 3485 76840
rect 8227 76839 8285 76840
rect 10435 76839 10493 76840
rect 17443 76839 17501 76840
rect 19267 76839 19325 76840
rect 5347 76796 5405 76797
rect 19372 76796 19412 76840
rect 1507 76756 1516 76796
rect 1556 76756 1565 76796
rect 1699 76756 1708 76796
rect 1748 76756 2540 76796
rect 3052 76756 3148 76796
rect 3188 76756 3197 76796
rect 4771 76756 4780 76796
rect 4820 76756 5356 76796
rect 5396 76756 5405 76796
rect 6307 76756 6316 76796
rect 6356 76756 10540 76796
rect 10580 76756 11360 76796
rect 14755 76756 14764 76796
rect 14804 76756 18124 76796
rect 18164 76756 18173 76796
rect 19363 76756 19372 76796
rect 19412 76756 19421 76796
rect 0 76712 80 76732
rect 1411 76712 1469 76713
rect 0 76672 1420 76712
rect 1460 76672 1469 76712
rect 0 76652 80 76672
rect 1411 76671 1469 76672
rect 2179 76712 2237 76713
rect 3052 76712 3092 76756
rect 5347 76755 5405 76756
rect 3235 76712 3293 76713
rect 10147 76712 10205 76713
rect 2179 76672 2188 76712
rect 2228 76672 3092 76712
rect 3150 76672 3244 76712
rect 3284 76672 3293 76712
rect 3715 76672 3724 76712
rect 3764 76672 4108 76712
rect 4148 76672 4157 76712
rect 7075 76672 7084 76712
rect 7124 76672 9196 76712
rect 9236 76672 9245 76712
rect 10062 76672 10156 76712
rect 10196 76672 10205 76712
rect 11320 76712 11360 76756
rect 11320 76672 11692 76712
rect 11732 76672 12364 76712
rect 12404 76672 12413 76712
rect 13411 76672 13420 76712
rect 13460 76672 14476 76712
rect 14516 76672 14668 76712
rect 14708 76672 18028 76712
rect 18068 76672 18077 76712
rect 2179 76671 2237 76672
rect 3235 76671 3293 76672
rect 10147 76671 10205 76672
rect 2083 76628 2141 76629
rect 2083 76588 2092 76628
rect 2132 76588 2188 76628
rect 2228 76588 2237 76628
rect 2371 76588 2380 76628
rect 2420 76588 2764 76628
rect 2804 76588 3052 76628
rect 3092 76588 3101 76628
rect 6211 76588 6220 76628
rect 6260 76588 8524 76628
rect 8564 76588 13324 76628
rect 13364 76588 13373 76628
rect 2083 76587 2141 76588
rect 2563 76544 2621 76545
rect 8323 76544 8381 76545
rect 16291 76544 16349 76545
rect 1891 76504 1900 76544
rect 1940 76504 2572 76544
rect 2612 76504 2621 76544
rect 4579 76504 4588 76544
rect 4628 76504 8332 76544
rect 8372 76504 8381 76544
rect 8899 76504 8908 76544
rect 8948 76504 14380 76544
rect 14420 76504 14429 76544
rect 16291 76504 16300 76544
rect 16340 76504 20140 76544
rect 20180 76504 20189 76544
rect 2563 76503 2621 76504
rect 8323 76503 8381 76504
rect 16291 76503 16349 76504
rect 2371 76460 2429 76461
rect 2371 76420 2380 76460
rect 2420 76420 13516 76460
rect 13556 76420 13565 76460
rect 2371 76419 2429 76420
rect 0 76376 80 76396
rect 2563 76376 2621 76377
rect 4771 76376 4829 76377
rect 8419 76376 8477 76377
rect 10156 76376 10196 76420
rect 0 76336 1612 76376
rect 1652 76336 1661 76376
rect 2563 76336 2572 76376
rect 2612 76336 4780 76376
rect 4820 76336 4829 76376
rect 4919 76336 4928 76376
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 5296 76336 5305 76376
rect 8334 76336 8428 76376
rect 8468 76336 8477 76376
rect 10147 76336 10156 76376
rect 10196 76336 10205 76376
rect 12163 76336 12172 76376
rect 12212 76336 12364 76376
rect 12404 76336 12413 76376
rect 20039 76336 20048 76376
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20416 76336 20425 76376
rect 0 76316 80 76336
rect 2563 76335 2621 76336
rect 4771 76335 4829 76336
rect 8419 76335 8477 76336
rect 18019 76292 18077 76293
rect 19651 76292 19709 76293
rect 4387 76252 4396 76292
rect 4436 76252 7468 76292
rect 7508 76252 7517 76292
rect 8323 76252 8332 76292
rect 8372 76252 15436 76292
rect 15476 76252 15485 76292
rect 18019 76252 18028 76292
rect 18068 76252 19660 76292
rect 19700 76252 19709 76292
rect 18019 76251 18077 76252
rect 19651 76251 19709 76252
rect 1795 76208 1853 76209
rect 6691 76208 6749 76209
rect 18403 76208 18461 76209
rect 1411 76168 1420 76208
rect 1460 76168 1804 76208
rect 1844 76168 1853 76208
rect 6606 76168 6700 76208
rect 6740 76168 6749 76208
rect 6883 76168 6892 76208
rect 6932 76168 7372 76208
rect 7412 76168 7421 76208
rect 7939 76168 7948 76208
rect 7988 76168 7997 76208
rect 18403 76168 18412 76208
rect 18452 76168 20044 76208
rect 20084 76168 20093 76208
rect 1795 76167 1853 76168
rect 6691 76167 6749 76168
rect 1411 76124 1469 76125
rect 7948 76124 7988 76168
rect 18403 76167 18461 76168
rect 1411 76084 1420 76124
rect 1460 76084 4972 76124
rect 5012 76084 5021 76124
rect 6787 76084 6796 76124
rect 6836 76084 7852 76124
rect 7892 76084 7901 76124
rect 7948 76084 9004 76124
rect 9044 76084 9676 76124
rect 9716 76084 9725 76124
rect 15427 76084 15436 76124
rect 15476 76084 15916 76124
rect 15956 76084 16108 76124
rect 16148 76084 16157 76124
rect 1411 76083 1469 76084
rect 0 76040 80 76060
rect 1804 76041 1844 76084
rect 1315 76040 1373 76041
rect 0 76000 1324 76040
rect 1364 76000 1373 76040
rect 0 75980 80 76000
rect 1315 75999 1373 76000
rect 1795 76040 1853 76041
rect 15523 76040 15581 76041
rect 1795 76000 1804 76040
rect 1844 76000 1884 76040
rect 4099 76000 4108 76040
rect 4148 76000 4876 76040
rect 4916 76000 4925 76040
rect 6220 76000 6644 76040
rect 7171 76000 7180 76040
rect 7220 76000 8044 76040
rect 8084 76000 8093 76040
rect 13411 76000 13420 76040
rect 13460 76000 13469 76040
rect 15523 76000 15532 76040
rect 15572 76000 15628 76040
rect 15668 76000 15677 76040
rect 17443 76000 17452 76040
rect 17492 76000 17836 76040
rect 17876 76000 18028 76040
rect 18068 76000 19852 76040
rect 19892 76000 19901 76040
rect 1795 75999 1853 76000
rect 6220 75956 6260 76000
rect 6604 75956 6644 76000
rect 13420 75956 13460 76000
rect 15523 75999 15581 76000
rect 1219 75916 1228 75956
rect 1268 75916 6260 75956
rect 6403 75916 6412 75956
rect 6452 75916 6461 75956
rect 6604 75916 10060 75956
rect 10100 75916 10109 75956
rect 11299 75916 11308 75956
rect 11348 75916 13460 75956
rect 13507 75916 13516 75956
rect 13556 75916 15052 75956
rect 15092 75916 15101 75956
rect 6412 75872 6452 75916
rect 4963 75832 4972 75872
rect 5012 75832 6356 75872
rect 6412 75832 7084 75872
rect 7124 75832 7948 75872
rect 7988 75832 7997 75872
rect 16675 75832 16684 75872
rect 16724 75832 16972 75872
rect 17012 75832 17021 75872
rect 1603 75748 1612 75788
rect 1652 75748 4588 75788
rect 4628 75748 4637 75788
rect 0 75704 80 75724
rect 6316 75704 6356 75832
rect 19939 75788 19997 75789
rect 11320 75748 19276 75788
rect 19316 75748 19948 75788
rect 19988 75748 19997 75788
rect 11320 75704 11360 75748
rect 19939 75747 19997 75748
rect 0 75664 6260 75704
rect 6316 75664 9868 75704
rect 9908 75664 11360 75704
rect 12643 75664 12652 75704
rect 12692 75664 13460 75704
rect 13891 75664 13900 75704
rect 13940 75664 14380 75704
rect 14420 75664 14429 75704
rect 18211 75664 18220 75704
rect 18260 75664 19660 75704
rect 19700 75664 19709 75704
rect 0 75644 80 75664
rect 163 75580 172 75620
rect 212 75580 2380 75620
rect 2420 75580 2429 75620
rect 3679 75580 3688 75620
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 4056 75580 4065 75620
rect 1891 75536 1949 75537
rect 1795 75496 1804 75536
rect 1844 75496 1900 75536
rect 1940 75496 1949 75536
rect 6220 75536 6260 75664
rect 13420 75621 13460 75664
rect 13411 75620 13469 75621
rect 6307 75580 6316 75620
rect 6356 75580 6604 75620
rect 6644 75580 6653 75620
rect 6787 75580 6796 75620
rect 6836 75580 11404 75620
rect 11444 75580 11980 75620
rect 12020 75580 12029 75620
rect 12163 75580 12172 75620
rect 12212 75580 12844 75620
rect 12884 75580 12893 75620
rect 13411 75580 13420 75620
rect 13460 75580 13996 75620
rect 14036 75580 14045 75620
rect 17347 75580 17356 75620
rect 17396 75580 17644 75620
rect 17684 75580 17693 75620
rect 18799 75580 18808 75620
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 19176 75580 19185 75620
rect 13411 75579 13469 75580
rect 7555 75536 7613 75537
rect 6220 75496 7564 75536
rect 7604 75496 9772 75536
rect 9812 75496 15340 75536
rect 15380 75496 15389 75536
rect 1891 75495 1949 75496
rect 7555 75495 7613 75496
rect 4291 75452 4349 75453
rect 1603 75412 1612 75452
rect 1652 75412 4300 75452
rect 4340 75412 4349 75452
rect 5923 75412 5932 75452
rect 5972 75412 8468 75452
rect 11203 75412 11212 75452
rect 11252 75412 11404 75452
rect 11444 75412 11453 75452
rect 11971 75412 11980 75452
rect 12020 75412 16876 75452
rect 16916 75412 16925 75452
rect 4291 75411 4349 75412
rect 0 75368 80 75388
rect 8428 75368 8468 75412
rect 0 75328 2476 75368
rect 2516 75328 8140 75368
rect 8180 75328 8332 75368
rect 8372 75328 8381 75368
rect 8428 75328 13516 75368
rect 13556 75328 13565 75368
rect 17251 75328 17260 75368
rect 17300 75328 18220 75368
rect 18260 75328 18269 75368
rect 0 75308 80 75328
rect 1411 75284 1469 75285
rect 1326 75244 1420 75284
rect 1460 75244 1469 75284
rect 1411 75243 1469 75244
rect 3331 75284 3389 75285
rect 17251 75284 17309 75285
rect 3331 75244 3340 75284
rect 3380 75244 4108 75284
rect 4148 75244 4588 75284
rect 4628 75244 4637 75284
rect 4867 75244 4876 75284
rect 4916 75244 6220 75284
rect 6260 75244 6269 75284
rect 11299 75244 11308 75284
rect 11348 75244 11788 75284
rect 11828 75244 11980 75284
rect 12020 75244 12029 75284
rect 13027 75244 13036 75284
rect 13076 75244 13612 75284
rect 13652 75244 13661 75284
rect 17155 75244 17164 75284
rect 17204 75244 17260 75284
rect 17300 75244 17309 75284
rect 3331 75243 3389 75244
rect 17251 75243 17309 75244
rect 2755 75200 2813 75201
rect 12547 75200 12605 75201
rect 15715 75200 15773 75201
rect 2670 75160 2764 75200
rect 2804 75160 2813 75200
rect 3235 75160 3244 75200
rect 3284 75160 3628 75200
rect 3668 75160 3677 75200
rect 4483 75160 4492 75200
rect 4532 75160 6508 75200
rect 6548 75160 6557 75200
rect 9379 75160 9388 75200
rect 9428 75160 11020 75200
rect 11060 75160 11069 75200
rect 12462 75160 12556 75200
rect 12596 75160 12605 75200
rect 15331 75160 15340 75200
rect 15380 75160 15724 75200
rect 15764 75160 15773 75200
rect 15907 75160 15916 75200
rect 15956 75160 16588 75200
rect 16628 75160 17740 75200
rect 17780 75160 17789 75200
rect 2755 75159 2813 75160
rect 12547 75159 12605 75160
rect 15715 75159 15773 75160
rect 3715 75076 3724 75116
rect 3764 75076 5452 75116
rect 5492 75076 7084 75116
rect 7124 75076 13804 75116
rect 13844 75076 13853 75116
rect 0 75032 80 75052
rect 1219 75032 1277 75033
rect 4099 75032 4157 75033
rect 18691 75032 18749 75033
rect 0 74992 1228 75032
rect 1268 74992 1277 75032
rect 2563 74992 2572 75032
rect 2612 74992 3436 75032
rect 3476 74992 3485 75032
rect 4099 74992 4108 75032
rect 4148 74992 4876 75032
rect 4916 74992 4925 75032
rect 11203 74992 11212 75032
rect 11252 74992 11788 75032
rect 11828 74992 11837 75032
rect 15523 74992 15532 75032
rect 15572 74992 15820 75032
rect 15860 74992 15869 75032
rect 17731 74992 17740 75032
rect 17780 74992 18412 75032
rect 18452 74992 18461 75032
rect 18691 74992 18700 75032
rect 18740 74992 20044 75032
rect 20084 74992 20093 75032
rect 0 74972 80 74992
rect 1219 74991 1277 74992
rect 4099 74991 4157 74992
rect 18691 74991 18749 74992
rect 451 74908 460 74948
rect 500 74908 3148 74948
rect 3188 74908 6508 74948
rect 6548 74908 7564 74948
rect 7604 74908 7613 74948
rect 7660 74908 13996 74948
rect 14036 74908 14045 74948
rect 7660 74864 7700 74908
rect 1123 74824 1132 74864
rect 1172 74824 1900 74864
rect 1940 74824 4492 74864
rect 4532 74824 4541 74864
rect 4919 74824 4928 74864
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 5296 74824 5305 74864
rect 7267 74824 7276 74864
rect 7316 74824 7700 74864
rect 9187 74864 9245 74865
rect 9187 74824 9196 74864
rect 9236 74824 12460 74864
rect 12500 74824 12509 74864
rect 20039 74824 20048 74864
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20416 74824 20425 74864
rect 9187 74823 9245 74824
rect 2851 74740 2860 74780
rect 2900 74740 3148 74780
rect 3188 74740 3197 74780
rect 14659 74740 14668 74780
rect 14708 74740 15052 74780
rect 15092 74740 15101 74780
rect 0 74696 80 74716
rect 0 74656 2284 74696
rect 2324 74656 2333 74696
rect 9763 74656 9772 74696
rect 9812 74656 10828 74696
rect 10868 74656 10877 74696
rect 11971 74656 11980 74696
rect 12020 74656 13900 74696
rect 13940 74656 13949 74696
rect 0 74636 80 74656
rect 7747 74612 7805 74613
rect 15427 74612 15485 74613
rect 7662 74572 7756 74612
rect 7796 74572 7805 74612
rect 9475 74572 9484 74612
rect 9524 74572 10060 74612
rect 10100 74572 14516 74612
rect 15139 74572 15148 74612
rect 15188 74572 15436 74612
rect 15476 74572 15485 74612
rect 20227 74572 20236 74612
rect 20276 74572 21292 74612
rect 21332 74572 21341 74612
rect 7747 74571 7805 74572
rect 2755 74528 2813 74529
rect 14476 74528 14516 74572
rect 15427 74571 15485 74572
rect 2755 74488 2764 74528
rect 2804 74488 6604 74528
rect 6644 74488 8044 74528
rect 8084 74488 8093 74528
rect 9571 74488 9580 74528
rect 9620 74488 10252 74528
rect 10292 74488 10301 74528
rect 12547 74488 12556 74528
rect 12596 74488 12844 74528
rect 12884 74488 12893 74528
rect 13123 74488 13132 74528
rect 13172 74488 13612 74528
rect 13652 74488 13661 74528
rect 14467 74488 14476 74528
rect 14516 74488 14525 74528
rect 16483 74488 16492 74528
rect 16532 74488 16972 74528
rect 17012 74488 17021 74528
rect 18019 74488 18028 74528
rect 18068 74488 18077 74528
rect 2755 74487 2813 74488
rect 3331 74444 3389 74445
rect 10723 74444 10781 74445
rect 17923 74444 17981 74445
rect 1507 74404 1516 74444
rect 1556 74404 2956 74444
rect 2996 74404 3005 74444
rect 3139 74404 3148 74444
rect 3188 74404 3340 74444
rect 3380 74404 4300 74444
rect 4340 74404 5356 74444
rect 5396 74404 5405 74444
rect 10637 74404 10732 74444
rect 10772 74404 11404 74444
rect 11444 74404 11453 74444
rect 17838 74404 17932 74444
rect 17972 74404 17981 74444
rect 3331 74403 3389 74404
rect 10723 74403 10781 74404
rect 17923 74403 17981 74404
rect 0 74360 80 74380
rect 1699 74360 1757 74361
rect 18028 74360 18068 74488
rect 0 74320 1708 74360
rect 1748 74320 1757 74360
rect 13987 74320 13996 74360
rect 14036 74320 16204 74360
rect 16244 74320 16253 74360
rect 18028 74320 19660 74360
rect 19700 74320 19709 74360
rect 0 74300 80 74320
rect 1699 74319 1757 74320
rect 3427 74276 3485 74277
rect 3331 74236 3340 74276
rect 3380 74236 3436 74276
rect 3476 74236 3485 74276
rect 3619 74236 3628 74276
rect 3668 74236 3677 74276
rect 5827 74236 5836 74276
rect 5876 74236 7852 74276
rect 7892 74236 10868 74276
rect 11011 74236 11020 74276
rect 11060 74236 16012 74276
rect 16052 74236 19084 74276
rect 19124 74236 19276 74276
rect 19316 74236 19325 74276
rect 3427 74235 3485 74236
rect 3628 74192 3668 74236
rect 10828 74192 10868 74236
rect 2851 74152 2860 74192
rect 2900 74152 7412 74192
rect 9475 74152 9484 74192
rect 9524 74152 9868 74192
rect 9908 74152 9917 74192
rect 10828 74152 12076 74192
rect 12116 74152 12125 74192
rect 3679 74068 3688 74108
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 4056 74068 4065 74108
rect 5635 74068 5644 74108
rect 5684 74068 5932 74108
rect 5972 74068 5981 74108
rect 0 74024 80 74044
rect 7372 74024 7412 74152
rect 16195 74108 16253 74109
rect 9283 74068 9292 74108
rect 9332 74068 11212 74108
rect 11252 74068 11261 74108
rect 11395 74068 11404 74108
rect 11444 74068 13708 74108
rect 13748 74068 16204 74108
rect 16244 74068 16253 74108
rect 18799 74068 18808 74108
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 19176 74068 19185 74108
rect 16195 74067 16253 74068
rect 14275 74024 14333 74025
rect 0 73984 2188 74024
rect 2228 73984 7276 74024
rect 7316 73984 7325 74024
rect 7372 73984 11020 74024
rect 11060 73984 11069 74024
rect 11320 73984 14284 74024
rect 14324 73984 14333 74024
rect 0 73964 80 73984
rect 11320 73940 11360 73984
rect 14275 73983 14333 73984
rect 2371 73900 2380 73940
rect 2420 73900 11360 73940
rect 13411 73900 13420 73940
rect 13460 73900 13900 73940
rect 13940 73900 13949 73940
rect 10435 73856 10493 73857
rect 3139 73816 3148 73856
rect 3188 73816 3532 73856
rect 3572 73816 3581 73856
rect 4771 73816 4780 73856
rect 4820 73816 5644 73856
rect 5684 73816 5693 73856
rect 9955 73816 9964 73856
rect 10004 73816 10156 73856
rect 10196 73816 10205 73856
rect 10350 73816 10444 73856
rect 10484 73816 10493 73856
rect 15331 73816 15340 73856
rect 15380 73816 15389 73856
rect 10435 73815 10493 73816
rect 15340 73772 15380 73816
rect 739 73732 748 73772
rect 788 73732 2540 73772
rect 5347 73732 5356 73772
rect 5396 73732 13708 73772
rect 13748 73732 14764 73772
rect 14804 73732 14813 73772
rect 15340 73732 16108 73772
rect 16148 73732 16157 73772
rect 0 73688 80 73708
rect 2500 73688 2540 73732
rect 8611 73688 8669 73689
rect 0 73648 1036 73688
rect 1076 73648 1085 73688
rect 2500 73648 3532 73688
rect 3572 73648 6604 73688
rect 6644 73648 6653 73688
rect 7075 73648 7084 73688
rect 7124 73648 7468 73688
rect 7508 73648 7660 73688
rect 7700 73648 7709 73688
rect 8131 73648 8140 73688
rect 8180 73648 8189 73688
rect 8419 73648 8428 73688
rect 8468 73648 8620 73688
rect 8660 73648 8669 73688
rect 0 73628 80 73648
rect 6883 73604 6941 73605
rect 8140 73604 8180 73648
rect 8611 73647 8669 73648
rect 9868 73648 10348 73688
rect 10388 73648 10397 73688
rect 10627 73648 10636 73688
rect 10676 73648 10828 73688
rect 10868 73648 10877 73688
rect 13123 73648 13132 73688
rect 13172 73648 13516 73688
rect 13556 73648 13565 73688
rect 18115 73648 18124 73688
rect 18164 73648 19756 73688
rect 19796 73648 19805 73688
rect 9868 73604 9908 73648
rect 2659 73564 2668 73604
rect 2708 73564 6892 73604
rect 6932 73564 8180 73604
rect 9859 73564 9868 73604
rect 9908 73564 9917 73604
rect 6883 73563 6941 73564
rect 7651 73520 7709 73521
rect 10156 73520 10196 73648
rect 12067 73564 12076 73604
rect 12116 73564 12940 73604
rect 12980 73564 16396 73604
rect 16436 73564 16445 73604
rect 6979 73480 6988 73520
rect 7028 73480 7372 73520
rect 7412 73480 7421 73520
rect 7566 73480 7660 73520
rect 7700 73480 7709 73520
rect 7843 73480 7852 73520
rect 7892 73480 8236 73520
rect 8276 73480 8285 73520
rect 10147 73480 10156 73520
rect 10196 73480 10205 73520
rect 13987 73480 13996 73520
rect 14036 73480 14284 73520
rect 14324 73480 14333 73520
rect 17827 73480 17836 73520
rect 17876 73480 18508 73520
rect 18548 73480 18557 73520
rect 7651 73479 7709 73480
rect 2947 73436 3005 73437
rect 2947 73396 2956 73436
rect 2996 73396 3340 73436
rect 3380 73396 3389 73436
rect 8131 73396 8140 73436
rect 8180 73396 8620 73436
rect 8660 73396 8669 73436
rect 18403 73396 18412 73436
rect 18452 73396 18700 73436
rect 18740 73396 18749 73436
rect 2947 73395 3005 73396
rect 0 73352 80 73372
rect 8227 73352 8285 73353
rect 0 73312 2540 73352
rect 4919 73312 4928 73352
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 5296 73312 5305 73352
rect 6691 73312 6700 73352
rect 6740 73312 7084 73352
rect 7124 73312 7133 73352
rect 8142 73312 8236 73352
rect 8276 73312 8285 73352
rect 9763 73312 9772 73352
rect 9812 73312 10540 73352
rect 10580 73312 10589 73352
rect 20039 73312 20048 73352
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20416 73312 20425 73352
rect 0 73292 80 73312
rect 2500 73268 2540 73312
rect 8227 73311 8285 73312
rect 10435 73268 10493 73269
rect 2500 73228 3340 73268
rect 3380 73228 3389 73268
rect 5635 73228 5644 73268
rect 5684 73228 9388 73268
rect 9428 73228 9676 73268
rect 9716 73228 9725 73268
rect 10350 73228 10444 73268
rect 10484 73228 10493 73268
rect 10435 73227 10493 73228
rect 643 73184 701 73185
rect 12451 73184 12509 73185
rect 643 73144 652 73184
rect 692 73144 1172 73184
rect 1219 73144 1228 73184
rect 1268 73144 1277 73184
rect 5644 73144 5932 73184
rect 5972 73144 5981 73184
rect 7555 73144 7564 73184
rect 7604 73144 7948 73184
rect 7988 73144 7997 73184
rect 10243 73144 10252 73184
rect 10292 73144 10676 73184
rect 643 73143 701 73144
rect 1132 73101 1172 73144
rect 1123 73100 1181 73101
rect 1123 73060 1132 73100
rect 1172 73060 1181 73100
rect 1123 73059 1181 73060
rect 0 73016 80 73036
rect 1228 73016 1268 73144
rect 3139 73100 3197 73101
rect 5644 73100 5684 73144
rect 10636 73101 10676 73144
rect 12172 73144 12460 73184
rect 12500 73144 12509 73184
rect 10627 73100 10685 73101
rect 3108 73060 3148 73100
rect 3188 73060 3197 73100
rect 5635 73060 5644 73100
rect 5684 73060 5693 73100
rect 10596 73060 10636 73100
rect 10676 73060 10685 73100
rect 3139 73059 3197 73060
rect 10627 73059 10685 73060
rect 2371 73016 2429 73017
rect 0 72976 1172 73016
rect 1228 72976 2380 73016
rect 2420 72976 2429 73016
rect 3148 73016 3188 73059
rect 10636 73016 10676 73059
rect 12172 73016 12212 73144
rect 12451 73143 12509 73144
rect 13507 73184 13565 73185
rect 13507 73144 13516 73184
rect 13556 73144 13804 73184
rect 13844 73144 13853 73184
rect 15235 73144 15244 73184
rect 15284 73144 17548 73184
rect 17588 73144 18124 73184
rect 18164 73144 18173 73184
rect 19843 73144 19852 73184
rect 19892 73144 20044 73184
rect 20084 73144 20093 73184
rect 13507 73143 13565 73144
rect 13507 73060 13516 73100
rect 13556 73060 13900 73100
rect 13940 73060 13949 73100
rect 17604 73060 17644 73100
rect 17684 73060 17693 73100
rect 13900 73016 13940 73060
rect 17644 73016 17684 73060
rect 3148 72976 3628 73016
rect 3668 72976 3677 73016
rect 4867 72976 4876 73016
rect 4916 72976 7756 73016
rect 7796 72976 7805 73016
rect 10243 72976 10252 73016
rect 10292 72976 10676 73016
rect 11320 72976 12212 73016
rect 12259 72976 12268 73016
rect 12308 72976 13612 73016
rect 13652 72976 13804 73016
rect 13844 72976 13853 73016
rect 13900 72976 14284 73016
rect 14324 72976 14333 73016
rect 17251 72976 17260 73016
rect 17300 72976 17684 73016
rect 0 72956 80 72976
rect 1132 72848 1172 72976
rect 2371 72975 2429 72976
rect 1315 72932 1373 72933
rect 6796 72932 6836 72976
rect 11320 72932 11360 72976
rect 1315 72892 1324 72932
rect 1364 72892 2540 72932
rect 6787 72892 6796 72932
rect 6836 72892 6876 72932
rect 7843 72892 7852 72932
rect 7892 72892 11360 72932
rect 12643 72892 12652 72932
rect 12692 72892 13132 72932
rect 13172 72892 13181 72932
rect 15907 72892 15916 72932
rect 15956 72892 16396 72932
rect 16436 72892 16445 72932
rect 16867 72892 16876 72932
rect 16916 72892 17452 72932
rect 17492 72892 17501 72932
rect 1315 72891 1373 72892
rect 2500 72848 2540 72892
rect 13507 72848 13565 72849
rect 1132 72808 1420 72848
rect 1460 72808 1469 72848
rect 2500 72808 4780 72848
rect 4820 72808 10540 72848
rect 10580 72808 10589 72848
rect 13422 72808 13516 72848
rect 13556 72808 13565 72848
rect 15427 72808 15436 72848
rect 15476 72808 15724 72848
rect 15764 72808 15773 72848
rect 17539 72808 17548 72848
rect 17588 72808 18124 72848
rect 18164 72808 18173 72848
rect 13507 72807 13565 72808
rect 19651 72764 19709 72765
rect 5251 72724 5260 72764
rect 5300 72724 6700 72764
rect 6740 72724 6749 72764
rect 19651 72724 19660 72764
rect 19700 72724 19852 72764
rect 19892 72724 19901 72764
rect 19651 72723 19709 72724
rect 0 72680 80 72700
rect 3235 72680 3293 72681
rect 0 72640 3244 72680
rect 3284 72640 9100 72680
rect 9140 72640 12844 72680
rect 12884 72640 12893 72680
rect 0 72620 80 72640
rect 3235 72639 3293 72640
rect 3679 72556 3688 72596
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 4056 72556 4065 72596
rect 18799 72556 18808 72596
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 19176 72556 19185 72596
rect 21424 72512 21504 72532
rect 5731 72472 5740 72512
rect 5780 72472 6124 72512
rect 6164 72472 6173 72512
rect 21091 72472 21100 72512
rect 21140 72472 21504 72512
rect 21424 72452 21504 72472
rect 9379 72428 9437 72429
rect 2467 72388 2476 72428
rect 2516 72388 2956 72428
rect 2996 72388 5836 72428
rect 5876 72388 5885 72428
rect 9294 72388 9388 72428
rect 9428 72388 11404 72428
rect 11444 72388 11453 72428
rect 11683 72388 11692 72428
rect 11732 72388 15340 72428
rect 15380 72388 15389 72428
rect 0 72344 80 72364
rect 3427 72344 3485 72345
rect 0 72304 2860 72344
rect 2900 72304 2909 72344
rect 3342 72304 3436 72344
rect 3476 72304 3485 72344
rect 4003 72304 4012 72344
rect 4052 72304 4300 72344
rect 4340 72304 4349 72344
rect 0 72284 80 72304
rect 3427 72303 3485 72304
rect 4291 72136 4300 72176
rect 4340 72136 5452 72176
rect 5492 72136 5501 72176
rect 451 72092 509 72093
rect 451 72052 460 72092
rect 500 72052 4876 72092
rect 4916 72052 4925 72092
rect 451 72051 509 72052
rect 0 72008 80 72028
rect 2659 72008 2717 72009
rect 0 71968 2668 72008
rect 2708 71968 2717 72008
rect 5251 71968 5260 72008
rect 5300 71968 5309 72008
rect 0 71948 80 71968
rect 2659 71967 2717 71968
rect 5260 71924 5300 71968
rect 259 71884 268 71924
rect 308 71884 5300 71924
rect 5836 71924 5876 72388
rect 9379 72387 9437 72388
rect 7171 72304 7180 72344
rect 7220 72304 15244 72344
rect 15284 72304 15293 72344
rect 11875 72260 11933 72261
rect 9187 72220 9196 72260
rect 9236 72220 9772 72260
rect 9812 72220 9821 72260
rect 11790 72220 11884 72260
rect 11924 72220 11933 72260
rect 11875 72219 11933 72220
rect 18403 72176 18461 72177
rect 21424 72176 21504 72196
rect 5923 72136 5932 72176
rect 5972 72136 6604 72176
rect 6644 72136 6653 72176
rect 10243 72136 10252 72176
rect 10292 72136 10828 72176
rect 10868 72136 10877 72176
rect 11683 72136 11692 72176
rect 11732 72136 13420 72176
rect 13460 72136 13469 72176
rect 14659 72136 14668 72176
rect 14708 72136 15052 72176
rect 15092 72136 15244 72176
rect 15284 72136 15293 72176
rect 18403 72136 18412 72176
rect 18452 72136 21504 72176
rect 18403 72135 18461 72136
rect 21424 72116 21504 72136
rect 19267 72092 19325 72093
rect 9667 72052 9676 72092
rect 9716 72052 10636 72092
rect 10676 72052 11116 72092
rect 11156 72052 11165 72092
rect 13987 72052 13996 72092
rect 14036 72052 14572 72092
rect 14612 72052 14621 72092
rect 18979 72052 18988 72092
rect 19028 72052 19276 72092
rect 19316 72052 19372 72092
rect 19412 72052 19440 72092
rect 19267 72051 19325 72052
rect 7939 72008 7997 72009
rect 17443 72008 17501 72009
rect 7747 71968 7756 72008
rect 7796 71968 7948 72008
rect 7988 71968 7997 72008
rect 10435 71968 10444 72008
rect 10484 71968 10828 72008
rect 10868 71968 11308 72008
rect 11348 71968 11360 72008
rect 13411 71968 13420 72008
rect 13460 71968 13804 72008
rect 13844 71968 13853 72008
rect 15427 71968 15436 72008
rect 15476 71968 16396 72008
rect 16436 71968 16445 72008
rect 17358 71968 17452 72008
rect 17492 71968 17501 72008
rect 7939 71967 7997 71968
rect 5836 71884 5932 71924
rect 5972 71884 5981 71924
rect 7651 71884 7660 71924
rect 7700 71884 7948 71924
rect 7988 71884 7997 71924
rect 3523 71840 3581 71841
rect 11203 71840 11261 71841
rect 1315 71800 1324 71840
rect 1364 71800 1804 71840
rect 1844 71800 1853 71840
rect 3235 71800 3244 71840
rect 3284 71800 3532 71840
rect 3572 71800 3581 71840
rect 4919 71800 4928 71840
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 5296 71800 5305 71840
rect 6019 71800 6028 71840
rect 6068 71800 7564 71840
rect 7604 71800 7613 71840
rect 9283 71800 9292 71840
rect 9332 71800 11212 71840
rect 11252 71800 11261 71840
rect 11320 71840 11360 71968
rect 17443 71967 17501 71968
rect 13027 71884 13036 71924
rect 13076 71884 14188 71924
rect 14228 71884 16780 71924
rect 16820 71884 16829 71924
rect 21424 71841 21504 71860
rect 12547 71840 12605 71841
rect 13219 71840 13277 71841
rect 21379 71840 21504 71841
rect 11320 71800 11788 71840
rect 11828 71800 11837 71840
rect 12355 71800 12364 71840
rect 12404 71800 12556 71840
rect 12596 71800 12605 71840
rect 13134 71800 13228 71840
rect 13268 71800 13277 71840
rect 13411 71800 13420 71840
rect 13460 71800 14228 71840
rect 20039 71800 20048 71840
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20416 71800 20425 71840
rect 21379 71800 21388 71840
rect 21428 71800 21504 71840
rect 3523 71799 3581 71800
rect 11203 71799 11261 71800
rect 12547 71799 12605 71800
rect 13219 71799 13277 71800
rect 10147 71756 10205 71757
rect 13795 71756 13853 71757
rect 14188 71756 14228 71800
rect 21379 71799 21504 71800
rect 21424 71780 21504 71799
rect 2563 71716 2572 71756
rect 2612 71716 2956 71756
rect 2996 71716 3005 71756
rect 3331 71716 3340 71756
rect 3380 71716 3532 71756
rect 3572 71716 3581 71756
rect 4387 71716 4396 71756
rect 4436 71716 4588 71756
rect 4628 71716 4637 71756
rect 5347 71716 5356 71756
rect 5396 71716 10156 71756
rect 10196 71716 10205 71756
rect 10147 71715 10205 71716
rect 11320 71716 13804 71756
rect 13844 71716 13853 71756
rect 14179 71716 14188 71756
rect 14228 71716 14237 71756
rect 0 71672 80 71692
rect 11320 71672 11360 71716
rect 13795 71715 13853 71716
rect 13411 71672 13469 71673
rect 0 71632 1364 71672
rect 1411 71632 1420 71672
rect 1460 71632 2092 71672
rect 2132 71632 8812 71672
rect 8852 71632 8861 71672
rect 10051 71632 10060 71672
rect 10100 71632 11360 71672
rect 13326 71632 13420 71672
rect 13460 71632 13469 71672
rect 0 71612 80 71632
rect 1324 71588 1364 71632
rect 13411 71631 13469 71632
rect 1315 71548 1324 71588
rect 1364 71548 1373 71588
rect 2563 71548 2572 71588
rect 2612 71548 3340 71588
rect 3380 71548 6068 71588
rect 7459 71548 7468 71588
rect 7508 71548 9100 71588
rect 9140 71548 9149 71588
rect 10339 71548 10348 71588
rect 10388 71548 10732 71588
rect 10772 71548 10781 71588
rect 12355 71548 12364 71588
rect 12404 71548 12652 71588
rect 12692 71548 12701 71588
rect 13987 71548 13996 71588
rect 14036 71548 14380 71588
rect 14420 71548 14429 71588
rect 6028 71504 6068 71548
rect 13315 71504 13373 71505
rect 14563 71504 14621 71505
rect 20803 71504 20861 71505
rect 21424 71504 21504 71524
rect 4291 71464 4300 71504
rect 4340 71464 4684 71504
rect 4724 71464 4733 71504
rect 6019 71464 6028 71504
rect 6068 71464 7372 71504
rect 7412 71464 7421 71504
rect 8515 71464 8524 71504
rect 8564 71464 8908 71504
rect 8948 71464 8957 71504
rect 9772 71464 12212 71504
rect 12259 71464 12268 71504
rect 12308 71464 13132 71504
rect 13172 71464 13181 71504
rect 13315 71464 13324 71504
rect 13364 71464 13458 71504
rect 14478 71464 14572 71504
rect 14612 71464 14621 71504
rect 15619 71464 15628 71504
rect 15668 71464 15820 71504
rect 15860 71464 17164 71504
rect 17204 71464 17452 71504
rect 17492 71464 19660 71504
rect 19700 71464 19709 71504
rect 20803 71464 20812 71504
rect 20852 71464 21504 71504
rect 1795 71380 1804 71420
rect 1844 71380 9676 71420
rect 9716 71380 9725 71420
rect 0 71336 80 71356
rect 1315 71336 1373 71337
rect 0 71296 1324 71336
rect 1364 71296 1373 71336
rect 0 71276 80 71296
rect 1315 71295 1373 71296
rect 4771 71336 4829 71337
rect 9772 71336 9812 71464
rect 12172 71420 12212 71464
rect 13315 71463 13373 71464
rect 14563 71463 14621 71464
rect 20803 71463 20861 71464
rect 21424 71444 21504 71464
rect 16195 71420 16253 71421
rect 12172 71380 15148 71420
rect 15188 71380 15724 71420
rect 15764 71380 15773 71420
rect 16110 71380 16204 71420
rect 16244 71380 16253 71420
rect 16195 71379 16253 71380
rect 17635 71336 17693 71337
rect 4771 71296 4780 71336
rect 4820 71296 4876 71336
rect 4916 71296 4925 71336
rect 5347 71296 5356 71336
rect 5396 71296 6220 71336
rect 6260 71296 6269 71336
rect 6883 71296 6892 71336
rect 6932 71296 9812 71336
rect 10531 71296 10540 71336
rect 10580 71296 15436 71336
rect 15476 71296 15485 71336
rect 15916 71296 17644 71336
rect 17684 71296 18604 71336
rect 18644 71296 18653 71336
rect 4771 71295 4829 71296
rect 4876 71252 4916 71296
rect 9763 71252 9821 71253
rect 15916 71252 15956 71296
rect 17635 71295 17693 71296
rect 19843 71252 19901 71253
rect 4003 71212 4012 71252
rect 4052 71212 4300 71252
rect 4340 71212 4349 71252
rect 4876 71212 9772 71252
rect 9812 71212 9821 71252
rect 10627 71212 10636 71252
rect 10676 71212 11308 71252
rect 11348 71212 11596 71252
rect 11636 71212 11645 71252
rect 12067 71212 12076 71252
rect 12116 71212 15956 71252
rect 16003 71212 16012 71252
rect 16052 71212 16492 71252
rect 16532 71212 16541 71252
rect 16588 71212 18316 71252
rect 18356 71212 19852 71252
rect 19892 71212 19901 71252
rect 9763 71211 9821 71212
rect 1795 71168 1853 71169
rect 13219 71168 13277 71169
rect 1411 71128 1420 71168
rect 1460 71128 1804 71168
rect 1844 71128 1853 71168
rect 3523 71128 3532 71168
rect 3572 71128 8468 71168
rect 8803 71128 8812 71168
rect 8852 71128 13228 71168
rect 13268 71128 13277 71168
rect 1795 71127 1853 71128
rect 8428 71084 8468 71128
rect 13219 71127 13277 71128
rect 13795 71168 13853 71169
rect 16588 71168 16628 71212
rect 19843 71211 19901 71212
rect 13795 71128 13804 71168
rect 13844 71128 16628 71168
rect 16771 71168 16829 71169
rect 21424 71168 21504 71188
rect 16771 71128 16780 71168
rect 16820 71128 21504 71168
rect 13795 71127 13853 71128
rect 16771 71127 16829 71128
rect 21424 71108 21504 71128
rect 14371 71084 14429 71085
rect 19555 71084 19613 71085
rect 3679 71044 3688 71084
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 4056 71044 4065 71084
rect 7651 71044 7660 71084
rect 7700 71044 8236 71084
rect 8276 71044 8285 71084
rect 8419 71044 8428 71084
rect 8468 71044 14380 71084
rect 14420 71044 14429 71084
rect 18799 71044 18808 71084
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 19176 71044 19185 71084
rect 19555 71044 19564 71084
rect 19604 71044 19756 71084
rect 19796 71044 19805 71084
rect 14371 71043 14429 71044
rect 19555 71043 19613 71044
rect 0 71000 80 71020
rect 0 70960 12076 71000
rect 12116 70960 12125 71000
rect 12355 70960 12364 71000
rect 12404 70960 12413 71000
rect 13315 70960 13324 71000
rect 13364 70960 16012 71000
rect 16052 70960 16061 71000
rect 17251 70960 17260 71000
rect 17300 70960 17548 71000
rect 17588 70960 19564 71000
rect 19604 70960 19613 71000
rect 0 70940 80 70960
rect 3523 70916 3581 70917
rect 7843 70916 7901 70917
rect 3523 70876 3532 70916
rect 3572 70876 4396 70916
rect 4436 70876 7852 70916
rect 7892 70876 7901 70916
rect 3523 70875 3581 70876
rect 7843 70875 7901 70876
rect 8611 70916 8669 70917
rect 12364 70916 12404 70960
rect 8611 70876 8620 70916
rect 8660 70876 8716 70916
rect 8756 70876 8765 70916
rect 8995 70876 9004 70916
rect 9044 70876 9388 70916
rect 9428 70876 10924 70916
rect 10964 70876 10973 70916
rect 11320 70876 11692 70916
rect 11732 70876 11741 70916
rect 11980 70876 12268 70916
rect 12308 70876 12317 70916
rect 12364 70876 14380 70916
rect 14420 70876 14429 70916
rect 14563 70876 14572 70916
rect 14612 70876 15052 70916
rect 15092 70876 15101 70916
rect 15235 70876 15244 70916
rect 15284 70876 15820 70916
rect 15860 70876 15869 70916
rect 8611 70875 8669 70876
rect 3331 70832 3389 70833
rect 5635 70832 5693 70833
rect 11320 70832 11360 70876
rect 2467 70792 2476 70832
rect 2516 70792 3340 70832
rect 3380 70792 4436 70832
rect 4483 70792 4492 70832
rect 4532 70792 4541 70832
rect 4771 70792 4780 70832
rect 4820 70792 5644 70832
rect 5684 70792 5693 70832
rect 9091 70792 9100 70832
rect 9140 70792 11360 70832
rect 3331 70791 3389 70792
rect 4396 70748 4436 70792
rect 4492 70748 4532 70792
rect 5635 70791 5693 70792
rect 6979 70748 7037 70749
rect 4387 70708 4396 70748
rect 4436 70708 4445 70748
rect 4492 70708 4916 70748
rect 6883 70708 6892 70748
rect 6932 70708 6988 70748
rect 7028 70708 7037 70748
rect 11980 70748 12020 70876
rect 15139 70832 15197 70833
rect 21424 70832 21504 70852
rect 12067 70792 12076 70832
rect 12116 70792 12460 70832
rect 12500 70792 12509 70832
rect 12739 70792 12748 70832
rect 12788 70792 13036 70832
rect 13076 70792 13085 70832
rect 15139 70792 15148 70832
rect 15188 70792 21504 70832
rect 15139 70791 15197 70792
rect 21424 70772 21504 70792
rect 19651 70748 19709 70749
rect 11980 70708 13748 70748
rect 14947 70708 14956 70748
rect 14996 70708 15148 70748
rect 15188 70708 15197 70748
rect 19566 70708 19660 70748
rect 19700 70708 19709 70748
rect 0 70664 80 70684
rect 4876 70664 4916 70708
rect 6979 70707 7037 70708
rect 7939 70664 7997 70665
rect 12547 70664 12605 70665
rect 13708 70664 13748 70708
rect 19651 70707 19709 70708
rect 0 70624 1036 70664
rect 1076 70624 1085 70664
rect 1219 70624 1228 70664
rect 1268 70624 2092 70664
rect 2132 70624 2380 70664
rect 2420 70624 2429 70664
rect 3043 70624 3052 70664
rect 3092 70624 3532 70664
rect 3572 70624 3581 70664
rect 4867 70624 4876 70664
rect 4916 70624 7948 70664
rect 7988 70624 7997 70664
rect 0 70604 80 70624
rect 7939 70623 7997 70624
rect 8044 70624 8332 70664
rect 8372 70624 8381 70664
rect 8803 70624 8812 70664
rect 8852 70624 9484 70664
rect 9524 70624 9533 70664
rect 10915 70624 10924 70664
rect 10964 70624 11500 70664
rect 11540 70624 11549 70664
rect 11779 70624 11788 70664
rect 11828 70624 12076 70664
rect 12116 70624 12125 70664
rect 12547 70624 12556 70664
rect 12596 70624 12844 70664
rect 12884 70624 12893 70664
rect 13708 70624 15244 70664
rect 15284 70624 15293 70664
rect 17923 70624 17932 70664
rect 17972 70624 17981 70664
rect 4291 70580 4349 70581
rect 8044 70580 8084 70624
rect 12547 70623 12605 70624
rect 8995 70580 9053 70581
rect 15043 70580 15101 70581
rect 15523 70580 15581 70581
rect 3139 70540 3148 70580
rect 3188 70540 3197 70580
rect 4206 70540 4300 70580
rect 4340 70540 4349 70580
rect 8035 70540 8044 70580
rect 8084 70540 8093 70580
rect 8995 70540 9004 70580
rect 9044 70540 10060 70580
rect 10100 70540 10109 70580
rect 10531 70540 10540 70580
rect 10580 70540 11116 70580
rect 11156 70540 11165 70580
rect 15043 70540 15052 70580
rect 15092 70540 15148 70580
rect 15188 70540 15197 70580
rect 15438 70540 15532 70580
rect 15572 70540 15581 70580
rect 17635 70540 17644 70580
rect 17684 70540 17693 70580
rect 3148 70496 3188 70540
rect 4291 70539 4349 70540
rect 8995 70539 9053 70540
rect 15043 70539 15101 70540
rect 15523 70539 15581 70540
rect 2371 70456 2380 70496
rect 2420 70456 2668 70496
rect 2708 70456 2717 70496
rect 3148 70456 4204 70496
rect 4244 70456 4253 70496
rect 4780 70456 12652 70496
rect 12692 70456 14188 70496
rect 14228 70456 14237 70496
rect 0 70328 80 70348
rect 0 70288 940 70328
rect 980 70288 989 70328
rect 0 70268 80 70288
rect 4780 70160 4820 70456
rect 7939 70372 7948 70412
rect 7988 70372 8428 70412
rect 8468 70372 8477 70412
rect 10147 70372 10156 70412
rect 10196 70372 10636 70412
rect 10676 70372 10685 70412
rect 11299 70372 11308 70412
rect 11348 70372 12076 70412
rect 12116 70372 12125 70412
rect 17644 70328 17684 70540
rect 17932 70496 17972 70624
rect 20707 70496 20765 70497
rect 21424 70496 21504 70516
rect 17932 70456 18124 70496
rect 18164 70456 18508 70496
rect 18548 70456 18557 70496
rect 19363 70456 19372 70496
rect 19412 70456 19948 70496
rect 19988 70456 19997 70496
rect 20707 70456 20716 70496
rect 20756 70456 21504 70496
rect 20707 70455 20765 70456
rect 21424 70436 21504 70456
rect 18211 70328 18269 70329
rect 4919 70288 4928 70328
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 5296 70288 5305 70328
rect 6307 70288 6316 70328
rect 6356 70288 16684 70328
rect 16724 70288 17452 70328
rect 17492 70288 17501 70328
rect 17644 70288 17836 70328
rect 17876 70288 17885 70328
rect 18211 70288 18220 70328
rect 18260 70288 18700 70328
rect 18740 70288 18749 70328
rect 20039 70288 20048 70328
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20416 70288 20425 70328
rect 18211 70287 18269 70288
rect 11299 70244 11357 70245
rect 11299 70204 11308 70244
rect 11348 70204 20524 70244
rect 20564 70204 20573 70244
rect 11299 70203 11357 70204
rect 5347 70160 5405 70161
rect 7171 70160 7229 70161
rect 11203 70160 11261 70161
rect 14563 70160 14621 70161
rect 17827 70160 17885 70161
rect 21424 70160 21504 70180
rect 172 70120 4820 70160
rect 5155 70120 5164 70160
rect 5204 70120 5356 70160
rect 5396 70120 5405 70160
rect 6595 70120 6604 70160
rect 6644 70120 6892 70160
rect 6932 70120 6941 70160
rect 7171 70120 7180 70160
rect 7220 70120 7756 70160
rect 7796 70120 7805 70160
rect 11118 70120 11212 70160
rect 11252 70120 11261 70160
rect 0 69992 80 70012
rect 0 69932 116 69992
rect 76 69908 116 69932
rect 172 69908 212 70120
rect 5347 70119 5405 70120
rect 7171 70119 7229 70120
rect 11203 70119 11261 70120
rect 11980 70120 14572 70160
rect 14612 70120 14621 70160
rect 15427 70120 15436 70160
rect 15476 70120 15572 70160
rect 7180 70076 7220 70119
rect 9475 70076 9533 70077
rect 11980 70076 12020 70120
rect 14563 70119 14621 70120
rect 4483 70036 4492 70076
rect 4532 70036 7220 70076
rect 7939 70036 7948 70076
rect 7988 70036 9484 70076
rect 9524 70036 9533 70076
rect 9475 70035 9533 70036
rect 11320 70036 11980 70076
rect 12020 70036 12029 70076
rect 14659 70036 14668 70076
rect 14708 70036 14956 70076
rect 14996 70036 15005 70076
rect 4291 69992 4349 69993
rect 11320 69992 11360 70036
rect 1315 69952 1324 69992
rect 1364 69952 4052 69992
rect 4012 69908 4052 69952
rect 4291 69952 4300 69992
rect 4340 69952 7276 69992
rect 7316 69952 7325 69992
rect 7555 69952 7564 69992
rect 7604 69952 8627 69992
rect 8667 69952 11360 69992
rect 11683 69952 11692 69992
rect 11732 69952 12076 69992
rect 12116 69952 12125 69992
rect 13219 69952 13228 69992
rect 13268 69952 13420 69992
rect 13460 69952 13469 69992
rect 14275 69952 14284 69992
rect 14324 69952 15340 69992
rect 15380 69952 15389 69992
rect 4291 69951 4349 69952
rect 11587 69908 11645 69909
rect 15532 69908 15572 70120
rect 17827 70120 17836 70160
rect 17876 70120 21504 70160
rect 17827 70119 17885 70120
rect 21424 70100 21504 70120
rect 19939 70076 19997 70077
rect 19854 70036 19948 70076
rect 19988 70036 19997 70076
rect 19939 70035 19997 70036
rect 18499 69992 18557 69993
rect 18499 69952 18508 69992
rect 18548 69952 18796 69992
rect 18836 69952 18845 69992
rect 18499 69951 18557 69952
rect 76 69868 212 69908
rect 4003 69868 4012 69908
rect 4052 69868 11444 69908
rect 11502 69868 11596 69908
rect 11636 69868 11645 69908
rect 15523 69868 15532 69908
rect 15572 69868 15581 69908
rect 15916 69868 16300 69908
rect 16340 69868 16349 69908
rect 11404 69824 11444 69868
rect 11587 69867 11645 69868
rect 14563 69824 14621 69825
rect 15916 69824 15956 69868
rect 19267 69824 19325 69825
rect 21424 69824 21504 69844
rect 11404 69784 14572 69824
rect 14612 69784 14621 69824
rect 15427 69784 15436 69824
rect 15476 69784 15956 69824
rect 16012 69784 19276 69824
rect 19316 69784 19325 69824
rect 19459 69784 19468 69824
rect 19508 69784 19852 69824
rect 19892 69784 19901 69824
rect 20140 69784 21504 69824
rect 14563 69783 14621 69784
rect 355 69700 364 69740
rect 404 69700 6316 69740
rect 6356 69700 6365 69740
rect 11299 69700 11308 69740
rect 11348 69700 11692 69740
rect 11732 69700 11741 69740
rect 11971 69700 11980 69740
rect 12020 69700 12172 69740
rect 12212 69700 12221 69740
rect 0 69656 80 69676
rect 16012 69656 16052 69784
rect 19267 69783 19325 69784
rect 16099 69740 16157 69741
rect 20140 69740 20180 69784
rect 21424 69764 21504 69784
rect 16099 69700 16108 69740
rect 16148 69700 20180 69740
rect 16099 69699 16157 69700
rect 0 69616 16052 69656
rect 16387 69616 16396 69656
rect 16436 69616 16876 69656
rect 16916 69616 16925 69656
rect 18019 69616 18028 69656
rect 18068 69616 18316 69656
rect 18356 69616 18365 69656
rect 0 69596 80 69616
rect 1411 69532 1420 69572
rect 1460 69532 1900 69572
rect 1940 69532 1949 69572
rect 3679 69532 3688 69572
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 4056 69532 4065 69572
rect 18799 69532 18808 69572
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 19176 69532 19185 69572
rect 20611 69488 20669 69489
rect 21424 69488 21504 69508
rect 2500 69448 16876 69488
rect 16916 69448 16925 69488
rect 20611 69448 20620 69488
rect 20660 69448 21504 69488
rect 2275 69404 2333 69405
rect 2500 69404 2540 69448
rect 20611 69447 20669 69448
rect 21424 69428 21504 69448
rect 1891 69364 1900 69404
rect 1940 69364 2284 69404
rect 2324 69364 2333 69404
rect 2275 69363 2333 69364
rect 2380 69364 2540 69404
rect 4099 69364 4108 69404
rect 4148 69364 4396 69404
rect 4436 69364 4445 69404
rect 7267 69364 7276 69404
rect 7316 69364 14764 69404
rect 14804 69364 14813 69404
rect 0 69320 80 69340
rect 2380 69320 2420 69364
rect 13603 69320 13661 69321
rect 0 69280 2420 69320
rect 6019 69280 6028 69320
rect 6068 69280 6700 69320
rect 6740 69280 7468 69320
rect 7508 69280 7517 69320
rect 9763 69280 9772 69320
rect 9812 69280 11212 69320
rect 11252 69280 13228 69320
rect 13268 69280 13277 69320
rect 13603 69280 13612 69320
rect 13652 69280 14092 69320
rect 14132 69280 14141 69320
rect 0 69260 80 69280
rect 13603 69279 13661 69280
rect 17635 69236 17693 69237
rect 2467 69196 2476 69236
rect 2516 69196 3052 69236
rect 3092 69196 4108 69236
rect 4148 69196 4492 69236
rect 4532 69196 7852 69236
rect 7892 69196 7901 69236
rect 8899 69196 8908 69236
rect 8948 69196 12844 69236
rect 12884 69196 12893 69236
rect 17635 69196 17644 69236
rect 17684 69196 17932 69236
rect 17972 69196 17981 69236
rect 17635 69195 17693 69196
rect 2083 69152 2141 69153
rect 2371 69152 2429 69153
rect 3139 69152 3197 69153
rect 21424 69152 21504 69172
rect 1219 69112 1228 69152
rect 1268 69112 2092 69152
rect 2132 69112 2380 69152
rect 2420 69112 2429 69152
rect 2659 69112 2668 69152
rect 2708 69112 3148 69152
rect 3188 69112 3197 69152
rect 4675 69112 4684 69152
rect 4724 69112 5548 69152
rect 5588 69112 6028 69152
rect 6068 69112 6077 69152
rect 8419 69112 8428 69152
rect 8468 69112 10348 69152
rect 10388 69112 10397 69152
rect 10819 69112 10828 69152
rect 10868 69112 12460 69152
rect 12500 69112 12509 69152
rect 14179 69112 14188 69152
rect 14228 69112 14476 69152
rect 14516 69112 14525 69152
rect 15907 69112 15916 69152
rect 15956 69112 16300 69152
rect 16340 69112 19180 69152
rect 19220 69112 19372 69152
rect 19412 69112 19421 69152
rect 20515 69112 20524 69152
rect 20564 69112 21504 69152
rect 2083 69111 2141 69112
rect 2371 69111 2429 69112
rect 3139 69111 3197 69112
rect 21424 69092 21504 69112
rect 19555 69068 19613 69069
rect 6883 69028 6892 69068
rect 6932 69028 8332 69068
rect 8372 69028 13420 69068
rect 13460 69028 13469 69068
rect 19459 69028 19468 69068
rect 19508 69028 19564 69068
rect 19604 69028 19613 69068
rect 19555 69027 19613 69028
rect 0 68984 80 69004
rect 163 68984 221 68985
rect 6883 68984 6941 68985
rect 19267 68984 19325 68985
rect 0 68944 172 68984
rect 212 68944 221 68984
rect 4099 68944 4108 68984
rect 4148 68944 4300 68984
rect 4340 68944 4349 68984
rect 6883 68944 6892 68984
rect 6932 68944 13804 68984
rect 13844 68944 13853 68984
rect 14659 68944 14668 68984
rect 14708 68944 16108 68984
rect 16148 68944 16157 68984
rect 19267 68944 19276 68984
rect 19316 68944 20044 68984
rect 20084 68944 20093 68984
rect 0 68924 80 68944
rect 163 68943 221 68944
rect 6883 68943 6941 68944
rect 19267 68943 19325 68944
rect 3235 68900 3293 68901
rect 2947 68860 2956 68900
rect 2996 68860 3244 68900
rect 3284 68860 3293 68900
rect 4195 68860 4204 68900
rect 4244 68860 5588 68900
rect 9379 68860 9388 68900
rect 9428 68860 9964 68900
rect 10004 68860 10013 68900
rect 10627 68860 10636 68900
rect 10676 68860 10828 68900
rect 10868 68860 10877 68900
rect 3235 68859 3293 68860
rect 5548 68816 5588 68860
rect 21424 68816 21504 68836
rect 4919 68776 4928 68816
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 5296 68776 5305 68816
rect 5539 68776 5548 68816
rect 5588 68776 5932 68816
rect 5972 68776 5981 68816
rect 20039 68776 20048 68816
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20416 68776 20425 68816
rect 20524 68776 21504 68816
rect 2851 68732 2909 68733
rect 3331 68732 3389 68733
rect 13795 68732 13853 68733
rect 20524 68732 20564 68776
rect 21424 68756 21504 68776
rect 2851 68692 2860 68732
rect 2900 68692 3340 68732
rect 3380 68692 11212 68732
rect 11252 68692 11261 68732
rect 11395 68692 11404 68732
rect 11444 68692 12556 68732
rect 12596 68692 12605 68732
rect 13795 68692 13804 68732
rect 13844 68692 20564 68732
rect 2851 68691 2909 68692
rect 3331 68691 3389 68692
rect 13795 68691 13853 68692
rect 0 68648 80 68668
rect 0 68608 15436 68648
rect 15476 68608 15485 68648
rect 19363 68608 19372 68648
rect 19412 68608 19660 68648
rect 19700 68608 19709 68648
rect 0 68588 80 68608
rect 2851 68564 2909 68565
rect 11875 68564 11933 68565
rect 2851 68524 2860 68564
rect 2900 68524 3436 68564
rect 3476 68524 3485 68564
rect 11320 68524 11884 68564
rect 11924 68524 11933 68564
rect 13219 68524 13228 68564
rect 13268 68524 14572 68564
rect 14612 68524 14621 68564
rect 2851 68523 2909 68524
rect 6307 68480 6365 68481
rect 6883 68480 6941 68481
rect 11320 68480 11360 68524
rect 11875 68523 11933 68524
rect 20899 68480 20957 68481
rect 21424 68480 21504 68500
rect 1699 68440 1708 68480
rect 1748 68440 2572 68480
rect 2612 68440 2621 68480
rect 2755 68440 2764 68480
rect 2804 68440 3340 68480
rect 3380 68440 3389 68480
rect 6307 68440 6316 68480
rect 6356 68440 6508 68480
rect 6548 68440 6892 68480
rect 6932 68440 6941 68480
rect 7267 68440 7276 68480
rect 7316 68440 10156 68480
rect 10196 68440 11360 68480
rect 14179 68440 14188 68480
rect 14228 68440 17164 68480
rect 17204 68440 17644 68480
rect 17684 68440 17693 68480
rect 20899 68440 20908 68480
rect 20948 68440 21504 68480
rect 6307 68439 6365 68440
rect 6883 68439 6941 68440
rect 20899 68439 20957 68440
rect 21424 68420 21504 68440
rect 1219 68356 1228 68396
rect 1268 68356 1516 68396
rect 1556 68356 1804 68396
rect 1844 68356 1853 68396
rect 8611 68356 8620 68396
rect 8660 68356 9868 68396
rect 9908 68356 9917 68396
rect 14275 68356 14284 68396
rect 14324 68356 14956 68396
rect 14996 68356 15005 68396
rect 0 68312 80 68332
rect 0 68272 13268 68312
rect 13315 68272 13324 68312
rect 13364 68272 13804 68312
rect 13844 68272 13853 68312
rect 0 68252 80 68272
rect 13228 68228 13268 68272
rect 2083 68188 2092 68228
rect 2132 68188 2668 68228
rect 2708 68188 2717 68228
rect 7747 68188 7756 68228
rect 7796 68188 9388 68228
rect 9428 68188 9772 68228
rect 9812 68188 9821 68228
rect 12355 68188 12364 68228
rect 12404 68188 13036 68228
rect 13076 68188 13085 68228
rect 13228 68188 18412 68228
rect 18452 68188 18461 68228
rect 21424 68144 21504 68164
rect 20611 68104 20620 68144
rect 20660 68104 21504 68144
rect 21424 68084 21504 68104
rect 3679 68020 3688 68060
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 4056 68020 4065 68060
rect 7939 68020 7948 68060
rect 7988 68020 8908 68060
rect 8948 68020 8957 68060
rect 9091 68020 9100 68060
rect 9140 68020 9964 68060
rect 10004 68020 10013 68060
rect 18799 68020 18808 68060
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 19176 68020 19185 68060
rect 0 67976 80 67996
rect 259 67976 317 67977
rect 13507 67976 13565 67977
rect 13987 67976 14045 67977
rect 0 67936 268 67976
rect 308 67936 317 67976
rect 5731 67936 5740 67976
rect 5780 67936 9292 67976
rect 9332 67936 9341 67976
rect 12355 67936 12364 67976
rect 12404 67936 12556 67976
rect 12596 67936 12605 67976
rect 13507 67936 13516 67976
rect 13556 67936 13996 67976
rect 14036 67936 14045 67976
rect 0 67916 80 67936
rect 259 67935 317 67936
rect 13507 67935 13565 67936
rect 13987 67935 14045 67936
rect 2500 67852 14764 67892
rect 14804 67852 14813 67892
rect 2500 67808 2540 67852
rect 5155 67808 5213 67809
rect 21424 67808 21504 67828
rect 67 67768 76 67808
rect 116 67768 2540 67808
rect 4483 67768 4492 67808
rect 4532 67768 4684 67808
rect 4724 67768 4733 67808
rect 5070 67768 5164 67808
rect 5204 67768 5213 67808
rect 5635 67768 5644 67808
rect 5684 67768 6124 67808
rect 6164 67768 6173 67808
rect 7651 67768 7660 67808
rect 7700 67768 8812 67808
rect 8852 67768 9484 67808
rect 9524 67768 9533 67808
rect 20899 67768 20908 67808
rect 20948 67768 21504 67808
rect 5155 67767 5213 67768
rect 21424 67748 21504 67768
rect 9091 67724 9149 67725
rect 2275 67684 2284 67724
rect 2324 67684 8428 67724
rect 8468 67684 8477 67724
rect 8995 67684 9004 67724
rect 9044 67684 9100 67724
rect 9140 67684 9149 67724
rect 9091 67683 9149 67684
rect 11587 67724 11645 67725
rect 18211 67724 18269 67725
rect 11587 67684 11596 67724
rect 11636 67684 11980 67724
rect 12020 67684 12029 67724
rect 12355 67684 12364 67724
rect 12404 67684 13612 67724
rect 13652 67684 13661 67724
rect 14851 67684 14860 67724
rect 14900 67684 18220 67724
rect 18260 67684 18269 67724
rect 11587 67683 11645 67684
rect 18211 67683 18269 67684
rect 0 67641 80 67660
rect 0 67640 125 67641
rect 0 67600 76 67640
rect 116 67600 125 67640
rect 0 67599 125 67600
rect 1027 67640 1085 67641
rect 5923 67640 5981 67641
rect 15907 67640 15965 67641
rect 1027 67600 1036 67640
rect 1076 67600 4780 67640
rect 4820 67600 4829 67640
rect 5251 67600 5260 67640
rect 5300 67600 5932 67640
rect 5972 67600 5981 67640
rect 7356 67600 7365 67640
rect 7405 67600 7414 67640
rect 7459 67600 7468 67640
rect 7508 67600 9868 67640
rect 9908 67600 9917 67640
rect 10147 67600 10156 67640
rect 10196 67600 10348 67640
rect 10388 67600 10397 67640
rect 11320 67600 15916 67640
rect 15956 67600 15965 67640
rect 17443 67600 17452 67640
rect 17492 67600 18028 67640
rect 18068 67600 18077 67640
rect 1027 67599 1085 67600
rect 0 67580 80 67599
rect 4780 67556 4820 67600
rect 5923 67599 5981 67600
rect 6403 67556 6461 67557
rect 4780 67516 6412 67556
rect 6452 67516 6461 67556
rect 7372 67556 7412 67600
rect 11320 67556 11360 67600
rect 15907 67599 15965 67600
rect 7372 67516 7508 67556
rect 8419 67516 8428 67556
rect 8468 67516 9580 67556
rect 9620 67516 11360 67556
rect 6403 67515 6461 67516
rect 7075 67432 7084 67472
rect 7124 67432 7372 67472
rect 7412 67432 7421 67472
rect 2659 67388 2717 67389
rect 7468 67388 7508 67516
rect 21424 67472 21504 67492
rect 9187 67432 9196 67472
rect 9236 67432 13228 67472
rect 13268 67432 13277 67472
rect 20140 67432 21504 67472
rect 17347 67388 17405 67389
rect 20140 67388 20180 67432
rect 21424 67412 21504 67432
rect 2659 67348 2668 67388
rect 2708 67348 7412 67388
rect 7468 67348 9676 67388
rect 9716 67348 9725 67388
rect 17347 67348 17356 67388
rect 17396 67348 20180 67388
rect 2659 67347 2717 67348
rect 0 67304 80 67324
rect 7372 67304 7412 67348
rect 17347 67347 17405 67348
rect 11203 67304 11261 67305
rect 0 67264 76 67304
rect 116 67264 125 67304
rect 4919 67264 4928 67304
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 5296 67264 5305 67304
rect 7372 67264 11212 67304
rect 11252 67264 18604 67304
rect 18644 67264 18653 67304
rect 20039 67264 20048 67304
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20416 67264 20425 67304
rect 0 67244 80 67264
rect 11203 67263 11261 67264
rect 2947 67180 2956 67220
rect 2996 67180 5204 67220
rect 7363 67180 7372 67220
rect 7412 67180 9772 67220
rect 9812 67180 9821 67220
rect 15907 67180 15916 67220
rect 15956 67180 16108 67220
rect 16148 67180 16157 67220
rect 19651 67180 19660 67220
rect 19700 67180 19852 67220
rect 19892 67180 19901 67220
rect 1507 67136 1565 67137
rect 5164 67136 5204 67180
rect 7651 67136 7709 67137
rect 21424 67136 21504 67156
rect 1507 67096 1516 67136
rect 1556 67096 4204 67136
rect 4244 67096 4253 67136
rect 5155 67096 5164 67136
rect 5204 67096 7660 67136
rect 7700 67096 7709 67136
rect 8611 67096 8620 67136
rect 8660 67096 8812 67136
rect 8852 67096 8861 67136
rect 8908 67096 9868 67136
rect 9908 67096 9917 67136
rect 12931 67096 12940 67136
rect 12980 67096 18124 67136
rect 18164 67096 18173 67136
rect 20707 67096 20716 67136
rect 20756 67096 21504 67136
rect 1507 67095 1565 67096
rect 7651 67095 7709 67096
rect 8908 67052 8948 67096
rect 21424 67076 21504 67096
rect 16195 67052 16253 67053
rect 19651 67052 19709 67053
rect 8419 67012 8428 67052
rect 8468 67012 8948 67052
rect 9283 67012 9292 67052
rect 9332 67012 12748 67052
rect 12788 67012 12797 67052
rect 16099 67012 16108 67052
rect 16148 67012 16204 67052
rect 16244 67012 16253 67052
rect 19566 67012 19660 67052
rect 19700 67012 19709 67052
rect 16195 67011 16253 67012
rect 19651 67011 19709 67012
rect 0 66968 80 66988
rect 16675 66968 16733 66969
rect 0 66928 5396 66968
rect 6499 66928 6508 66968
rect 6548 66928 6844 66968
rect 6884 66928 9484 66968
rect 9524 66928 9533 66968
rect 12259 66928 12268 66968
rect 12308 66928 12556 66968
rect 12596 66928 12605 66968
rect 16590 66928 16684 66968
rect 16724 66928 16733 66968
rect 0 66908 80 66928
rect 5356 66884 5396 66928
rect 16675 66927 16733 66928
rect 5356 66844 7564 66884
rect 7604 66844 7613 66884
rect 8812 66844 9196 66884
rect 9236 66844 9245 66884
rect 9292 66844 10540 66884
rect 10580 66844 10589 66884
rect 11683 66844 11692 66884
rect 11732 66844 12076 66884
rect 12116 66844 12125 66884
rect 14860 66844 17068 66884
rect 17108 66844 18988 66884
rect 19028 66844 19037 66884
rect 835 66800 893 66801
rect 7267 66800 7325 66801
rect 8812 66800 8852 66844
rect 9292 66800 9332 66844
rect 14860 66800 14900 66844
rect 19747 66800 19805 66801
rect 21424 66800 21504 66820
rect 835 66760 844 66800
rect 884 66760 1132 66800
rect 1172 66760 1181 66800
rect 3523 66760 3532 66800
rect 3572 66760 4108 66800
rect 4148 66760 6508 66800
rect 6548 66760 6557 66800
rect 6604 66760 7276 66800
rect 7316 66760 7325 66800
rect 8131 66760 8140 66800
rect 8180 66760 8620 66800
rect 8660 66760 8669 66800
rect 8803 66760 8812 66800
rect 8852 66760 8861 66800
rect 9283 66760 9292 66800
rect 9332 66760 9341 66800
rect 9571 66760 9580 66800
rect 9620 66760 10636 66800
rect 10676 66760 10685 66800
rect 14851 66760 14860 66800
rect 14900 66760 14909 66800
rect 15427 66760 15436 66800
rect 15476 66760 16012 66800
rect 16052 66760 16061 66800
rect 19747 66760 19756 66800
rect 19796 66760 20524 66800
rect 20564 66760 20573 66800
rect 20995 66760 21004 66800
rect 21044 66760 21504 66800
rect 835 66759 893 66760
rect 1795 66716 1853 66717
rect 6604 66716 6644 66760
rect 7267 66759 7325 66760
rect 19747 66759 19805 66760
rect 21424 66740 21504 66760
rect 1795 66676 1804 66716
rect 1844 66676 6644 66716
rect 6691 66716 6749 66717
rect 8899 66716 8957 66717
rect 6691 66676 6700 66716
rect 6740 66676 8908 66716
rect 8948 66676 8957 66716
rect 1795 66675 1853 66676
rect 6691 66675 6749 66676
rect 8899 66675 8957 66676
rect 9091 66716 9149 66717
rect 9091 66676 9100 66716
rect 9140 66676 13228 66716
rect 13268 66676 13277 66716
rect 9091 66675 9149 66676
rect 0 66632 80 66652
rect 0 66592 8524 66632
rect 8564 66592 8573 66632
rect 10531 66592 10540 66632
rect 10580 66592 11116 66632
rect 11156 66592 11165 66632
rect 12643 66592 12652 66632
rect 12692 66592 13036 66632
rect 13076 66592 13085 66632
rect 0 66572 80 66592
rect 931 66508 940 66548
rect 980 66508 2380 66548
rect 2420 66508 2429 66548
rect 3679 66508 3688 66548
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 4056 66508 4065 66548
rect 6595 66508 6604 66548
rect 6644 66508 7084 66548
rect 7124 66508 7133 66548
rect 2275 66464 2333 66465
rect 7555 66464 7613 66465
rect 8323 66464 8381 66465
rect 1027 66424 1036 66464
rect 1076 66424 2284 66464
rect 2324 66424 2333 66464
rect 5731 66424 5740 66464
rect 5780 66424 6508 66464
rect 6548 66424 6557 66464
rect 7555 66424 7564 66464
rect 7604 66424 8332 66464
rect 8372 66424 8381 66464
rect 2275 66423 2333 66424
rect 7555 66423 7613 66424
rect 8323 66423 8381 66424
rect 7267 66380 7325 66381
rect 4579 66340 4588 66380
rect 4628 66340 6700 66380
rect 6740 66340 7276 66380
rect 7316 66340 7325 66380
rect 7267 66339 7325 66340
rect 0 66296 80 66316
rect 0 66256 76 66296
rect 116 66256 125 66296
rect 1411 66256 1420 66296
rect 1460 66256 8468 66296
rect 0 66236 80 66256
rect 1987 66172 1996 66212
rect 2036 66172 5068 66212
rect 5108 66172 6412 66212
rect 6452 66172 6461 66212
rect 7075 66172 7084 66212
rect 7124 66172 7164 66212
rect 3331 66128 3389 66129
rect 7084 66128 7124 66172
rect 3246 66088 3340 66128
rect 3380 66088 4204 66128
rect 4244 66088 4253 66128
rect 5923 66088 5932 66128
rect 5972 66088 7468 66128
rect 7508 66088 7517 66128
rect 3331 66087 3389 66088
rect 6979 66044 7037 66045
rect 2500 66004 6988 66044
rect 7028 66004 7037 66044
rect 8428 66044 8468 66256
rect 8524 66212 8564 66592
rect 10627 66508 10636 66548
rect 10676 66508 11020 66548
rect 11060 66508 12460 66548
rect 12500 66508 12509 66548
rect 18799 66508 18808 66548
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 19176 66508 19185 66548
rect 14179 66464 14237 66465
rect 21424 66464 21504 66484
rect 8611 66424 8620 66464
rect 8660 66424 11360 66464
rect 11320 66380 11360 66424
rect 14179 66424 14188 66464
rect 14228 66424 21504 66464
rect 14179 66423 14237 66424
rect 21424 66404 21504 66424
rect 18499 66380 18557 66381
rect 11320 66340 12364 66380
rect 12404 66340 12413 66380
rect 13219 66340 13228 66380
rect 13268 66340 18508 66380
rect 18548 66340 18557 66380
rect 18499 66339 18557 66340
rect 8995 66256 9004 66296
rect 9044 66256 9484 66296
rect 9524 66256 9533 66296
rect 17635 66256 17644 66296
rect 17684 66256 17932 66296
rect 17972 66256 17981 66296
rect 8524 66172 18220 66212
rect 18260 66172 18269 66212
rect 18979 66172 18988 66212
rect 19028 66172 19756 66212
rect 19796 66172 19805 66212
rect 21424 66128 21504 66148
rect 14083 66088 14092 66128
rect 14132 66088 15724 66128
rect 15764 66088 17164 66128
rect 17204 66088 19468 66128
rect 19508 66088 19517 66128
rect 20515 66088 20524 66128
rect 20564 66088 21504 66128
rect 21424 66068 21504 66088
rect 17059 66044 17117 66045
rect 8428 66004 10828 66044
rect 10868 66004 11212 66044
rect 11252 66004 11261 66044
rect 17059 66004 17068 66044
rect 17108 66004 20812 66044
rect 20852 66004 20861 66044
rect 0 65960 80 65980
rect 2500 65960 2540 66004
rect 6979 66003 7037 66004
rect 17059 66003 17117 66004
rect 8323 65960 8381 65961
rect 0 65920 2540 65960
rect 4483 65920 4492 65960
rect 4532 65920 4780 65960
rect 4820 65920 4829 65960
rect 5827 65920 5836 65960
rect 5876 65920 6508 65960
rect 6548 65920 6557 65960
rect 6979 65920 6988 65960
rect 7028 65920 7756 65960
rect 7796 65920 7805 65960
rect 8323 65920 8332 65960
rect 8372 65920 16684 65960
rect 16724 65920 18316 65960
rect 18356 65920 18365 65960
rect 0 65900 80 65920
rect 8323 65919 8381 65920
rect 7171 65876 7229 65877
rect 6787 65836 6796 65876
rect 6836 65836 7180 65876
rect 7220 65836 7229 65876
rect 14563 65836 14572 65876
rect 14612 65836 14860 65876
rect 14900 65836 14909 65876
rect 7171 65835 7229 65836
rect 7267 65792 7325 65793
rect 21424 65792 21504 65812
rect 4919 65752 4928 65792
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 5296 65752 5305 65792
rect 7182 65752 7276 65792
rect 7316 65752 7325 65792
rect 20039 65752 20048 65792
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20416 65752 20425 65792
rect 20803 65752 20812 65792
rect 20852 65752 21504 65792
rect 7267 65751 7325 65752
rect 21424 65732 21504 65752
rect 1411 65708 1469 65709
rect 1411 65668 1420 65708
rect 1460 65668 7756 65708
rect 7796 65668 7805 65708
rect 12355 65668 12364 65708
rect 12404 65668 12844 65708
rect 12884 65668 15532 65708
rect 15572 65668 19756 65708
rect 19796 65668 19805 65708
rect 1411 65667 1469 65668
rect 0 65624 80 65644
rect 3139 65624 3197 65625
rect 0 65584 1516 65624
rect 1556 65584 1565 65624
rect 2851 65584 2860 65624
rect 2900 65584 3148 65624
rect 3188 65584 3197 65624
rect 6307 65584 6316 65624
rect 6356 65584 6836 65624
rect 0 65564 80 65584
rect 3139 65583 3197 65584
rect 6796 65540 6836 65584
rect 6796 65500 9100 65540
rect 9140 65500 9149 65540
rect 15235 65500 15244 65540
rect 15284 65500 16012 65540
rect 16052 65500 16061 65540
rect 18115 65500 18124 65540
rect 18164 65500 19372 65540
rect 19412 65500 19421 65540
rect 3331 65456 3389 65457
rect 9379 65456 9437 65457
rect 11587 65456 11645 65457
rect 2563 65416 2572 65456
rect 2612 65416 2956 65456
rect 2996 65416 3005 65456
rect 3052 65416 3340 65456
rect 3380 65416 3436 65456
rect 3476 65416 3485 65456
rect 7075 65416 7084 65456
rect 7124 65416 7564 65456
rect 7604 65416 7613 65456
rect 9294 65416 9388 65456
rect 9428 65416 9437 65456
rect 11502 65416 11596 65456
rect 11636 65416 11645 65456
rect 1699 65372 1757 65373
rect 3052 65372 3092 65416
rect 3331 65415 3389 65416
rect 9379 65415 9437 65416
rect 11587 65415 11645 65416
rect 11971 65456 12029 65457
rect 15523 65456 15581 65457
rect 21424 65456 21504 65476
rect 11971 65416 11980 65456
rect 12020 65416 12172 65456
rect 12212 65416 12221 65456
rect 13900 65416 15340 65456
rect 15380 65416 15389 65456
rect 15523 65416 15532 65456
rect 15572 65416 21504 65456
rect 11971 65415 12029 65416
rect 13900 65372 13940 65416
rect 15523 65415 15581 65416
rect 21424 65396 21504 65416
rect 1699 65332 1708 65372
rect 1748 65332 3092 65372
rect 3331 65332 3340 65372
rect 3380 65332 3389 65372
rect 3523 65332 3532 65372
rect 3572 65332 5644 65372
rect 5684 65332 5693 65372
rect 6499 65332 6508 65372
rect 6548 65332 13940 65372
rect 14755 65332 14764 65372
rect 14804 65332 17548 65372
rect 17588 65332 17597 65372
rect 1699 65331 1757 65332
rect 0 65288 80 65308
rect 3340 65288 3380 65332
rect 16579 65288 16637 65289
rect 0 65248 3148 65288
rect 3188 65248 3380 65288
rect 5827 65248 5836 65288
rect 5876 65248 8044 65288
rect 8084 65248 8093 65288
rect 9667 65248 9676 65288
rect 9716 65248 10252 65288
rect 10292 65248 10301 65288
rect 10435 65248 10444 65288
rect 10484 65248 11308 65288
rect 11348 65248 11357 65288
rect 11596 65248 14380 65288
rect 14420 65248 14429 65288
rect 16579 65248 16588 65288
rect 16628 65248 16684 65288
rect 16724 65248 16733 65288
rect 0 65228 80 65248
rect 11596 65204 11636 65248
rect 16579 65247 16637 65248
rect 739 65164 748 65204
rect 788 65164 2540 65204
rect 2500 65120 2540 65164
rect 3628 65164 11636 65204
rect 13219 65204 13277 65205
rect 17155 65204 17213 65205
rect 13219 65164 13228 65204
rect 13268 65164 14764 65204
rect 14804 65164 14813 65204
rect 17155 65164 17164 65204
rect 17204 65164 19180 65204
rect 19220 65164 19229 65204
rect 3628 65120 3668 65164
rect 13219 65163 13277 65164
rect 17155 65163 17213 65164
rect 14467 65120 14525 65121
rect 21187 65120 21245 65121
rect 21424 65120 21504 65140
rect 2500 65080 3668 65120
rect 4675 65080 4684 65120
rect 4724 65080 7948 65120
rect 7988 65080 7997 65120
rect 9187 65080 9196 65120
rect 9236 65080 9580 65120
rect 9620 65080 9629 65120
rect 10627 65080 10636 65120
rect 10676 65080 10924 65120
rect 10964 65080 10973 65120
rect 14179 65080 14188 65120
rect 14228 65080 14476 65120
rect 14516 65080 14525 65120
rect 14947 65080 14956 65120
rect 14996 65080 17932 65120
rect 17972 65080 17981 65120
rect 21187 65080 21196 65120
rect 21236 65080 21504 65120
rect 14467 65079 14525 65080
rect 21187 65079 21245 65080
rect 21424 65060 21504 65080
rect 3679 64996 3688 65036
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 4056 64996 4065 65036
rect 5731 64996 5740 65036
rect 5780 64996 6220 65036
rect 6260 64996 6269 65036
rect 6403 64996 6412 65036
rect 6452 64996 9004 65036
rect 9044 64996 9053 65036
rect 13027 64996 13036 65036
rect 13076 64996 18412 65036
rect 18452 64996 18604 65036
rect 18644 64996 18653 65036
rect 18799 64996 18808 65036
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 19176 64996 19185 65036
rect 19276 64996 20620 65036
rect 20660 64996 20669 65036
rect 0 64952 80 64972
rect 14947 64952 15005 64953
rect 19276 64952 19316 64996
rect 0 64912 2188 64952
rect 2228 64912 2237 64952
rect 3235 64912 3244 64952
rect 3284 64912 3532 64952
rect 3572 64912 3581 64952
rect 6115 64912 6124 64952
rect 6164 64912 10540 64952
rect 10580 64912 10589 64952
rect 14947 64912 14956 64952
rect 14996 64912 19316 64952
rect 19372 64912 20524 64952
rect 20564 64912 20573 64952
rect 0 64892 80 64912
rect 14947 64911 15005 64912
rect 12547 64868 12605 64869
rect 19372 64868 19412 64912
rect 20515 64868 20573 64869
rect 12547 64828 12556 64868
rect 12596 64828 19412 64868
rect 19843 64828 19852 64868
rect 19892 64828 20524 64868
rect 20564 64828 20573 64868
rect 12547 64827 12605 64828
rect 20515 64827 20573 64828
rect 20995 64784 21053 64785
rect 21424 64784 21504 64804
rect 3139 64744 3148 64784
rect 3188 64744 6412 64784
rect 6452 64744 6461 64784
rect 7267 64744 7276 64784
rect 7316 64744 7325 64784
rect 20995 64744 21004 64784
rect 21044 64744 21504 64784
rect 2659 64700 2717 64701
rect 2574 64660 2668 64700
rect 2708 64660 2717 64700
rect 3331 64660 3340 64700
rect 3380 64660 3628 64700
rect 3668 64660 3677 64700
rect 5443 64660 5452 64700
rect 5492 64660 5932 64700
rect 5972 64660 5981 64700
rect 2659 64659 2717 64660
rect 0 64616 80 64636
rect 2179 64616 2237 64617
rect 0 64576 2188 64616
rect 2228 64576 2237 64616
rect 4483 64576 4492 64616
rect 4532 64576 6316 64616
rect 6356 64576 7084 64616
rect 7124 64576 7133 64616
rect 0 64556 80 64576
rect 2179 64575 2237 64576
rect 2467 64532 2525 64533
rect 7276 64532 7316 64744
rect 20995 64743 21053 64744
rect 21424 64724 21504 64744
rect 15715 64700 15773 64701
rect 8899 64660 8908 64700
rect 8948 64660 9580 64700
rect 9620 64660 9629 64700
rect 15715 64660 15724 64700
rect 15764 64660 21004 64700
rect 21044 64660 21053 64700
rect 15715 64659 15773 64660
rect 7555 64616 7613 64617
rect 19939 64616 19997 64617
rect 7555 64576 7564 64616
rect 7604 64576 7852 64616
rect 7892 64576 7901 64616
rect 8515 64576 8524 64616
rect 8564 64576 9292 64616
rect 9332 64576 9868 64616
rect 9908 64576 9917 64616
rect 10014 64576 10023 64616
rect 10063 64576 10348 64616
rect 10388 64576 10397 64616
rect 10819 64576 10828 64616
rect 10868 64576 13900 64616
rect 13940 64576 15724 64616
rect 15764 64576 16492 64616
rect 16532 64576 16541 64616
rect 19843 64576 19852 64616
rect 19892 64576 19948 64616
rect 19988 64576 19997 64616
rect 7555 64575 7613 64576
rect 19939 64575 19997 64576
rect 2467 64492 2476 64532
rect 2516 64492 3820 64532
rect 3860 64492 3869 64532
rect 5251 64492 5260 64532
rect 5300 64492 7660 64532
rect 7700 64492 7709 64532
rect 9091 64492 9100 64532
rect 9140 64492 10924 64532
rect 10964 64492 10973 64532
rect 11395 64492 11404 64532
rect 11444 64492 14476 64532
rect 14516 64492 18316 64532
rect 18356 64492 18365 64532
rect 2467 64491 2525 64492
rect 6307 64448 6365 64449
rect 8131 64448 8189 64449
rect 5443 64408 5452 64448
rect 5492 64408 5740 64448
rect 5780 64408 5789 64448
rect 6307 64408 6316 64448
rect 6356 64408 7508 64448
rect 7843 64408 7852 64448
rect 7892 64408 8140 64448
rect 8180 64408 8189 64448
rect 6307 64407 6365 64408
rect 1027 64364 1085 64365
rect 6019 64364 6077 64365
rect 6883 64364 6941 64365
rect 7468 64364 7508 64408
rect 8131 64407 8189 64408
rect 11011 64448 11069 64449
rect 13219 64448 13277 64449
rect 19267 64448 19325 64449
rect 21424 64448 21504 64468
rect 11011 64408 11020 64448
rect 11060 64408 13228 64448
rect 13268 64408 13277 64448
rect 15523 64408 15532 64448
rect 15572 64408 15916 64448
rect 15956 64408 15965 64448
rect 19182 64408 19276 64448
rect 19316 64408 19325 64448
rect 19651 64408 19660 64448
rect 19700 64408 20044 64448
rect 20084 64408 20093 64448
rect 20611 64408 20620 64448
rect 20660 64408 21504 64448
rect 11011 64407 11069 64408
rect 13219 64407 13277 64408
rect 19267 64407 19325 64408
rect 21424 64388 21504 64408
rect 16387 64364 16445 64365
rect 1027 64324 1036 64364
rect 1076 64324 4588 64364
rect 4628 64324 4637 64364
rect 6019 64324 6028 64364
rect 6068 64324 6220 64364
rect 6260 64324 6269 64364
rect 6403 64324 6412 64364
rect 6452 64324 6892 64364
rect 6932 64324 6941 64364
rect 7459 64324 7468 64364
rect 7508 64324 7517 64364
rect 9091 64324 9100 64364
rect 9140 64324 10252 64364
rect 10292 64324 10301 64364
rect 11779 64324 11788 64364
rect 11828 64324 12500 64364
rect 12739 64324 12748 64364
rect 12788 64324 16108 64364
rect 16148 64324 16396 64364
rect 16436 64324 16445 64364
rect 1027 64323 1085 64324
rect 6019 64323 6077 64324
rect 6883 64323 6941 64324
rect 0 64280 80 64300
rect 8515 64280 8573 64281
rect 0 64240 460 64280
rect 500 64240 509 64280
rect 4919 64240 4928 64280
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 5296 64240 5305 64280
rect 7267 64240 7276 64280
rect 7316 64240 7564 64280
rect 7604 64240 7613 64280
rect 8419 64240 8428 64280
rect 8468 64240 8524 64280
rect 8564 64240 8573 64280
rect 0 64220 80 64240
rect 8515 64239 8573 64240
rect 9091 64280 9149 64281
rect 11491 64280 11549 64281
rect 12460 64280 12500 64324
rect 16387 64323 16445 64324
rect 15811 64280 15869 64281
rect 9091 64240 9100 64280
rect 9140 64240 10060 64280
rect 10100 64240 10109 64280
rect 11406 64240 11500 64280
rect 11540 64240 11549 64280
rect 12420 64240 12460 64280
rect 12500 64240 12509 64280
rect 12643 64240 12652 64280
rect 12692 64240 12844 64280
rect 12884 64240 12893 64280
rect 15726 64240 15820 64280
rect 15860 64240 15869 64280
rect 20039 64240 20048 64280
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20416 64240 20425 64280
rect 9091 64239 9149 64240
rect 11491 64239 11549 64240
rect 15811 64239 15869 64240
rect 17251 64196 17309 64197
rect 3811 64156 3820 64196
rect 3860 64156 9388 64196
rect 9428 64156 11020 64196
rect 11060 64156 11069 64196
rect 17251 64156 17260 64196
rect 17300 64156 20812 64196
rect 20852 64156 20861 64196
rect 17251 64155 17309 64156
rect 17923 64112 17981 64113
rect 21424 64112 21504 64132
rect 8227 64072 8236 64112
rect 8276 64072 9772 64112
rect 9812 64072 9821 64112
rect 11491 64072 11500 64112
rect 11540 64072 12076 64112
rect 12116 64072 12125 64112
rect 12355 64072 12364 64112
rect 12404 64072 16300 64112
rect 16340 64072 16349 64112
rect 17923 64072 17932 64112
rect 17972 64072 21504 64112
rect 17923 64071 17981 64072
rect 21424 64052 21504 64072
rect 1411 63988 1420 64028
rect 1460 63988 1996 64028
rect 2036 63988 2045 64028
rect 2659 63988 2668 64028
rect 2708 63988 5068 64028
rect 5108 63988 5117 64028
rect 12835 63988 12844 64028
rect 12884 63988 13708 64028
rect 13748 63988 13757 64028
rect 0 63944 80 63964
rect 5827 63944 5885 63945
rect 17539 63944 17597 63945
rect 0 63904 2572 63944
rect 2612 63904 2621 63944
rect 5742 63904 5836 63944
rect 5876 63904 5885 63944
rect 6019 63904 6028 63944
rect 6068 63904 8044 63944
rect 8084 63904 8093 63944
rect 8323 63904 8332 63944
rect 8372 63904 8716 63944
rect 8756 63904 9388 63944
rect 9428 63904 9437 63944
rect 10147 63904 10156 63944
rect 10196 63904 10444 63944
rect 10484 63904 10493 63944
rect 11587 63904 11596 63944
rect 11636 63904 13516 63944
rect 13556 63904 14668 63944
rect 14708 63904 14717 63944
rect 17539 63904 17548 63944
rect 17588 63904 20180 63944
rect 0 63884 80 63904
rect 2500 63860 2540 63904
rect 5827 63903 5885 63904
rect 17539 63903 17597 63904
rect 10531 63860 10589 63861
rect 20140 63860 20180 63904
rect 2500 63820 8428 63860
rect 8468 63820 8477 63860
rect 10531 63820 10540 63860
rect 10580 63820 16300 63860
rect 16340 63820 19372 63860
rect 19412 63820 19421 63860
rect 20140 63820 20908 63860
rect 20948 63820 20957 63860
rect 10531 63819 10589 63820
rect 10540 63776 10580 63819
rect 14275 63776 14333 63777
rect 21424 63776 21504 63796
rect 1411 63736 1420 63776
rect 1460 63736 1612 63776
rect 1652 63736 1661 63776
rect 4579 63736 4588 63776
rect 4628 63736 5932 63776
rect 5972 63736 5981 63776
rect 7747 63736 7756 63776
rect 7796 63736 10580 63776
rect 11011 63736 11020 63776
rect 11060 63736 12748 63776
rect 12788 63736 12797 63776
rect 14275 63736 14284 63776
rect 14324 63736 14476 63776
rect 14516 63736 14525 63776
rect 15724 63736 20716 63776
rect 20756 63736 20765 63776
rect 21187 63736 21196 63776
rect 21236 63736 21504 63776
rect 14275 63735 14333 63736
rect 1315 63652 1324 63692
rect 1364 63652 3820 63692
rect 3860 63652 3869 63692
rect 4771 63652 4780 63692
rect 4820 63652 5260 63692
rect 5300 63652 5309 63692
rect 5443 63652 5452 63692
rect 5492 63652 7276 63692
rect 7316 63652 9964 63692
rect 10004 63652 10828 63692
rect 10868 63652 10877 63692
rect 13315 63652 13324 63692
rect 13364 63652 13708 63692
rect 13748 63652 13757 63692
rect 0 63608 80 63628
rect 0 63568 4492 63608
rect 4532 63568 4541 63608
rect 0 63548 80 63568
rect 7468 63524 7508 63652
rect 10819 63608 10877 63609
rect 15724 63608 15764 63736
rect 21424 63716 21504 63736
rect 19939 63652 19948 63692
rect 19988 63652 20812 63692
rect 20852 63652 20861 63692
rect 8515 63568 8524 63608
rect 8564 63568 10772 63608
rect 8323 63524 8381 63525
rect 8515 63524 8573 63525
rect 10732 63524 10772 63568
rect 10819 63568 10828 63608
rect 10868 63568 15764 63608
rect 18211 63608 18269 63609
rect 18211 63568 18220 63608
rect 18260 63568 18604 63608
rect 18644 63568 18653 63608
rect 10819 63567 10877 63568
rect 18211 63567 18269 63568
rect 3679 63484 3688 63524
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 4056 63484 4065 63524
rect 7459 63484 7468 63524
rect 7508 63484 7517 63524
rect 8323 63484 8332 63524
rect 8372 63484 8524 63524
rect 8564 63484 10676 63524
rect 10732 63484 11596 63524
rect 11636 63484 11645 63524
rect 18307 63484 18316 63524
rect 18356 63484 18700 63524
rect 18740 63484 18749 63524
rect 18799 63484 18808 63524
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 19176 63484 19185 63524
rect 8323 63483 8381 63484
rect 8515 63483 8573 63484
rect 835 63440 893 63441
rect 10636 63440 10676 63484
rect 19267 63440 19325 63441
rect 21424 63440 21504 63460
rect 835 63400 844 63440
rect 884 63400 6988 63440
rect 7028 63400 7037 63440
rect 9964 63400 10580 63440
rect 10636 63400 14900 63440
rect 17731 63400 17740 63440
rect 17780 63400 17932 63440
rect 17972 63400 17981 63440
rect 19267 63400 19276 63440
rect 19316 63400 21504 63440
rect 835 63399 893 63400
rect 0 63272 80 63292
rect 451 63272 509 63273
rect 0 63232 460 63272
rect 500 63232 509 63272
rect 0 63212 80 63232
rect 451 63231 509 63232
rect 1411 63272 1469 63273
rect 1987 63272 2045 63273
rect 9379 63272 9437 63273
rect 1411 63232 1420 63272
rect 1460 63232 1516 63272
rect 1556 63232 1565 63272
rect 1891 63232 1900 63272
rect 1940 63232 1996 63272
rect 2036 63232 2045 63272
rect 2851 63232 2860 63272
rect 2900 63232 4684 63272
rect 4724 63232 4733 63272
rect 6403 63232 6412 63272
rect 6452 63232 6892 63272
rect 6932 63232 6941 63272
rect 9379 63232 9388 63272
rect 9428 63232 9484 63272
rect 9524 63232 9533 63272
rect 1411 63231 1469 63232
rect 1987 63231 2045 63232
rect 9379 63231 9437 63232
rect 3427 63188 3485 63189
rect 8515 63188 8573 63189
rect 9964 63188 10004 63400
rect 10339 63356 10397 63357
rect 10254 63316 10348 63356
rect 10388 63316 10397 63356
rect 10540 63356 10580 63400
rect 14860 63356 14900 63400
rect 19267 63399 19325 63400
rect 21424 63380 21504 63400
rect 10540 63316 11884 63356
rect 11924 63316 11933 63356
rect 14851 63316 14860 63356
rect 14900 63316 19756 63356
rect 19796 63316 19805 63356
rect 10339 63315 10397 63316
rect 10243 63272 10301 63273
rect 10158 63232 10252 63272
rect 10292 63232 10301 63272
rect 10243 63231 10301 63232
rect 11320 63232 12364 63272
rect 12404 63232 12413 63272
rect 15523 63232 15532 63272
rect 15572 63232 15724 63272
rect 15764 63232 15773 63272
rect 16867 63232 16876 63272
rect 16916 63232 18412 63272
rect 18452 63232 18461 63272
rect 11320 63188 11360 63232
rect 1699 63148 1708 63188
rect 1748 63148 2572 63188
rect 2612 63148 2621 63188
rect 3427 63148 3436 63188
rect 3476 63148 6508 63188
rect 6548 63148 6557 63188
rect 8515 63148 8524 63188
rect 8564 63148 9868 63188
rect 9908 63148 10004 63188
rect 10339 63148 10348 63188
rect 10388 63148 10732 63188
rect 10772 63148 11360 63188
rect 18019 63148 18028 63188
rect 18068 63148 18220 63188
rect 18260 63148 18269 63188
rect 3427 63147 3485 63148
rect 8515 63147 8573 63148
rect 4387 63104 4445 63105
rect 6019 63104 6077 63105
rect 18499 63104 18557 63105
rect 21424 63104 21504 63124
rect 4195 63064 4204 63104
rect 4244 63064 4396 63104
rect 4436 63064 4445 63104
rect 5059 63064 5068 63104
rect 5108 63064 6028 63104
rect 6068 63064 6077 63104
rect 7651 63064 7660 63104
rect 7700 63064 9292 63104
rect 9332 63064 9341 63104
rect 9763 63064 9772 63104
rect 9812 63064 10156 63104
rect 10196 63064 10205 63104
rect 10627 63064 10636 63104
rect 10676 63064 11308 63104
rect 11348 63064 11357 63104
rect 11875 63064 11884 63104
rect 11924 63064 14092 63104
rect 14132 63064 14141 63104
rect 15715 63064 15724 63104
rect 15764 63064 16204 63104
rect 16244 63064 16253 63104
rect 18499 63064 18508 63104
rect 18548 63064 18988 63104
rect 19028 63064 19037 63104
rect 20995 63064 21004 63104
rect 21044 63064 21504 63104
rect 4387 63063 4445 63064
rect 6019 63063 6077 63064
rect 9292 63020 9332 63064
rect 18499 63063 18557 63064
rect 21424 63044 21504 63064
rect 16963 63020 17021 63021
rect 931 62980 940 63020
rect 980 62980 2284 63020
rect 2324 62980 2333 63020
rect 2659 62980 2668 63020
rect 2708 62980 3148 63020
rect 3188 62980 3197 63020
rect 4291 62980 4300 63020
rect 4340 62980 6604 63020
rect 6644 62980 6653 63020
rect 8419 62980 8428 63020
rect 8468 62980 8812 63020
rect 8852 62980 8861 63020
rect 9292 62980 10252 63020
rect 10292 62980 10301 63020
rect 12451 62980 12460 63020
rect 12500 62980 13996 63020
rect 14036 62980 15916 63020
rect 15956 62980 15965 63020
rect 16483 62980 16492 63020
rect 16532 62980 16972 63020
rect 17012 62980 17021 63020
rect 16963 62979 17021 62980
rect 0 62936 80 62956
rect 7747 62936 7805 62937
rect 0 62896 212 62936
rect 0 62876 80 62896
rect 172 62768 212 62896
rect 1420 62896 7756 62936
rect 7796 62896 7805 62936
rect 451 62852 509 62853
rect 1420 62852 1460 62896
rect 7747 62895 7805 62896
rect 451 62812 460 62852
rect 500 62812 1460 62852
rect 1507 62812 1516 62852
rect 1556 62812 2188 62852
rect 2228 62812 8716 62852
rect 8756 62812 8765 62852
rect 11875 62812 11884 62852
rect 11924 62812 12076 62852
rect 12116 62812 12125 62852
rect 451 62811 509 62812
rect 5347 62768 5405 62769
rect 21424 62768 21504 62788
rect 172 62728 1420 62768
rect 1460 62728 1469 62768
rect 4919 62728 4928 62768
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 5296 62728 5305 62768
rect 5347 62728 5356 62768
rect 5396 62728 5452 62768
rect 5492 62728 5501 62768
rect 5731 62728 5740 62768
rect 5780 62728 6316 62768
rect 6356 62728 6365 62768
rect 11491 62728 11500 62768
rect 11540 62728 12172 62768
rect 12212 62728 12221 62768
rect 20039 62728 20048 62768
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20416 62728 20425 62768
rect 20515 62728 20524 62768
rect 20564 62728 21504 62768
rect 5347 62727 5405 62728
rect 21424 62708 21504 62728
rect 4291 62684 4349 62685
rect 5827 62684 5885 62685
rect 9955 62684 10013 62685
rect 1228 62644 2956 62684
rect 2996 62644 3005 62684
rect 4291 62644 4300 62684
rect 4340 62644 4396 62684
rect 4436 62644 4445 62684
rect 5742 62644 5836 62684
rect 5876 62644 5885 62684
rect 9475 62644 9484 62684
rect 9524 62644 9964 62684
rect 10004 62644 10013 62684
rect 0 62600 80 62620
rect 1228 62600 1268 62644
rect 4291 62643 4349 62644
rect 5827 62643 5885 62644
rect 9955 62643 10013 62644
rect 10060 62644 19660 62684
rect 19700 62644 19709 62684
rect 8611 62600 8669 62601
rect 10060 62600 10100 62644
rect 14563 62600 14621 62601
rect 16867 62600 16925 62601
rect 0 62560 1268 62600
rect 2467 62560 2476 62600
rect 2516 62560 5068 62600
rect 5108 62560 5117 62600
rect 7555 62560 7564 62600
rect 7604 62560 7756 62600
rect 7796 62560 7805 62600
rect 8611 62560 8620 62600
rect 8660 62560 10100 62600
rect 10819 62560 10828 62600
rect 10868 62560 11116 62600
rect 11156 62560 11165 62600
rect 14563 62560 14572 62600
rect 14612 62560 16108 62600
rect 16148 62560 16157 62600
rect 16782 62560 16876 62600
rect 16916 62560 16925 62600
rect 0 62540 80 62560
rect 8611 62559 8669 62560
rect 14563 62559 14621 62560
rect 16867 62559 16925 62560
rect 1699 62516 1757 62517
rect 9955 62516 10013 62517
rect 1699 62476 1708 62516
rect 1748 62476 2540 62516
rect 3043 62476 3052 62516
rect 3092 62476 3340 62516
rect 3380 62476 3389 62516
rect 4003 62476 4012 62516
rect 4052 62476 8620 62516
rect 8660 62476 8669 62516
rect 8995 62476 9004 62516
rect 9044 62476 9292 62516
rect 9332 62476 9341 62516
rect 9870 62476 9964 62516
rect 10004 62476 10013 62516
rect 1699 62475 1757 62476
rect 2500 62432 2540 62476
rect 9955 62475 10013 62476
rect 10060 62476 15532 62516
rect 15572 62476 15581 62516
rect 20140 62476 21292 62516
rect 21332 62476 21341 62516
rect 10060 62432 10100 62476
rect 2500 62392 10100 62432
rect 10156 62392 19892 62432
rect 10156 62348 10196 62392
rect 15331 62348 15389 62349
rect 19852 62348 19892 62392
rect 2563 62308 2572 62348
rect 2612 62308 3052 62348
rect 3092 62308 3101 62348
rect 3811 62308 3820 62348
rect 3860 62308 7084 62348
rect 7124 62308 7133 62348
rect 7267 62308 7276 62348
rect 7316 62308 10196 62348
rect 10243 62308 10252 62348
rect 10292 62308 10444 62348
rect 10484 62308 12364 62348
rect 12404 62308 15340 62348
rect 15380 62308 15389 62348
rect 19843 62308 19852 62348
rect 19892 62308 19901 62348
rect 15331 62307 15389 62308
rect 0 62264 80 62284
rect 20140 62264 20180 62476
rect 20227 62432 20285 62433
rect 21424 62432 21504 62452
rect 20227 62392 20236 62432
rect 20276 62392 21504 62432
rect 20227 62391 20285 62392
rect 21424 62372 21504 62392
rect 0 62224 1228 62264
rect 1268 62224 1277 62264
rect 3907 62224 3916 62264
rect 3956 62224 4108 62264
rect 4148 62224 15340 62264
rect 15380 62224 15389 62264
rect 15436 62224 20180 62264
rect 0 62204 80 62224
rect 15436 62180 15476 62224
rect 2755 62140 2764 62180
rect 2804 62140 4492 62180
rect 4532 62140 4541 62180
rect 6499 62140 6508 62180
rect 6548 62140 7276 62180
rect 7316 62140 7325 62180
rect 7939 62140 7948 62180
rect 7988 62140 8236 62180
rect 8276 62140 8285 62180
rect 12163 62140 12172 62180
rect 12212 62140 12556 62180
rect 12596 62140 12605 62180
rect 13507 62140 13516 62180
rect 13556 62140 15476 62180
rect 21424 62096 21504 62116
rect 3427 62056 3436 62096
rect 3476 62056 4588 62096
rect 4628 62056 4637 62096
rect 7075 62056 7084 62096
rect 7124 62056 12940 62096
rect 12980 62056 12989 62096
rect 13699 62056 13708 62096
rect 13748 62056 21504 62096
rect 21424 62036 21504 62056
rect 3235 62012 3293 62013
rect 3235 61972 3244 62012
rect 3284 61972 3532 62012
rect 3572 61972 3581 62012
rect 3679 61972 3688 62012
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 4056 61972 4065 62012
rect 9667 61972 9676 62012
rect 9716 61972 16780 62012
rect 16820 61972 16829 62012
rect 18799 61972 18808 62012
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 19176 61972 19185 62012
rect 3235 61971 3293 61972
rect 0 61928 80 61948
rect 3427 61928 3485 61929
rect 4387 61928 4445 61929
rect 11203 61928 11261 61929
rect 0 61888 172 61928
rect 212 61888 221 61928
rect 3427 61888 3436 61928
rect 3476 61888 4204 61928
rect 4244 61888 4253 61928
rect 4302 61888 4396 61928
rect 4436 61888 4445 61928
rect 10723 61888 10732 61928
rect 10772 61888 11212 61928
rect 11252 61888 11261 61928
rect 13315 61888 13324 61928
rect 13364 61888 20524 61928
rect 20564 61888 20573 61928
rect 0 61868 80 61888
rect 3427 61887 3485 61888
rect 4387 61887 4445 61888
rect 11203 61887 11261 61888
rect 4579 61844 4637 61845
rect 17635 61844 17693 61845
rect 4579 61804 4588 61844
rect 4628 61804 13036 61844
rect 13076 61804 13085 61844
rect 13891 61804 13900 61844
rect 13940 61804 14476 61844
rect 14516 61804 14525 61844
rect 16195 61804 16204 61844
rect 16244 61804 17644 61844
rect 17684 61804 17693 61844
rect 4579 61803 4637 61804
rect 17635 61803 17693 61804
rect 1123 61760 1181 61761
rect 4291 61760 4349 61761
rect 11491 61760 11549 61761
rect 11971 61760 12029 61761
rect 21424 61760 21504 61780
rect 1027 61720 1036 61760
rect 1076 61720 1132 61760
rect 1172 61720 1181 61760
rect 4206 61720 4300 61760
rect 4340 61720 4349 61760
rect 11107 61720 11116 61760
rect 11156 61720 11252 61760
rect 11299 61720 11308 61760
rect 11348 61720 11500 61760
rect 11540 61720 11549 61760
rect 11886 61720 11980 61760
rect 12020 61720 12029 61760
rect 16099 61720 16108 61760
rect 16148 61720 21504 61760
rect 1123 61719 1181 61720
rect 4291 61719 4349 61720
rect 643 61676 701 61677
rect 4195 61676 4253 61677
rect 11212 61676 11252 61720
rect 11491 61719 11549 61720
rect 11971 61719 12029 61720
rect 21424 61700 21504 61720
rect 643 61636 652 61676
rect 692 61636 4204 61676
rect 4244 61636 4253 61676
rect 9571 61636 9580 61676
rect 9620 61636 10156 61676
rect 10196 61636 11156 61676
rect 11212 61636 14860 61676
rect 14900 61636 14909 61676
rect 16291 61636 16300 61676
rect 16340 61636 19756 61676
rect 19796 61636 19805 61676
rect 643 61635 701 61636
rect 4195 61635 4253 61636
rect 0 61592 80 61612
rect 2755 61592 2813 61593
rect 0 61552 2764 61592
rect 2804 61552 2813 61592
rect 0 61532 80 61552
rect 2755 61551 2813 61552
rect 3235 61592 3293 61593
rect 11116 61592 11156 61636
rect 19459 61592 19517 61593
rect 3235 61552 3244 61592
rect 3284 61552 3628 61592
rect 3668 61552 3677 61592
rect 6499 61552 6508 61592
rect 6548 61552 6892 61592
rect 6932 61552 6941 61592
rect 7459 61552 7468 61592
rect 7508 61552 7660 61592
rect 7700 61552 7709 61592
rect 8803 61552 8812 61592
rect 8852 61552 11020 61592
rect 11060 61552 11069 61592
rect 11116 61552 12268 61592
rect 12308 61552 16684 61592
rect 16724 61552 16733 61592
rect 17539 61552 17548 61592
rect 17588 61552 17597 61592
rect 19459 61552 19468 61592
rect 19508 61552 19564 61592
rect 19604 61552 19613 61592
rect 3235 61551 3293 61552
rect 15619 61508 15677 61509
rect 8899 61468 8908 61508
rect 8948 61468 9388 61508
rect 9428 61468 11116 61508
rect 11156 61468 11165 61508
rect 13987 61468 13996 61508
rect 14036 61468 14476 61508
rect 14516 61468 14525 61508
rect 15139 61468 15148 61508
rect 15188 61468 15628 61508
rect 15668 61468 15677 61508
rect 17548 61508 17588 61552
rect 19459 61551 19517 61552
rect 19843 61508 19901 61509
rect 17548 61468 18220 61508
rect 18260 61468 19372 61508
rect 19412 61468 19421 61508
rect 19843 61468 19852 61508
rect 19892 61468 20044 61508
rect 20084 61468 20093 61508
rect 15619 61467 15677 61468
rect 10627 61424 10685 61425
rect 17620 61424 17660 61468
rect 19843 61467 19901 61468
rect 20707 61424 20765 61425
rect 21424 61424 21504 61444
rect 3331 61384 3340 61424
rect 3380 61384 3628 61424
rect 3668 61384 4588 61424
rect 4628 61384 6124 61424
rect 6164 61384 6173 61424
rect 8812 61384 10636 61424
rect 10676 61384 10685 61424
rect 11011 61384 11020 61424
rect 11060 61384 11788 61424
rect 11828 61384 15916 61424
rect 15956 61384 15965 61424
rect 17443 61384 17452 61424
rect 17492 61384 17660 61424
rect 19939 61384 19948 61424
rect 19988 61384 20716 61424
rect 20756 61384 20765 61424
rect 8812 61340 8852 61384
rect 10627 61383 10685 61384
rect 20707 61383 20765 61384
rect 20812 61384 21504 61424
rect 643 61300 652 61340
rect 692 61300 8852 61340
rect 10147 61300 10156 61340
rect 10196 61300 16300 61340
rect 16340 61300 16349 61340
rect 0 61256 80 61276
rect 13219 61256 13277 61257
rect 0 61216 1516 61256
rect 1556 61216 1565 61256
rect 4919 61216 4928 61256
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 5296 61216 5305 61256
rect 6019 61216 6028 61256
rect 6068 61216 10868 61256
rect 0 61196 80 61216
rect 10828 61172 10868 61216
rect 11320 61216 11404 61256
rect 11444 61216 11453 61256
rect 12163 61216 12172 61256
rect 12212 61216 12460 61256
rect 12500 61216 12509 61256
rect 13219 61216 13228 61256
rect 13268 61216 13420 61256
rect 13460 61216 15340 61256
rect 15380 61216 15389 61256
rect 20039 61216 20048 61256
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20416 61216 20425 61256
rect 11320 61172 11360 61216
rect 13219 61215 13277 61216
rect 14851 61172 14909 61173
rect 20812 61172 20852 61384
rect 21424 61364 21504 61384
rect 3139 61132 3148 61172
rect 3188 61132 4780 61172
rect 4820 61132 7660 61172
rect 7700 61132 7709 61172
rect 10060 61132 10444 61172
rect 10484 61132 10493 61172
rect 10828 61132 11360 61172
rect 11779 61132 11788 61172
rect 11828 61132 12844 61172
rect 12884 61132 12893 61172
rect 14766 61132 14860 61172
rect 14900 61132 14909 61172
rect 15043 61132 15052 61172
rect 15092 61132 20852 61172
rect 6019 61088 6077 61089
rect 7555 61088 7613 61089
rect 172 61048 3244 61088
rect 3284 61048 3293 61088
rect 6019 61048 6028 61088
rect 6068 61048 6412 61088
rect 6452 61048 7564 61088
rect 7604 61048 7613 61088
rect 7747 61048 7756 61088
rect 7796 61048 8140 61088
rect 8180 61048 9772 61088
rect 9812 61048 9821 61088
rect 0 60920 80 60940
rect 172 60920 212 61048
rect 6019 61047 6077 61048
rect 7555 61047 7613 61048
rect 9187 61004 9245 61005
rect 835 60964 844 61004
rect 884 60964 9196 61004
rect 9236 60964 9245 61004
rect 9187 60963 9245 60964
rect 7555 60920 7613 60921
rect 8131 60920 8189 60921
rect 10060 60920 10100 61132
rect 14851 61131 14909 61132
rect 21424 61088 21504 61108
rect 12739 61048 12748 61088
rect 12788 61048 14228 61088
rect 14947 61048 14956 61088
rect 14996 61048 15436 61088
rect 15476 61048 15485 61088
rect 19747 61048 19756 61088
rect 19796 61048 21504 61088
rect 14188 61004 14228 61048
rect 21424 61028 21504 61048
rect 10243 60964 10252 61004
rect 10292 60964 10540 61004
rect 10580 60964 10589 61004
rect 10636 60964 14092 61004
rect 14132 60964 14141 61004
rect 14188 60964 16972 61004
rect 17012 60964 17021 61004
rect 0 60880 212 60920
rect 1603 60880 1612 60920
rect 1652 60880 1900 60920
rect 1940 60880 1949 60920
rect 2500 60880 3532 60920
rect 3572 60880 5164 60920
rect 5204 60880 7180 60920
rect 7220 60880 7229 60920
rect 7555 60880 7564 60920
rect 7604 60880 8140 60920
rect 8180 60880 8524 60920
rect 8564 60880 8573 60920
rect 8899 60880 8908 60920
rect 8948 60880 8957 60920
rect 10051 60880 10060 60920
rect 10100 60880 10109 60920
rect 0 60860 80 60880
rect 2500 60836 2540 60880
rect 7555 60879 7613 60880
rect 8131 60879 8189 60880
rect 8908 60836 8948 60880
rect 10636 60836 10676 60964
rect 14563 60880 14572 60920
rect 14612 60880 15532 60920
rect 15572 60880 15581 60920
rect 17347 60880 17356 60920
rect 17396 60880 17548 60920
rect 17588 60880 19276 60920
rect 19316 60880 19325 60920
rect 1315 60796 1324 60836
rect 1364 60796 2540 60836
rect 6883 60796 6892 60836
rect 6932 60796 7468 60836
rect 7508 60796 7517 60836
rect 8908 60796 9868 60836
rect 9908 60796 10676 60836
rect 13027 60796 13036 60836
rect 13076 60796 14476 60836
rect 14516 60796 14525 60836
rect 18499 60796 18508 60836
rect 18548 60796 20044 60836
rect 20084 60796 20093 60836
rect 21424 60752 21504 60772
rect 7171 60712 7180 60752
rect 7220 60712 13612 60752
rect 13652 60712 13661 60752
rect 14083 60712 14092 60752
rect 14132 60712 16244 60752
rect 17155 60712 17164 60752
rect 17204 60712 21504 60752
rect 6979 60668 7037 60669
rect 16204 60668 16244 60712
rect 21424 60692 21504 60712
rect 3043 60628 3052 60668
rect 3092 60628 4300 60668
rect 4340 60628 4349 60668
rect 4963 60628 4972 60668
rect 5012 60628 6316 60668
rect 6356 60628 6365 60668
rect 6979 60628 6988 60668
rect 7028 60628 11020 60668
rect 11060 60628 11069 60668
rect 11116 60628 12788 60668
rect 13027 60628 13036 60668
rect 13076 60628 14996 60668
rect 16195 60628 16204 60668
rect 16244 60628 16253 60668
rect 20227 60628 20236 60668
rect 20276 60628 20716 60668
rect 20756 60628 20765 60668
rect 6979 60627 7037 60628
rect 0 60584 80 60604
rect 7555 60584 7613 60585
rect 11116 60584 11156 60628
rect 0 60544 268 60584
rect 308 60544 317 60584
rect 1699 60544 1708 60584
rect 1748 60544 5492 60584
rect 0 60524 80 60544
rect 5452 60500 5492 60544
rect 7555 60544 7564 60584
rect 7604 60544 7852 60584
rect 7892 60544 7901 60584
rect 9763 60544 9772 60584
rect 9812 60544 11156 60584
rect 12748 60584 12788 60628
rect 14956 60584 14996 60628
rect 12748 60544 13228 60584
rect 13268 60544 14900 60584
rect 14956 60544 15017 60584
rect 15057 60544 15244 60584
rect 15284 60544 15293 60584
rect 7555 60543 7613 60544
rect 13315 60500 13373 60501
rect 14860 60500 14900 60544
rect 3331 60460 3340 60500
rect 3380 60460 3532 60500
rect 3572 60460 3581 60500
rect 3679 60460 3688 60500
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 4056 60460 4065 60500
rect 5452 60460 8332 60500
rect 8372 60460 8381 60500
rect 8515 60460 8524 60500
rect 8564 60460 13268 60500
rect 13228 60416 13268 60460
rect 13315 60460 13324 60500
rect 13364 60460 13804 60500
rect 13844 60460 13853 60500
rect 14083 60460 14092 60500
rect 14132 60460 14764 60500
rect 14804 60460 14813 60500
rect 14860 60460 16876 60500
rect 16916 60460 16925 60500
rect 18799 60460 18808 60500
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 19176 60460 19185 60500
rect 13315 60459 13373 60460
rect 14851 60416 14909 60417
rect 21424 60416 21504 60436
rect 2083 60376 2092 60416
rect 2132 60376 12268 60416
rect 12308 60376 12317 60416
rect 13228 60376 13900 60416
rect 13940 60376 14476 60416
rect 14516 60376 14525 60416
rect 14851 60376 14860 60416
rect 14900 60376 14956 60416
rect 14996 60376 15005 60416
rect 17539 60376 17548 60416
rect 17588 60376 21504 60416
rect 14851 60375 14909 60376
rect 21424 60356 21504 60376
rect 13219 60332 13277 60333
rect 2947 60292 2956 60332
rect 2996 60292 4780 60332
rect 4820 60292 4829 60332
rect 4876 60292 12500 60332
rect 12643 60292 12652 60332
rect 12692 60292 13228 60332
rect 13268 60292 18892 60332
rect 18932 60292 18941 60332
rect 0 60248 80 60268
rect 4876 60248 4916 60292
rect 0 60208 364 60248
rect 404 60208 413 60248
rect 2755 60208 2764 60248
rect 2804 60208 3244 60248
rect 3284 60208 3293 60248
rect 3340 60208 4916 60248
rect 6019 60248 6077 60249
rect 7747 60248 7805 60249
rect 6019 60208 6028 60248
rect 6068 60208 6700 60248
rect 6740 60208 6749 60248
rect 7651 60208 7660 60248
rect 7700 60208 7756 60248
rect 7796 60208 7805 60248
rect 10723 60208 10732 60248
rect 10772 60208 11212 60248
rect 11252 60208 11261 60248
rect 11587 60208 11596 60248
rect 11636 60208 11645 60248
rect 0 60188 80 60208
rect 3340 60165 3380 60208
rect 6019 60207 6077 60208
rect 7747 60207 7805 60208
rect 3331 60164 3389 60165
rect 11011 60164 11069 60165
rect 11203 60164 11261 60165
rect 3331 60124 3340 60164
rect 3380 60124 3389 60164
rect 4099 60124 4108 60164
rect 4148 60124 7084 60164
rect 7124 60124 7133 60164
rect 10926 60124 11020 60164
rect 11060 60124 11069 60164
rect 11118 60124 11127 60164
rect 11167 60124 11212 60164
rect 11252 60124 11261 60164
rect 3331 60123 3389 60124
rect 11011 60123 11069 60124
rect 11203 60123 11261 60124
rect 4099 60080 4157 60081
rect 11596 60080 11636 60208
rect 12067 60080 12125 60081
rect 3811 60040 3820 60080
rect 3860 60040 4108 60080
rect 4148 60040 4157 60080
rect 6211 60040 6220 60080
rect 6260 60040 6700 60080
rect 6740 60040 12076 60080
rect 12116 60040 12125 60080
rect 4099 60039 4157 60040
rect 12067 60039 12125 60040
rect 12460 59996 12500 60292
rect 13219 60291 13277 60292
rect 15907 60248 15965 60249
rect 15907 60208 15916 60248
rect 15956 60208 18412 60248
rect 18452 60208 18461 60248
rect 15907 60207 15965 60208
rect 12643 60124 12652 60164
rect 12692 60124 17356 60164
rect 17396 60124 17405 60164
rect 21424 60080 21504 60100
rect 12547 60040 12556 60080
rect 12596 60040 13228 60080
rect 13268 60040 13900 60080
rect 13940 60040 13949 60080
rect 14092 60040 14860 60080
rect 14900 60040 14909 60080
rect 16771 60040 16780 60080
rect 16820 60040 21504 60080
rect 14092 59996 14132 60040
rect 3619 59956 3628 59996
rect 3668 59956 4300 59996
rect 4340 59956 6988 59996
rect 7028 59956 11596 59996
rect 11636 59956 11788 59996
rect 11828 59956 11837 59996
rect 12460 59956 14132 59996
rect 0 59912 80 59932
rect 4099 59912 4157 59913
rect 11116 59912 11156 59956
rect 12451 59912 12509 59913
rect 12643 59912 12701 59913
rect 14380 59912 14420 60040
rect 21424 60020 21504 60040
rect 15811 59912 15869 59913
rect 0 59872 2540 59912
rect 0 59852 80 59872
rect 2500 59828 2540 59872
rect 4099 59872 4108 59912
rect 4148 59872 7660 59912
rect 7700 59872 7709 59912
rect 11107 59872 11116 59912
rect 11156 59872 11165 59912
rect 12451 59872 12460 59912
rect 12500 59872 12652 59912
rect 12692 59872 12701 59912
rect 14371 59872 14380 59912
rect 14420 59872 14429 59912
rect 15811 59872 15820 59912
rect 15860 59872 16108 59912
rect 16148 59872 16157 59912
rect 19555 59872 19564 59912
rect 19604 59872 20908 59912
rect 20948 59872 20957 59912
rect 4099 59871 4157 59872
rect 7660 59828 7700 59872
rect 12451 59871 12509 59872
rect 12643 59871 12701 59872
rect 15811 59871 15869 59872
rect 11203 59828 11261 59829
rect 19939 59828 19997 59829
rect 2500 59788 5396 59828
rect 7660 59788 10636 59828
rect 10676 59788 11212 59828
rect 11252 59788 11261 59828
rect 14947 59788 14956 59828
rect 14996 59788 19948 59828
rect 19988 59788 19997 59828
rect 5356 59744 5396 59788
rect 11203 59787 11261 59788
rect 19939 59787 19997 59788
rect 11971 59744 12029 59745
rect 21424 59744 21504 59764
rect 4919 59704 4928 59744
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 5296 59704 5305 59744
rect 5356 59704 5836 59744
rect 5876 59704 10444 59744
rect 10484 59704 10493 59744
rect 11971 59704 11980 59744
rect 12020 59704 12364 59744
rect 12404 59704 12413 59744
rect 14275 59704 14284 59744
rect 14324 59704 14476 59744
rect 14516 59704 14525 59744
rect 16387 59704 16396 59744
rect 16436 59704 16780 59744
rect 16820 59704 16829 59744
rect 20039 59704 20048 59744
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20416 59704 20425 59744
rect 20803 59704 20812 59744
rect 20852 59704 21504 59744
rect 11971 59703 12029 59704
rect 21424 59684 21504 59704
rect 7267 59660 7325 59661
rect 7267 59620 7276 59660
rect 7316 59620 7372 59660
rect 7412 59620 7421 59660
rect 8515 59620 8524 59660
rect 8564 59620 9964 59660
rect 10004 59620 10013 59660
rect 10243 59620 10252 59660
rect 10292 59620 11212 59660
rect 11252 59620 19756 59660
rect 19796 59620 19805 59660
rect 7267 59619 7325 59620
rect 0 59576 80 59596
rect 0 59536 8428 59576
rect 8468 59536 8477 59576
rect 8611 59536 8620 59576
rect 8660 59536 11980 59576
rect 12020 59536 12029 59576
rect 12835 59536 12844 59576
rect 12884 59536 13036 59576
rect 13076 59536 13085 59576
rect 14659 59536 14668 59576
rect 14708 59536 15244 59576
rect 15284 59536 15293 59576
rect 15907 59536 15916 59576
rect 15956 59536 16396 59576
rect 16436 59536 16445 59576
rect 0 59516 80 59536
rect 11779 59492 11837 59493
rect 19555 59492 19613 59493
rect 11694 59452 11788 59492
rect 11828 59452 11837 59492
rect 14467 59452 14476 59492
rect 14516 59452 16588 59492
rect 16628 59452 16637 59492
rect 19470 59452 19564 59492
rect 19604 59452 19613 59492
rect 11779 59451 11837 59452
rect 19555 59451 19613 59452
rect 4579 59408 4637 59409
rect 14659 59408 14717 59409
rect 19267 59408 19325 59409
rect 21424 59408 21504 59428
rect 4494 59368 4588 59408
rect 4628 59368 6220 59408
rect 6260 59368 6412 59408
rect 6452 59368 6461 59408
rect 8323 59368 8332 59408
rect 8372 59368 8620 59408
rect 8660 59368 8669 59408
rect 10531 59368 10540 59408
rect 10580 59368 11020 59408
rect 11060 59368 11069 59408
rect 12643 59368 12652 59408
rect 12692 59368 14092 59408
rect 14132 59368 14141 59408
rect 14574 59368 14668 59408
rect 14708 59368 14717 59408
rect 18211 59368 18220 59408
rect 18260 59368 19276 59408
rect 19316 59368 19325 59408
rect 4579 59367 4637 59368
rect 14659 59367 14717 59368
rect 19267 59367 19325 59368
rect 21292 59368 21504 59408
rect 4195 59324 4253 59325
rect 3715 59284 3724 59324
rect 3764 59284 4204 59324
rect 4244 59284 4253 59324
rect 4195 59283 4253 59284
rect 4387 59324 4445 59325
rect 4387 59284 4396 59324
rect 4436 59284 4530 59324
rect 4771 59284 4780 59324
rect 4820 59284 5164 59324
rect 5204 59284 5213 59324
rect 5347 59284 5356 59324
rect 5396 59284 14476 59324
rect 14516 59284 14525 59324
rect 14572 59284 19756 59324
rect 19796 59284 19805 59324
rect 4387 59283 4445 59284
rect 0 59240 80 59260
rect 3139 59240 3197 59241
rect 6883 59240 6941 59241
rect 8515 59240 8573 59241
rect 0 59200 748 59240
rect 788 59200 797 59240
rect 3139 59200 3148 59240
rect 3188 59200 4972 59240
rect 5012 59200 5021 59240
rect 6787 59200 6796 59240
rect 6836 59200 6892 59240
rect 6932 59200 7180 59240
rect 7220 59200 7229 59240
rect 7276 59200 8524 59240
rect 8564 59200 8573 59240
rect 0 59180 80 59200
rect 3139 59199 3197 59200
rect 6883 59199 6941 59200
rect 7276 59156 7316 59200
rect 8515 59199 8573 59200
rect 9091 59240 9149 59241
rect 14572 59240 14612 59284
rect 14851 59240 14909 59241
rect 9091 59200 9100 59240
rect 9140 59200 9484 59240
rect 9524 59200 9533 59240
rect 10147 59200 10156 59240
rect 10196 59200 10732 59240
rect 10772 59200 11020 59240
rect 11060 59200 11069 59240
rect 11971 59200 11980 59240
rect 12020 59200 14572 59240
rect 14612 59200 14621 59240
rect 14851 59200 14860 59240
rect 14900 59200 16684 59240
rect 16724 59200 16733 59240
rect 17155 59200 17164 59240
rect 17204 59200 20180 59240
rect 9091 59199 9149 59200
rect 14851 59199 14909 59200
rect 20140 59156 20180 59200
rect 21292 59156 21332 59368
rect 21424 59348 21504 59368
rect 2659 59116 2668 59156
rect 2708 59116 4204 59156
rect 4244 59116 4253 59156
rect 6403 59116 6412 59156
rect 6452 59116 7316 59156
rect 17539 59116 17548 59156
rect 17588 59116 17597 59156
rect 19747 59116 19756 59156
rect 19796 59116 19948 59156
rect 19988 59116 19997 59156
rect 20140 59116 21332 59156
rect 12259 59072 12317 59073
rect 17548 59072 17588 59116
rect 21424 59072 21504 59092
rect 12259 59032 12268 59072
rect 12308 59032 13516 59072
rect 13556 59032 13565 59072
rect 17548 59032 21504 59072
rect 12259 59031 12317 59032
rect 21424 59012 21504 59032
rect 259 58988 317 58989
rect 259 58948 268 58988
rect 308 58948 2540 58988
rect 3679 58948 3688 58988
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 4056 58948 4065 58988
rect 6115 58948 6124 58988
rect 6164 58948 6508 58988
rect 6548 58948 6557 58988
rect 7459 58948 7468 58988
rect 7508 58948 15340 58988
rect 15380 58948 15389 58988
rect 18799 58948 18808 58988
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 19176 58948 19185 58988
rect 259 58947 317 58948
rect 0 58904 80 58924
rect 2500 58904 2540 58948
rect 0 58864 940 58904
rect 980 58864 989 58904
rect 2500 58864 6988 58904
rect 7028 58864 7037 58904
rect 0 58844 80 58864
rect 7468 58820 7508 58948
rect 14083 58904 14141 58905
rect 8899 58864 8908 58904
rect 8948 58864 9580 58904
rect 9620 58864 11308 58904
rect 11348 58864 11357 58904
rect 13699 58864 13708 58904
rect 13748 58864 14092 58904
rect 14132 58864 14141 58904
rect 14083 58863 14141 58864
rect 1411 58780 1420 58820
rect 1460 58780 2540 58820
rect 3331 58780 3340 58820
rect 3380 58780 3628 58820
rect 3668 58780 3677 58820
rect 3724 58780 7508 58820
rect 11011 58780 11020 58820
rect 11060 58780 11404 58820
rect 11444 58780 11453 58820
rect 2500 58736 2540 58780
rect 3724 58736 3764 58780
rect 10339 58736 10397 58737
rect 21424 58736 21504 58756
rect 2500 58696 3764 58736
rect 6211 58696 6220 58736
rect 6260 58696 10348 58736
rect 10388 58696 13708 58736
rect 13748 58696 13757 58736
rect 18595 58696 18604 58736
rect 18644 58696 19796 58736
rect 19843 58696 19852 58736
rect 19892 58696 21504 58736
rect 10339 58695 10397 58696
rect 8323 58652 8381 58653
rect 8515 58652 8573 58653
rect 19267 58652 19325 58653
rect 19756 58652 19796 58696
rect 21424 58676 21504 58696
rect 6307 58612 6316 58652
rect 6356 58612 8332 58652
rect 8372 58612 8524 58652
rect 8564 58612 8573 58652
rect 15331 58612 15340 58652
rect 15380 58612 17260 58652
rect 17300 58612 17309 58652
rect 19267 58612 19276 58652
rect 19316 58612 19660 58652
rect 19700 58612 19709 58652
rect 19756 58612 20044 58652
rect 20084 58612 20093 58652
rect 8323 58611 8381 58612
rect 8515 58611 8573 58612
rect 19267 58611 19325 58612
rect 0 58568 80 58588
rect 15715 58568 15773 58569
rect 0 58528 1324 58568
rect 1364 58528 1373 58568
rect 3043 58528 3052 58568
rect 3092 58528 3436 58568
rect 3476 58528 3485 58568
rect 4675 58528 4684 58568
rect 4724 58528 11212 58568
rect 11252 58528 12364 58568
rect 12404 58528 12413 58568
rect 15715 58528 15724 58568
rect 15764 58528 17644 58568
rect 17684 58528 18124 58568
rect 18164 58528 18173 58568
rect 0 58508 80 58528
rect 15715 58527 15773 58528
rect 8131 58484 8189 58485
rect 8707 58484 8765 58485
rect 4291 58444 4300 58484
rect 4340 58444 5932 58484
rect 5972 58444 5981 58484
rect 6787 58444 6796 58484
rect 6836 58444 7372 58484
rect 7412 58444 7421 58484
rect 7555 58444 7564 58484
rect 7604 58444 8140 58484
rect 8180 58444 8716 58484
rect 8756 58444 9292 58484
rect 9332 58444 9341 58484
rect 10435 58444 10444 58484
rect 10484 58444 10828 58484
rect 10868 58444 10877 58484
rect 8131 58443 8189 58444
rect 8707 58443 8765 58444
rect 21424 58400 21504 58420
rect 2500 58360 9676 58400
rect 9716 58360 9725 58400
rect 10051 58360 10060 58400
rect 10100 58360 12748 58400
rect 12788 58360 12797 58400
rect 17443 58360 17452 58400
rect 17492 58360 21504 58400
rect 0 58232 80 58252
rect 2500 58232 2540 58360
rect 21424 58340 21504 58360
rect 4099 58316 4157 58317
rect 4014 58276 4108 58316
rect 4148 58276 4157 58316
rect 4099 58275 4157 58276
rect 0 58192 2540 58232
rect 4919 58192 4928 58232
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 5296 58192 5305 58232
rect 5923 58192 5932 58232
rect 5972 58192 7468 58232
rect 7508 58192 8908 58232
rect 8948 58192 8957 58232
rect 20039 58192 20048 58232
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20416 58192 20425 58232
rect 0 58172 80 58192
rect 12355 58148 12413 58149
rect 12355 58108 12364 58148
rect 12404 58108 16684 58148
rect 16724 58108 16733 58148
rect 12355 58107 12413 58108
rect 19843 58064 19901 58065
rect 21424 58064 21504 58084
rect 3619 58024 3628 58064
rect 3668 58024 7412 58064
rect 8035 58024 8044 58064
rect 8084 58024 8716 58064
rect 8756 58024 8765 58064
rect 12643 58024 12652 58064
rect 12692 58024 13132 58064
rect 13172 58024 13181 58064
rect 15724 58024 17356 58064
rect 17396 58024 17405 58064
rect 19843 58024 19852 58064
rect 19892 58024 21504 58064
rect 7372 57980 7412 58024
rect 8227 57980 8285 57981
rect 15724 57980 15764 58024
rect 19843 58023 19901 58024
rect 21424 58004 21504 58024
rect 16483 57980 16541 57981
rect 17635 57980 17693 57981
rect 2659 57940 2668 57980
rect 2708 57940 2956 57980
rect 2996 57940 4300 57980
rect 4340 57940 4349 57980
rect 4483 57940 4492 57980
rect 4532 57940 5068 57980
rect 5108 57940 5117 57980
rect 7372 57940 8236 57980
rect 8276 57940 8285 57980
rect 11395 57940 11404 57980
rect 11444 57940 11484 57980
rect 12739 57940 12748 57980
rect 12788 57940 13324 57980
rect 13364 57940 13373 57980
rect 13699 57940 13708 57980
rect 13748 57940 15764 57980
rect 16398 57940 16492 57980
rect 16532 57940 16541 57980
rect 17539 57940 17548 57980
rect 17588 57940 17644 57980
rect 17684 57940 19276 57980
rect 19316 57940 19325 57980
rect 8227 57939 8285 57940
rect 0 57896 80 57916
rect 1315 57896 1373 57897
rect 4195 57896 4253 57897
rect 8131 57896 8189 57897
rect 11404 57896 11444 57940
rect 15724 57896 15764 57940
rect 16483 57939 16541 57940
rect 17635 57939 17693 57940
rect 0 57856 1324 57896
rect 1364 57856 1373 57896
rect 4003 57856 4012 57896
rect 4052 57856 4204 57896
rect 4244 57856 4253 57896
rect 8035 57856 8044 57896
rect 8084 57856 8140 57896
rect 8180 57856 8189 57896
rect 8419 57856 8428 57896
rect 8468 57856 8908 57896
rect 8948 57856 8957 57896
rect 9283 57856 9292 57896
rect 9332 57856 13132 57896
rect 13172 57856 13181 57896
rect 15715 57856 15724 57896
rect 15764 57856 15773 57896
rect 17059 57856 17068 57896
rect 17108 57856 19084 57896
rect 19124 57856 19133 57896
rect 0 57836 80 57856
rect 1315 57855 1373 57856
rect 4195 57855 4253 57856
rect 8131 57855 8189 57856
rect 1507 57772 1516 57812
rect 1556 57772 5356 57812
rect 5396 57772 5405 57812
rect 8995 57772 9004 57812
rect 9044 57772 9388 57812
rect 9428 57772 9437 57812
rect 12355 57772 12364 57812
rect 12404 57772 14092 57812
rect 14132 57772 14141 57812
rect 17827 57772 17836 57812
rect 17876 57772 20180 57812
rect 3235 57728 3293 57729
rect 4579 57728 4637 57729
rect 15331 57728 15389 57729
rect 20140 57728 20180 57772
rect 21424 57728 21504 57748
rect 3235 57688 3244 57728
rect 3284 57688 3532 57728
rect 3572 57688 3581 57728
rect 4291 57688 4300 57728
rect 4340 57688 4588 57728
rect 4628 57688 4637 57728
rect 15312 57688 15340 57728
rect 15380 57688 15436 57728
rect 15476 57688 16588 57728
rect 16628 57688 16972 57728
rect 17012 57688 17021 57728
rect 20140 57688 21504 57728
rect 3235 57687 3293 57688
rect 4579 57687 4637 57688
rect 15331 57687 15389 57688
rect 21424 57668 21504 57688
rect 5635 57604 5644 57644
rect 5684 57604 11360 57644
rect 15523 57604 15532 57644
rect 15572 57604 15724 57644
rect 15764 57604 15773 57644
rect 17347 57604 17356 57644
rect 17396 57604 17836 57644
rect 17876 57604 17885 57644
rect 0 57560 80 57580
rect 11320 57560 11360 57604
rect 11491 57560 11549 57561
rect 0 57520 1420 57560
rect 1460 57520 1469 57560
rect 2083 57520 2092 57560
rect 2132 57520 9964 57560
rect 10004 57520 10013 57560
rect 11320 57520 11500 57560
rect 11540 57520 11549 57560
rect 0 57500 80 57520
rect 11491 57519 11549 57520
rect 11779 57560 11837 57561
rect 11779 57520 11788 57560
rect 11828 57520 17932 57560
rect 17972 57520 17981 57560
rect 11779 57519 11837 57520
rect 7651 57476 7709 57477
rect 3679 57436 3688 57476
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 4056 57436 4065 57476
rect 7566 57436 7660 57476
rect 7700 57436 7709 57476
rect 8419 57436 8428 57476
rect 8468 57436 8812 57476
rect 8852 57436 8861 57476
rect 9379 57436 9388 57476
rect 9428 57436 11308 57476
rect 11348 57436 15916 57476
rect 15956 57436 15965 57476
rect 18799 57436 18808 57476
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 19176 57436 19185 57476
rect 7651 57435 7709 57436
rect 13987 57392 14045 57393
rect 6787 57352 6796 57392
rect 6836 57352 12556 57392
rect 12596 57352 12605 57392
rect 13902 57352 13996 57392
rect 14036 57352 14045 57392
rect 13987 57351 14045 57352
rect 20707 57392 20765 57393
rect 21424 57392 21504 57412
rect 20707 57352 20716 57392
rect 20756 57352 21504 57392
rect 20707 57351 20765 57352
rect 21424 57332 21504 57352
rect 7267 57308 7325 57309
rect 1699 57268 1708 57308
rect 1748 57268 7276 57308
rect 7316 57268 19756 57308
rect 19796 57268 19805 57308
rect 7267 57267 7325 57268
rect 0 57224 80 57244
rect 3427 57224 3485 57225
rect 6979 57224 7037 57225
rect 0 57184 1228 57224
rect 1268 57184 1277 57224
rect 3427 57184 3436 57224
rect 3476 57184 3628 57224
rect 3668 57184 3677 57224
rect 3811 57184 3820 57224
rect 3860 57184 6988 57224
rect 7028 57184 7037 57224
rect 0 57164 80 57184
rect 3427 57183 3485 57184
rect 6979 57183 7037 57184
rect 7747 57224 7805 57225
rect 7747 57184 7756 57224
rect 7796 57184 9388 57224
rect 9428 57184 11020 57224
rect 11060 57184 11069 57224
rect 12259 57184 12268 57224
rect 12308 57184 14092 57224
rect 14132 57184 14141 57224
rect 15052 57184 15148 57224
rect 15188 57184 15197 57224
rect 16195 57184 16204 57224
rect 16244 57184 16780 57224
rect 16820 57184 16829 57224
rect 7747 57183 7805 57184
rect 1699 57100 1708 57140
rect 1748 57100 7948 57140
rect 7988 57100 7997 57140
rect 8044 57100 14612 57140
rect 8044 57056 8084 57100
rect 14572 57056 14612 57100
rect 15052 57056 15092 57184
rect 16003 57100 16012 57140
rect 16052 57100 16876 57140
rect 16916 57100 16925 57140
rect 21424 57056 21504 57076
rect 7267 57016 7276 57056
rect 7316 57016 8084 57056
rect 8131 57016 8140 57056
rect 8180 57016 8332 57056
rect 8372 57016 8381 57056
rect 9763 57016 9772 57056
rect 9812 57016 10156 57056
rect 10196 57016 10205 57056
rect 11011 57016 11020 57056
rect 11060 57016 13420 57056
rect 13460 57016 13469 57056
rect 14563 57016 14572 57056
rect 14612 57016 14621 57056
rect 15043 57016 15052 57056
rect 15092 57016 15101 57056
rect 15715 57016 15724 57056
rect 15764 57016 16492 57056
rect 16532 57016 16541 57056
rect 16963 57016 16972 57056
rect 17012 57016 17260 57056
rect 17300 57016 17309 57056
rect 19939 57016 19948 57056
rect 19988 57016 19997 57056
rect 20707 57016 20716 57056
rect 20756 57016 21504 57056
rect 11779 56972 11837 56973
rect 19948 56972 19988 57016
rect 21424 56996 21504 57016
rect 2755 56932 2764 56972
rect 2804 56932 5260 56972
rect 5300 56932 5309 56972
rect 6979 56932 6988 56972
rect 7028 56932 11788 56972
rect 11828 56932 11837 56972
rect 12067 56932 12076 56972
rect 12116 56932 12268 56972
rect 12308 56932 12317 56972
rect 15139 56932 15148 56972
rect 15188 56932 15436 56972
rect 15476 56932 15485 56972
rect 19747 56932 19756 56972
rect 19796 56932 19988 56972
rect 11779 56931 11837 56932
rect 0 56888 80 56908
rect 0 56848 1900 56888
rect 1940 56848 1949 56888
rect 2500 56848 15244 56888
rect 15284 56848 15293 56888
rect 19555 56848 19564 56888
rect 19604 56848 20812 56888
rect 20852 56848 20861 56888
rect 0 56828 80 56848
rect 2500 56804 2540 56848
rect 13699 56804 13757 56805
rect 1699 56764 1708 56804
rect 1748 56764 2540 56804
rect 6979 56764 6988 56804
rect 7028 56764 7276 56804
rect 7316 56764 7325 56804
rect 7651 56764 7660 56804
rect 7700 56764 8428 56804
rect 8468 56764 8477 56804
rect 11491 56764 11500 56804
rect 11540 56764 11980 56804
rect 12020 56764 13612 56804
rect 13652 56764 13708 56804
rect 13748 56764 13757 56804
rect 19843 56764 19852 56804
rect 19892 56764 20756 56804
rect 13699 56763 13757 56764
rect 7939 56720 7997 56721
rect 12355 56720 12413 56721
rect 20716 56720 20756 56764
rect 21424 56720 21504 56740
rect 4919 56680 4928 56720
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 5296 56680 5305 56720
rect 7939 56680 7948 56720
rect 7988 56680 8140 56720
rect 8180 56680 8524 56720
rect 8564 56680 8573 56720
rect 11299 56680 11308 56720
rect 11348 56680 11596 56720
rect 11636 56680 11645 56720
rect 12259 56680 12268 56720
rect 12308 56680 12364 56720
rect 12404 56680 12413 56720
rect 13411 56680 13420 56720
rect 13460 56680 14956 56720
rect 14996 56680 15005 56720
rect 16195 56680 16204 56720
rect 16244 56680 16780 56720
rect 16820 56680 16829 56720
rect 20039 56680 20048 56720
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20416 56680 20425 56720
rect 20716 56680 21504 56720
rect 7939 56679 7997 56680
rect 12355 56679 12413 56680
rect 21424 56660 21504 56680
rect 8707 56636 8765 56637
rect 14755 56636 14813 56637
rect 2467 56596 2476 56636
rect 2516 56596 6412 56636
rect 6452 56596 6461 56636
rect 7747 56596 7756 56636
rect 7796 56596 8716 56636
rect 8756 56596 9772 56636
rect 9812 56596 9821 56636
rect 11395 56596 11404 56636
rect 11444 56596 11924 56636
rect 13987 56596 13996 56636
rect 14036 56596 14764 56636
rect 14804 56596 14813 56636
rect 15331 56596 15340 56636
rect 15380 56596 15724 56636
rect 15764 56596 15773 56636
rect 16963 56596 16972 56636
rect 17012 56596 17644 56636
rect 17684 56596 17693 56636
rect 8707 56595 8765 56596
rect 0 56552 80 56572
rect 11884 56552 11924 56596
rect 14755 56595 14813 56596
rect 15715 56552 15773 56553
rect 0 56512 10060 56552
rect 10100 56512 10109 56552
rect 11299 56512 11308 56552
rect 11348 56512 11788 56552
rect 11828 56512 11837 56552
rect 11884 56512 14092 56552
rect 14132 56512 14141 56552
rect 15043 56512 15052 56552
rect 15092 56512 15724 56552
rect 15764 56512 15773 56552
rect 0 56492 80 56512
rect 15715 56511 15773 56512
rect 3043 56428 3052 56468
rect 3092 56428 3628 56468
rect 3668 56428 3677 56468
rect 5155 56428 5164 56468
rect 5204 56428 5836 56468
rect 5876 56428 5885 56468
rect 10339 56428 10348 56468
rect 10388 56428 11212 56468
rect 11252 56428 11261 56468
rect 12547 56428 12556 56468
rect 12596 56428 14860 56468
rect 14900 56428 14909 56468
rect 19747 56428 19756 56468
rect 19796 56428 20180 56468
rect 20140 56384 20180 56428
rect 21424 56384 21504 56404
rect 2947 56344 2956 56384
rect 2996 56344 3436 56384
rect 3476 56344 3485 56384
rect 4675 56344 4684 56384
rect 4724 56344 7084 56384
rect 7124 56344 7133 56384
rect 9571 56344 9580 56384
rect 9620 56344 11884 56384
rect 11924 56344 11933 56384
rect 14275 56344 14284 56384
rect 14324 56344 15340 56384
rect 15380 56344 15389 56384
rect 16579 56344 16588 56384
rect 16628 56344 17836 56384
rect 17876 56344 17885 56384
rect 19363 56344 19372 56384
rect 19412 56344 19421 56384
rect 20140 56344 21504 56384
rect 16963 56300 17021 56301
rect 19372 56300 19412 56344
rect 21424 56324 21504 56344
rect 4195 56260 4204 56300
rect 4244 56260 5836 56300
rect 5876 56260 5885 56300
rect 6403 56260 6412 56300
rect 6452 56260 15820 56300
rect 15860 56260 16012 56300
rect 16052 56260 16061 56300
rect 16963 56260 16972 56300
rect 17012 56260 17740 56300
rect 17780 56260 19412 56300
rect 16963 56259 17021 56260
rect 0 56216 80 56236
rect 2755 56216 2813 56217
rect 14755 56216 14813 56217
rect 0 56176 2764 56216
rect 2804 56176 2813 56216
rect 6691 56176 6700 56216
rect 6740 56176 11308 56216
rect 11348 56176 11357 56216
rect 11491 56176 11500 56216
rect 11540 56176 11692 56216
rect 11732 56176 11741 56216
rect 12355 56176 12364 56216
rect 12404 56176 12556 56216
rect 12596 56176 12605 56216
rect 14083 56176 14092 56216
rect 14132 56176 14764 56216
rect 14804 56176 14813 56216
rect 15235 56176 15244 56216
rect 15284 56176 15628 56216
rect 15668 56176 17356 56216
rect 17396 56176 17405 56216
rect 18691 56176 18700 56216
rect 18740 56176 19372 56216
rect 19412 56176 19421 56216
rect 0 56156 80 56176
rect 2755 56175 2813 56176
rect 14755 56175 14813 56176
rect 13987 56132 14045 56133
rect 14563 56132 14621 56133
rect 19939 56132 19997 56133
rect 3331 56092 3340 56132
rect 3380 56092 3724 56132
rect 3764 56092 3773 56132
rect 4099 56092 4108 56132
rect 4148 56092 4492 56132
rect 4532 56092 4541 56132
rect 9571 56092 9580 56132
rect 9620 56092 9772 56132
rect 9812 56092 9821 56132
rect 13987 56092 13996 56132
rect 14036 56092 14284 56132
rect 14324 56092 14333 56132
rect 14563 56092 14572 56132
rect 14612 56092 17644 56132
rect 17684 56092 17693 56132
rect 18124 56092 19756 56132
rect 19796 56092 19805 56132
rect 19854 56092 19948 56132
rect 19988 56092 19997 56132
rect 13987 56091 14045 56092
rect 14563 56091 14621 56092
rect 18124 56048 18164 56092
rect 19939 56091 19997 56092
rect 21424 56048 21504 56068
rect 1315 56008 1324 56048
rect 1364 56008 1996 56048
rect 2036 56008 4628 56048
rect 8227 56008 8236 56048
rect 8276 56008 10252 56048
rect 10292 56008 10301 56048
rect 11788 56008 18124 56048
rect 18164 56008 18173 56048
rect 19651 56008 19660 56048
rect 19700 56008 21504 56048
rect 4588 55964 4628 56008
rect 11491 55964 11549 55965
rect 11788 55964 11828 56008
rect 21424 55988 21504 56008
rect 3679 55924 3688 55964
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 4056 55924 4065 55964
rect 4588 55924 11116 55964
rect 11156 55924 11165 55964
rect 11491 55924 11500 55964
rect 11540 55924 11788 55964
rect 11828 55924 11837 55964
rect 12547 55924 12556 55964
rect 12596 55924 14764 55964
rect 14804 55924 17164 55964
rect 17204 55924 17213 55964
rect 18799 55924 18808 55964
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 19176 55924 19185 55964
rect 11491 55923 11549 55924
rect 0 55880 80 55900
rect 0 55840 12940 55880
rect 12980 55840 12989 55880
rect 0 55820 80 55840
rect 3043 55756 3052 55796
rect 3092 55756 9484 55796
rect 9524 55756 9533 55796
rect 10243 55756 10252 55796
rect 10292 55756 15820 55796
rect 15860 55756 18604 55796
rect 18644 55756 19756 55796
rect 19796 55756 19805 55796
rect 3235 55712 3293 55713
rect 8707 55712 8765 55713
rect 13411 55712 13469 55713
rect 21424 55712 21504 55732
rect 172 55672 2540 55712
rect 3150 55672 3244 55712
rect 3284 55672 3293 55712
rect 8622 55672 8716 55712
rect 8756 55672 8765 55712
rect 10531 55672 10540 55712
rect 10580 55672 11020 55712
rect 11060 55672 11069 55712
rect 11320 55672 13420 55712
rect 13460 55672 13469 55712
rect 0 55544 80 55564
rect 172 55544 212 55672
rect 2500 55628 2540 55672
rect 3235 55671 3293 55672
rect 8707 55671 8765 55672
rect 11320 55628 11360 55672
rect 13411 55671 13469 55672
rect 16876 55672 17452 55712
rect 17492 55672 18124 55712
rect 18164 55672 18173 55712
rect 20515 55672 20524 55712
rect 20564 55672 21504 55712
rect 12643 55628 12701 55629
rect 16876 55628 16916 55672
rect 21424 55652 21504 55672
rect 17635 55628 17693 55629
rect 2500 55588 11360 55628
rect 12163 55588 12172 55628
rect 12212 55588 12364 55628
rect 12404 55588 12413 55628
rect 12643 55588 12652 55628
rect 12692 55588 16916 55628
rect 16963 55588 16972 55628
rect 17012 55588 17644 55628
rect 17684 55588 18700 55628
rect 18740 55588 18749 55628
rect 12643 55587 12701 55588
rect 17635 55587 17693 55588
rect 7651 55544 7709 55545
rect 11587 55544 11645 55545
rect 14083 55544 14141 55545
rect 16963 55544 17021 55545
rect 0 55504 212 55544
rect 3139 55504 3148 55544
rect 3188 55504 7084 55544
rect 7124 55504 7133 55544
rect 7651 55504 7660 55544
rect 7700 55504 7756 55544
rect 7796 55504 7805 55544
rect 8323 55504 8332 55544
rect 8372 55504 8381 55544
rect 11502 55504 11596 55544
rect 11636 55504 11645 55544
rect 11779 55504 11788 55544
rect 11828 55504 12404 55544
rect 0 55484 80 55504
rect 7651 55503 7709 55504
rect 1476 55420 1516 55460
rect 1556 55420 1565 55460
rect 5443 55420 5452 55460
rect 5492 55420 5740 55460
rect 5780 55420 5789 55460
rect 7908 55420 7948 55460
rect 7988 55420 7997 55460
rect 1516 55376 1556 55420
rect 7948 55376 7988 55420
rect 8332 55376 8372 55504
rect 11587 55503 11645 55504
rect 12364 55460 12404 55504
rect 14083 55504 14092 55544
rect 14132 55504 14476 55544
rect 14516 55504 14525 55544
rect 15523 55504 15532 55544
rect 15572 55504 15668 55544
rect 14083 55503 14141 55504
rect 13411 55460 13469 55461
rect 12355 55420 12364 55460
rect 12404 55420 12413 55460
rect 12931 55420 12940 55460
rect 12980 55420 12989 55460
rect 13411 55420 13420 55460
rect 13460 55420 13556 55460
rect 643 55336 652 55376
rect 692 55336 1556 55376
rect 2659 55336 2668 55376
rect 2708 55336 4204 55376
rect 4244 55336 4253 55376
rect 7948 55336 8236 55376
rect 8276 55336 8285 55376
rect 8332 55336 8660 55376
rect 8515 55292 8573 55293
rect 547 55252 556 55292
rect 596 55252 5452 55292
rect 5492 55252 5501 55292
rect 8323 55252 8332 55292
rect 8372 55252 8524 55292
rect 8564 55252 8573 55292
rect 8515 55251 8573 55252
rect 0 55208 80 55228
rect 8620 55208 8660 55336
rect 12940 55292 12980 55420
rect 13411 55419 13469 55420
rect 13516 55376 13556 55420
rect 15628 55376 15668 55504
rect 16963 55504 16972 55544
rect 17012 55504 17068 55544
rect 17108 55504 17117 55544
rect 19372 55504 19564 55544
rect 19604 55504 19613 55544
rect 20035 55504 20044 55544
rect 20084 55504 20180 55544
rect 16963 55503 17021 55504
rect 19372 55460 19412 55504
rect 20140 55460 20180 55504
rect 15972 55420 16012 55460
rect 16052 55420 16061 55460
rect 19363 55420 19372 55460
rect 19412 55420 19421 55460
rect 20140 55420 20756 55460
rect 16012 55376 16052 55420
rect 13507 55336 13516 55376
rect 13556 55336 13565 55376
rect 14467 55336 14476 55376
rect 14516 55336 15668 55376
rect 15811 55336 15820 55376
rect 15860 55336 16052 55376
rect 20716 55376 20756 55420
rect 21424 55376 21504 55396
rect 20716 55336 21504 55376
rect 21424 55316 21504 55336
rect 13699 55292 13757 55293
rect 15331 55292 15389 55293
rect 12940 55252 13420 55292
rect 13460 55252 13469 55292
rect 13699 55252 13708 55292
rect 13748 55252 15340 55292
rect 15380 55252 15389 55292
rect 13699 55251 13757 55252
rect 15331 55251 15389 55252
rect 16003 55292 16061 55293
rect 18115 55292 18173 55293
rect 16003 55252 16012 55292
rect 16052 55252 18124 55292
rect 18164 55252 18173 55292
rect 16003 55251 16061 55252
rect 18115 55251 18173 55252
rect 16387 55208 16445 55209
rect 0 55168 940 55208
rect 980 55168 989 55208
rect 1603 55168 1612 55208
rect 1652 55168 3532 55208
rect 3572 55168 3581 55208
rect 4919 55168 4928 55208
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 5296 55168 5305 55208
rect 8515 55168 8524 55208
rect 8564 55168 8660 55208
rect 13996 55168 16396 55208
rect 16436 55168 16445 55208
rect 17251 55168 17260 55208
rect 17300 55168 17836 55208
rect 17876 55168 17885 55208
rect 20039 55168 20048 55208
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20416 55168 20425 55208
rect 0 55148 80 55168
rect 2083 55084 2092 55124
rect 2132 55084 8044 55124
rect 8084 55084 8093 55124
rect 1315 55000 1324 55040
rect 1364 55000 10156 55040
rect 10196 55000 10205 55040
rect 7747 54956 7805 54957
rect 2179 54916 2188 54956
rect 2228 54916 2476 54956
rect 2516 54916 2525 54956
rect 3619 54916 3628 54956
rect 3668 54916 6604 54956
rect 6644 54916 6796 54956
rect 6836 54916 6845 54956
rect 7662 54916 7756 54956
rect 7796 54916 7805 54956
rect 9667 54916 9676 54956
rect 9716 54916 11308 54956
rect 11348 54916 11357 54956
rect 7747 54915 7805 54916
rect 0 54872 80 54892
rect 1411 54872 1469 54873
rect 13996 54872 14036 55168
rect 16387 55167 16445 55168
rect 14083 55124 14141 55125
rect 16003 55124 16061 55125
rect 14083 55084 14092 55124
rect 14132 55084 14572 55124
rect 14612 55084 14621 55124
rect 16003 55084 16012 55124
rect 16052 55084 16108 55124
rect 16148 55084 16157 55124
rect 18883 55084 18892 55124
rect 18932 55084 19276 55124
rect 19316 55084 19325 55124
rect 14083 55083 14141 55084
rect 16003 55083 16061 55084
rect 19939 55040 19997 55041
rect 21424 55040 21504 55060
rect 14371 55000 14380 55040
rect 14420 55000 14429 55040
rect 14947 55000 14956 55040
rect 14996 55000 15916 55040
rect 15956 55000 15965 55040
rect 16483 55000 16492 55040
rect 16532 55000 17068 55040
rect 17108 55000 17117 55040
rect 19939 55000 19948 55040
rect 19988 55000 21504 55040
rect 14083 54956 14141 54957
rect 14380 54956 14420 55000
rect 19939 54999 19997 55000
rect 21424 54980 21504 55000
rect 14083 54916 14092 54956
rect 14132 54916 14420 54956
rect 15331 54916 15340 54956
rect 15380 54916 16108 54956
rect 16148 54916 16157 54956
rect 19267 54916 19276 54956
rect 19316 54916 19564 54956
rect 19604 54916 19613 54956
rect 14083 54915 14141 54916
rect 14467 54872 14525 54873
rect 0 54832 1420 54872
rect 1460 54832 1469 54872
rect 4675 54832 4684 54872
rect 4724 54832 14036 54872
rect 14382 54832 14476 54872
rect 14516 54832 14525 54872
rect 0 54812 80 54832
rect 1411 54831 1469 54832
rect 14467 54831 14525 54832
rect 14668 54832 18412 54872
rect 18452 54832 18461 54872
rect 14668 54789 14708 54832
rect 11491 54788 11549 54789
rect 14659 54788 14717 54789
rect 15331 54788 15389 54789
rect 16387 54788 16445 54789
rect 2500 54748 11500 54788
rect 11540 54748 11549 54788
rect 14083 54748 14092 54788
rect 14132 54748 14668 54788
rect 14708 54748 14717 54788
rect 14851 54748 14860 54788
rect 14900 54748 14909 54788
rect 15331 54748 15340 54788
rect 15380 54748 15436 54788
rect 15476 54748 15485 54788
rect 16387 54748 16396 54788
rect 16436 54748 19756 54788
rect 19796 54748 19805 54788
rect 19939 54748 19948 54788
rect 19988 54748 19997 54788
rect 2500 54704 2540 54748
rect 11491 54747 11549 54748
rect 14659 54747 14717 54748
rect 8131 54704 8189 54705
rect 14860 54704 14900 54748
rect 15331 54747 15389 54748
rect 16387 54747 16445 54748
rect 1795 54664 1804 54704
rect 1844 54664 2540 54704
rect 2947 54664 2956 54704
rect 2996 54664 3340 54704
rect 3380 54664 3389 54704
rect 3523 54664 3532 54704
rect 3572 54664 3860 54704
rect 3427 54620 3485 54621
rect 3820 54620 3860 54664
rect 8131 54664 8140 54704
rect 8180 54664 14900 54704
rect 16579 54704 16637 54705
rect 19948 54704 19988 54748
rect 21424 54704 21504 54724
rect 16579 54664 16588 54704
rect 16628 54664 18892 54704
rect 18932 54664 18941 54704
rect 19948 54664 21504 54704
rect 8131 54663 8189 54664
rect 16579 54663 16637 54664
rect 21424 54644 21504 54664
rect 12451 54620 12509 54621
rect 1891 54580 1900 54620
rect 1940 54580 2380 54620
rect 2420 54580 2429 54620
rect 2500 54580 3436 54620
rect 3476 54580 3724 54620
rect 3764 54580 3773 54620
rect 3820 54580 12460 54620
rect 12500 54580 12509 54620
rect 0 54536 80 54556
rect 1603 54536 1661 54537
rect 0 54496 1612 54536
rect 1652 54496 1661 54536
rect 0 54476 80 54496
rect 1603 54495 1661 54496
rect 547 54452 605 54453
rect 2500 54452 2540 54580
rect 3427 54579 3485 54580
rect 12451 54579 12509 54580
rect 6115 54496 6124 54536
rect 6164 54496 6892 54536
rect 6932 54496 6941 54536
rect 7651 54496 7660 54536
rect 7700 54496 8140 54536
rect 8180 54496 8189 54536
rect 6019 54452 6077 54453
rect 547 54412 556 54452
rect 596 54412 2540 54452
rect 3679 54412 3688 54452
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 4056 54412 4065 54452
rect 6019 54412 6028 54452
rect 6068 54412 6316 54452
rect 6356 54412 6365 54452
rect 16003 54412 16012 54452
rect 16052 54412 16300 54452
rect 16340 54412 16349 54452
rect 16483 54412 16492 54452
rect 16532 54412 17164 54452
rect 17204 54412 17213 54452
rect 18799 54412 18808 54452
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 19176 54412 19185 54452
rect 547 54411 605 54412
rect 6019 54411 6077 54412
rect 8131 54368 8189 54369
rect 21424 54368 21504 54388
rect 2563 54328 2572 54368
rect 2612 54328 3860 54368
rect 8046 54328 8140 54368
rect 8180 54328 8189 54368
rect 17827 54328 17836 54368
rect 17876 54328 21504 54368
rect 3820 54284 3860 54328
rect 8131 54327 8189 54328
rect 21424 54308 21504 54328
rect 2500 54244 2860 54284
rect 2900 54244 2909 54284
rect 3811 54244 3820 54284
rect 3860 54244 3869 54284
rect 11971 54244 11980 54284
rect 12020 54244 12268 54284
rect 12308 54244 12317 54284
rect 14371 54244 14380 54284
rect 14420 54244 14668 54284
rect 14708 54244 14717 54284
rect 15907 54244 15916 54284
rect 15956 54244 16300 54284
rect 16340 54244 16349 54284
rect 0 54200 80 54220
rect 2500 54200 2540 54244
rect 13987 54200 14045 54201
rect 16099 54200 16157 54201
rect 19651 54200 19709 54201
rect 0 54160 2540 54200
rect 2659 54160 2668 54200
rect 2708 54160 4012 54200
rect 4052 54160 4061 54200
rect 11299 54160 11308 54200
rect 11348 54160 12844 54200
rect 12884 54160 12893 54200
rect 13987 54160 13996 54200
rect 14036 54160 14188 54200
rect 14228 54160 14237 54200
rect 16099 54160 16108 54200
rect 16148 54160 17740 54200
rect 17780 54160 17789 54200
rect 19555 54160 19564 54200
rect 19604 54160 19660 54200
rect 19700 54160 19709 54200
rect 0 54140 80 54160
rect 13987 54159 14045 54160
rect 16099 54159 16157 54160
rect 19651 54159 19709 54160
rect 20515 54200 20573 54201
rect 20515 54160 20524 54200
rect 20564 54160 21292 54200
rect 21332 54160 21341 54200
rect 20515 54159 20573 54160
rect 2467 54116 2525 54117
rect 2755 54116 2813 54117
rect 11491 54116 11549 54117
rect 2467 54076 2476 54116
rect 2516 54076 2764 54116
rect 2804 54076 2813 54116
rect 2467 54075 2525 54076
rect 2755 54075 2813 54076
rect 3244 54076 9868 54116
rect 9908 54076 9917 54116
rect 11472 54076 11500 54116
rect 11540 54076 11596 54116
rect 11636 54076 17644 54116
rect 17684 54076 17693 54116
rect 19651 54076 19660 54116
rect 19700 54076 19709 54116
rect 2371 54032 2429 54033
rect 3244 54032 3284 54076
rect 11491 54075 11549 54076
rect 7651 54032 7709 54033
rect 8323 54032 8381 54033
rect 10819 54032 10877 54033
rect 16963 54032 17021 54033
rect 1411 53992 1420 54032
rect 1460 53992 1469 54032
rect 2371 53992 2380 54032
rect 2420 53992 3284 54032
rect 3331 53992 3340 54032
rect 3380 53992 5644 54032
rect 5684 53992 6124 54032
rect 6164 53992 7564 54032
rect 7604 53992 7660 54032
rect 7700 53992 7728 54032
rect 8323 53992 8332 54032
rect 8372 53992 8524 54032
rect 8564 53992 8573 54032
rect 8707 53992 8716 54032
rect 8756 53992 10828 54032
rect 10868 53992 10877 54032
rect 14467 53992 14476 54032
rect 14516 53992 16108 54032
rect 16148 53992 16157 54032
rect 16878 53992 16972 54032
rect 17012 53992 19084 54032
rect 19124 53992 19276 54032
rect 19316 53992 19325 54032
rect 0 53864 80 53884
rect 0 53824 212 53864
rect 0 53804 80 53824
rect 172 53696 212 53824
rect 1420 53780 1460 53992
rect 2371 53991 2429 53992
rect 7651 53991 7709 53992
rect 8323 53991 8381 53992
rect 10819 53991 10877 53992
rect 16963 53991 17021 53992
rect 19660 53948 19700 54076
rect 21424 54032 21504 54052
rect 20227 53992 20236 54032
rect 20276 53992 21504 54032
rect 21424 53972 21504 53992
rect 2083 53908 2092 53948
rect 2132 53908 10060 53948
rect 10100 53908 10109 53948
rect 11107 53908 11116 53948
rect 11156 53908 11404 53948
rect 11444 53908 11453 53948
rect 13219 53908 13228 53948
rect 13268 53908 19700 53948
rect 8611 53824 8620 53864
rect 8660 53824 14764 53864
rect 14804 53824 14813 53864
rect 18883 53824 18892 53864
rect 18932 53824 20044 53864
rect 20084 53824 20093 53864
rect 17539 53780 17597 53781
rect 19363 53780 19421 53781
rect 1420 53740 5780 53780
rect 7075 53740 7084 53780
rect 7124 53740 8716 53780
rect 8756 53740 8765 53780
rect 11395 53740 11404 53780
rect 11444 53740 14860 53780
rect 14900 53740 14909 53780
rect 17539 53740 17548 53780
rect 17588 53740 19372 53780
rect 19412 53740 19421 53780
rect 19747 53740 19756 53780
rect 19796 53740 20564 53780
rect 5740 53696 5780 53740
rect 17539 53739 17597 53740
rect 19363 53739 19421 53740
rect 14275 53696 14333 53697
rect 20524 53696 20564 53740
rect 21424 53696 21504 53716
rect 172 53656 2540 53696
rect 4919 53656 4928 53696
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 5296 53656 5305 53696
rect 5731 53656 5740 53696
rect 5780 53656 5789 53696
rect 7843 53656 7852 53696
rect 7892 53656 8524 53696
rect 8564 53656 8573 53696
rect 11107 53656 11116 53696
rect 11156 53656 11308 53696
rect 11348 53656 11357 53696
rect 12643 53656 12652 53696
rect 12692 53656 12844 53696
rect 12884 53656 12893 53696
rect 14275 53656 14284 53696
rect 14324 53656 18028 53696
rect 18068 53656 18316 53696
rect 18356 53656 18365 53696
rect 20039 53656 20048 53696
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20416 53656 20425 53696
rect 20524 53656 21504 53696
rect 2500 53612 2540 53656
rect 14275 53655 14333 53656
rect 21424 53636 21504 53656
rect 16387 53612 16445 53613
rect 2500 53572 11252 53612
rect 16195 53572 16204 53612
rect 16244 53572 16396 53612
rect 16436 53572 16445 53612
rect 0 53528 80 53548
rect 3235 53528 3293 53529
rect 8707 53528 8765 53529
rect 11212 53528 11252 53572
rect 16387 53571 16445 53572
rect 12739 53528 12797 53529
rect 0 53488 3244 53528
rect 3284 53488 3293 53528
rect 8622 53488 8716 53528
rect 8756 53488 8765 53528
rect 11203 53488 11212 53528
rect 11252 53488 11261 53528
rect 12067 53488 12076 53528
rect 12116 53488 12748 53528
rect 12788 53488 12797 53528
rect 0 53468 80 53488
rect 3235 53487 3293 53488
rect 8707 53487 8765 53488
rect 12739 53487 12797 53488
rect 14947 53528 15005 53529
rect 14947 53488 14956 53528
rect 14996 53488 19180 53528
rect 19220 53488 19229 53528
rect 14947 53487 15005 53488
rect 1507 53404 1516 53444
rect 1556 53404 1565 53444
rect 3523 53404 3532 53444
rect 3572 53404 4012 53444
rect 4052 53404 4061 53444
rect 5827 53404 5836 53444
rect 5876 53404 6028 53444
rect 6068 53404 14476 53444
rect 14516 53404 14525 53444
rect 15427 53404 15436 53444
rect 15476 53404 16588 53444
rect 16628 53404 16637 53444
rect 19939 53404 19948 53444
rect 19988 53404 20180 53444
rect 1516 53360 1556 53404
rect 4387 53360 4445 53361
rect 20140 53360 20180 53404
rect 21424 53360 21504 53380
rect 76 53320 1556 53360
rect 2563 53320 2572 53360
rect 2612 53320 4396 53360
rect 4436 53320 13228 53360
rect 13268 53320 13277 53360
rect 13699 53320 13708 53360
rect 13748 53320 14668 53360
rect 14708 53320 15628 53360
rect 15668 53320 15677 53360
rect 19075 53320 19084 53360
rect 19124 53320 19564 53360
rect 19604 53320 19613 53360
rect 20140 53320 21504 53360
rect 76 53212 116 53320
rect 4387 53319 4445 53320
rect 21424 53300 21504 53320
rect 11491 53276 11549 53277
rect 13219 53276 13277 53277
rect 14275 53276 14333 53277
rect 1891 53236 1900 53276
rect 1940 53236 5740 53276
rect 5780 53236 5789 53276
rect 9859 53236 9868 53276
rect 9908 53236 9917 53276
rect 11203 53236 11212 53276
rect 11252 53236 11500 53276
rect 11540 53236 11549 53276
rect 12163 53236 12172 53276
rect 12212 53236 13228 53276
rect 13268 53236 13324 53276
rect 13364 53236 13373 53276
rect 14190 53236 14284 53276
rect 14324 53236 14333 53276
rect 15715 53236 15724 53276
rect 15764 53236 16108 53276
rect 16148 53236 16157 53276
rect 19939 53236 19948 53276
rect 19988 53236 19997 53276
rect 0 53152 116 53212
rect 0 53132 80 53152
rect 9868 53108 9908 53236
rect 11491 53235 11549 53236
rect 13219 53235 13277 53236
rect 14275 53235 14333 53236
rect 11107 53192 11165 53193
rect 12451 53192 12509 53193
rect 14083 53192 14141 53193
rect 19948 53192 19988 53236
rect 11107 53152 11116 53192
rect 11156 53152 11308 53192
rect 11348 53152 11357 53192
rect 12451 53152 12460 53192
rect 12500 53152 12652 53192
rect 12692 53152 12701 53192
rect 14083 53152 14092 53192
rect 14132 53152 14188 53192
rect 14228 53152 14237 53192
rect 14851 53152 14860 53192
rect 14900 53152 19988 53192
rect 11107 53151 11165 53152
rect 12451 53151 12509 53152
rect 14083 53151 14141 53152
rect 8611 53068 8620 53108
rect 8660 53068 18892 53108
rect 18932 53068 18941 53108
rect 4579 53024 4637 53025
rect 12739 53024 12797 53025
rect 15043 53024 15101 53025
rect 21424 53024 21504 53044
rect 4494 52984 4588 53024
rect 4628 52984 11884 53024
rect 11924 52984 11933 53024
rect 12739 52984 12748 53024
rect 12788 52984 13612 53024
rect 13652 52984 13661 53024
rect 15043 52984 15052 53024
rect 15092 52984 16876 53024
rect 16916 52984 16925 53024
rect 19843 52984 19852 53024
rect 19892 52984 21504 53024
rect 4579 52983 4637 52984
rect 12739 52983 12797 52984
rect 15043 52983 15101 52984
rect 21424 52964 21504 52984
rect 17731 52940 17789 52941
rect 19843 52940 19901 52941
rect 3679 52900 3688 52940
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 4056 52900 4065 52940
rect 5059 52900 5068 52940
rect 5108 52900 5356 52940
rect 5396 52900 7564 52940
rect 7604 52900 9100 52940
rect 9140 52900 9149 52940
rect 11011 52900 11020 52940
rect 11060 52900 13804 52940
rect 13844 52900 17588 52940
rect 17635 52900 17644 52940
rect 17684 52900 17740 52940
rect 17780 52900 17789 52940
rect 18799 52900 18808 52940
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 19176 52900 19185 52940
rect 19651 52900 19660 52940
rect 19700 52900 19852 52940
rect 19892 52900 19901 52940
rect 0 52856 80 52876
rect 13219 52856 13277 52857
rect 15619 52856 15677 52857
rect 17548 52856 17588 52900
rect 17731 52899 17789 52900
rect 19843 52899 19901 52900
rect 19948 52900 21100 52940
rect 21140 52900 21149 52940
rect 19948 52857 19988 52900
rect 19939 52856 19997 52857
rect 0 52816 1804 52856
rect 1844 52816 1853 52856
rect 1987 52816 1996 52856
rect 2036 52816 4972 52856
rect 5012 52816 5021 52856
rect 7843 52816 7852 52856
rect 7892 52816 9484 52856
rect 9524 52816 9772 52856
rect 9812 52816 9821 52856
rect 13219 52816 13228 52856
rect 13268 52816 15052 52856
rect 15092 52816 15101 52856
rect 15523 52816 15532 52856
rect 15572 52816 15628 52856
rect 15668 52816 15677 52856
rect 17539 52816 17548 52856
rect 17588 52816 17597 52856
rect 19939 52816 19948 52856
rect 19988 52816 19997 52856
rect 0 52796 80 52816
rect 13219 52815 13277 52816
rect 15619 52815 15677 52816
rect 19939 52815 19997 52816
rect 20140 52816 20716 52856
rect 20756 52816 20765 52856
rect 5059 52772 5117 52773
rect 19459 52772 19517 52773
rect 20140 52772 20180 52816
rect 2563 52732 2572 52772
rect 2612 52732 3244 52772
rect 3284 52732 3293 52772
rect 3811 52732 3820 52772
rect 3860 52732 4492 52772
rect 4532 52732 4541 52772
rect 5059 52732 5068 52772
rect 5108 52732 5452 52772
rect 5492 52732 5501 52772
rect 19459 52732 19468 52772
rect 19508 52732 20180 52772
rect 5059 52731 5117 52732
rect 19459 52731 19517 52732
rect 21424 52688 21504 52708
rect 1507 52648 1516 52688
rect 1556 52648 4684 52688
rect 4724 52648 11116 52688
rect 11156 52648 11165 52688
rect 14371 52648 14380 52688
rect 14420 52648 14860 52688
rect 14900 52648 15244 52688
rect 15284 52648 15293 52688
rect 18979 52648 18988 52688
rect 19028 52648 19468 52688
rect 19508 52648 19517 52688
rect 20131 52648 20140 52688
rect 20180 52648 21504 52688
rect 21424 52628 21504 52648
rect 7843 52604 7901 52605
rect 7843 52564 7852 52604
rect 7892 52564 19756 52604
rect 19796 52564 19805 52604
rect 7843 52563 7901 52564
rect 0 52520 80 52540
rect 6883 52520 6941 52521
rect 0 52480 1612 52520
rect 1652 52480 1661 52520
rect 3331 52480 3340 52520
rect 3380 52480 4204 52520
rect 4244 52480 4253 52520
rect 6595 52480 6604 52520
rect 6644 52480 6892 52520
rect 6932 52480 6941 52520
rect 7171 52480 7180 52520
rect 7220 52480 9388 52520
rect 9428 52480 11020 52520
rect 11060 52480 11069 52520
rect 11320 52480 12940 52520
rect 12980 52480 12989 52520
rect 13315 52480 13324 52520
rect 13364 52480 15244 52520
rect 15284 52480 15293 52520
rect 15715 52480 15724 52520
rect 15764 52480 15916 52520
rect 15956 52480 15965 52520
rect 0 52460 80 52480
rect 6883 52479 6941 52480
rect 6892 52436 6932 52479
rect 11320 52436 11360 52480
rect 4291 52396 4300 52436
rect 4340 52396 4492 52436
rect 4532 52396 4541 52436
rect 6892 52396 8716 52436
rect 8756 52396 11360 52436
rect 13507 52396 13516 52436
rect 13556 52396 14188 52436
rect 14228 52396 15052 52436
rect 15092 52396 15101 52436
rect 17155 52396 17164 52436
rect 17204 52396 17452 52436
rect 17492 52396 17501 52436
rect 1603 52352 1661 52353
rect 16579 52352 16637 52353
rect 19459 52352 19517 52353
rect 21424 52352 21504 52372
rect 1518 52312 1612 52352
rect 1652 52312 1661 52352
rect 6595 52312 6604 52352
rect 6644 52312 8428 52352
rect 8468 52312 8477 52352
rect 8899 52312 8908 52352
rect 8948 52312 15148 52352
rect 15188 52312 16588 52352
rect 16628 52312 16637 52352
rect 19171 52312 19180 52352
rect 19220 52312 19468 52352
rect 19508 52312 19517 52352
rect 19939 52312 19948 52352
rect 19988 52312 21504 52352
rect 1603 52311 1661 52312
rect 16579 52311 16637 52312
rect 19459 52311 19517 52312
rect 21424 52292 21504 52312
rect 11683 52268 11741 52269
rect 16099 52268 16157 52269
rect 11683 52228 11692 52268
rect 11732 52228 11980 52268
rect 12020 52228 12029 52268
rect 16014 52228 16108 52268
rect 16148 52228 16157 52268
rect 11683 52227 11741 52228
rect 16099 52227 16157 52228
rect 0 52184 80 52204
rect 10531 52184 10589 52185
rect 0 52144 2380 52184
rect 2420 52144 2429 52184
rect 4919 52144 4928 52184
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 5296 52144 5305 52184
rect 6211 52144 6220 52184
rect 6260 52144 6508 52184
rect 6548 52144 6557 52184
rect 10531 52144 10540 52184
rect 10580 52144 19372 52184
rect 19412 52144 19421 52184
rect 20039 52144 20048 52184
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20416 52144 20425 52184
rect 0 52124 80 52144
rect 10531 52143 10589 52144
rect 2371 52100 2429 52101
rect 2947 52100 3005 52101
rect 15715 52100 15773 52101
rect 16483 52100 16541 52101
rect 2371 52060 2380 52100
rect 2420 52060 2956 52100
rect 2996 52060 3005 52100
rect 11683 52060 11692 52100
rect 11732 52060 13036 52100
rect 13076 52060 13085 52100
rect 15715 52060 15724 52100
rect 15764 52060 16012 52100
rect 16052 52060 16061 52100
rect 16483 52060 16492 52100
rect 16532 52060 16684 52100
rect 16724 52060 16733 52100
rect 2371 52059 2429 52060
rect 2947 52059 3005 52060
rect 15715 52059 15773 52060
rect 16483 52059 16541 52060
rect 21424 52016 21504 52036
rect 5059 51976 5068 52016
rect 5108 51976 9292 52016
rect 9332 51976 9341 52016
rect 10531 51976 10540 52016
rect 10580 51976 12844 52016
rect 12884 51976 13804 52016
rect 13844 51976 13853 52016
rect 16771 51976 16780 52016
rect 16820 51976 17164 52016
rect 17204 51976 17213 52016
rect 19555 51976 19564 52016
rect 19604 51976 21504 52016
rect 21424 51956 21504 51976
rect 16579 51932 16637 51933
rect 20899 51932 20957 51933
rect 2371 51892 2380 51932
rect 2420 51892 8236 51932
rect 8276 51892 8285 51932
rect 11107 51892 11116 51932
rect 11156 51892 14572 51932
rect 14612 51892 15724 51932
rect 15764 51892 15773 51932
rect 16483 51892 16492 51932
rect 16532 51892 16588 51932
rect 16628 51892 16637 51932
rect 19075 51892 19084 51932
rect 19124 51892 20908 51932
rect 20948 51892 20957 51932
rect 16579 51891 16637 51892
rect 20899 51891 20957 51892
rect 0 51848 80 51868
rect 0 51808 1708 51848
rect 1748 51808 1757 51848
rect 3811 51808 3820 51848
rect 3860 51808 10636 51848
rect 10676 51808 10685 51848
rect 11011 51808 11020 51848
rect 11060 51808 14092 51848
rect 14132 51808 14141 51848
rect 14851 51808 14860 51848
rect 14900 51808 18412 51848
rect 18452 51808 18461 51848
rect 0 51788 80 51808
rect 1891 51764 1949 51765
rect 6019 51764 6077 51765
rect 163 51724 172 51764
rect 212 51724 1076 51764
rect 1507 51724 1516 51764
rect 1556 51724 1900 51764
rect 1940 51724 2092 51764
rect 2132 51724 2141 51764
rect 2755 51724 2764 51764
rect 2804 51724 3532 51764
rect 3572 51724 4396 51764
rect 4436 51724 4445 51764
rect 5934 51724 6028 51764
rect 6068 51724 6077 51764
rect 931 51680 989 51681
rect 739 51640 748 51680
rect 788 51640 940 51680
rect 980 51640 989 51680
rect 1036 51680 1076 51724
rect 1891 51723 1949 51724
rect 6019 51723 6077 51724
rect 8323 51764 8381 51765
rect 13411 51764 13469 51765
rect 16963 51764 17021 51765
rect 8323 51724 8332 51764
rect 8372 51724 10444 51764
rect 10484 51724 10493 51764
rect 13411 51724 13420 51764
rect 13460 51724 13516 51764
rect 13556 51724 13565 51764
rect 15043 51724 15052 51764
rect 15092 51724 15820 51764
rect 15860 51724 15869 51764
rect 16099 51724 16108 51764
rect 16148 51724 16188 51764
rect 16291 51724 16300 51764
rect 16340 51724 16972 51764
rect 17012 51724 17021 51764
rect 8323 51723 8381 51724
rect 13411 51723 13469 51724
rect 16108 51680 16148 51724
rect 16963 51723 17021 51724
rect 18499 51764 18557 51765
rect 18499 51724 18508 51764
rect 18548 51724 19756 51764
rect 19796 51724 19805 51764
rect 18499 51723 18557 51724
rect 21424 51680 21504 51700
rect 1036 51640 1556 51680
rect 2947 51640 2956 51680
rect 2996 51640 4108 51680
rect 4148 51640 4157 51680
rect 7747 51640 7756 51680
rect 7796 51640 8236 51680
rect 8276 51640 10060 51680
rect 10100 51640 10109 51680
rect 10819 51640 10828 51680
rect 10868 51640 12076 51680
rect 12116 51640 12125 51680
rect 13795 51640 13804 51680
rect 13844 51640 14572 51680
rect 14612 51640 14860 51680
rect 14900 51640 14909 51680
rect 15139 51640 15148 51680
rect 15188 51640 16780 51680
rect 16820 51640 16829 51680
rect 19555 51640 19564 51680
rect 19604 51640 20084 51680
rect 20131 51640 20140 51680
rect 20180 51640 21504 51680
rect 931 51639 989 51640
rect 1516 51596 1556 51640
rect 20044 51596 20084 51640
rect 21424 51620 21504 51640
rect 1507 51556 1516 51596
rect 1556 51556 1565 51596
rect 7939 51556 7948 51596
rect 7988 51556 8620 51596
rect 8660 51556 8669 51596
rect 9283 51556 9292 51596
rect 9332 51556 10252 51596
rect 10292 51556 10301 51596
rect 12259 51556 12268 51596
rect 12308 51556 16108 51596
rect 16148 51556 16157 51596
rect 20044 51556 21140 51596
rect 0 51512 80 51532
rect 19555 51512 19613 51513
rect 20995 51512 21053 51513
rect 0 51472 1996 51512
rect 2036 51472 2045 51512
rect 5827 51472 5836 51512
rect 5876 51472 6124 51512
rect 6164 51472 6173 51512
rect 14083 51472 14092 51512
rect 14132 51472 14476 51512
rect 14516 51472 14525 51512
rect 19555 51472 19564 51512
rect 19604 51472 21004 51512
rect 21044 51472 21053 51512
rect 0 51452 80 51472
rect 19555 51471 19613 51472
rect 20995 51471 21053 51472
rect 3679 51388 3688 51428
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 4056 51388 4065 51428
rect 18799 51388 18808 51428
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 19176 51388 19185 51428
rect 163 51344 221 51345
rect 15043 51344 15101 51345
rect 21100 51344 21140 51556
rect 21424 51344 21504 51364
rect 163 51304 172 51344
rect 212 51304 5836 51344
rect 5876 51304 5885 51344
rect 11491 51304 11500 51344
rect 11540 51304 11828 51344
rect 163 51303 221 51304
rect 11788 51260 11828 51304
rect 15043 51304 15052 51344
rect 15092 51304 15340 51344
rect 15380 51304 15389 51344
rect 21100 51304 21504 51344
rect 15043 51303 15101 51304
rect 21424 51284 21504 51304
rect 7843 51220 7852 51260
rect 7892 51220 8524 51260
rect 8564 51220 8716 51260
rect 8756 51220 8765 51260
rect 11779 51220 11788 51260
rect 11828 51220 11837 51260
rect 15427 51220 15436 51260
rect 15476 51220 16204 51260
rect 16244 51220 16253 51260
rect 0 51176 80 51196
rect 4387 51176 4445 51177
rect 4579 51176 4637 51177
rect 0 51136 1324 51176
rect 1364 51136 1373 51176
rect 4302 51136 4396 51176
rect 4436 51136 4445 51176
rect 4494 51136 4588 51176
rect 4628 51136 4637 51176
rect 4771 51136 4780 51176
rect 4820 51136 7660 51176
rect 7700 51136 12692 51176
rect 12739 51136 12748 51176
rect 12788 51136 13708 51176
rect 13748 51136 13757 51176
rect 14755 51136 14764 51176
rect 14804 51136 15052 51176
rect 15092 51136 15101 51176
rect 0 51116 80 51136
rect 4387 51135 4445 51136
rect 4579 51135 4637 51136
rect 12652 51092 12692 51136
rect 3043 51052 3052 51092
rect 3092 51052 11404 51092
rect 11444 51052 11453 51092
rect 11779 51052 11788 51092
rect 11828 51052 12172 51092
rect 12212 51052 12221 51092
rect 12652 51052 16300 51092
rect 16340 51052 16349 51092
rect 21424 51008 21504 51028
rect 3235 50968 3244 51008
rect 3284 50968 3532 51008
rect 3572 50968 4492 51008
rect 4532 50968 4541 51008
rect 5923 50968 5932 51008
rect 5972 50968 6412 51008
rect 6452 50968 7660 51008
rect 7700 50968 11360 51008
rect 12067 50968 12076 51008
rect 12116 50968 13996 51008
rect 14036 50968 14045 51008
rect 14179 50968 14188 51008
rect 14228 50968 14956 51008
rect 14996 50968 15005 51008
rect 15523 50968 15532 51008
rect 15572 50968 15724 51008
rect 15764 50968 15773 51008
rect 17539 50968 17548 51008
rect 17588 50968 19564 51008
rect 19604 50968 19613 51008
rect 20131 50968 20140 51008
rect 20180 50968 21504 51008
rect 4099 50924 4157 50925
rect 10339 50924 10397 50925
rect 547 50884 556 50924
rect 596 50884 844 50924
rect 884 50884 893 50924
rect 4099 50884 4108 50924
rect 4148 50884 4204 50924
rect 4244 50884 4253 50924
rect 4387 50884 4396 50924
rect 4436 50884 5068 50924
rect 5108 50884 5117 50924
rect 10254 50884 10348 50924
rect 10388 50884 11212 50924
rect 11252 50884 11261 50924
rect 4099 50883 4157 50884
rect 10339 50883 10397 50884
rect 0 50840 80 50860
rect 11320 50840 11360 50968
rect 21424 50948 21504 50968
rect 19267 50924 19325 50925
rect 16291 50884 16300 50924
rect 16340 50884 19276 50924
rect 19316 50884 19325 50924
rect 19267 50883 19325 50884
rect 0 50800 8428 50840
rect 8468 50800 8477 50840
rect 11320 50800 18316 50840
rect 18356 50800 18365 50840
rect 0 50780 80 50800
rect 4387 50756 4445 50757
rect 6019 50756 6077 50757
rect 4387 50716 4396 50756
rect 4436 50716 5548 50756
rect 5588 50716 6028 50756
rect 6068 50716 7756 50756
rect 7796 50716 7805 50756
rect 8611 50716 8620 50756
rect 8660 50716 12268 50756
rect 12308 50716 12317 50756
rect 15715 50716 15724 50756
rect 15764 50716 17356 50756
rect 17396 50716 17548 50756
rect 17588 50716 17597 50756
rect 4387 50715 4445 50716
rect 6019 50715 6077 50716
rect 11683 50672 11741 50673
rect 21424 50672 21504 50692
rect 4919 50632 4928 50672
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 5296 50632 5305 50672
rect 11598 50632 11692 50672
rect 11732 50632 11741 50672
rect 20039 50632 20048 50672
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20416 50632 20425 50672
rect 20716 50632 21504 50672
rect 11683 50631 11741 50632
rect 20716 50588 20756 50632
rect 21424 50612 21504 50632
rect 10051 50548 10060 50588
rect 10100 50548 10636 50588
rect 10676 50548 11404 50588
rect 11444 50548 11453 50588
rect 11971 50548 11980 50588
rect 12020 50548 12364 50588
rect 12404 50548 12413 50588
rect 13987 50548 13996 50588
rect 14036 50548 15052 50588
rect 15092 50548 15101 50588
rect 19939 50548 19948 50588
rect 19988 50548 20756 50588
rect 0 50504 80 50524
rect 0 50464 1804 50504
rect 1844 50464 1853 50504
rect 2467 50464 2476 50504
rect 2516 50464 2540 50504
rect 5443 50464 5452 50504
rect 5492 50464 5740 50504
rect 5780 50464 5789 50504
rect 17731 50464 17740 50504
rect 17780 50464 18028 50504
rect 18068 50464 18077 50504
rect 0 50444 80 50464
rect 2500 50420 2540 50464
rect 17731 50420 17789 50421
rect 2500 50380 3956 50420
rect 10147 50380 10156 50420
rect 10196 50380 11212 50420
rect 11252 50380 11261 50420
rect 16579 50380 16588 50420
rect 16628 50380 17164 50420
rect 17204 50380 17213 50420
rect 17635 50380 17644 50420
rect 17684 50380 17740 50420
rect 17780 50380 17789 50420
rect 3916 50336 3956 50380
rect 17731 50379 17789 50380
rect 19267 50336 19325 50337
rect 21424 50336 21504 50356
rect 2659 50296 2668 50336
rect 2708 50296 3148 50336
rect 3188 50296 3197 50336
rect 3907 50296 3916 50336
rect 3956 50296 6124 50336
rect 6164 50296 7180 50336
rect 7220 50296 7229 50336
rect 7939 50296 7948 50336
rect 7988 50296 9004 50336
rect 9044 50296 9053 50336
rect 9187 50296 9196 50336
rect 9236 50296 9868 50336
rect 9908 50296 10348 50336
rect 10388 50296 10397 50336
rect 10819 50296 10828 50336
rect 10868 50296 11116 50336
rect 11156 50296 11165 50336
rect 12931 50296 12940 50336
rect 12980 50296 14380 50336
rect 14420 50296 14429 50336
rect 15907 50296 15916 50336
rect 15956 50296 16204 50336
rect 16244 50296 16253 50336
rect 16963 50296 16972 50336
rect 17012 50296 17932 50336
rect 17972 50296 17981 50336
rect 19171 50296 19180 50336
rect 19220 50296 19276 50336
rect 19316 50296 19325 50336
rect 19555 50296 19564 50336
rect 19604 50296 21504 50336
rect 1699 50252 1757 50253
rect 1614 50212 1708 50252
rect 1748 50212 1757 50252
rect 4291 50212 4300 50252
rect 4340 50212 4876 50252
rect 4916 50212 4925 50252
rect 1699 50211 1757 50212
rect 0 50168 80 50188
rect 5932 50168 5972 50296
rect 9004 50252 9044 50296
rect 19267 50295 19325 50296
rect 21424 50276 21504 50296
rect 9004 50212 9772 50252
rect 9812 50212 9821 50252
rect 13027 50212 13036 50252
rect 13076 50212 13085 50252
rect 13219 50212 13228 50252
rect 13268 50212 13516 50252
rect 13556 50212 13565 50252
rect 13036 50168 13076 50212
rect 0 50128 2860 50168
rect 2900 50128 2909 50168
rect 5923 50128 5932 50168
rect 5972 50128 5981 50168
rect 13036 50128 13420 50168
rect 13460 50128 13469 50168
rect 13795 50128 13804 50168
rect 13844 50128 14188 50168
rect 14228 50128 14237 50168
rect 16099 50128 16108 50168
rect 16148 50128 16396 50168
rect 16436 50128 16445 50168
rect 0 50108 80 50128
rect 10051 50044 10060 50084
rect 10100 50044 11884 50084
rect 11924 50044 14284 50084
rect 14324 50044 14333 50084
rect 14563 50044 14572 50084
rect 14612 50044 18604 50084
rect 18644 50044 18653 50084
rect 67 50000 125 50001
rect 21424 50000 21504 50020
rect 67 49960 76 50000
rect 116 49960 2476 50000
rect 2516 49960 2525 50000
rect 8323 49960 8332 50000
rect 8372 49960 15764 50000
rect 67 49959 125 49960
rect 1603 49876 1612 49916
rect 1652 49876 1996 49916
rect 2036 49876 2045 49916
rect 3679 49876 3688 49916
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 4056 49876 4065 49916
rect 8899 49876 8908 49916
rect 8948 49876 12596 49916
rect 12643 49876 12652 49916
rect 12692 49876 13036 49916
rect 13076 49876 13085 49916
rect 0 49832 80 49852
rect 12556 49832 12596 49876
rect 15724 49832 15764 49960
rect 20140 49960 21504 50000
rect 20140 49917 20180 49960
rect 21424 49940 21504 49960
rect 20131 49916 20189 49917
rect 18799 49876 18808 49916
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 19176 49876 19185 49916
rect 20131 49876 20140 49916
rect 20180 49876 20189 49916
rect 20131 49875 20189 49876
rect 0 49792 1516 49832
rect 1556 49792 1565 49832
rect 8131 49792 8140 49832
rect 8180 49792 8428 49832
rect 8468 49792 9484 49832
rect 9524 49792 10060 49832
rect 10100 49792 10109 49832
rect 12556 49792 14572 49832
rect 14612 49792 14621 49832
rect 15724 49792 21388 49832
rect 21428 49792 21437 49832
rect 0 49772 80 49792
rect 1891 49748 1949 49749
rect 15619 49748 15677 49749
rect 1891 49708 1900 49748
rect 1940 49708 2540 49748
rect 4099 49708 4108 49748
rect 4148 49708 4684 49748
rect 4724 49708 4733 49748
rect 5635 49708 5644 49748
rect 5684 49708 5932 49748
rect 5972 49708 5981 49748
rect 8515 49708 8524 49748
rect 8564 49708 15628 49748
rect 15668 49708 15677 49748
rect 1891 49707 1949 49708
rect 2500 49664 2540 49708
rect 15619 49707 15677 49708
rect 10435 49664 10493 49665
rect 20707 49664 20765 49665
rect 21424 49664 21504 49684
rect 2500 49624 6700 49664
rect 6740 49624 10444 49664
rect 10484 49624 10493 49664
rect 11971 49624 11980 49664
rect 12020 49624 16340 49664
rect 10435 49623 10493 49624
rect 16300 49580 16340 49624
rect 20707 49624 20716 49664
rect 20756 49624 21504 49664
rect 20707 49623 20765 49624
rect 21424 49604 21504 49624
rect 1411 49540 1420 49580
rect 1460 49540 9004 49580
rect 9044 49540 11156 49580
rect 16291 49540 16300 49580
rect 16340 49540 16349 49580
rect 0 49496 80 49516
rect 9667 49496 9725 49497
rect 0 49456 1900 49496
rect 1940 49456 1949 49496
rect 4579 49456 4588 49496
rect 4628 49456 6028 49496
rect 6068 49456 9484 49496
rect 9524 49456 9676 49496
rect 9716 49456 9725 49496
rect 9859 49456 9868 49496
rect 9908 49456 10540 49496
rect 10580 49456 11020 49496
rect 11060 49456 11069 49496
rect 0 49436 80 49456
rect 9667 49455 9725 49456
rect 11116 49412 11156 49540
rect 13603 49456 13612 49496
rect 13652 49456 13804 49496
rect 13844 49456 13996 49496
rect 14036 49456 14045 49496
rect 14275 49456 14284 49496
rect 14324 49456 16588 49496
rect 16628 49456 19084 49496
rect 19124 49456 19133 49496
rect 10147 49372 10156 49412
rect 10196 49372 10828 49412
rect 10868 49372 10877 49412
rect 11116 49372 18124 49412
rect 18164 49372 18173 49412
rect 18499 49372 18508 49412
rect 18548 49372 18557 49412
rect 18508 49328 18548 49372
rect 1699 49288 1708 49328
rect 1748 49288 4492 49328
rect 4532 49288 4541 49328
rect 5827 49288 5836 49328
rect 5876 49288 18548 49328
rect 18595 49328 18653 49329
rect 20515 49328 20573 49329
rect 21424 49328 21504 49348
rect 18595 49288 18604 49328
rect 18644 49288 20524 49328
rect 20564 49288 20573 49328
rect 21379 49288 21388 49328
rect 21428 49288 21504 49328
rect 18595 49287 18653 49288
rect 20515 49287 20573 49288
rect 21424 49268 21504 49288
rect 13699 49244 13757 49245
rect 3811 49204 3820 49244
rect 3860 49204 5644 49244
rect 5684 49204 5693 49244
rect 8995 49204 9004 49244
rect 9044 49204 11212 49244
rect 11252 49204 11261 49244
rect 13603 49204 13612 49244
rect 13652 49204 13708 49244
rect 13748 49204 13757 49244
rect 13699 49203 13757 49204
rect 14467 49244 14525 49245
rect 14467 49204 14476 49244
rect 14516 49204 14764 49244
rect 14804 49204 14813 49244
rect 14467 49203 14525 49204
rect 0 49160 80 49180
rect 10435 49160 10493 49161
rect 0 49120 1324 49160
rect 1364 49120 1373 49160
rect 4919 49120 4928 49160
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 5296 49120 5305 49160
rect 9475 49120 9484 49160
rect 9524 49120 9772 49160
rect 9812 49120 9821 49160
rect 10435 49120 10444 49160
rect 10484 49120 11020 49160
rect 11060 49120 11069 49160
rect 11395 49120 11404 49160
rect 11444 49120 13996 49160
rect 14036 49120 14045 49160
rect 16387 49120 16396 49160
rect 16436 49120 17740 49160
rect 17780 49120 17789 49160
rect 18115 49120 18124 49160
rect 18164 49120 18412 49160
rect 18452 49120 18461 49160
rect 20039 49120 20048 49160
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20416 49120 20425 49160
rect 0 49100 80 49120
rect 10435 49119 10493 49120
rect 7171 49036 7180 49076
rect 7220 49036 7564 49076
rect 7604 49036 7613 49076
rect 7939 49036 7948 49076
rect 7988 49036 9676 49076
rect 9716 49036 9725 49076
rect 10627 49036 10636 49076
rect 10676 49036 10685 49076
rect 16483 49036 16492 49076
rect 16532 49036 17068 49076
rect 17108 49036 17117 49076
rect 10636 48992 10676 49036
rect 14659 48992 14717 48993
rect 15715 48992 15773 48993
rect 21424 48992 21504 49012
rect 8227 48952 8236 48992
rect 8276 48952 10676 48992
rect 14574 48952 14668 48992
rect 14708 48952 15724 48992
rect 15764 48952 18316 48992
rect 18356 48952 18365 48992
rect 21283 48952 21292 48992
rect 21332 48952 21504 48992
rect 14659 48951 14717 48952
rect 15715 48951 15773 48952
rect 21424 48932 21504 48952
rect 2572 48868 10676 48908
rect 11203 48868 11212 48908
rect 11252 48868 13172 48908
rect 0 48824 80 48844
rect 2572 48824 2612 48868
rect 10339 48824 10397 48825
rect 10636 48824 10676 48868
rect 13132 48824 13172 48868
rect 13219 48824 13277 48825
rect 16579 48824 16637 48825
rect 0 48784 1612 48824
rect 1652 48784 1661 48824
rect 2563 48784 2572 48824
rect 2612 48784 2621 48824
rect 3331 48784 3340 48824
rect 3380 48784 5356 48824
rect 5396 48784 6508 48824
rect 6548 48784 6796 48824
rect 6836 48784 6845 48824
rect 8035 48784 8044 48824
rect 8084 48784 9388 48824
rect 9428 48784 9437 48824
rect 10254 48784 10348 48824
rect 10388 48784 10397 48824
rect 10627 48784 10636 48824
rect 10676 48784 11360 48824
rect 11587 48784 11596 48824
rect 11636 48784 11884 48824
rect 11924 48784 11933 48824
rect 13123 48784 13132 48824
rect 13172 48784 13228 48824
rect 13268 48784 13277 48824
rect 14371 48784 14380 48824
rect 14420 48784 15052 48824
rect 15092 48784 15101 48824
rect 15523 48784 15532 48824
rect 15572 48784 15916 48824
rect 15956 48784 15965 48824
rect 16494 48784 16588 48824
rect 16628 48784 16637 48824
rect 0 48764 80 48784
rect 10339 48783 10397 48784
rect 11320 48740 11360 48784
rect 13219 48783 13277 48784
rect 16579 48783 16637 48784
rect 15715 48740 15773 48741
rect 4195 48700 4204 48740
rect 4244 48700 4780 48740
rect 4820 48700 8428 48740
rect 8468 48700 11212 48740
rect 11252 48700 11261 48740
rect 11320 48700 11980 48740
rect 12020 48700 12029 48740
rect 15630 48700 15724 48740
rect 15764 48700 15773 48740
rect 15715 48699 15773 48700
rect 20899 48656 20957 48657
rect 21424 48656 21504 48676
rect 2467 48616 2476 48656
rect 2516 48616 16012 48656
rect 16052 48616 16061 48656
rect 20899 48616 20908 48656
rect 20948 48616 21504 48656
rect 20899 48615 20957 48616
rect 21424 48596 21504 48616
rect 4003 48532 4012 48572
rect 4052 48532 4300 48572
rect 4340 48532 4349 48572
rect 14275 48532 14284 48572
rect 14324 48532 14572 48572
rect 14612 48532 14621 48572
rect 0 48488 80 48508
rect 1987 48488 2045 48489
rect 0 48448 1996 48488
rect 2036 48448 2045 48488
rect 0 48428 80 48448
rect 1987 48447 2045 48448
rect 3679 48364 3688 48404
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 4056 48364 4065 48404
rect 4771 48364 4780 48404
rect 4820 48364 6316 48404
rect 6356 48364 11788 48404
rect 11828 48364 11837 48404
rect 16483 48364 16492 48404
rect 16532 48364 16972 48404
rect 17012 48364 18124 48404
rect 18164 48364 18173 48404
rect 18799 48364 18808 48404
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 19176 48364 19185 48404
rect 21424 48320 21504 48340
rect 7651 48280 7660 48320
rect 7700 48280 10252 48320
rect 10292 48280 11360 48320
rect 17251 48280 17260 48320
rect 17300 48280 21504 48320
rect 11320 48236 11360 48280
rect 21424 48260 21504 48280
rect 19459 48236 19517 48237
rect 6019 48196 6028 48236
rect 6068 48196 6316 48236
rect 6356 48196 6604 48236
rect 6644 48196 6653 48236
rect 11320 48196 11596 48236
rect 11636 48196 12172 48236
rect 12212 48196 12221 48236
rect 19267 48196 19276 48236
rect 19316 48196 19468 48236
rect 19508 48196 19517 48236
rect 19459 48195 19517 48196
rect 0 48152 80 48172
rect 3139 48152 3197 48153
rect 0 48112 3148 48152
rect 3188 48112 3197 48152
rect 7171 48112 7180 48152
rect 7220 48112 11360 48152
rect 11875 48112 11884 48152
rect 11924 48112 21332 48152
rect 0 48092 80 48112
rect 3139 48111 3197 48112
rect 8707 48068 8765 48069
rect 1699 48028 1708 48068
rect 1748 48028 7948 48068
rect 7988 48028 7997 48068
rect 8622 48028 8716 48068
rect 8756 48028 8765 48068
rect 8707 48027 8765 48028
rect 3139 47984 3197 47985
rect 3139 47944 3148 47984
rect 3188 47944 3244 47984
rect 3284 47944 3293 47984
rect 6403 47944 6412 47984
rect 6452 47944 7180 47984
rect 7220 47944 7229 47984
rect 8227 47944 8236 47984
rect 8276 47944 8620 47984
rect 8660 47944 8669 47984
rect 8803 47944 8812 47984
rect 8852 47944 10924 47984
rect 10964 47944 10973 47984
rect 3139 47943 3197 47944
rect 11320 47900 11360 48112
rect 13987 48028 13996 48068
rect 14036 48028 14380 48068
rect 14420 48028 16588 48068
rect 16628 48028 16637 48068
rect 21292 47984 21332 48112
rect 21424 47984 21504 48004
rect 13603 47944 13612 47984
rect 13652 47944 13804 47984
rect 13844 47944 13853 47984
rect 15907 47944 15916 47984
rect 15956 47944 16492 47984
rect 16532 47944 17260 47984
rect 17300 47944 17309 47984
rect 17827 47944 17836 47984
rect 17876 47944 19372 47984
rect 19412 47944 19421 47984
rect 21292 47944 21504 47984
rect 21424 47924 21504 47944
rect 18499 47900 18557 47901
rect 1795 47860 1804 47900
rect 1844 47860 4492 47900
rect 4532 47860 4541 47900
rect 6307 47860 6316 47900
rect 6356 47860 11212 47900
rect 11252 47860 11261 47900
rect 11308 47860 18508 47900
rect 18548 47860 18557 47900
rect 0 47816 80 47836
rect 0 47776 1420 47816
rect 1460 47776 1469 47816
rect 3811 47776 3820 47816
rect 3860 47776 4108 47816
rect 4148 47776 6988 47816
rect 7028 47776 7037 47816
rect 0 47756 80 47776
rect 2083 47692 2092 47732
rect 2132 47692 9868 47732
rect 9908 47692 9917 47732
rect 11308 47648 11348 47860
rect 18499 47859 18557 47860
rect 15427 47776 15436 47816
rect 15476 47776 16108 47816
rect 16148 47776 16157 47816
rect 16291 47776 16300 47816
rect 16340 47776 16972 47816
rect 17012 47776 17021 47816
rect 16291 47732 16349 47733
rect 16291 47692 16300 47732
rect 16340 47692 20564 47732
rect 16291 47691 16349 47692
rect 20524 47648 20564 47692
rect 21424 47648 21504 47668
rect 4919 47608 4928 47648
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 5296 47608 5305 47648
rect 6019 47608 6028 47648
rect 6068 47608 7660 47648
rect 7700 47608 7709 47648
rect 11011 47608 11020 47648
rect 11060 47608 11348 47648
rect 20039 47608 20048 47648
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20416 47608 20425 47648
rect 20524 47608 21504 47648
rect 21424 47588 21504 47608
rect 18307 47524 18316 47564
rect 18356 47524 19372 47564
rect 19412 47524 19421 47564
rect 0 47480 80 47500
rect 0 47440 1900 47480
rect 1940 47440 1949 47480
rect 2179 47440 2188 47480
rect 2228 47440 12076 47480
rect 12116 47440 12125 47480
rect 14947 47440 14956 47480
rect 14996 47440 18892 47480
rect 18932 47440 18941 47480
rect 0 47420 80 47440
rect 3331 47356 3340 47396
rect 3380 47356 3820 47396
rect 3860 47356 3869 47396
rect 6979 47356 6988 47396
rect 7028 47356 7276 47396
rect 7316 47356 11404 47396
rect 11444 47356 11453 47396
rect 13507 47356 13516 47396
rect 13556 47356 16300 47396
rect 16340 47356 16349 47396
rect 20035 47356 20044 47396
rect 20084 47356 21292 47396
rect 21332 47356 21341 47396
rect 1891 47312 1949 47313
rect 4099 47312 4157 47313
rect 16579 47312 16637 47313
rect 20707 47312 20765 47313
rect 21424 47312 21504 47332
rect 1806 47272 1900 47312
rect 1940 47272 1949 47312
rect 3907 47272 3916 47312
rect 3956 47272 4108 47312
rect 4148 47272 4157 47312
rect 4291 47272 4300 47312
rect 4340 47272 7700 47312
rect 10147 47272 10156 47312
rect 10196 47272 10924 47312
rect 10964 47272 10973 47312
rect 12259 47272 12268 47312
rect 12308 47272 14188 47312
rect 14228 47272 14237 47312
rect 14467 47272 14476 47312
rect 14516 47272 16492 47312
rect 16532 47272 16588 47312
rect 16628 47272 16637 47312
rect 17923 47272 17932 47312
rect 17972 47272 18316 47312
rect 18356 47272 18365 47312
rect 18499 47272 18508 47312
rect 18548 47272 18796 47312
rect 18836 47272 18845 47312
rect 19555 47272 19564 47312
rect 19604 47272 20716 47312
rect 20756 47272 20765 47312
rect 20899 47272 20908 47312
rect 20948 47272 21504 47312
rect 1891 47271 1949 47272
rect 4099 47271 4157 47272
rect 7660 47228 7700 47272
rect 10819 47228 10877 47229
rect 1699 47188 1708 47228
rect 1748 47188 7564 47228
rect 7604 47188 7613 47228
rect 7660 47188 10828 47228
rect 10868 47188 10877 47228
rect 10924 47228 10964 47272
rect 14476 47228 14516 47272
rect 16579 47271 16637 47272
rect 20707 47271 20765 47272
rect 21424 47252 21504 47272
rect 10924 47188 14516 47228
rect 10819 47187 10877 47188
rect 0 47144 80 47164
rect 8323 47144 8381 47145
rect 0 47104 652 47144
rect 692 47104 701 47144
rect 6595 47104 6604 47144
rect 6644 47104 8332 47144
rect 8372 47104 10060 47144
rect 10100 47104 10109 47144
rect 11683 47104 11692 47144
rect 11732 47104 19316 47144
rect 0 47084 80 47104
rect 8323 47103 8381 47104
rect 7843 47060 7901 47061
rect 7843 47020 7852 47060
rect 7892 47020 12940 47060
rect 12980 47020 12989 47060
rect 18700 47020 18892 47060
rect 18932 47020 18941 47060
rect 7843 47019 7901 47020
rect 2851 46936 2860 46976
rect 2900 46936 10444 46976
rect 10484 46936 10493 46976
rect 13411 46892 13469 46893
rect 3679 46852 3688 46892
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 4056 46852 4065 46892
rect 9763 46852 9772 46892
rect 9812 46852 9964 46892
rect 10004 46852 10013 46892
rect 12931 46852 12940 46892
rect 12980 46852 13420 46892
rect 13460 46852 13469 46892
rect 13411 46851 13469 46852
rect 0 46808 80 46828
rect 0 46768 2284 46808
rect 2324 46768 2333 46808
rect 4387 46768 4396 46808
rect 4436 46768 8428 46808
rect 8468 46768 8716 46808
rect 8756 46768 8765 46808
rect 16579 46768 16588 46808
rect 16628 46768 17164 46808
rect 17204 46768 17213 46808
rect 0 46748 80 46768
rect 1123 46724 1181 46725
rect 18700 46724 18740 47020
rect 18799 46852 18808 46892
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 19176 46852 19185 46892
rect 19276 46808 19316 47104
rect 21424 46976 21504 46996
rect 19939 46936 19948 46976
rect 19988 46936 21504 46976
rect 21424 46916 21504 46936
rect 19276 46768 20180 46808
rect 940 46684 1132 46724
rect 1172 46684 1181 46724
rect 940 46641 980 46684
rect 1123 46683 1181 46684
rect 2500 46684 3148 46724
rect 3188 46684 3197 46724
rect 7660 46684 9676 46724
rect 9716 46684 9964 46724
rect 10004 46684 10013 46724
rect 18700 46684 18988 46724
rect 19028 46684 19037 46724
rect 931 46640 989 46641
rect 2500 46640 2540 46684
rect 7660 46640 7700 46684
rect 20140 46640 20180 46768
rect 21424 46640 21504 46660
rect 931 46600 940 46640
rect 980 46600 989 46640
rect 2467 46600 2476 46640
rect 2516 46600 2540 46640
rect 7620 46600 7660 46640
rect 7700 46600 7709 46640
rect 20140 46600 21504 46640
rect 931 46599 989 46600
rect 21424 46580 21504 46600
rect 2755 46556 2813 46557
rect 2755 46516 2764 46556
rect 2804 46516 3052 46556
rect 3092 46516 3101 46556
rect 3427 46516 3436 46556
rect 3476 46516 5548 46556
rect 5588 46516 5597 46556
rect 2755 46515 2813 46516
rect 0 46472 80 46492
rect 6883 46472 6941 46473
rect 0 46432 3244 46472
rect 3284 46432 3293 46472
rect 6403 46432 6412 46472
rect 6452 46432 6892 46472
rect 6932 46432 6941 46472
rect 0 46412 80 46432
rect 6883 46431 6941 46432
rect 10531 46472 10589 46473
rect 11875 46472 11933 46473
rect 15715 46472 15773 46473
rect 10531 46432 10540 46472
rect 10580 46432 10924 46472
rect 10964 46432 10973 46472
rect 11875 46432 11884 46472
rect 11924 46432 13132 46472
rect 13172 46432 13181 46472
rect 14947 46432 14956 46472
rect 14996 46432 15724 46472
rect 15764 46432 16972 46472
rect 17012 46432 17356 46472
rect 17396 46432 17405 46472
rect 10531 46431 10589 46432
rect 11875 46431 11933 46432
rect 15715 46431 15773 46432
rect 7747 46388 7805 46389
rect 1411 46348 1420 46388
rect 1460 46348 7756 46388
rect 7796 46348 7805 46388
rect 10243 46348 10252 46388
rect 10292 46348 15724 46388
rect 15764 46348 15773 46388
rect 7747 46347 7805 46348
rect 9763 46304 9821 46305
rect 21424 46304 21504 46324
rect 1315 46264 1324 46304
rect 1364 46264 9004 46304
rect 9044 46264 9053 46304
rect 9763 46264 9772 46304
rect 9812 46264 21504 46304
rect 9763 46263 9821 46264
rect 21424 46244 21504 46264
rect 3331 46180 3340 46220
rect 3380 46180 5356 46220
rect 5396 46180 6028 46220
rect 6068 46180 6077 46220
rect 12547 46180 12556 46220
rect 12596 46180 13228 46220
rect 13268 46180 13277 46220
rect 0 46136 80 46156
rect 0 46096 1516 46136
rect 1556 46096 1565 46136
rect 4919 46096 4928 46136
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 5296 46096 5305 46136
rect 11395 46096 11404 46136
rect 11444 46096 19372 46136
rect 19412 46096 19421 46136
rect 20039 46096 20048 46136
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20416 46096 20425 46136
rect 0 46076 80 46096
rect 11779 46012 11788 46052
rect 11828 46012 12172 46052
rect 12212 46012 17452 46052
rect 17492 46012 17836 46052
rect 17876 46012 17885 46052
rect 21424 45968 21504 45988
rect 7756 45928 13748 45968
rect 18403 45928 18412 45968
rect 18452 45928 18796 45968
rect 18836 45928 18845 45968
rect 20803 45928 20812 45968
rect 20852 45928 21504 45968
rect 7756 45884 7796 45928
rect 2500 45844 2860 45884
rect 2900 45844 2909 45884
rect 6115 45844 6124 45884
rect 6164 45844 7756 45884
rect 7796 45844 7805 45884
rect 8131 45844 8140 45884
rect 8180 45844 10252 45884
rect 10292 45844 10301 45884
rect 0 45800 80 45820
rect 2500 45800 2540 45844
rect 7843 45800 7901 45801
rect 13708 45800 13748 45928
rect 21424 45908 21504 45928
rect 19459 45844 19468 45884
rect 19508 45844 19756 45884
rect 19796 45844 19805 45884
rect 0 45760 2540 45800
rect 4099 45760 4108 45800
rect 4148 45760 4396 45800
rect 4436 45760 7852 45800
rect 7892 45760 8716 45800
rect 8756 45760 8765 45800
rect 13699 45760 13708 45800
rect 13748 45760 13757 45800
rect 17347 45760 17356 45800
rect 17396 45760 18700 45800
rect 18740 45760 18749 45800
rect 0 45740 80 45760
rect 7843 45759 7901 45760
rect 6403 45676 6412 45716
rect 6452 45676 19756 45716
rect 19796 45676 19805 45716
rect 21424 45632 21504 45652
rect 1987 45592 1996 45632
rect 2036 45592 10348 45632
rect 10388 45592 10924 45632
rect 10964 45592 10973 45632
rect 17347 45592 17356 45632
rect 17396 45592 21504 45632
rect 21424 45572 21504 45592
rect 12547 45548 12605 45549
rect 19939 45548 19997 45549
rect 2500 45508 2668 45548
rect 2708 45508 2717 45548
rect 12547 45508 12556 45548
rect 12596 45508 19564 45548
rect 19604 45508 19613 45548
rect 19854 45508 19948 45548
rect 19988 45508 19997 45548
rect 0 45464 80 45484
rect 2500 45464 2540 45508
rect 12547 45507 12605 45508
rect 19939 45507 19997 45508
rect 0 45424 2540 45464
rect 3532 45424 7276 45464
rect 7316 45424 7660 45464
rect 7700 45424 7709 45464
rect 18691 45424 18700 45464
rect 18740 45424 19756 45464
rect 19796 45424 19805 45464
rect 0 45404 80 45424
rect 3532 45380 3572 45424
rect 8131 45380 8189 45381
rect 11971 45380 12029 45381
rect 1603 45340 1612 45380
rect 1652 45340 2380 45380
rect 2420 45340 3572 45380
rect 3679 45340 3688 45380
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 4056 45340 4065 45380
rect 4771 45340 4780 45380
rect 4820 45340 7084 45380
rect 7124 45340 7133 45380
rect 7363 45340 7372 45380
rect 7412 45340 8140 45380
rect 8180 45340 8189 45380
rect 11587 45340 11596 45380
rect 11636 45340 11980 45380
rect 12020 45340 12029 45380
rect 16195 45340 16204 45380
rect 16244 45340 16972 45380
rect 17012 45340 17021 45380
rect 18799 45340 18808 45380
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 19176 45340 19185 45380
rect 7084 45296 7124 45340
rect 8131 45339 8189 45340
rect 11971 45339 12029 45340
rect 17155 45296 17213 45297
rect 21424 45296 21504 45316
rect 7084 45256 8908 45296
rect 8948 45256 9196 45296
rect 9236 45256 9245 45296
rect 9955 45256 9964 45296
rect 10004 45256 11500 45296
rect 11540 45256 11692 45296
rect 11732 45256 13420 45296
rect 13460 45256 13469 45296
rect 17155 45256 17164 45296
rect 17204 45256 21504 45296
rect 17155 45255 17213 45256
rect 21424 45236 21504 45256
rect 15907 45212 15965 45213
rect 2755 45172 2764 45212
rect 2804 45172 3916 45212
rect 3956 45172 3965 45212
rect 15907 45172 15916 45212
rect 15956 45172 18316 45212
rect 18356 45172 18365 45212
rect 15907 45171 15965 45172
rect 0 45128 80 45148
rect 10531 45128 10589 45129
rect 0 45088 1516 45128
rect 1556 45088 1565 45128
rect 6883 45088 6892 45128
rect 6932 45088 9716 45128
rect 10435 45088 10444 45128
rect 10484 45088 10540 45128
rect 10580 45088 10589 45128
rect 0 45068 80 45088
rect 1795 45004 1804 45044
rect 1844 45004 9580 45044
rect 9620 45004 9629 45044
rect 7939 44960 7997 44961
rect 9676 44960 9716 45088
rect 10531 45087 10589 45088
rect 16099 45044 16157 45045
rect 16003 45004 16012 45044
rect 16052 45004 16108 45044
rect 16148 45004 16157 45044
rect 16099 45003 16157 45004
rect 10627 44960 10685 44961
rect 18499 44960 18557 44961
rect 3235 44920 3244 44960
rect 3284 44920 5644 44960
rect 5684 44920 5836 44960
rect 5876 44920 5885 44960
rect 7854 44920 7948 44960
rect 7988 44920 8236 44960
rect 8276 44920 8285 44960
rect 9676 44920 10636 44960
rect 10676 44920 10685 44960
rect 18414 44920 18508 44960
rect 18548 44920 18557 44960
rect 7939 44919 7997 44920
rect 10627 44919 10685 44920
rect 18499 44919 18557 44920
rect 20131 44960 20189 44961
rect 21424 44960 21504 44980
rect 20131 44920 20140 44960
rect 20180 44920 21504 44960
rect 20131 44919 20189 44920
rect 21424 44900 21504 44920
rect 8323 44876 8381 44877
rect 2083 44836 2092 44876
rect 2132 44836 5452 44876
rect 5492 44836 5501 44876
rect 8238 44836 8332 44876
rect 8372 44836 8620 44876
rect 8660 44836 8669 44876
rect 8323 44835 8381 44836
rect 0 44792 80 44812
rect 4099 44792 4157 44793
rect 0 44752 1612 44792
rect 1652 44752 1661 44792
rect 3811 44752 3820 44792
rect 3860 44752 4108 44792
rect 4148 44752 12652 44792
rect 12692 44752 12701 44792
rect 0 44732 80 44752
rect 4099 44751 4157 44752
rect 10915 44708 10973 44709
rect 10915 44668 10924 44708
rect 10964 44668 17932 44708
rect 17972 44668 17981 44708
rect 10915 44667 10973 44668
rect 21424 44624 21504 44644
rect 4919 44584 4928 44624
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 5296 44584 5305 44624
rect 20039 44584 20048 44624
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20416 44584 20425 44624
rect 20707 44584 20716 44624
rect 20756 44584 21504 44624
rect 21424 44564 21504 44584
rect 13795 44540 13853 44541
rect 6892 44500 11884 44540
rect 11924 44500 11933 44540
rect 13795 44500 13804 44540
rect 13844 44500 18316 44540
rect 18356 44500 18365 44540
rect 0 44456 80 44476
rect 0 44416 1228 44456
rect 1268 44416 1277 44456
rect 4291 44416 4300 44456
rect 4340 44416 4876 44456
rect 4916 44416 4925 44456
rect 0 44396 80 44416
rect 2467 44332 2476 44372
rect 2516 44332 5548 44372
rect 5588 44332 5597 44372
rect 3427 44248 3436 44288
rect 3476 44248 3820 44288
rect 3860 44248 3869 44288
rect 6892 44204 6932 44500
rect 13795 44499 13853 44500
rect 10147 44456 10205 44457
rect 10147 44416 10156 44456
rect 10196 44416 18124 44456
rect 18164 44416 18173 44456
rect 10147 44415 10205 44416
rect 21424 44288 21504 44308
rect 9379 44248 9388 44288
rect 9428 44248 9964 44288
rect 10004 44248 10013 44288
rect 12067 44248 12076 44288
rect 12116 44248 12748 44288
rect 12788 44248 13228 44288
rect 13268 44248 13277 44288
rect 15043 44248 15052 44288
rect 15092 44248 15476 44288
rect 16195 44248 16204 44288
rect 16244 44248 19852 44288
rect 19892 44248 19901 44288
rect 20515 44248 20524 44288
rect 20564 44248 21504 44288
rect 1795 44164 1804 44204
rect 1844 44164 6932 44204
rect 8227 44204 8285 44205
rect 12451 44204 12509 44205
rect 15043 44204 15101 44205
rect 15436 44204 15476 44248
rect 21424 44228 21504 44248
rect 8227 44164 8236 44204
rect 8276 44164 12460 44204
rect 12500 44164 12509 44204
rect 12643 44164 12652 44204
rect 12692 44164 13036 44204
rect 13076 44164 13085 44204
rect 15043 44164 15052 44204
rect 15092 44164 15148 44204
rect 15188 44164 15197 44204
rect 15427 44164 15436 44204
rect 15476 44164 15485 44204
rect 8227 44163 8285 44164
rect 12451 44163 12509 44164
rect 15043 44163 15101 44164
rect 0 44120 80 44140
rect 17347 44120 17405 44121
rect 0 44080 14956 44120
rect 14996 44080 15005 44120
rect 17262 44080 17356 44120
rect 17396 44080 17405 44120
rect 19555 44080 19564 44120
rect 19604 44080 20620 44120
rect 20660 44080 20669 44120
rect 0 44060 80 44080
rect 17347 44079 17405 44080
rect 19459 44036 19517 44037
rect 19459 43996 19468 44036
rect 19508 43996 19756 44036
rect 19796 43996 19805 44036
rect 19459 43995 19517 43996
rect 21424 43952 21504 43972
rect 17539 43912 17548 43952
rect 17588 43912 21504 43952
rect 21424 43892 21504 43912
rect 3679 43828 3688 43868
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 4056 43828 4065 43868
rect 18799 43828 18808 43868
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 19176 43828 19185 43868
rect 0 43784 80 43804
rect 2083 43784 2141 43785
rect 0 43744 1612 43784
rect 1652 43744 1661 43784
rect 2083 43744 2092 43784
rect 2132 43744 19756 43784
rect 19796 43744 19805 43784
rect 0 43724 80 43744
rect 2083 43743 2141 43744
rect 2467 43700 2525 43701
rect 6883 43700 6941 43701
rect 18403 43700 18461 43701
rect 19747 43700 19805 43701
rect 2467 43660 2476 43700
rect 2516 43660 6412 43700
rect 6452 43660 6461 43700
rect 6883 43660 6892 43700
rect 6932 43660 7084 43700
rect 7124 43660 7133 43700
rect 13411 43660 13420 43700
rect 13460 43660 17740 43700
rect 17780 43660 17789 43700
rect 18403 43660 18412 43700
rect 18452 43660 18796 43700
rect 18836 43660 18845 43700
rect 19747 43660 19756 43700
rect 19796 43660 19948 43700
rect 19988 43660 19997 43700
rect 21292 43660 21428 43700
rect 2467 43659 2525 43660
rect 6883 43659 6941 43660
rect 18403 43659 18461 43660
rect 19747 43659 19805 43660
rect 172 43576 13132 43616
rect 13172 43576 13181 43616
rect 0 43448 80 43468
rect 0 43388 116 43448
rect 76 43364 116 43388
rect 172 43364 212 43576
rect 4771 43532 4829 43533
rect 4771 43492 4780 43532
rect 4820 43492 9388 43532
rect 9428 43492 9437 43532
rect 10915 43492 10924 43532
rect 10964 43492 17548 43532
rect 17588 43492 17597 43532
rect 4771 43491 4829 43492
rect 21292 43448 21332 43660
rect 21388 43636 21428 43660
rect 21388 43576 21504 43636
rect 21424 43556 21504 43576
rect 2467 43408 2476 43448
rect 2516 43408 3436 43448
rect 3476 43408 3485 43448
rect 6307 43408 6316 43448
rect 6356 43408 6604 43448
rect 6644 43408 6653 43448
rect 6787 43408 6796 43448
rect 6836 43408 8236 43448
rect 8276 43408 8285 43448
rect 15235 43408 15244 43448
rect 15284 43408 16204 43448
rect 16244 43408 16253 43448
rect 17443 43408 17452 43448
rect 17492 43408 21332 43448
rect 2179 43364 2237 43365
rect 76 43324 212 43364
rect 2094 43324 2188 43364
rect 2228 43324 6932 43364
rect 7171 43324 7180 43364
rect 7220 43324 7372 43364
rect 7412 43324 7421 43364
rect 8419 43324 8428 43364
rect 8468 43324 18604 43364
rect 18644 43324 18653 43364
rect 2179 43323 2237 43324
rect 4099 43280 4157 43281
rect 4003 43240 4012 43280
rect 4052 43240 4108 43280
rect 4148 43240 4157 43280
rect 6892 43280 6932 43324
rect 12355 43280 12413 43281
rect 20899 43280 20957 43281
rect 21424 43280 21504 43300
rect 6892 43240 11360 43280
rect 4099 43239 4157 43240
rect 7363 43196 7421 43197
rect 11320 43196 11360 43240
rect 12355 43240 12364 43280
rect 12404 43240 19180 43280
rect 19220 43240 19229 43280
rect 20899 43240 20908 43280
rect 20948 43240 21504 43280
rect 12355 43239 12413 43240
rect 20899 43239 20957 43240
rect 21424 43220 21504 43240
rect 18595 43196 18653 43197
rect 2083 43156 2092 43196
rect 2132 43156 3916 43196
rect 3956 43156 3965 43196
rect 6883 43156 6892 43196
rect 6932 43156 7372 43196
rect 7412 43156 7421 43196
rect 7939 43156 7948 43196
rect 7988 43156 8524 43196
rect 8564 43156 8573 43196
rect 11320 43156 18604 43196
rect 18644 43156 19372 43196
rect 19412 43156 19421 43196
rect 7363 43155 7421 43156
rect 18595 43155 18653 43156
rect 0 43112 80 43132
rect 0 43072 3724 43112
rect 3764 43072 3773 43112
rect 4919 43072 4928 43112
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 5296 43072 5305 43112
rect 5347 43072 5356 43112
rect 5396 43072 8428 43112
rect 8468 43072 8477 43112
rect 20039 43072 20048 43112
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20416 43072 20425 43112
rect 0 43052 80 43072
rect 2371 43028 2429 43029
rect 6211 43028 6269 43029
rect 2371 42988 2380 43028
rect 2420 42988 3532 43028
rect 3572 42988 5548 43028
rect 5588 42988 5597 43028
rect 6211 42988 6220 43028
rect 6260 42988 11360 43028
rect 2371 42987 2429 42988
rect 6211 42987 6269 42988
rect 11320 42944 11360 42988
rect 21424 42944 21504 42964
rect 3715 42904 3724 42944
rect 3764 42904 6644 42944
rect 6979 42904 6988 42944
rect 7028 42904 7372 42944
rect 7412 42904 7421 42944
rect 11320 42904 18124 42944
rect 18164 42904 18173 42944
rect 20899 42904 20908 42944
rect 20948 42904 21504 42944
rect 6499 42860 6557 42861
rect 3139 42820 3148 42860
rect 3188 42820 4684 42860
rect 4724 42820 4733 42860
rect 5635 42820 5644 42860
rect 5684 42820 6508 42860
rect 6548 42820 6557 42860
rect 6604 42860 6644 42904
rect 21424 42884 21504 42904
rect 14179 42860 14237 42861
rect 20035 42860 20093 42861
rect 21187 42860 21245 42861
rect 6604 42820 11692 42860
rect 11732 42820 11741 42860
rect 14179 42820 14188 42860
rect 14228 42820 18988 42860
rect 19028 42820 19037 42860
rect 20035 42820 20044 42860
rect 20084 42820 21196 42860
rect 21236 42820 21245 42860
rect 6499 42819 6557 42820
rect 14179 42819 14237 42820
rect 20035 42819 20093 42820
rect 21187 42819 21245 42820
rect 0 42776 80 42796
rect 1315 42776 1373 42777
rect 2467 42776 2525 42777
rect 16579 42776 16637 42777
rect 21379 42776 21437 42777
rect 0 42736 1324 42776
rect 1364 42736 2476 42776
rect 2516 42736 2525 42776
rect 2755 42736 2764 42776
rect 2804 42736 3436 42776
rect 3476 42736 3485 42776
rect 3619 42736 3628 42776
rect 3668 42736 3916 42776
rect 3956 42736 4108 42776
rect 4148 42736 4157 42776
rect 4483 42736 4492 42776
rect 4532 42736 5012 42776
rect 7267 42736 7276 42776
rect 7316 42736 8428 42776
rect 8468 42736 8477 42776
rect 8707 42736 8716 42776
rect 8756 42736 9100 42776
rect 9140 42736 9149 42776
rect 12067 42736 12076 42776
rect 12116 42736 12748 42776
rect 12788 42736 14092 42776
rect 14132 42736 14380 42776
rect 14420 42736 14429 42776
rect 16579 42736 16588 42776
rect 16628 42736 17932 42776
rect 17972 42736 17981 42776
rect 19555 42736 19564 42776
rect 19604 42736 21388 42776
rect 21428 42736 21437 42776
rect 0 42716 80 42736
rect 1315 42735 1373 42736
rect 2467 42735 2525 42736
rect 3436 42692 3476 42736
rect 4972 42692 5012 42736
rect 16579 42735 16637 42736
rect 21379 42735 21437 42736
rect 8515 42692 8573 42693
rect 3436 42652 4876 42692
rect 4916 42652 4925 42692
rect 4972 42652 8524 42692
rect 8564 42652 8573 42692
rect 8515 42651 8573 42652
rect 10915 42692 10973 42693
rect 10915 42652 10924 42692
rect 10964 42652 11308 42692
rect 11348 42652 11357 42692
rect 13123 42652 13132 42692
rect 13172 42652 17164 42692
rect 17204 42652 17213 42692
rect 17347 42652 17356 42692
rect 17396 42652 18796 42692
rect 18836 42652 18845 42692
rect 10915 42651 10973 42652
rect 9667 42608 9725 42609
rect 15139 42608 15197 42609
rect 16771 42608 16829 42609
rect 17923 42608 17981 42609
rect 4195 42568 4204 42608
rect 4244 42568 4396 42608
rect 4436 42568 4445 42608
rect 6700 42568 7180 42608
rect 7220 42568 7229 42608
rect 9187 42568 9196 42608
rect 9236 42568 9388 42608
rect 9428 42568 9437 42608
rect 9667 42568 9676 42608
rect 9716 42568 11500 42608
rect 11540 42568 11549 42608
rect 15054 42568 15148 42608
rect 15188 42568 15197 42608
rect 16686 42568 16780 42608
rect 16820 42568 16829 42608
rect 17838 42568 17932 42608
rect 17972 42568 17981 42608
rect 6700 42524 6740 42568
rect 9667 42567 9725 42568
rect 15139 42567 15197 42568
rect 16771 42567 16829 42568
rect 17923 42567 17981 42568
rect 20995 42608 21053 42609
rect 21424 42608 21504 42628
rect 20995 42568 21004 42608
rect 21044 42568 21504 42608
rect 20995 42567 21053 42568
rect 21424 42548 21504 42568
rect 17539 42524 17597 42525
rect 19939 42524 19997 42525
rect 3043 42484 3052 42524
rect 3092 42484 3244 42524
rect 3284 42484 3293 42524
rect 6691 42484 6700 42524
rect 6740 42484 6749 42524
rect 6979 42484 6988 42524
rect 7028 42484 9100 42524
rect 9140 42484 9149 42524
rect 17539 42484 17548 42524
rect 17588 42484 19372 42524
rect 19412 42484 19421 42524
rect 19854 42484 19948 42524
rect 19988 42484 19997 42524
rect 17539 42483 17597 42484
rect 19939 42483 19997 42484
rect 0 42440 80 42460
rect 11107 42440 11165 42441
rect 0 42400 5260 42440
rect 5300 42400 5452 42440
rect 5492 42400 5501 42440
rect 7171 42400 7180 42440
rect 7220 42400 7372 42440
rect 7412 42400 7421 42440
rect 8227 42400 8236 42440
rect 8276 42400 11116 42440
rect 11156 42400 11165 42440
rect 11299 42400 11308 42440
rect 11348 42400 12460 42440
rect 12500 42400 17260 42440
rect 17300 42400 17309 42440
rect 17635 42400 17644 42440
rect 17684 42400 18604 42440
rect 18644 42400 18653 42440
rect 19276 42400 21004 42440
rect 21044 42400 21053 42440
rect 0 42380 80 42400
rect 11107 42399 11165 42400
rect 17251 42356 17309 42357
rect 1795 42316 1804 42356
rect 1844 42316 3572 42356
rect 3679 42316 3688 42356
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 4056 42316 4065 42356
rect 6499 42316 6508 42356
rect 6548 42316 7660 42356
rect 7700 42316 11692 42356
rect 11732 42316 11741 42356
rect 17251 42316 17260 42356
rect 17300 42316 18220 42356
rect 18260 42316 18269 42356
rect 18799 42316 18808 42356
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 19176 42316 19185 42356
rect 0 42104 80 42124
rect 3532 42104 3572 42316
rect 17251 42315 17309 42316
rect 19276 42272 19316 42400
rect 21424 42272 21504 42292
rect 5251 42232 5260 42272
rect 5300 42232 7220 42272
rect 7843 42232 7852 42272
rect 7892 42232 8428 42272
rect 8468 42232 8477 42272
rect 8524 42232 13132 42272
rect 13172 42232 13181 42272
rect 13228 42232 18260 42272
rect 4195 42188 4253 42189
rect 4483 42188 4541 42189
rect 7180 42188 7220 42232
rect 8524 42189 8564 42232
rect 7843 42188 7901 42189
rect 8515 42188 8573 42189
rect 13228 42188 13268 42232
rect 15523 42188 15581 42189
rect 17827 42188 17885 42189
rect 4195 42148 4204 42188
rect 4244 42148 4396 42188
rect 4436 42148 4492 42188
rect 4532 42148 4876 42188
rect 4916 42148 6988 42188
rect 7028 42148 7037 42188
rect 7180 42148 7852 42188
rect 7892 42148 8236 42188
rect 8276 42148 8285 42188
rect 8515 42148 8524 42188
rect 8564 42148 8573 42188
rect 11107 42148 11116 42188
rect 11156 42148 13268 42188
rect 15139 42148 15148 42188
rect 15188 42148 15532 42188
rect 15572 42148 15581 42188
rect 17742 42148 17836 42188
rect 17876 42148 17885 42188
rect 4195 42147 4253 42148
rect 4483 42147 4541 42148
rect 7843 42147 7901 42148
rect 8515 42147 8573 42148
rect 15523 42147 15581 42148
rect 17827 42147 17885 42148
rect 18220 42104 18260 42232
rect 18988 42232 19316 42272
rect 19852 42232 20948 42272
rect 20995 42232 21004 42272
rect 21044 42232 21504 42272
rect 18988 42188 19028 42232
rect 19363 42188 19421 42189
rect 18979 42148 18988 42188
rect 19028 42148 19037 42188
rect 19278 42148 19372 42188
rect 19412 42148 19421 42188
rect 19363 42147 19421 42148
rect 0 42064 3476 42104
rect 3532 42064 18124 42104
rect 18164 42064 18173 42104
rect 18220 42064 19756 42104
rect 19796 42064 19805 42104
rect 0 42044 80 42064
rect 3436 42020 3476 42064
rect 7747 42020 7805 42021
rect 10339 42020 10397 42021
rect 2755 41980 2764 42020
rect 2804 41980 2956 42020
rect 2996 41980 3005 42020
rect 3436 41980 5260 42020
rect 5300 41980 5309 42020
rect 5539 41980 5548 42020
rect 5588 41980 6892 42020
rect 6932 41980 7756 42020
rect 7796 41980 10348 42020
rect 10388 41980 10397 42020
rect 11491 41980 11500 42020
rect 11540 41980 19180 42020
rect 19220 41980 19229 42020
rect 7747 41979 7805 41980
rect 10339 41979 10397 41980
rect 3235 41936 3293 41937
rect 11011 41936 11069 41937
rect 13699 41936 13757 41937
rect 19852 41936 19892 42232
rect 20803 42188 20861 42189
rect 20131 42148 20140 42188
rect 20180 42148 20812 42188
rect 20852 42148 20861 42188
rect 20908 42188 20948 42232
rect 21424 42212 21504 42232
rect 20908 42148 21100 42188
rect 21140 42148 21149 42188
rect 20803 42147 20861 42148
rect 3043 41896 3052 41936
rect 3092 41896 3244 41936
rect 3284 41896 3293 41936
rect 3619 41896 3628 41936
rect 3668 41896 4588 41936
rect 4628 41896 4637 41936
rect 6307 41896 6316 41936
rect 6356 41896 6508 41936
rect 6548 41896 6557 41936
rect 6691 41896 6700 41936
rect 6740 41896 7276 41936
rect 7316 41896 7564 41936
rect 7604 41896 7613 41936
rect 7747 41896 7756 41936
rect 7796 41896 8044 41936
rect 8084 41896 8093 41936
rect 11011 41896 11020 41936
rect 11060 41896 11116 41936
rect 11156 41896 11165 41936
rect 13123 41896 13132 41936
rect 13172 41896 13708 41936
rect 13748 41896 15820 41936
rect 15860 41896 15869 41936
rect 16771 41896 16780 41936
rect 16820 41896 16829 41936
rect 16876 41896 19892 41936
rect 21292 41980 21428 42020
rect 3235 41895 3293 41896
rect 11011 41895 11069 41896
rect 13699 41895 13757 41896
rect 9763 41852 9821 41853
rect 10243 41852 10301 41853
rect 16780 41852 16820 41896
rect 2947 41812 2956 41852
rect 2996 41812 4012 41852
rect 4052 41812 4061 41852
rect 7171 41812 7180 41852
rect 7220 41812 8236 41852
rect 8276 41812 8285 41852
rect 9763 41812 9772 41852
rect 9812 41812 9868 41852
rect 9908 41812 9917 41852
rect 10243 41812 10252 41852
rect 10292 41812 11212 41852
rect 11252 41812 11261 41852
rect 13507 41812 13516 41852
rect 13556 41812 16820 41852
rect 9763 41811 9821 41812
rect 10243 41811 10301 41812
rect 0 41768 80 41788
rect 7171 41768 7229 41769
rect 7651 41768 7709 41769
rect 8707 41768 8765 41769
rect 14284 41768 14324 41812
rect 16876 41768 16916 41896
rect 20140 41812 21196 41852
rect 21236 41812 21245 41852
rect 0 41728 5356 41768
rect 5396 41728 5405 41768
rect 6979 41728 6988 41768
rect 7028 41728 7180 41768
rect 7220 41728 7229 41768
rect 7566 41728 7660 41768
rect 7700 41728 7709 41768
rect 7843 41728 7852 41768
rect 7892 41728 8140 41768
rect 8180 41728 8189 41768
rect 8622 41728 8716 41768
rect 8756 41728 8765 41768
rect 9091 41728 9100 41768
rect 9140 41728 9428 41768
rect 9475 41728 9484 41768
rect 9524 41728 10540 41768
rect 10580 41728 10589 41768
rect 14275 41728 14284 41768
rect 14324 41728 14364 41768
rect 16387 41728 16396 41768
rect 16436 41728 16916 41768
rect 17155 41768 17213 41769
rect 20140 41768 20180 41812
rect 17155 41728 17164 41768
rect 17204 41728 19564 41768
rect 19604 41728 19613 41768
rect 19747 41728 19756 41768
rect 19796 41728 20180 41768
rect 0 41708 80 41728
rect 7171 41727 7229 41728
rect 7651 41727 7709 41728
rect 8707 41727 8765 41728
rect 6115 41644 6124 41684
rect 6164 41644 7276 41684
rect 7316 41644 7325 41684
rect 7459 41644 7468 41684
rect 7508 41644 8276 41684
rect 9283 41644 9292 41684
rect 9332 41644 9341 41684
rect 8236 41600 8276 41644
rect 8899 41600 8957 41601
rect 9292 41600 9332 41644
rect 4919 41560 4928 41600
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 5296 41560 5305 41600
rect 6595 41560 6604 41600
rect 6644 41560 7756 41600
rect 7796 41560 7805 41600
rect 8227 41560 8236 41600
rect 8276 41560 8285 41600
rect 8332 41560 8716 41600
rect 8756 41560 8765 41600
rect 8899 41560 8908 41600
rect 8948 41560 9004 41600
rect 9044 41560 9053 41600
rect 9196 41560 9332 41600
rect 9388 41600 9428 41728
rect 17155 41727 17213 41728
rect 10435 41684 10493 41685
rect 21292 41684 21332 41980
rect 21388 41956 21428 41980
rect 21388 41896 21504 41956
rect 21424 41876 21504 41896
rect 10051 41644 10060 41684
rect 10100 41644 10444 41684
rect 10484 41644 10493 41684
rect 11299 41644 11308 41684
rect 11348 41644 21332 41684
rect 10435 41643 10493 41644
rect 16387 41600 16445 41601
rect 21424 41600 21504 41620
rect 9388 41560 9676 41600
rect 9716 41560 9725 41600
rect 10243 41560 10252 41600
rect 10292 41560 10636 41600
rect 10676 41560 10685 41600
rect 12739 41560 12748 41600
rect 12788 41560 13612 41600
rect 13652 41560 13661 41600
rect 13987 41560 13996 41600
rect 14036 41560 14956 41600
rect 14996 41560 15005 41600
rect 16387 41560 16396 41600
rect 16436 41560 16876 41600
rect 16916 41560 16925 41600
rect 17827 41560 17836 41600
rect 17876 41560 19948 41600
rect 19988 41560 19997 41600
rect 20039 41560 20048 41600
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20416 41560 20425 41600
rect 21091 41560 21100 41600
rect 21140 41560 21504 41600
rect 4291 41516 4349 41517
rect 8332 41516 8372 41560
rect 8899 41559 8957 41560
rect 4003 41476 4012 41516
rect 4052 41476 4300 41516
rect 4340 41476 4349 41516
rect 4291 41475 4349 41476
rect 6412 41476 8332 41516
rect 8372 41476 8381 41516
rect 8524 41476 8908 41516
rect 8948 41476 8957 41516
rect 0 41432 80 41452
rect 1987 41432 2045 41433
rect 6412 41432 6452 41476
rect 6883 41432 6941 41433
rect 0 41392 1996 41432
rect 2036 41392 2045 41432
rect 2275 41392 2284 41432
rect 2324 41392 3820 41432
rect 3860 41392 4684 41432
rect 4724 41392 4733 41432
rect 4867 41392 4876 41432
rect 4916 41392 5836 41432
rect 5876 41392 6412 41432
rect 6452 41392 6461 41432
rect 6883 41392 6892 41432
rect 6932 41392 7372 41432
rect 7412 41392 7508 41432
rect 7555 41392 7564 41432
rect 7604 41392 8044 41432
rect 8084 41392 8428 41432
rect 8468 41392 8477 41432
rect 0 41372 80 41392
rect 1987 41391 2045 41392
rect 6883 41391 6941 41392
rect 7468 41348 7508 41392
rect 8524 41348 8564 41476
rect 9196 41432 9236 41560
rect 16387 41559 16445 41560
rect 21424 41540 21504 41560
rect 9763 41516 9821 41517
rect 17827 41516 17885 41517
rect 9763 41476 9772 41516
rect 9812 41476 11156 41516
rect 14179 41476 14188 41516
rect 14228 41476 14860 41516
rect 14900 41476 14909 41516
rect 15907 41476 15916 41516
rect 15956 41476 16588 41516
rect 16628 41476 16637 41516
rect 17731 41476 17740 41516
rect 17780 41476 17836 41516
rect 17876 41476 17885 41516
rect 9763 41475 9821 41476
rect 8611 41392 8620 41432
rect 8660 41392 9236 41432
rect 9283 41392 9292 41432
rect 9332 41392 11020 41432
rect 11060 41392 11069 41432
rect 2563 41308 2572 41348
rect 2612 41308 3436 41348
rect 3476 41308 4204 41348
rect 4244 41308 4253 41348
rect 5539 41308 5548 41348
rect 5588 41308 7412 41348
rect 7468 41308 7948 41348
rect 7988 41308 8332 41348
rect 8372 41308 8564 41348
rect 9763 41308 9772 41348
rect 9812 41308 9964 41348
rect 10004 41308 10013 41348
rect 10723 41308 10732 41348
rect 10772 41308 11060 41348
rect 7372 41264 7412 41308
rect 9964 41264 10004 41308
rect 1219 41224 1228 41264
rect 1268 41224 1612 41264
rect 1652 41224 1661 41264
rect 2659 41224 2668 41264
rect 2708 41224 2860 41264
rect 2900 41224 3340 41264
rect 3380 41224 4396 41264
rect 4436 41224 4445 41264
rect 4771 41224 4780 41264
rect 4820 41224 7316 41264
rect 7372 41224 7892 41264
rect 8707 41224 8716 41264
rect 8756 41224 9004 41264
rect 9044 41224 9053 41264
rect 9187 41224 9196 41264
rect 9236 41224 9868 41264
rect 9908 41224 9917 41264
rect 9964 41224 10252 41264
rect 10292 41224 10444 41264
rect 10484 41224 10493 41264
rect 10915 41224 10924 41264
rect 10964 41224 10973 41264
rect 4099 41180 4157 41181
rect 1987 41140 1996 41180
rect 2036 41140 3724 41180
rect 3764 41140 3773 41180
rect 3907 41140 3916 41180
rect 3956 41140 4108 41180
rect 4148 41140 4157 41180
rect 4099 41139 4157 41140
rect 0 41096 80 41116
rect 4675 41096 4733 41097
rect 6883 41096 6941 41097
rect 0 41056 1900 41096
rect 1940 41056 1949 41096
rect 3811 41056 3820 41096
rect 3860 41056 4108 41096
rect 4148 41056 4157 41096
rect 4590 41056 4684 41096
rect 4724 41056 4733 41096
rect 6691 41056 6700 41096
rect 6740 41056 6892 41096
rect 6932 41056 6941 41096
rect 7276 41096 7316 41224
rect 7852 41096 7892 41224
rect 10924 41180 10964 41224
rect 11020 41180 11060 41308
rect 9283 41140 9292 41180
rect 9332 41140 10964 41180
rect 11011 41140 11020 41180
rect 11060 41140 11069 41180
rect 8899 41096 8957 41097
rect 7276 41056 7372 41096
rect 7412 41056 7421 41096
rect 7852 41056 8908 41096
rect 8948 41056 11060 41096
rect 0 41036 80 41056
rect 4675 41055 4733 41056
rect 6883 41055 6941 41056
rect 8899 41055 8957 41056
rect 7651 41012 7709 41013
rect 9187 41012 9245 41013
rect 3139 40972 3148 41012
rect 3188 40972 7660 41012
rect 7700 40972 9196 41012
rect 9236 40972 9245 41012
rect 9571 40972 9580 41012
rect 9620 40972 9772 41012
rect 9812 40972 9821 41012
rect 7651 40971 7709 40972
rect 9187 40971 9245 40972
rect 3427 40928 3485 40929
rect 8803 40928 8861 40929
rect 3427 40888 3436 40928
rect 3476 40888 4340 40928
rect 3427 40887 3485 40888
rect 3679 40804 3688 40844
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 4056 40804 4065 40844
rect 0 40760 80 40780
rect 4195 40760 4253 40761
rect 0 40720 4204 40760
rect 4244 40720 4253 40760
rect 4300 40760 4340 40888
rect 5932 40888 8428 40928
rect 8468 40888 8620 40928
rect 8660 40888 8669 40928
rect 8803 40888 8812 40928
rect 8852 40888 10964 40928
rect 5932 40844 5972 40888
rect 8803 40887 8861 40888
rect 4483 40804 4492 40844
rect 4532 40804 5932 40844
rect 5972 40804 5981 40844
rect 6499 40804 6508 40844
rect 6548 40804 6892 40844
rect 6932 40804 10828 40844
rect 10868 40804 10877 40844
rect 8707 40760 8765 40761
rect 10924 40760 10964 40888
rect 11020 40844 11060 41056
rect 11116 40928 11156 41476
rect 17827 41475 17885 41476
rect 15043 41432 15101 41433
rect 20611 41432 20669 41433
rect 13699 41392 13708 41432
rect 13748 41392 15052 41432
rect 15092 41392 15101 41432
rect 15523 41392 15532 41432
rect 15572 41392 18316 41432
rect 18356 41392 18365 41432
rect 20227 41392 20236 41432
rect 20276 41392 20620 41432
rect 20660 41392 20669 41432
rect 15043 41391 15101 41392
rect 20611 41391 20669 41392
rect 14371 41308 14380 41348
rect 14420 41308 14668 41348
rect 14708 41308 14717 41348
rect 17635 41308 17644 41348
rect 17684 41308 18508 41348
rect 18548 41308 18557 41348
rect 21424 41264 21504 41284
rect 11203 41224 11212 41264
rect 11252 41224 19564 41264
rect 19604 41224 19613 41264
rect 21187 41224 21196 41264
rect 21236 41224 21504 41264
rect 21424 41204 21504 41224
rect 15235 41140 15244 41180
rect 15284 41140 15436 41180
rect 15476 41140 16972 41180
rect 17012 41140 17164 41180
rect 17204 41140 17213 41180
rect 17923 41140 17932 41180
rect 17972 41140 18796 41180
rect 18836 41140 18845 41180
rect 20035 41140 20044 41180
rect 20084 41140 20093 41180
rect 12643 41096 12701 41097
rect 20044 41096 20084 41140
rect 12643 41056 12652 41096
rect 12692 41056 20084 41096
rect 12643 41055 12701 41056
rect 14851 41012 14909 41013
rect 13411 40972 13420 41012
rect 13460 40972 14668 41012
rect 14708 40972 14717 41012
rect 14851 40972 14860 41012
rect 14900 40972 17740 41012
rect 17780 40972 17789 41012
rect 17836 40972 19180 41012
rect 19220 40972 19229 41012
rect 19363 40972 19372 41012
rect 19412 40972 19660 41012
rect 19700 40972 19709 41012
rect 14851 40971 14909 40972
rect 16099 40928 16157 40929
rect 11116 40888 13652 40928
rect 13699 40888 13708 40928
rect 13748 40888 14860 40928
rect 14900 40888 14909 40928
rect 16014 40888 16108 40928
rect 16148 40888 16157 40928
rect 13612 40844 13652 40888
rect 16099 40887 16157 40888
rect 17836 40844 17876 40972
rect 21424 40928 21504 40948
rect 11020 40804 12556 40844
rect 12596 40804 12605 40844
rect 13612 40804 14380 40844
rect 14420 40804 17876 40844
rect 18124 40888 21504 40928
rect 4300 40720 6316 40760
rect 6356 40720 7604 40760
rect 0 40700 80 40720
rect 4195 40719 4253 40720
rect 6499 40676 6557 40677
rect 7564 40676 7604 40720
rect 8707 40720 8716 40760
rect 8756 40720 10060 40760
rect 10100 40720 10109 40760
rect 10924 40720 17836 40760
rect 17876 40720 17885 40760
rect 8707 40719 8765 40720
rect 9187 40676 9245 40677
rect 10915 40676 10973 40677
rect 13507 40676 13565 40677
rect 18124 40676 18164 40888
rect 21424 40868 21504 40888
rect 18799 40804 18808 40844
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 19176 40804 19185 40844
rect 2947 40636 2956 40676
rect 2996 40636 4780 40676
rect 4820 40636 4829 40676
rect 6499 40636 6508 40676
rect 6548 40636 6988 40676
rect 7028 40636 7037 40676
rect 7459 40636 7468 40676
rect 7508 40636 7517 40676
rect 7564 40636 8276 40676
rect 8323 40636 8332 40676
rect 8372 40636 8908 40676
rect 8948 40636 8957 40676
rect 9187 40636 9196 40676
rect 9236 40636 9676 40676
rect 9716 40636 9725 40676
rect 9955 40636 9964 40676
rect 10004 40636 10444 40676
rect 10484 40636 10493 40676
rect 10830 40636 10924 40676
rect 10964 40636 10973 40676
rect 13315 40636 13324 40676
rect 13364 40636 13516 40676
rect 13556 40636 13565 40676
rect 15427 40636 15436 40676
rect 15476 40636 15764 40676
rect 16099 40636 16108 40676
rect 16148 40636 16157 40676
rect 17443 40636 17452 40676
rect 17492 40636 18164 40676
rect 18211 40636 18220 40676
rect 18260 40636 19276 40676
rect 19316 40636 19325 40676
rect 6499 40635 6557 40636
rect 7363 40592 7421 40593
rect 2851 40552 2860 40592
rect 2900 40552 3916 40592
rect 3956 40552 3965 40592
rect 4291 40552 4300 40592
rect 4340 40552 4684 40592
rect 4724 40552 4733 40592
rect 5251 40552 5260 40592
rect 5300 40552 7372 40592
rect 7412 40552 7421 40592
rect 7468 40592 7508 40636
rect 8236 40593 8276 40636
rect 9187 40635 9245 40636
rect 10915 40635 10973 40636
rect 13507 40635 13565 40636
rect 8227 40592 8285 40593
rect 13219 40592 13277 40593
rect 15724 40592 15764 40636
rect 7468 40552 7852 40592
rect 7892 40552 7901 40592
rect 8227 40552 8236 40592
rect 8276 40552 8285 40592
rect 9091 40552 9100 40592
rect 9140 40552 9868 40592
rect 9908 40552 9917 40592
rect 10051 40552 10060 40592
rect 10100 40552 10348 40592
rect 10388 40552 10397 40592
rect 12643 40552 12652 40592
rect 12692 40552 13228 40592
rect 13268 40552 13277 40592
rect 13507 40552 13516 40592
rect 13556 40552 15340 40592
rect 15380 40552 15389 40592
rect 15715 40552 15724 40592
rect 15764 40552 15773 40592
rect 7363 40551 7421 40552
rect 8227 40551 8285 40552
rect 13219 40551 13277 40552
rect 2947 40508 3005 40509
rect 3427 40508 3485 40509
rect 6883 40508 6941 40509
rect 2947 40468 2956 40508
rect 2996 40468 3436 40508
rect 3476 40468 3628 40508
rect 3668 40468 3677 40508
rect 4099 40468 4108 40508
rect 4148 40468 4396 40508
rect 4436 40468 4445 40508
rect 5347 40468 5356 40508
rect 5396 40468 6892 40508
rect 6932 40468 6941 40508
rect 2947 40467 3005 40468
rect 3427 40467 3485 40468
rect 6883 40467 6941 40468
rect 7171 40508 7229 40509
rect 11491 40508 11549 40509
rect 16108 40508 16148 40636
rect 20611 40592 20669 40593
rect 21424 40592 21504 40612
rect 20611 40552 20620 40592
rect 20660 40552 21504 40592
rect 20611 40551 20669 40552
rect 21424 40532 21504 40552
rect 7171 40468 7180 40508
rect 7220 40468 7276 40508
rect 7316 40468 7325 40508
rect 7651 40468 7660 40508
rect 7700 40468 8524 40508
rect 8564 40468 8573 40508
rect 8899 40468 8908 40508
rect 8948 40468 10252 40508
rect 10292 40468 10301 40508
rect 11406 40468 11500 40508
rect 11540 40468 11549 40508
rect 15811 40468 15820 40508
rect 15860 40468 16148 40508
rect 7171 40467 7229 40468
rect 11491 40467 11549 40468
rect 0 40424 80 40444
rect 10339 40424 10397 40425
rect 0 40384 2228 40424
rect 2275 40384 2284 40424
rect 2324 40384 2572 40424
rect 2612 40384 2860 40424
rect 2900 40384 4148 40424
rect 4195 40384 4204 40424
rect 4244 40384 4588 40424
rect 4628 40384 4637 40424
rect 5731 40384 5740 40424
rect 5780 40384 6068 40424
rect 6787 40384 6796 40424
rect 6836 40384 7468 40424
rect 7508 40384 7517 40424
rect 7939 40384 7948 40424
rect 7988 40384 8812 40424
rect 8852 40384 8861 40424
rect 9283 40384 9292 40424
rect 9332 40384 9341 40424
rect 9475 40384 9484 40424
rect 9524 40384 10156 40424
rect 10196 40384 10205 40424
rect 10339 40384 10348 40424
rect 10388 40384 10482 40424
rect 11320 40384 19948 40424
rect 19988 40384 19997 40424
rect 0 40364 80 40384
rect 2188 40340 2228 40384
rect 3331 40340 3389 40341
rect 2188 40300 3340 40340
rect 3380 40300 3389 40340
rect 4108 40340 4148 40384
rect 6028 40340 6068 40384
rect 9292 40340 9332 40384
rect 10339 40383 10397 40384
rect 11320 40340 11360 40384
rect 14083 40340 14141 40341
rect 4108 40300 4972 40340
rect 5012 40300 5356 40340
rect 5396 40300 5405 40340
rect 6019 40300 6028 40340
rect 6068 40300 6077 40340
rect 7267 40300 7276 40340
rect 7316 40300 9332 40340
rect 10252 40300 11360 40340
rect 13998 40300 14092 40340
rect 14132 40300 14141 40340
rect 3331 40299 3389 40300
rect 8899 40256 8957 40257
rect 10252 40256 10292 40300
rect 14083 40299 14141 40300
rect 14275 40340 14333 40341
rect 15043 40340 15101 40341
rect 19459 40340 19517 40341
rect 14275 40300 14284 40340
rect 14324 40300 15052 40340
rect 15092 40300 16108 40340
rect 16148 40300 16300 40340
rect 16340 40300 16349 40340
rect 19374 40300 19468 40340
rect 19508 40300 19517 40340
rect 14275 40299 14333 40300
rect 15043 40299 15101 40300
rect 19459 40299 19517 40300
rect 21424 40256 21504 40276
rect 2659 40216 2668 40256
rect 2708 40216 3532 40256
rect 3572 40216 3581 40256
rect 3628 40216 5740 40256
rect 5780 40216 8236 40256
rect 8276 40216 8285 40256
rect 8899 40216 8908 40256
rect 8948 40216 9004 40256
rect 9044 40216 9053 40256
rect 9283 40216 9292 40256
rect 9332 40216 9580 40256
rect 9620 40216 9629 40256
rect 10243 40216 10252 40256
rect 10292 40216 10301 40256
rect 13699 40216 13708 40256
rect 13748 40216 19220 40256
rect 20515 40216 20524 40256
rect 20564 40216 21504 40256
rect 3628 40172 3668 40216
rect 8899 40215 8957 40216
rect 19180 40172 19220 40216
rect 21424 40196 21504 40216
rect 2947 40132 2956 40172
rect 2996 40132 3668 40172
rect 4492 40132 7852 40172
rect 7892 40132 10636 40172
rect 10676 40132 10685 40172
rect 13603 40132 13612 40172
rect 13652 40132 16588 40172
rect 16628 40132 16780 40172
rect 16820 40132 16829 40172
rect 17059 40132 17068 40172
rect 17108 40132 17452 40172
rect 17492 40132 17501 40172
rect 19171 40132 19180 40172
rect 19220 40132 19229 40172
rect 0 40088 80 40108
rect 4492 40088 4532 40132
rect 4780 40088 4820 40132
rect 16099 40088 16157 40089
rect 0 40048 1708 40088
rect 1748 40048 1757 40088
rect 3139 40048 3148 40088
rect 3188 40048 4532 40088
rect 4771 40048 4780 40088
rect 4820 40048 4860 40088
rect 4919 40048 4928 40088
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 5296 40048 5305 40088
rect 8035 40048 8044 40088
rect 8084 40048 8428 40088
rect 8468 40048 8477 40088
rect 8899 40048 8908 40088
rect 8948 40048 9484 40088
rect 9524 40048 9533 40088
rect 11320 40048 16108 40088
rect 16148 40048 16157 40088
rect 20039 40048 20048 40088
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20416 40048 20425 40088
rect 0 40028 80 40048
rect 2083 39964 2092 40004
rect 2132 39964 7700 40004
rect 7747 39964 7756 40004
rect 7796 39964 10732 40004
rect 10772 39964 10781 40004
rect 7660 39920 7700 39964
rect 7843 39920 7901 39921
rect 8227 39920 8285 39921
rect 11320 39920 11360 40048
rect 16099 40047 16157 40048
rect 13027 39964 13036 40004
rect 13076 39964 13516 40004
rect 13556 39964 13565 40004
rect 13996 39964 15148 40004
rect 15188 39964 15197 40004
rect 15715 39964 15724 40004
rect 15764 39964 18124 40004
rect 18164 39964 18173 40004
rect 13996 39920 14036 39964
rect 14179 39920 14237 39921
rect 17923 39920 17981 39921
rect 21424 39920 21504 39940
rect 2467 39880 2476 39920
rect 2516 39880 3340 39920
rect 3380 39880 6644 39920
rect 6691 39880 6700 39920
rect 6740 39880 7276 39920
rect 7316 39880 7325 39920
rect 7651 39880 7660 39920
rect 7700 39880 7709 39920
rect 7843 39880 7852 39920
rect 7892 39880 7948 39920
rect 7988 39880 7997 39920
rect 8227 39880 8236 39920
rect 8276 39880 8332 39920
rect 8372 39880 8381 39920
rect 8515 39880 8524 39920
rect 8564 39880 11360 39920
rect 12556 39880 13132 39920
rect 13172 39880 14036 39920
rect 14094 39880 14188 39920
rect 14228 39880 14237 39920
rect 14467 39880 14476 39920
rect 14516 39880 14764 39920
rect 14804 39880 14813 39920
rect 15235 39880 15244 39920
rect 15284 39880 15476 39920
rect 6604 39836 6644 39880
rect 7843 39879 7901 39880
rect 8227 39879 8285 39880
rect 3811 39796 3820 39836
rect 3860 39796 4972 39836
rect 5012 39796 5021 39836
rect 6604 39796 8372 39836
rect 8419 39796 8428 39836
rect 8468 39796 10540 39836
rect 10580 39796 10589 39836
rect 0 39752 80 39772
rect 4291 39752 4349 39753
rect 4675 39752 4733 39753
rect 8332 39752 8372 39796
rect 8707 39752 8765 39753
rect 0 39712 556 39752
rect 596 39712 605 39752
rect 4291 39712 4300 39752
rect 4340 39712 4492 39752
rect 4532 39712 4541 39752
rect 4675 39712 4684 39752
rect 4724 39712 4876 39752
rect 4916 39712 4925 39752
rect 5164 39712 6508 39752
rect 6548 39712 6557 39752
rect 6883 39712 6892 39752
rect 6932 39712 7372 39752
rect 7412 39712 7421 39752
rect 8332 39712 8716 39752
rect 8756 39712 8765 39752
rect 0 39692 80 39712
rect 4291 39711 4349 39712
rect 4675 39711 4733 39712
rect 5164 39668 5204 39712
rect 8707 39711 8765 39712
rect 9772 39712 10348 39752
rect 10388 39712 10397 39752
rect 9772 39668 9812 39712
rect 2476 39628 5204 39668
rect 5251 39628 5260 39668
rect 5300 39628 8524 39668
rect 8564 39628 8573 39668
rect 9187 39628 9196 39668
rect 9236 39628 9716 39668
rect 9763 39628 9772 39668
rect 9812 39628 9821 39668
rect 2476 39584 2516 39628
rect 8899 39584 8957 39585
rect 9676 39584 9716 39628
rect 12556 39584 12596 39880
rect 14179 39879 14237 39880
rect 14275 39796 14284 39836
rect 14324 39796 14708 39836
rect 12739 39712 12748 39752
rect 12788 39712 13132 39752
rect 13172 39712 13324 39752
rect 13364 39712 14188 39752
rect 14228 39712 14237 39752
rect 12931 39628 12940 39668
rect 12980 39628 14380 39668
rect 14420 39628 14429 39668
rect 14668 39584 14708 39796
rect 15436 39752 15476 39880
rect 17923 39880 17932 39920
rect 17972 39880 18412 39920
rect 18452 39880 18461 39920
rect 19843 39880 19852 39920
rect 19892 39880 21004 39920
rect 21044 39880 21053 39920
rect 21100 39880 21504 39920
rect 17923 39879 17981 39880
rect 21100 39836 21140 39880
rect 21424 39860 21504 39880
rect 17731 39796 17740 39836
rect 17780 39796 18114 39836
rect 18154 39796 18163 39836
rect 20611 39796 20620 39836
rect 20660 39796 21140 39836
rect 15427 39712 15436 39752
rect 15476 39712 15485 39752
rect 21424 39584 21504 39604
rect 2467 39544 2476 39584
rect 2516 39544 2525 39584
rect 6979 39544 6988 39584
rect 7028 39544 8908 39584
rect 8948 39544 9580 39584
rect 9620 39544 9629 39584
rect 9676 39544 9868 39584
rect 9908 39544 9917 39584
rect 12547 39544 12556 39584
rect 12596 39544 12605 39584
rect 13411 39544 13420 39584
rect 13460 39544 14476 39584
rect 14516 39544 14525 39584
rect 14659 39544 14668 39584
rect 14708 39544 14717 39584
rect 15139 39544 15148 39584
rect 15188 39544 15532 39584
rect 15572 39544 15581 39584
rect 20131 39544 20140 39584
rect 20180 39544 21504 39584
rect 8899 39543 8957 39544
rect 21424 39524 21504 39544
rect 19363 39500 19421 39501
rect 4003 39460 4012 39500
rect 4052 39460 9716 39500
rect 13027 39460 13036 39500
rect 13076 39460 13804 39500
rect 13844 39460 14380 39500
rect 14420 39460 14429 39500
rect 19171 39460 19180 39500
rect 19220 39460 19372 39500
rect 19412 39460 19421 39500
rect 0 39416 80 39436
rect 1603 39416 1661 39417
rect 2083 39416 2141 39417
rect 4012 39416 4052 39460
rect 0 39376 1612 39416
rect 1652 39376 2092 39416
rect 2132 39376 2141 39416
rect 2371 39376 2380 39416
rect 2420 39376 4052 39416
rect 6883 39416 6941 39417
rect 8803 39416 8861 39417
rect 6883 39376 6892 39416
rect 6932 39376 8140 39416
rect 8180 39376 8812 39416
rect 8852 39376 8861 39416
rect 0 39356 80 39376
rect 1603 39375 1661 39376
rect 2083 39375 2141 39376
rect 6883 39375 6941 39376
rect 8803 39375 8861 39376
rect 9676 39332 9716 39460
rect 19363 39459 19421 39460
rect 10252 39376 12268 39416
rect 12308 39376 12317 39416
rect 10252 39332 10292 39376
rect 12547 39332 12605 39333
rect 13699 39332 13757 39333
rect 3679 39292 3688 39332
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 4056 39292 4065 39332
rect 6499 39292 6508 39332
rect 6548 39292 7564 39332
rect 7604 39292 7613 39332
rect 9667 39292 9676 39332
rect 9716 39292 10292 39332
rect 11299 39292 11308 39332
rect 11348 39292 12556 39332
rect 12596 39292 12605 39332
rect 13614 39292 13708 39332
rect 13748 39292 13757 39332
rect 13987 39292 13996 39332
rect 14036 39292 14284 39332
rect 14324 39292 14333 39332
rect 18799 39292 18808 39332
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 19176 39292 19185 39332
rect 7564 39248 7604 39292
rect 12547 39291 12605 39292
rect 13699 39291 13757 39292
rect 9763 39248 9821 39249
rect 10243 39248 10301 39249
rect 7564 39208 9772 39248
rect 9812 39208 9821 39248
rect 10158 39208 10252 39248
rect 10292 39208 10301 39248
rect 9763 39207 9821 39208
rect 10243 39207 10301 39208
rect 20707 39248 20765 39249
rect 21424 39248 21504 39268
rect 20707 39208 20716 39248
rect 20756 39208 21504 39248
rect 20707 39207 20765 39208
rect 21424 39188 21504 39208
rect 14179 39164 14237 39165
rect 18211 39164 18269 39165
rect 2179 39124 2188 39164
rect 2228 39124 2540 39164
rect 7651 39124 7660 39164
rect 7700 39124 14188 39164
rect 14228 39124 14860 39164
rect 14900 39124 14909 39164
rect 17539 39124 17548 39164
rect 17588 39124 17597 39164
rect 18211 39124 18220 39164
rect 18260 39124 19084 39164
rect 19124 39124 19468 39164
rect 19508 39124 19517 39164
rect 0 39080 80 39100
rect 2371 39080 2429 39081
rect 0 39040 2380 39080
rect 2420 39040 2429 39080
rect 2500 39080 2540 39124
rect 14179 39123 14237 39124
rect 6211 39080 6269 39081
rect 7171 39080 7229 39081
rect 10147 39080 10205 39081
rect 17548 39080 17588 39124
rect 18211 39123 18269 39124
rect 2500 39040 5356 39080
rect 5396 39040 6220 39080
rect 6260 39040 6892 39080
rect 6932 39040 6941 39080
rect 7171 39040 7180 39080
rect 7220 39040 10156 39080
rect 10196 39040 10205 39080
rect 12259 39040 12268 39080
rect 12308 39040 15340 39080
rect 15380 39040 15389 39080
rect 16291 39040 16300 39080
rect 16340 39040 17588 39080
rect 17827 39040 17836 39080
rect 17876 39040 18508 39080
rect 18548 39040 18557 39080
rect 0 39020 80 39040
rect 2371 39039 2429 39040
rect 6211 39039 6269 39040
rect 7171 39039 7229 39040
rect 10147 39039 10205 39040
rect 3043 38996 3101 38997
rect 4099 38996 4157 38997
rect 3043 38956 3052 38996
rect 3092 38956 3148 38996
rect 3188 38956 3197 38996
rect 3532 38956 4108 38996
rect 4148 38956 4157 38996
rect 4387 38956 4396 38996
rect 4436 38956 4876 38996
rect 4916 38956 7756 38996
rect 7796 38956 7805 38996
rect 11875 38956 11884 38996
rect 11924 38956 13228 38996
rect 13268 38956 13277 38996
rect 16300 38956 19468 38996
rect 19508 38956 19517 38996
rect 3043 38955 3101 38956
rect 2755 38872 2764 38912
rect 2804 38872 3052 38912
rect 3092 38872 3101 38912
rect 3532 38828 3572 38956
rect 4099 38955 4157 38956
rect 4771 38912 4829 38913
rect 3619 38872 3628 38912
rect 3668 38872 4780 38912
rect 4820 38872 6412 38912
rect 6452 38872 7852 38912
rect 7892 38872 7901 38912
rect 8323 38872 8332 38912
rect 8372 38872 8620 38912
rect 8660 38872 8669 38912
rect 9763 38872 9772 38912
rect 9812 38872 10732 38912
rect 10772 38872 11980 38912
rect 12020 38872 12029 38912
rect 12355 38872 12364 38912
rect 12404 38872 12844 38912
rect 12884 38872 12893 38912
rect 14563 38872 14572 38912
rect 14612 38872 14956 38912
rect 14996 38872 15005 38912
rect 4771 38871 4829 38872
rect 16300 38829 16340 38956
rect 18211 38912 18269 38913
rect 19459 38912 19517 38913
rect 21424 38912 21504 38932
rect 16963 38872 16972 38912
rect 17012 38872 18220 38912
rect 18260 38872 18269 38912
rect 18403 38872 18412 38912
rect 18452 38872 18796 38912
rect 18836 38872 18845 38912
rect 18979 38872 18988 38912
rect 19028 38872 19468 38912
rect 19508 38872 19517 38912
rect 2659 38788 2668 38828
rect 2708 38788 3572 38828
rect 4195 38828 4253 38829
rect 7459 38828 7517 38829
rect 13219 38828 13277 38829
rect 16291 38828 16349 38829
rect 17644 38828 17684 38872
rect 18211 38871 18269 38872
rect 19459 38871 19517 38872
rect 20140 38872 21504 38912
rect 19267 38828 19325 38829
rect 4195 38788 4204 38828
rect 4244 38788 6932 38828
rect 6979 38788 6988 38828
rect 7028 38788 7468 38828
rect 7508 38788 7517 38828
rect 4195 38787 4253 38788
rect 0 38744 80 38764
rect 6892 38744 6932 38788
rect 7459 38787 7517 38788
rect 8620 38788 9964 38828
rect 10004 38788 10013 38828
rect 13134 38788 13228 38828
rect 13268 38788 13277 38828
rect 15235 38788 15244 38828
rect 15284 38788 16300 38828
rect 16340 38788 16349 38828
rect 17635 38788 17644 38828
rect 17684 38788 17724 38828
rect 18595 38788 18604 38828
rect 18644 38788 18892 38828
rect 18932 38788 19276 38828
rect 19316 38788 19325 38828
rect 8620 38744 8660 38788
rect 13219 38787 13277 38788
rect 16291 38787 16349 38788
rect 19267 38787 19325 38788
rect 0 38704 4204 38744
rect 4244 38704 4253 38744
rect 6892 38704 8660 38744
rect 8707 38744 8765 38745
rect 20140 38744 20180 38872
rect 21424 38852 21504 38872
rect 8707 38704 8716 38744
rect 8756 38704 13132 38744
rect 13172 38704 13181 38744
rect 16483 38704 16492 38744
rect 16532 38704 20180 38744
rect 0 38684 80 38704
rect 8707 38703 8765 38704
rect 4483 38660 4541 38661
rect 3523 38620 3532 38660
rect 3572 38620 4492 38660
rect 4532 38620 7468 38660
rect 7508 38620 7517 38660
rect 11020 38620 11212 38660
rect 11252 38620 11261 38660
rect 11395 38620 11404 38660
rect 11444 38620 11788 38660
rect 11828 38620 11837 38660
rect 13795 38620 13804 38660
rect 13844 38620 18124 38660
rect 18164 38620 18316 38660
rect 18356 38620 18508 38660
rect 18548 38620 18557 38660
rect 4483 38619 4541 38620
rect 11020 38576 11060 38620
rect 11404 38576 11444 38620
rect 21424 38576 21504 38596
rect 4919 38536 4928 38576
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 5296 38536 5305 38576
rect 6019 38536 6028 38576
rect 6068 38536 10540 38576
rect 10580 38536 11060 38576
rect 11107 38536 11116 38576
rect 11156 38536 11444 38576
rect 13123 38536 13132 38576
rect 13172 38536 18700 38576
rect 18740 38536 18749 38576
rect 20039 38536 20048 38576
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20416 38536 20425 38576
rect 20620 38536 21504 38576
rect 1411 38492 1469 38493
rect 1315 38452 1324 38492
rect 1364 38452 1420 38492
rect 1460 38452 1469 38492
rect 1411 38451 1469 38452
rect 3331 38492 3389 38493
rect 19747 38492 19805 38493
rect 20620 38492 20660 38536
rect 21424 38516 21504 38536
rect 3331 38452 3340 38492
rect 3380 38452 9292 38492
rect 9332 38452 10828 38492
rect 10868 38452 17836 38492
rect 17876 38452 17885 38492
rect 19747 38452 19756 38492
rect 19796 38452 20660 38492
rect 3331 38451 3389 38452
rect 19747 38451 19805 38452
rect 0 38408 80 38428
rect 4675 38408 4733 38409
rect 5827 38408 5885 38409
rect 12547 38408 12605 38409
rect 19555 38408 19613 38409
rect 0 38368 4684 38408
rect 4724 38368 4733 38408
rect 5539 38368 5548 38408
rect 5588 38368 5836 38408
rect 5876 38368 5885 38408
rect 9955 38368 9964 38408
rect 10004 38368 11360 38408
rect 12451 38368 12460 38408
rect 12500 38368 12556 38408
rect 12596 38368 15244 38408
rect 15284 38368 15724 38408
rect 15764 38368 15773 38408
rect 19470 38368 19564 38408
rect 19604 38368 19613 38408
rect 0 38348 80 38368
rect 4675 38367 4733 38368
rect 5827 38367 5885 38368
rect 10243 38324 10301 38325
rect 1315 38284 1324 38324
rect 1364 38284 1804 38324
rect 1844 38284 1853 38324
rect 4771 38284 4780 38324
rect 4820 38284 10252 38324
rect 10292 38284 10301 38324
rect 11320 38324 11360 38368
rect 12547 38367 12605 38368
rect 19555 38367 19613 38368
rect 12643 38324 12701 38325
rect 13411 38324 13469 38325
rect 20803 38324 20861 38325
rect 11320 38284 12652 38324
rect 12692 38284 13420 38324
rect 13460 38284 13469 38324
rect 13987 38284 13996 38324
rect 14036 38284 20812 38324
rect 20852 38284 20861 38324
rect 10243 38283 10301 38284
rect 12643 38283 12701 38284
rect 13411 38283 13469 38284
rect 20803 38283 20861 38284
rect 17827 38240 17885 38241
rect 19843 38240 19901 38241
rect 21424 38240 21504 38260
rect 1891 38200 1900 38240
rect 1940 38200 3916 38240
rect 3956 38200 3965 38240
rect 5155 38200 5164 38240
rect 5204 38200 6796 38240
rect 6836 38200 6845 38240
rect 10339 38200 10348 38240
rect 10388 38200 11212 38240
rect 11252 38200 11261 38240
rect 11683 38200 11692 38240
rect 11732 38200 13900 38240
rect 13940 38200 14668 38240
rect 14708 38200 14717 38240
rect 17742 38200 17836 38240
rect 17876 38200 17885 38240
rect 18307 38200 18316 38240
rect 18356 38200 18604 38240
rect 18644 38200 18653 38240
rect 19843 38200 19852 38240
rect 19892 38200 21504 38240
rect 17827 38199 17885 38200
rect 19843 38199 19901 38200
rect 21424 38180 21504 38200
rect 1987 38156 2045 38157
rect 2371 38156 2429 38157
rect 10243 38156 10301 38157
rect 1987 38116 1996 38156
rect 2036 38116 2380 38156
rect 2420 38116 5548 38156
rect 5588 38116 6220 38156
rect 6260 38116 6269 38156
rect 10243 38116 10252 38156
rect 10292 38116 11884 38156
rect 11924 38116 11933 38156
rect 13123 38116 13132 38156
rect 13172 38116 19756 38156
rect 19796 38116 19805 38156
rect 1987 38115 2045 38116
rect 2371 38115 2429 38116
rect 10243 38115 10301 38116
rect 0 38072 80 38092
rect 2659 38072 2717 38073
rect 19939 38072 19997 38073
rect 0 38032 212 38072
rect 0 38012 80 38032
rect 172 37904 212 38032
rect 2659 38032 2668 38072
rect 2708 38032 2956 38072
rect 2996 38032 3005 38072
rect 3907 38032 3916 38072
rect 3956 38032 7660 38072
rect 7700 38032 7709 38072
rect 10627 38032 10636 38072
rect 10676 38032 11308 38072
rect 11348 38032 11357 38072
rect 13795 38032 13804 38072
rect 13844 38032 14092 38072
rect 14132 38032 14141 38072
rect 19854 38032 19948 38072
rect 19988 38032 19997 38072
rect 2659 38031 2717 38032
rect 19939 38031 19997 38032
rect 10531 37948 10540 37988
rect 10580 37948 19372 37988
rect 19412 37948 19421 37988
rect 9667 37904 9725 37905
rect 21424 37904 21504 37924
rect 172 37864 9676 37904
rect 9716 37864 9725 37904
rect 9667 37863 9725 37864
rect 10732 37864 15436 37904
rect 15476 37864 15485 37904
rect 19267 37864 19276 37904
rect 19316 37864 21504 37904
rect 3679 37780 3688 37820
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 4056 37780 4065 37820
rect 6180 37780 6220 37820
rect 6260 37780 6269 37820
rect 0 37736 80 37756
rect 1219 37736 1277 37737
rect 6019 37736 6077 37737
rect 0 37696 1228 37736
rect 1268 37696 1277 37736
rect 5443 37696 5452 37736
rect 5492 37696 6028 37736
rect 6068 37696 6077 37736
rect 6220 37736 6260 37780
rect 10732 37736 10772 37864
rect 21424 37844 21504 37864
rect 16260 37780 16300 37820
rect 16340 37780 16349 37820
rect 18799 37780 18808 37820
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 19176 37780 19185 37820
rect 6220 37696 10772 37736
rect 16300 37736 16340 37780
rect 16300 37696 16876 37736
rect 16916 37696 16925 37736
rect 0 37676 80 37696
rect 1219 37695 1277 37696
rect 6019 37695 6077 37696
rect 3811 37652 3869 37653
rect 20611 37652 20669 37653
rect 2851 37612 2860 37652
rect 2900 37612 3148 37652
rect 3188 37612 3820 37652
rect 3860 37612 3869 37652
rect 5827 37612 5836 37652
rect 5876 37612 8716 37652
rect 8756 37612 8765 37652
rect 14467 37612 14476 37652
rect 14516 37612 20620 37652
rect 20660 37612 20669 37652
rect 3811 37611 3869 37612
rect 20611 37611 20669 37612
rect 5347 37568 5405 37569
rect 21424 37568 21504 37588
rect 2563 37528 2572 37568
rect 2612 37528 3340 37568
rect 3380 37528 3389 37568
rect 5347 37528 5356 37568
rect 5396 37528 5740 37568
rect 5780 37528 5789 37568
rect 6787 37528 6796 37568
rect 6836 37528 7948 37568
rect 7988 37528 9580 37568
rect 9620 37528 11596 37568
rect 11636 37528 12076 37568
rect 12116 37528 12125 37568
rect 13132 37528 15148 37568
rect 15188 37528 15197 37568
rect 16675 37528 16684 37568
rect 16724 37528 21504 37568
rect 5347 37527 5405 37528
rect 6307 37484 6365 37485
rect 13132 37484 13172 37528
rect 21424 37508 21504 37528
rect 6307 37444 6316 37484
rect 6356 37444 8332 37484
rect 8372 37444 13172 37484
rect 13219 37444 13228 37484
rect 13268 37444 16012 37484
rect 16052 37444 16061 37484
rect 6307 37443 6365 37444
rect 0 37400 80 37420
rect 3235 37400 3293 37401
rect 0 37360 1228 37400
rect 1268 37360 1277 37400
rect 3235 37360 3244 37400
rect 3284 37360 3532 37400
rect 3572 37360 3581 37400
rect 4003 37360 4012 37400
rect 4052 37360 4396 37400
rect 4436 37360 4445 37400
rect 6019 37360 6028 37400
rect 6068 37360 6412 37400
rect 6452 37360 6461 37400
rect 8707 37360 8716 37400
rect 8756 37360 13324 37400
rect 13364 37360 13373 37400
rect 15235 37360 15244 37400
rect 15284 37360 15916 37400
rect 15956 37360 15965 37400
rect 18691 37360 18700 37400
rect 18740 37360 19756 37400
rect 19796 37360 19805 37400
rect 0 37340 80 37360
rect 3235 37359 3293 37360
rect 4099 37316 4157 37317
rect 5635 37316 5693 37317
rect 9187 37316 9245 37317
rect 16195 37316 16253 37317
rect 4014 37276 4108 37316
rect 4148 37276 4157 37316
rect 4483 37276 4492 37316
rect 4532 37276 5644 37316
rect 5684 37276 5693 37316
rect 4099 37275 4157 37276
rect 5635 37275 5693 37276
rect 6124 37276 7412 37316
rect 7459 37276 7468 37316
rect 7508 37276 9196 37316
rect 9236 37276 9245 37316
rect 12835 37276 12844 37316
rect 12884 37276 13228 37316
rect 13268 37276 13277 37316
rect 16195 37276 16204 37316
rect 16244 37276 20180 37316
rect 6124 37232 6164 37276
rect 2851 37192 2860 37232
rect 2900 37192 6164 37232
rect 6211 37192 6220 37232
rect 6260 37192 7084 37232
rect 7124 37192 7133 37232
rect 7372 37148 7412 37276
rect 9187 37275 9245 37276
rect 16195 37275 16253 37276
rect 20140 37232 20180 37276
rect 21424 37232 21504 37252
rect 8131 37192 8140 37232
rect 8180 37192 8332 37232
rect 8372 37192 8381 37232
rect 18307 37192 18316 37232
rect 18356 37192 18892 37232
rect 18932 37192 18941 37232
rect 20140 37192 21504 37232
rect 21424 37172 21504 37192
rect 7939 37148 7997 37149
rect 15715 37148 15773 37149
rect 1315 37108 1324 37148
rect 1364 37108 6740 37148
rect 7372 37108 7468 37148
rect 7508 37108 7517 37148
rect 7939 37108 7948 37148
rect 7988 37108 15724 37148
rect 15764 37108 15773 37148
rect 0 37064 80 37084
rect 6700 37064 6740 37108
rect 7939 37107 7997 37108
rect 15715 37107 15773 37108
rect 17059 37148 17117 37149
rect 17059 37108 17068 37148
rect 17108 37108 21332 37148
rect 17059 37107 17117 37108
rect 11203 37064 11261 37065
rect 0 37024 3148 37064
rect 3188 37024 3197 37064
rect 4919 37024 4928 37064
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 5296 37024 5305 37064
rect 6403 37024 6412 37064
rect 6452 37024 6461 37064
rect 6691 37024 6700 37064
rect 6740 37024 7796 37064
rect 0 37004 80 37024
rect 6412 36980 6452 37024
rect 7756 36980 7796 37024
rect 11203 37024 11212 37064
rect 11252 37024 17660 37064
rect 20039 37024 20048 37064
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20416 37024 20425 37064
rect 11203 37023 11261 37024
rect 17620 36980 17660 37024
rect 6412 36940 7660 36980
rect 7700 36940 7709 36980
rect 7756 36940 11360 36980
rect 15427 36940 15436 36980
rect 15476 36940 15628 36980
rect 15668 36940 15677 36980
rect 17620 36940 20180 36980
rect 6979 36896 7037 36897
rect 11320 36896 11360 36940
rect 1411 36856 1420 36896
rect 1460 36856 1804 36896
rect 1844 36856 1853 36896
rect 4291 36856 4300 36896
rect 4340 36856 5452 36896
rect 5492 36856 5501 36896
rect 5548 36856 6740 36896
rect 6787 36856 6796 36896
rect 6836 36856 6988 36896
rect 7028 36856 7037 36896
rect 7555 36856 7564 36896
rect 7604 36856 8140 36896
rect 8180 36856 8189 36896
rect 11320 36856 15052 36896
rect 15092 36856 17068 36896
rect 17108 36856 18124 36896
rect 18164 36856 18173 36896
rect 739 36812 797 36813
rect 5548 36812 5588 36856
rect 6700 36812 6740 36856
rect 6979 36855 7037 36856
rect 739 36772 748 36812
rect 788 36772 4012 36812
rect 4052 36772 4061 36812
rect 4483 36772 4492 36812
rect 4532 36772 5588 36812
rect 6211 36772 6220 36812
rect 6260 36772 6604 36812
rect 6644 36772 6653 36812
rect 6700 36772 11788 36812
rect 11828 36772 14284 36812
rect 14324 36772 14333 36812
rect 14563 36772 14572 36812
rect 14612 36772 16684 36812
rect 16724 36772 16733 36812
rect 739 36771 797 36772
rect 0 36728 80 36748
rect 5827 36728 5885 36729
rect 19363 36728 19421 36729
rect 0 36688 1420 36728
rect 1460 36688 1469 36728
rect 4099 36688 4108 36728
rect 4148 36688 5260 36728
rect 5300 36688 5740 36728
rect 5780 36688 5836 36728
rect 5876 36688 5904 36728
rect 6307 36688 6316 36728
rect 6356 36688 7276 36728
rect 7316 36688 7325 36728
rect 11971 36688 11980 36728
rect 12020 36688 12748 36728
rect 12788 36688 12797 36728
rect 13603 36688 13612 36728
rect 13652 36688 15724 36728
rect 15764 36688 15773 36728
rect 19278 36688 19372 36728
rect 19412 36688 19421 36728
rect 20140 36728 20180 36940
rect 21292 36896 21332 37108
rect 21424 36896 21504 36916
rect 21292 36856 21504 36896
rect 21424 36836 21504 36856
rect 20140 36688 21332 36728
rect 0 36668 80 36688
rect 5827 36687 5885 36688
rect 19363 36687 19421 36688
rect 12739 36644 12797 36645
rect 5635 36604 5644 36644
rect 5684 36604 7756 36644
rect 7796 36604 7805 36644
rect 8899 36604 8908 36644
rect 8948 36604 11360 36644
rect 9091 36560 9149 36561
rect 11320 36560 11360 36604
rect 12739 36604 12748 36644
rect 12788 36604 12844 36644
rect 12884 36604 12893 36644
rect 13315 36604 13324 36644
rect 13364 36604 13373 36644
rect 14083 36604 14092 36644
rect 14132 36604 15820 36644
rect 15860 36604 16108 36644
rect 16148 36604 16157 36644
rect 17347 36604 17356 36644
rect 17396 36604 21100 36644
rect 21140 36604 21149 36644
rect 12739 36603 12797 36604
rect 13324 36560 13364 36604
rect 16675 36560 16733 36561
rect 19267 36560 19325 36561
rect 2659 36520 2668 36560
rect 2708 36520 4588 36560
rect 4628 36520 4637 36560
rect 5443 36520 5452 36560
rect 5492 36520 6356 36560
rect 6316 36476 6356 36520
rect 9091 36520 9100 36560
rect 9140 36520 9676 36560
rect 9716 36520 9725 36560
rect 11320 36520 13036 36560
rect 13076 36520 13364 36560
rect 15523 36520 15532 36560
rect 15572 36520 16300 36560
rect 16340 36520 16349 36560
rect 16675 36520 16684 36560
rect 16724 36520 17452 36560
rect 17492 36520 17501 36560
rect 17923 36520 17932 36560
rect 17972 36520 18508 36560
rect 18548 36520 18557 36560
rect 18787 36520 18796 36560
rect 18836 36520 19276 36560
rect 19316 36520 19325 36560
rect 21292 36560 21332 36688
rect 21424 36560 21504 36580
rect 21292 36520 21504 36560
rect 9091 36519 9149 36520
rect 16675 36519 16733 36520
rect 19267 36519 19325 36520
rect 21424 36500 21504 36520
rect 6307 36436 6316 36476
rect 6356 36436 6365 36476
rect 6595 36436 6604 36476
rect 6644 36436 11692 36476
rect 11732 36436 12460 36476
rect 12500 36436 12509 36476
rect 0 36392 80 36412
rect 2755 36392 2813 36393
rect 10435 36392 10493 36393
rect 0 36352 1324 36392
rect 1364 36352 2764 36392
rect 2804 36352 2813 36392
rect 4195 36352 4204 36392
rect 4244 36352 9908 36392
rect 0 36332 80 36352
rect 2755 36351 2813 36352
rect 9868 36308 9908 36352
rect 10435 36352 10444 36392
rect 10484 36352 21004 36392
rect 21044 36352 21053 36392
rect 10435 36351 10493 36352
rect 18403 36308 18461 36309
rect 3679 36268 3688 36308
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 4056 36268 4065 36308
rect 6019 36268 6028 36308
rect 6068 36268 6700 36308
rect 6740 36268 6749 36308
rect 9283 36268 9292 36308
rect 9332 36268 9484 36308
rect 9524 36268 9533 36308
rect 9868 36268 10348 36308
rect 10388 36268 10397 36308
rect 11395 36268 11404 36308
rect 11444 36268 16972 36308
rect 17012 36268 17021 36308
rect 17539 36268 17548 36308
rect 17588 36268 18412 36308
rect 18452 36268 18461 36308
rect 18799 36268 18808 36308
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 19176 36268 19185 36308
rect 19459 36268 19468 36308
rect 19508 36268 20852 36308
rect 18403 36267 18461 36268
rect 9859 36224 9917 36225
rect 20812 36224 20852 36268
rect 21424 36224 21504 36244
rect 9859 36184 9868 36224
rect 9908 36184 20716 36224
rect 20756 36184 20765 36224
rect 20812 36184 21504 36224
rect 9859 36183 9917 36184
rect 21424 36164 21504 36184
rect 5443 36100 5452 36140
rect 5492 36100 5836 36140
rect 5876 36100 5885 36140
rect 6403 36100 6412 36140
rect 6452 36100 6988 36140
rect 7028 36100 7037 36140
rect 8419 36100 8428 36140
rect 8468 36100 9868 36140
rect 9908 36100 9917 36140
rect 10819 36100 10828 36140
rect 10868 36100 11404 36140
rect 11444 36100 11453 36140
rect 14755 36100 14764 36140
rect 14804 36100 14956 36140
rect 14996 36100 15005 36140
rect 0 36056 80 36076
rect 9379 36056 9437 36057
rect 17059 36056 17117 36057
rect 0 36016 6604 36056
rect 6644 36016 6653 36056
rect 9379 36016 9388 36056
rect 9428 36016 17068 36056
rect 17108 36016 17117 36056
rect 0 35996 80 36016
rect 9379 36015 9437 36016
rect 17059 36015 17117 36016
rect 8524 35932 9292 35972
rect 9332 35932 9580 35972
rect 9620 35932 9629 35972
rect 9859 35932 9868 35972
rect 9908 35932 12364 35972
rect 12404 35932 12413 35972
rect 15724 35932 20812 35972
rect 20852 35932 20861 35972
rect 7843 35888 7901 35889
rect 5923 35848 5932 35888
rect 5972 35848 7564 35888
rect 7604 35848 7613 35888
rect 7747 35848 7756 35888
rect 7796 35848 7852 35888
rect 7892 35848 7901 35888
rect 7843 35847 7901 35848
rect 8524 35804 8564 35932
rect 8611 35888 8669 35889
rect 15724 35888 15764 35932
rect 8611 35848 8620 35888
rect 8660 35848 15764 35888
rect 17443 35888 17501 35889
rect 21424 35888 21504 35908
rect 17443 35848 17452 35888
rect 17492 35848 21504 35888
rect 8611 35847 8669 35848
rect 17443 35847 17501 35848
rect 21424 35828 21504 35848
rect 6691 35764 6700 35804
rect 6740 35764 8564 35804
rect 10339 35764 10348 35804
rect 10388 35764 18220 35804
rect 18260 35764 18508 35804
rect 18548 35764 18557 35804
rect 19747 35764 19756 35804
rect 19796 35764 19805 35804
rect 0 35720 80 35740
rect 7459 35720 7517 35721
rect 11011 35720 11069 35721
rect 0 35680 4492 35720
rect 4532 35680 4541 35720
rect 5251 35680 5260 35720
rect 5300 35680 5644 35720
rect 5684 35680 5693 35720
rect 6595 35680 6604 35720
rect 6644 35680 7468 35720
rect 7508 35680 8428 35720
rect 8468 35680 8477 35720
rect 9187 35680 9196 35720
rect 9236 35680 11020 35720
rect 11060 35680 11069 35720
rect 0 35660 80 35680
rect 7459 35679 7517 35680
rect 11011 35679 11069 35680
rect 11212 35636 11252 35764
rect 19756 35720 19796 35764
rect 12259 35680 12268 35720
rect 12308 35680 12844 35720
rect 12884 35680 12893 35720
rect 14467 35680 14476 35720
rect 14516 35680 14860 35720
rect 14900 35680 14909 35720
rect 15619 35680 15628 35720
rect 15668 35680 16492 35720
rect 16532 35680 16541 35720
rect 18115 35680 18124 35720
rect 18164 35680 19796 35720
rect 6979 35596 6988 35636
rect 7028 35596 7372 35636
rect 7412 35596 7421 35636
rect 11203 35596 11212 35636
rect 11252 35596 11261 35636
rect 11320 35596 16876 35636
rect 16916 35596 16925 35636
rect 5827 35552 5885 35553
rect 11320 35552 11360 35596
rect 21424 35552 21504 35572
rect 4919 35512 4928 35552
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 5296 35512 5305 35552
rect 5827 35512 5836 35552
rect 5876 35512 11360 35552
rect 20039 35512 20048 35552
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20416 35512 20425 35552
rect 21292 35512 21504 35552
rect 5827 35511 5885 35512
rect 4003 35428 4012 35468
rect 4052 35428 13132 35468
rect 13172 35428 13420 35468
rect 13460 35428 13469 35468
rect 16291 35428 16300 35468
rect 16340 35428 16876 35468
rect 16916 35428 17260 35468
rect 17300 35428 17452 35468
rect 17492 35428 18124 35468
rect 18164 35428 18173 35468
rect 0 35384 80 35404
rect 4012 35384 4052 35428
rect 8419 35384 8477 35385
rect 21292 35384 21332 35512
rect 21424 35492 21504 35512
rect 0 35344 4052 35384
rect 5443 35344 5452 35384
rect 5492 35344 5932 35384
rect 5972 35344 7180 35384
rect 7220 35344 7229 35384
rect 8419 35344 8428 35384
rect 8468 35344 21332 35384
rect 0 35324 80 35344
rect 8419 35343 8477 35344
rect 3523 35300 3581 35301
rect 8611 35300 8669 35301
rect 9667 35300 9725 35301
rect 19747 35300 19805 35301
rect 3523 35260 3532 35300
rect 3572 35260 3724 35300
rect 3764 35260 3773 35300
rect 6019 35260 6028 35300
rect 6068 35260 7468 35300
rect 7508 35260 7517 35300
rect 8526 35260 8620 35300
rect 8660 35260 8669 35300
rect 9582 35260 9676 35300
rect 9716 35260 9725 35300
rect 3523 35259 3581 35260
rect 8611 35259 8669 35260
rect 9667 35259 9725 35260
rect 17620 35260 17932 35300
rect 17972 35260 17981 35300
rect 19747 35260 19756 35300
rect 19796 35260 19852 35300
rect 19892 35260 19901 35300
rect 16867 35216 16925 35217
rect 17620 35216 17660 35260
rect 19747 35259 19805 35260
rect 21424 35216 21504 35236
rect 1987 35176 1996 35216
rect 2036 35176 2668 35216
rect 2708 35176 2717 35216
rect 2947 35176 2956 35216
rect 2996 35176 5260 35216
rect 5300 35176 5309 35216
rect 5443 35176 5452 35216
rect 5492 35176 6124 35216
rect 6164 35176 6173 35216
rect 6403 35176 6412 35216
rect 6452 35176 7084 35216
rect 7124 35176 7133 35216
rect 8995 35176 9004 35216
rect 9044 35176 10444 35216
rect 10484 35176 10924 35216
rect 10964 35176 10973 35216
rect 16867 35176 16876 35216
rect 16916 35176 17068 35216
rect 17108 35176 17117 35216
rect 17347 35176 17356 35216
rect 17396 35176 17660 35216
rect 17731 35176 17740 35216
rect 17780 35176 18508 35216
rect 18548 35176 19756 35216
rect 19796 35176 19805 35216
rect 21292 35176 21504 35216
rect 10924 35132 10964 35176
rect 16867 35175 16925 35176
rect 12739 35132 12797 35133
rect 21292 35132 21332 35176
rect 21424 35156 21504 35176
rect 5827 35092 5836 35132
rect 5876 35092 6316 35132
rect 6356 35092 6365 35132
rect 10924 35092 12076 35132
rect 12116 35092 12125 35132
rect 12654 35092 12748 35132
rect 12788 35092 12797 35132
rect 12739 35091 12797 35092
rect 14668 35092 17260 35132
rect 17300 35092 17836 35132
rect 17876 35092 17885 35132
rect 20236 35092 21332 35132
rect 0 35048 80 35068
rect 0 35008 2860 35048
rect 2900 35008 2909 35048
rect 6211 35008 6220 35048
rect 6260 35008 10348 35048
rect 10388 35008 10397 35048
rect 12835 35008 12844 35048
rect 12884 35008 13132 35048
rect 13172 35008 13181 35048
rect 0 34988 80 35008
rect 14668 34964 14708 35092
rect 16876 35048 16916 35092
rect 16867 35008 16876 35048
rect 16916 35008 16956 35048
rect 1795 34924 1804 34964
rect 1844 34924 2036 34964
rect 4963 34924 4972 34964
rect 5012 34924 14708 34964
rect 14755 34964 14813 34965
rect 14755 34924 14764 34964
rect 14804 34924 20180 34964
rect 1996 34880 2036 34924
rect 14755 34923 14813 34924
rect 11203 34880 11261 34881
rect 15619 34880 15677 34881
rect 1987 34840 1996 34880
rect 2036 34840 2045 34880
rect 5251 34840 5260 34880
rect 5300 34840 5644 34880
rect 5684 34840 5693 34880
rect 6595 34840 6604 34880
rect 6644 34840 7660 34880
rect 7700 34840 7709 34880
rect 11011 34840 11020 34880
rect 11060 34840 11212 34880
rect 11252 34840 11261 34880
rect 12259 34840 12268 34880
rect 12308 34840 12556 34880
rect 12596 34840 15628 34880
rect 15668 34840 15677 34880
rect 11203 34839 11261 34840
rect 15619 34839 15677 34840
rect 18403 34880 18461 34881
rect 20140 34880 20180 34924
rect 20236 34880 20276 35092
rect 21424 34880 21504 34900
rect 18403 34840 18412 34880
rect 18452 34840 19316 34880
rect 20140 34840 20276 34880
rect 20332 34840 21504 34880
rect 18403 34839 18461 34840
rect 16867 34796 16925 34797
rect 19276 34796 19316 34840
rect 20332 34796 20372 34840
rect 21424 34820 21504 34840
rect 3679 34756 3688 34796
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 4056 34756 4065 34796
rect 6211 34756 6220 34796
rect 6260 34756 11404 34796
rect 11444 34756 11453 34796
rect 11500 34756 14476 34796
rect 14516 34756 14525 34796
rect 16867 34756 16876 34796
rect 16916 34756 17068 34796
rect 17108 34756 17117 34796
rect 18799 34756 18808 34796
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 19176 34756 19185 34796
rect 19276 34756 20372 34796
rect 0 34712 80 34732
rect 2179 34712 2237 34713
rect 6883 34712 6941 34713
rect 11500 34712 11540 34756
rect 16867 34755 16925 34756
rect 20611 34712 20669 34713
rect 0 34672 2188 34712
rect 2228 34672 2237 34712
rect 3235 34672 3244 34712
rect 3284 34672 3532 34712
rect 3572 34672 3581 34712
rect 5539 34672 5548 34712
rect 5588 34672 5836 34712
rect 5876 34672 5885 34712
rect 6691 34672 6700 34712
rect 6740 34672 6892 34712
rect 6932 34672 6941 34712
rect 8899 34672 8908 34712
rect 8948 34672 11540 34712
rect 12547 34672 12556 34712
rect 12596 34672 12748 34712
rect 12788 34672 12797 34712
rect 19939 34672 19948 34712
rect 19988 34672 20620 34712
rect 20660 34672 20669 34712
rect 0 34652 80 34672
rect 2179 34671 2237 34672
rect 6883 34671 6941 34672
rect 20611 34671 20669 34672
rect 8803 34628 8861 34629
rect 20707 34628 20765 34629
rect 1315 34588 1324 34628
rect 1364 34588 4492 34628
rect 4532 34588 4541 34628
rect 6499 34588 6508 34628
rect 6548 34588 8812 34628
rect 8852 34588 8861 34628
rect 11011 34588 11020 34628
rect 11060 34588 20716 34628
rect 20756 34588 20765 34628
rect 8803 34587 8861 34588
rect 20707 34587 20765 34588
rect 21424 34544 21504 34564
rect 5443 34504 5452 34544
rect 5492 34504 6316 34544
rect 6356 34504 7180 34544
rect 7220 34504 7229 34544
rect 13603 34504 13612 34544
rect 13652 34504 13661 34544
rect 20707 34504 20716 34544
rect 20756 34504 21504 34544
rect 13612 34460 13652 34504
rect 21424 34484 21504 34504
rect 4003 34420 4012 34460
rect 4052 34420 13556 34460
rect 13612 34420 13804 34460
rect 13844 34420 13853 34460
rect 0 34376 80 34396
rect 7747 34376 7805 34377
rect 12355 34376 12413 34377
rect 13411 34376 13469 34377
rect 0 34336 1612 34376
rect 1652 34336 4204 34376
rect 4244 34336 4972 34376
rect 5012 34336 5021 34376
rect 5827 34336 5836 34376
rect 5876 34336 7084 34376
rect 7124 34336 7133 34376
rect 7555 34336 7564 34376
rect 7604 34336 7756 34376
rect 7796 34336 8524 34376
rect 8564 34336 8573 34376
rect 8803 34336 8812 34376
rect 8852 34336 9004 34376
rect 9044 34336 9053 34376
rect 9763 34336 9772 34376
rect 9812 34336 9964 34376
rect 10004 34336 10013 34376
rect 12270 34336 12364 34376
rect 12404 34336 13420 34376
rect 13460 34336 13469 34376
rect 13516 34376 13556 34420
rect 21379 34376 21437 34377
rect 13516 34336 13844 34376
rect 14179 34336 14188 34376
rect 14228 34336 14668 34376
rect 14708 34336 15820 34376
rect 15860 34336 17740 34376
rect 17780 34336 17789 34376
rect 19651 34336 19660 34376
rect 19700 34336 21388 34376
rect 21428 34336 21437 34376
rect 0 34316 80 34336
rect 7747 34335 7805 34336
rect 12355 34335 12413 34336
rect 13411 34335 13469 34336
rect 6691 34292 6749 34293
rect 6606 34252 6700 34292
rect 6740 34252 6749 34292
rect 6691 34251 6749 34252
rect 7363 34292 7421 34293
rect 13804 34292 13844 34336
rect 21379 34335 21437 34336
rect 16771 34292 16829 34293
rect 7363 34252 7372 34292
rect 7412 34252 7660 34292
rect 7700 34252 13708 34292
rect 13748 34252 13757 34292
rect 13804 34252 16780 34292
rect 16820 34252 16829 34292
rect 19555 34252 19564 34292
rect 19604 34252 20908 34292
rect 20948 34252 20957 34292
rect 7363 34251 7421 34252
rect 16771 34251 16829 34252
rect 10531 34208 10589 34209
rect 11299 34208 11357 34209
rect 21424 34208 21504 34228
rect 2851 34168 2860 34208
rect 2900 34168 5396 34208
rect 6019 34168 6028 34208
rect 6068 34168 6796 34208
rect 6836 34168 6845 34208
rect 6892 34168 10540 34208
rect 10580 34168 10636 34208
rect 10676 34168 10685 34208
rect 11299 34168 11308 34208
rect 11348 34168 21504 34208
rect 1411 34124 1469 34125
rect 460 34084 1420 34124
rect 1460 34084 4012 34124
rect 4052 34084 4061 34124
rect 0 34040 80 34060
rect 460 34040 500 34084
rect 1411 34083 1469 34084
rect 4675 34040 4733 34041
rect 5356 34040 5396 34168
rect 6019 34124 6077 34125
rect 6892 34124 6932 34168
rect 10531 34167 10589 34168
rect 11299 34167 11357 34168
rect 21424 34148 21504 34168
rect 6019 34084 6028 34124
rect 6068 34084 6220 34124
rect 6260 34084 6269 34124
rect 6316 34084 6932 34124
rect 7171 34084 7180 34124
rect 7220 34084 15860 34124
rect 6019 34083 6077 34084
rect 6316 34040 6356 34084
rect 8515 34040 8573 34041
rect 15820 34040 15860 34084
rect 16771 34040 16829 34041
rect 17155 34040 17213 34041
rect 0 34000 500 34040
rect 547 34000 556 34040
rect 596 34000 1804 34040
rect 1844 34000 4684 34040
rect 4724 34000 4733 34040
rect 4919 34000 4928 34040
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 5296 34000 5305 34040
rect 5356 34000 6356 34040
rect 6499 34000 6508 34040
rect 6548 34000 7564 34040
rect 7604 34000 7613 34040
rect 8515 34000 8524 34040
rect 8564 34000 8716 34040
rect 8756 34000 8765 34040
rect 8995 34000 9004 34040
rect 9044 34000 9292 34040
rect 9332 34000 9341 34040
rect 12643 34000 12652 34040
rect 12692 34000 13612 34040
rect 13652 34000 14188 34040
rect 14228 34000 14237 34040
rect 15811 34000 15820 34040
rect 15860 34000 15869 34040
rect 16771 34000 16780 34040
rect 16820 34000 17164 34040
rect 17204 34000 17213 34040
rect 17635 34000 17644 34040
rect 17684 34000 17932 34040
rect 17972 34000 17981 34040
rect 18403 34000 18412 34040
rect 18452 34000 18700 34040
rect 18740 34000 18749 34040
rect 20039 34000 20048 34040
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20416 34000 20425 34040
rect 0 33980 80 34000
rect 4675 33999 4733 34000
rect 8515 33999 8573 34000
rect 16771 33999 16829 34000
rect 17155 33999 17213 34000
rect 14467 33956 14525 33957
rect 1411 33916 1420 33956
rect 1460 33916 2476 33956
rect 2516 33916 11500 33956
rect 11540 33916 11549 33956
rect 11596 33916 14476 33956
rect 14516 33916 17660 33956
rect 4003 33872 4061 33873
rect 8227 33872 8285 33873
rect 11596 33872 11636 33916
rect 14467 33915 14525 33916
rect 17620 33872 17660 33916
rect 21424 33872 21504 33892
rect 3918 33832 4012 33872
rect 4052 33832 4061 33872
rect 6115 33832 6124 33872
rect 6164 33832 7468 33872
rect 7508 33832 7517 33872
rect 8142 33832 8236 33872
rect 8276 33832 8285 33872
rect 11395 33832 11404 33872
rect 11444 33832 11636 33872
rect 12643 33832 12652 33872
rect 12692 33832 13516 33872
rect 13556 33832 13565 33872
rect 15715 33832 15724 33872
rect 15764 33832 16204 33872
rect 16244 33832 16253 33872
rect 17620 33832 18932 33872
rect 20803 33832 20812 33872
rect 20852 33832 21504 33872
rect 4003 33831 4061 33832
rect 8227 33831 8285 33832
rect 18892 33788 18932 33832
rect 21424 33812 21504 33832
rect 2467 33748 2476 33788
rect 2516 33748 3052 33788
rect 3092 33748 3101 33788
rect 5731 33748 5740 33788
rect 5780 33748 6508 33788
rect 6548 33748 7660 33788
rect 7700 33748 7709 33788
rect 8419 33748 8428 33788
rect 8468 33748 8716 33788
rect 8756 33748 8765 33788
rect 11011 33748 11020 33788
rect 11060 33748 17644 33788
rect 17684 33748 17693 33788
rect 18883 33748 18892 33788
rect 18932 33748 19468 33788
rect 19508 33748 19517 33788
rect 0 33704 80 33724
rect 1987 33704 2045 33705
rect 0 33664 1996 33704
rect 2036 33664 2045 33704
rect 0 33644 80 33664
rect 1987 33663 2045 33664
rect 2179 33704 2237 33705
rect 8419 33704 8477 33705
rect 11011 33704 11069 33705
rect 16579 33704 16637 33705
rect 2179 33664 2188 33704
rect 2228 33664 4300 33704
rect 4340 33664 4349 33704
rect 6019 33664 6028 33704
rect 6068 33664 7276 33704
rect 7316 33664 7852 33704
rect 7892 33664 7901 33704
rect 8419 33664 8428 33704
rect 8468 33664 11020 33704
rect 11060 33664 11069 33704
rect 2179 33663 2237 33664
rect 8419 33663 8477 33664
rect 11011 33663 11069 33664
rect 11320 33664 13324 33704
rect 13364 33664 13940 33704
rect 13987 33664 13996 33704
rect 14036 33664 14668 33704
rect 14708 33664 14717 33704
rect 16494 33664 16588 33704
rect 16628 33664 16637 33704
rect 6403 33620 6461 33621
rect 11320 33620 11360 33664
rect 13900 33620 13940 33664
rect 16579 33663 16637 33664
rect 1123 33580 1132 33620
rect 1172 33580 6412 33620
rect 6452 33580 6461 33620
rect 6403 33579 6461 33580
rect 6604 33580 11360 33620
rect 11491 33580 11500 33620
rect 11540 33580 13420 33620
rect 13460 33580 13469 33620
rect 13900 33580 19564 33620
rect 19604 33580 19613 33620
rect 2755 33536 2813 33537
rect 6604 33536 6644 33580
rect 8419 33536 8477 33537
rect 9091 33536 9149 33537
rect 739 33496 748 33536
rect 788 33496 1036 33536
rect 1076 33496 1085 33536
rect 2755 33496 2764 33536
rect 2804 33496 6548 33536
rect 6595 33496 6604 33536
rect 6644 33496 6653 33536
rect 7756 33496 8428 33536
rect 8468 33496 8477 33536
rect 8803 33496 8812 33536
rect 8852 33496 9100 33536
rect 9140 33496 9149 33536
rect 2755 33495 2813 33496
rect 4675 33452 4733 33453
rect 6508 33452 6548 33496
rect 7756 33452 7796 33496
rect 8419 33495 8477 33496
rect 9091 33495 9149 33496
rect 18499 33536 18557 33537
rect 21424 33536 21504 33556
rect 18499 33496 18508 33536
rect 18548 33496 19084 33536
rect 19124 33496 19133 33536
rect 21283 33496 21292 33536
rect 21332 33496 21504 33536
rect 18499 33495 18557 33496
rect 21424 33476 21504 33496
rect 8227 33452 8285 33453
rect 3139 33412 3148 33452
rect 3188 33412 3820 33452
rect 3860 33412 3869 33452
rect 4675 33412 4684 33452
rect 4724 33412 4820 33452
rect 6508 33412 7796 33452
rect 7843 33412 7852 33452
rect 7892 33412 8236 33452
rect 8276 33412 8285 33452
rect 4675 33411 4733 33412
rect 0 33368 80 33388
rect 4780 33368 4820 33412
rect 8227 33411 8285 33412
rect 8332 33412 11360 33452
rect 16675 33412 16684 33452
rect 16724 33412 17356 33452
rect 17396 33412 17405 33452
rect 8332 33368 8372 33412
rect 8803 33368 8861 33369
rect 9955 33368 10013 33369
rect 10147 33368 10205 33369
rect 0 33328 4588 33368
rect 4628 33328 4637 33368
rect 4780 33328 8372 33368
rect 8718 33328 8812 33368
rect 8852 33328 8861 33368
rect 9379 33328 9388 33368
rect 9428 33328 9772 33368
rect 9812 33328 9821 33368
rect 9955 33328 9964 33368
rect 10004 33328 10156 33368
rect 10196 33328 10205 33368
rect 11320 33368 11360 33412
rect 11320 33328 16588 33368
rect 16628 33328 16637 33368
rect 0 33308 80 33328
rect 8803 33327 8861 33328
rect 9955 33327 10013 33328
rect 10147 33327 10205 33328
rect 3679 33244 3688 33284
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 4056 33244 4065 33284
rect 6595 33244 6604 33284
rect 6644 33244 11020 33284
rect 11060 33244 11069 33284
rect 18799 33244 18808 33284
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 19176 33244 19185 33284
rect 20035 33244 20044 33284
rect 20084 33244 20524 33284
rect 20564 33244 20573 33284
rect 21424 33200 21504 33220
rect 643 33160 652 33200
rect 692 33160 1132 33200
rect 1172 33160 1181 33200
rect 8035 33160 8044 33200
rect 8084 33160 8236 33200
rect 8276 33160 8285 33200
rect 8419 33160 8428 33200
rect 8468 33160 8620 33200
rect 8660 33160 8669 33200
rect 9379 33160 9388 33200
rect 9428 33160 12268 33200
rect 12308 33160 12317 33200
rect 14467 33160 14476 33200
rect 14516 33160 21504 33200
rect 21424 33140 21504 33160
rect 6979 33076 6988 33116
rect 7028 33076 7948 33116
rect 7988 33076 7997 33116
rect 9859 33076 9868 33116
rect 9908 33076 10156 33116
rect 10196 33076 10205 33116
rect 17923 33076 17932 33116
rect 17972 33076 19180 33116
rect 19220 33076 19229 33116
rect 0 33032 80 33052
rect 4675 33032 4733 33033
rect 8611 33032 8669 33033
rect 9379 33032 9437 33033
rect 13699 33032 13757 33033
rect 15235 33032 15293 33033
rect 0 32992 172 33032
rect 212 32992 221 33032
rect 2500 32992 4684 33032
rect 4724 32992 7316 33032
rect 8526 32992 8620 33032
rect 8660 32992 8669 33032
rect 9187 32992 9196 33032
rect 9236 32992 9388 33032
rect 9428 32992 9437 33032
rect 9571 32992 9580 33032
rect 9620 32992 13708 33032
rect 13748 32992 13757 33032
rect 14371 32992 14380 33032
rect 14420 32992 14764 33032
rect 14804 32992 14813 33032
rect 15150 32992 15244 33032
rect 15284 32992 15293 33032
rect 0 32972 80 32992
rect 2500 32948 2540 32992
rect 4675 32991 4733 32992
rect 7276 32948 7316 32992
rect 8611 32991 8669 32992
rect 9379 32991 9437 32992
rect 13699 32991 13757 32992
rect 15235 32991 15293 32992
rect 18499 32948 18557 32949
rect 1315 32908 1324 32948
rect 1364 32908 1708 32948
rect 1748 32908 2540 32948
rect 5923 32908 5932 32948
rect 5972 32908 7180 32948
rect 7220 32908 7229 32948
rect 7276 32908 10580 32948
rect 10627 32908 10636 32948
rect 10676 32908 11596 32948
rect 11636 32908 12268 32948
rect 12308 32908 12317 32948
rect 13411 32908 13420 32948
rect 13460 32908 18508 32948
rect 18548 32908 18557 32948
rect 3235 32864 3293 32865
rect 10540 32864 10580 32908
rect 18499 32907 18557 32908
rect 17923 32864 17981 32865
rect 21424 32864 21504 32884
rect 3216 32824 3244 32864
rect 3284 32824 3340 32864
rect 3380 32824 5836 32864
rect 5876 32824 5885 32864
rect 6499 32824 6508 32864
rect 6548 32824 7372 32864
rect 7412 32824 7421 32864
rect 7468 32824 9388 32864
rect 9428 32824 9437 32864
rect 10540 32824 16012 32864
rect 16052 32824 17932 32864
rect 17972 32824 17981 32864
rect 21091 32824 21100 32864
rect 21140 32824 21504 32864
rect 3235 32823 3293 32824
rect 6883 32780 6941 32781
rect 7468 32780 7508 32824
rect 17923 32823 17981 32824
rect 21424 32804 21504 32824
rect 8515 32780 8573 32781
rect 9379 32780 9437 32781
rect 14659 32780 14717 32781
rect 15523 32780 15581 32781
rect 4483 32740 4492 32780
rect 4532 32740 6836 32780
rect 0 32696 80 32716
rect 5827 32696 5885 32697
rect 6796 32696 6836 32740
rect 6883 32740 6892 32780
rect 6932 32740 7084 32780
rect 7124 32740 7133 32780
rect 7180 32740 7508 32780
rect 8131 32740 8140 32780
rect 8180 32740 8524 32780
rect 8564 32740 8573 32780
rect 8707 32740 8716 32780
rect 8756 32740 9388 32780
rect 9428 32740 9772 32780
rect 9812 32740 9821 32780
rect 10051 32740 10060 32780
rect 10100 32740 10348 32780
rect 10388 32740 10397 32780
rect 14659 32740 14668 32780
rect 14708 32740 15532 32780
rect 15572 32740 15581 32780
rect 18787 32740 18796 32780
rect 18836 32740 19468 32780
rect 19508 32740 19517 32780
rect 6883 32739 6941 32740
rect 7180 32696 7220 32740
rect 8515 32739 8573 32740
rect 9379 32739 9437 32740
rect 14659 32739 14717 32740
rect 15523 32739 15581 32740
rect 7459 32696 7517 32697
rect 10531 32696 10589 32697
rect 11491 32696 11549 32697
rect 0 32656 5780 32696
rect 0 32636 80 32656
rect 5740 32528 5780 32656
rect 5827 32656 5836 32696
rect 5876 32656 5932 32696
rect 5972 32656 5981 32696
rect 6796 32656 7220 32696
rect 7374 32656 7468 32696
rect 7508 32656 7517 32696
rect 5827 32655 5885 32656
rect 7459 32655 7517 32656
rect 7564 32656 9292 32696
rect 9332 32656 9341 32696
rect 10531 32656 10540 32696
rect 10580 32656 10732 32696
rect 10772 32656 10781 32696
rect 11011 32656 11020 32696
rect 11060 32656 11500 32696
rect 11540 32656 14572 32696
rect 14612 32656 14621 32696
rect 7564 32528 7604 32656
rect 10531 32655 10589 32656
rect 11491 32655 11549 32656
rect 8995 32572 9004 32612
rect 9044 32572 9676 32612
rect 9716 32572 9725 32612
rect 13891 32572 13900 32612
rect 13940 32572 20660 32612
rect 20620 32528 20660 32572
rect 21424 32528 21504 32548
rect 4919 32488 4928 32528
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 5296 32488 5305 32528
rect 5740 32488 7604 32528
rect 9091 32488 9100 32528
rect 9140 32488 9388 32528
rect 9428 32488 9437 32528
rect 20039 32488 20048 32528
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20416 32488 20425 32528
rect 20620 32488 21504 32528
rect 21424 32468 21504 32488
rect 547 32404 556 32444
rect 596 32404 14092 32444
rect 14132 32404 14141 32444
rect 0 32360 80 32380
rect 7747 32360 7805 32361
rect 15139 32360 15197 32361
rect 0 32320 7756 32360
rect 7796 32320 7805 32360
rect 8419 32320 8428 32360
rect 8468 32320 9100 32360
rect 9140 32320 9580 32360
rect 9620 32320 9629 32360
rect 15043 32320 15052 32360
rect 15092 32320 15148 32360
rect 15188 32320 15197 32360
rect 0 32300 80 32320
rect 7747 32319 7805 32320
rect 15139 32319 15197 32320
rect 3523 32276 3581 32277
rect 8515 32276 8573 32277
rect 3523 32236 3532 32276
rect 3572 32236 3724 32276
rect 3764 32236 3773 32276
rect 6604 32236 8524 32276
rect 8564 32236 8573 32276
rect 12163 32236 12172 32276
rect 12212 32236 12460 32276
rect 12500 32236 12509 32276
rect 19459 32236 19468 32276
rect 19508 32236 20180 32276
rect 3523 32235 3581 32236
rect 3043 32192 3101 32193
rect 67 32152 76 32192
rect 116 32152 2092 32192
rect 2132 32152 2141 32192
rect 2958 32152 3052 32192
rect 3092 32152 3101 32192
rect 3043 32151 3101 32152
rect 1891 32108 1949 32109
rect 1891 32068 1900 32108
rect 1940 32068 2572 32108
rect 2612 32068 2621 32108
rect 1891 32067 1949 32068
rect 0 32024 80 32044
rect 6604 32024 6644 32236
rect 8515 32235 8573 32236
rect 11011 32192 11069 32193
rect 15043 32192 15101 32193
rect 8515 32152 8524 32192
rect 8564 32152 9292 32192
rect 9332 32152 9341 32192
rect 9667 32152 9676 32192
rect 9716 32152 10156 32192
rect 10196 32152 10205 32192
rect 11011 32152 11020 32192
rect 11060 32152 11980 32192
rect 12020 32152 13900 32192
rect 13940 32152 13949 32192
rect 14958 32152 15052 32192
rect 15092 32152 15101 32192
rect 20140 32192 20180 32236
rect 21424 32192 21504 32212
rect 20140 32152 21504 32192
rect 11011 32151 11069 32152
rect 7555 32108 7613 32109
rect 13900 32108 13940 32152
rect 15043 32151 15101 32152
rect 21424 32132 21504 32152
rect 7555 32068 7564 32108
rect 7604 32068 12556 32108
rect 12596 32068 12605 32108
rect 13900 32068 14284 32108
rect 14324 32068 16300 32108
rect 16340 32068 16349 32108
rect 18307 32068 18316 32108
rect 18356 32068 18604 32108
rect 18644 32068 18653 32108
rect 7555 32067 7613 32068
rect 0 31984 6644 32024
rect 6883 31984 6892 32024
rect 6932 31984 12940 32024
rect 12980 31984 13132 32024
rect 13172 31984 13181 32024
rect 0 31964 80 31984
rect 5635 31940 5693 31941
rect 11299 31940 11357 31941
rect 5635 31900 5644 31940
rect 5684 31900 6988 31940
rect 7028 31900 8908 31940
rect 8948 31900 11308 31940
rect 11348 31900 11357 31940
rect 5635 31899 5693 31900
rect 11299 31899 11357 31900
rect 1603 31856 1661 31857
rect 4579 31856 4637 31857
rect 21424 31856 21504 31876
rect 1603 31816 1612 31856
rect 1652 31816 4588 31856
rect 4628 31816 5740 31856
rect 5780 31816 5789 31856
rect 6787 31816 6796 31856
rect 6836 31816 14036 31856
rect 20803 31816 20812 31856
rect 20852 31816 21504 31856
rect 1603 31815 1661 31816
rect 4579 31815 4637 31816
rect 9859 31772 9917 31773
rect 3679 31732 3688 31772
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 4056 31732 4065 31772
rect 9859 31732 9868 31772
rect 9908 31732 10060 31772
rect 10100 31732 10109 31772
rect 9859 31731 9917 31732
rect 0 31688 80 31708
rect 0 31648 2476 31688
rect 2516 31648 5644 31688
rect 5684 31648 8044 31688
rect 8084 31648 10156 31688
rect 10196 31648 10348 31688
rect 10388 31648 10397 31688
rect 0 31628 80 31648
rect 13996 31604 14036 31816
rect 21424 31796 21504 31816
rect 18799 31732 18808 31772
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 19176 31732 19185 31772
rect 15235 31688 15293 31689
rect 15235 31648 15244 31688
rect 15284 31648 15340 31688
rect 15380 31648 15389 31688
rect 15235 31647 15293 31648
rect 2275 31564 2284 31604
rect 2324 31564 2668 31604
rect 2708 31564 2717 31604
rect 5539 31564 5548 31604
rect 5588 31564 6740 31604
rect 6979 31564 6988 31604
rect 7028 31564 10636 31604
rect 10676 31564 10685 31604
rect 13987 31564 13996 31604
rect 14036 31564 15724 31604
rect 15764 31564 15773 31604
rect 6700 31520 6740 31564
rect 14563 31520 14621 31521
rect 17539 31520 17597 31521
rect 2563 31480 2572 31520
rect 2612 31480 2860 31520
rect 2900 31480 2909 31520
rect 5443 31480 5452 31520
rect 5492 31480 6604 31520
rect 6644 31480 6653 31520
rect 6700 31480 6796 31520
rect 6836 31480 6845 31520
rect 14563 31480 14572 31520
rect 14612 31480 17548 31520
rect 17588 31480 17597 31520
rect 14563 31479 14621 31480
rect 17539 31479 17597 31480
rect 20611 31520 20669 31521
rect 21424 31520 21504 31540
rect 20611 31480 20620 31520
rect 20660 31480 21504 31520
rect 20611 31479 20669 31480
rect 21424 31460 21504 31480
rect 1603 31436 1661 31437
rect 14179 31436 14237 31437
rect 14659 31436 14717 31437
rect 18499 31436 18557 31437
rect 1518 31396 1612 31436
rect 1652 31396 1661 31436
rect 1603 31395 1661 31396
rect 4204 31396 4684 31436
rect 4724 31396 4733 31436
rect 5635 31396 5644 31436
rect 5684 31396 6412 31436
rect 6452 31396 6461 31436
rect 14179 31396 14188 31436
rect 14228 31396 14668 31436
rect 14708 31396 14717 31436
rect 17251 31396 17260 31436
rect 17300 31396 17452 31436
rect 17492 31396 17972 31436
rect 0 31352 80 31372
rect 4204 31353 4244 31396
rect 14179 31395 14237 31396
rect 14659 31395 14717 31396
rect 4195 31352 4253 31353
rect 11491 31352 11549 31353
rect 17635 31352 17693 31353
rect 17932 31352 17972 31396
rect 18499 31396 18508 31436
rect 18548 31396 18988 31436
rect 19028 31396 19037 31436
rect 18499 31395 18557 31396
rect 0 31312 2956 31352
rect 2996 31312 3005 31352
rect 3427 31312 3436 31352
rect 3476 31312 3485 31352
rect 3907 31312 3916 31352
rect 3956 31312 4204 31352
rect 4244 31312 4253 31352
rect 4387 31312 4396 31352
rect 4436 31312 6508 31352
rect 6548 31312 7276 31352
rect 7316 31312 7325 31352
rect 8611 31312 8620 31352
rect 8660 31312 9292 31352
rect 9332 31312 9341 31352
rect 11299 31312 11308 31352
rect 11348 31312 11500 31352
rect 11540 31312 11549 31352
rect 11971 31312 11980 31352
rect 12020 31312 12652 31352
rect 12692 31312 13228 31352
rect 13268 31312 17644 31352
rect 17684 31312 17693 31352
rect 17923 31312 17932 31352
rect 17972 31312 18124 31352
rect 18164 31312 18173 31352
rect 0 31292 80 31312
rect 2371 31228 2380 31268
rect 2420 31228 2860 31268
rect 2900 31228 2909 31268
rect 3436 31184 3476 31312
rect 4195 31311 4253 31312
rect 11491 31311 11549 31312
rect 17635 31311 17693 31312
rect 5731 31268 5789 31269
rect 6499 31268 6557 31269
rect 8419 31268 8477 31269
rect 5059 31228 5068 31268
rect 5108 31228 5740 31268
rect 5780 31228 5789 31268
rect 6115 31228 6124 31268
rect 6164 31228 6508 31268
rect 6548 31228 8428 31268
rect 8468 31228 8477 31268
rect 5731 31227 5789 31228
rect 6499 31227 6557 31228
rect 8419 31227 8477 31228
rect 8707 31268 8765 31269
rect 8707 31228 8716 31268
rect 8756 31228 18508 31268
rect 18548 31228 18557 31268
rect 8707 31227 8765 31228
rect 7747 31184 7805 31185
rect 1699 31144 1708 31184
rect 1748 31144 3476 31184
rect 7651 31144 7660 31184
rect 7700 31144 7756 31184
rect 7796 31144 7805 31184
rect 7747 31143 7805 31144
rect 8899 31184 8957 31185
rect 21424 31184 21504 31204
rect 8899 31144 8908 31184
rect 8948 31144 9292 31184
rect 9332 31144 9341 31184
rect 14755 31144 14764 31184
rect 14804 31144 15148 31184
rect 15188 31144 15197 31184
rect 20131 31144 20140 31184
rect 20180 31144 20716 31184
rect 20756 31144 20765 31184
rect 20908 31144 21504 31184
rect 8899 31143 8957 31144
rect 2947 31060 2956 31100
rect 2996 31060 3148 31100
rect 3188 31060 3197 31100
rect 0 31016 80 31036
rect 13507 31016 13565 31017
rect 0 30976 364 31016
rect 404 30976 413 31016
rect 3811 30976 3820 31016
rect 3860 30976 4684 31016
rect 4724 30976 4733 31016
rect 4919 30976 4928 31016
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 5296 30976 5305 31016
rect 5827 30976 5836 31016
rect 5876 30976 6028 31016
rect 6068 30976 6077 31016
rect 6595 30976 6604 31016
rect 6644 30976 13036 31016
rect 13076 30976 13085 31016
rect 13315 30976 13324 31016
rect 13364 30976 13516 31016
rect 13556 30976 13565 31016
rect 16291 30976 16300 31016
rect 16340 30976 16684 31016
rect 16724 30976 16733 31016
rect 20039 30976 20048 31016
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20416 30976 20425 31016
rect 0 30956 80 30976
rect 13507 30975 13565 30976
rect 20908 30932 20948 31144
rect 21424 31124 21504 31144
rect 931 30892 940 30932
rect 980 30892 7124 30932
rect 11491 30892 11500 30932
rect 11540 30892 20948 30932
rect 4771 30808 4780 30848
rect 4820 30808 5260 30848
rect 5300 30808 5309 30848
rect 3043 30724 3052 30764
rect 3092 30724 3340 30764
rect 3380 30724 3389 30764
rect 0 30680 80 30700
rect 0 30640 1268 30680
rect 5539 30640 5548 30680
rect 5588 30640 5740 30680
rect 5780 30640 5789 30680
rect 6115 30640 6124 30680
rect 6164 30640 7028 30680
rect 0 30620 80 30640
rect 1228 30428 1268 30640
rect 2755 30596 2813 30597
rect 2659 30556 2668 30596
rect 2708 30556 2764 30596
rect 2804 30556 2813 30596
rect 3331 30556 3340 30596
rect 3380 30556 3532 30596
rect 3572 30556 3581 30596
rect 3811 30556 3820 30596
rect 3860 30556 6220 30596
rect 6260 30556 6836 30596
rect 2755 30555 2813 30556
rect 2467 30472 2476 30512
rect 2516 30472 2860 30512
rect 2900 30472 4492 30512
rect 4532 30472 5068 30512
rect 5108 30472 6124 30512
rect 6164 30472 6173 30512
rect 2755 30428 2813 30429
rect 6796 30428 6836 30556
rect 6988 30512 7028 30640
rect 7084 30596 7124 30892
rect 21424 30848 21504 30868
rect 13219 30808 13228 30848
rect 13268 30808 13516 30848
rect 13556 30808 13565 30848
rect 16483 30808 16492 30848
rect 16532 30808 21504 30848
rect 21424 30788 21504 30808
rect 9667 30764 9725 30765
rect 9667 30724 9676 30764
rect 9716 30724 9868 30764
rect 9908 30724 9917 30764
rect 17443 30724 17452 30764
rect 17492 30724 19276 30764
rect 19316 30724 19325 30764
rect 9667 30723 9725 30724
rect 7843 30680 7901 30681
rect 11011 30680 11069 30681
rect 15139 30680 15197 30681
rect 18595 30680 18653 30681
rect 7843 30640 7852 30680
rect 7892 30640 8236 30680
rect 8276 30640 8524 30680
rect 8564 30640 8573 30680
rect 8899 30640 8908 30680
rect 8948 30640 9484 30680
rect 9524 30640 10540 30680
rect 10580 30640 11020 30680
rect 11060 30640 11116 30680
rect 11156 30640 11165 30680
rect 11395 30640 11404 30680
rect 11444 30640 13132 30680
rect 13172 30640 13181 30680
rect 13891 30640 13900 30680
rect 13940 30640 14860 30680
rect 14900 30640 14909 30680
rect 15139 30640 15148 30680
rect 15188 30640 15244 30680
rect 15284 30640 15293 30680
rect 16483 30640 16492 30680
rect 16532 30640 17260 30680
rect 17300 30640 17309 30680
rect 18595 30640 18604 30680
rect 18644 30640 18796 30680
rect 18836 30640 18845 30680
rect 19651 30640 19660 30680
rect 19700 30640 21196 30680
rect 21236 30640 21245 30680
rect 7843 30639 7901 30640
rect 11011 30639 11069 30640
rect 15139 30639 15197 30640
rect 18595 30639 18653 30640
rect 7084 30556 11360 30596
rect 11491 30556 11500 30596
rect 11540 30556 11980 30596
rect 12020 30556 12029 30596
rect 12643 30556 12652 30596
rect 12692 30556 13612 30596
rect 13652 30556 15628 30596
rect 15668 30556 15677 30596
rect 19363 30556 19372 30596
rect 19412 30556 20044 30596
rect 20084 30556 20093 30596
rect 11320 30512 11360 30556
rect 14563 30512 14621 30513
rect 21424 30512 21504 30532
rect 6988 30472 9620 30512
rect 10723 30472 10732 30512
rect 10772 30472 11212 30512
rect 11252 30472 11261 30512
rect 11320 30472 14572 30512
rect 14612 30472 14621 30512
rect 16387 30472 16396 30512
rect 16436 30472 16972 30512
rect 17012 30472 17021 30512
rect 19459 30472 19468 30512
rect 19508 30472 21504 30512
rect 7747 30428 7805 30429
rect 9580 30428 9620 30472
rect 14563 30471 14621 30472
rect 21424 30452 21504 30472
rect 1228 30388 2764 30428
rect 2804 30388 6740 30428
rect 6796 30388 7756 30428
rect 7796 30388 7805 30428
rect 8803 30388 8812 30428
rect 8852 30388 9484 30428
rect 9524 30388 9533 30428
rect 9580 30388 11596 30428
rect 11636 30388 12268 30428
rect 12308 30388 12317 30428
rect 2755 30387 2813 30388
rect 0 30344 80 30364
rect 6700 30344 6740 30388
rect 7747 30387 7805 30388
rect 14659 30344 14717 30345
rect 0 30304 2572 30344
rect 2612 30304 6604 30344
rect 6644 30304 6653 30344
rect 6700 30304 14668 30344
rect 14708 30304 14717 30344
rect 0 30284 80 30304
rect 14659 30303 14717 30304
rect 5635 30260 5693 30261
rect 6499 30260 6557 30261
rect 14371 30260 14429 30261
rect 3679 30220 3688 30260
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 4056 30220 4065 30260
rect 5539 30220 5548 30260
rect 5588 30220 5644 30260
rect 5684 30220 5693 30260
rect 6414 30220 6508 30260
rect 6548 30220 6557 30260
rect 6787 30220 6796 30260
rect 6836 30220 7276 30260
rect 7316 30220 8812 30260
rect 8852 30220 8861 30260
rect 9187 30220 9196 30260
rect 9236 30220 9484 30260
rect 9524 30220 9533 30260
rect 11107 30220 11116 30260
rect 11156 30220 12652 30260
rect 12692 30220 12701 30260
rect 14371 30220 14380 30260
rect 14420 30220 16628 30260
rect 18799 30220 18808 30260
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 19176 30220 19185 30260
rect 5635 30219 5693 30220
rect 6499 30219 6557 30220
rect 14371 30219 14429 30220
rect 2083 30176 2141 30177
rect 2083 30136 2092 30176
rect 2132 30136 6700 30176
rect 6740 30136 14860 30176
rect 14900 30136 14909 30176
rect 2083 30135 2141 30136
rect 16588 30092 16628 30220
rect 21424 30176 21504 30196
rect 16771 30136 16780 30176
rect 16820 30136 21504 30176
rect 21424 30116 21504 30136
rect 19747 30092 19805 30093
rect 14371 30052 14380 30092
rect 14420 30052 14572 30092
rect 14612 30052 15916 30092
rect 15956 30052 15965 30092
rect 16588 30052 19756 30092
rect 19796 30052 19805 30092
rect 19747 30051 19805 30052
rect 0 30008 80 30028
rect 13507 30008 13565 30009
rect 0 29968 1420 30008
rect 1460 29968 1469 30008
rect 3139 29968 3148 30008
rect 3188 29968 3628 30008
rect 3668 29968 3677 30008
rect 13507 29968 13516 30008
rect 13556 29968 13708 30008
rect 13748 29968 13757 30008
rect 14179 29968 14188 30008
rect 14228 29968 20180 30008
rect 0 29948 80 29968
rect 13507 29967 13565 29968
rect 2947 29924 3005 29925
rect 6883 29924 6941 29925
rect 2862 29884 2956 29924
rect 2996 29884 6892 29924
rect 6932 29884 6941 29924
rect 7555 29884 7564 29924
rect 7604 29884 10636 29924
rect 10676 29884 11020 29924
rect 11060 29884 11069 29924
rect 12931 29884 12940 29924
rect 12980 29884 13516 29924
rect 13556 29884 14476 29924
rect 14516 29884 14525 29924
rect 2947 29883 3005 29884
rect 6883 29883 6941 29884
rect 4291 29840 4349 29841
rect 2500 29800 4300 29840
rect 4340 29800 4349 29840
rect 2500 29756 2540 29800
rect 4291 29799 4349 29800
rect 6307 29840 6365 29841
rect 12739 29840 12797 29841
rect 20140 29840 20180 29968
rect 21424 29840 21504 29860
rect 6307 29800 6316 29840
rect 6356 29800 8044 29840
rect 8084 29800 8093 29840
rect 12739 29800 12748 29840
rect 12788 29800 13036 29840
rect 13076 29800 15244 29840
rect 15284 29800 15293 29840
rect 15619 29800 15628 29840
rect 15668 29800 19372 29840
rect 19412 29800 19421 29840
rect 20140 29800 21504 29840
rect 6307 29799 6365 29800
rect 12739 29799 12797 29800
rect 21424 29780 21504 29800
rect 9859 29756 9917 29757
rect 1315 29716 1324 29756
rect 1364 29716 2540 29756
rect 2851 29716 2860 29756
rect 2900 29716 9868 29756
rect 9908 29716 9917 29756
rect 13411 29716 13420 29756
rect 13460 29716 14188 29756
rect 14228 29716 14237 29756
rect 17740 29716 18604 29756
rect 18644 29716 18653 29756
rect 9859 29715 9917 29716
rect 0 29672 80 29692
rect 4099 29672 4157 29673
rect 14179 29672 14237 29673
rect 17740 29672 17780 29716
rect 0 29632 1228 29672
rect 1268 29632 1277 29672
rect 4014 29632 4108 29672
rect 4148 29632 4157 29672
rect 5731 29632 5740 29672
rect 5780 29632 7852 29672
rect 7892 29632 7901 29672
rect 14179 29632 14188 29672
rect 14228 29632 17780 29672
rect 17827 29632 17836 29672
rect 17876 29632 18124 29672
rect 18164 29632 18173 29672
rect 0 29612 80 29632
rect 4099 29631 4157 29632
rect 14179 29631 14237 29632
rect 3427 29548 3436 29588
rect 3476 29548 12940 29588
rect 12980 29548 12989 29588
rect 13123 29548 13132 29588
rect 13172 29548 14764 29588
rect 14804 29548 14813 29588
rect 21424 29504 21504 29524
rect 4919 29464 4928 29504
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 5296 29464 5305 29504
rect 6595 29464 6604 29504
rect 6644 29464 6892 29504
rect 6932 29464 6941 29504
rect 7843 29464 7852 29504
rect 7892 29464 10060 29504
rect 10100 29464 10109 29504
rect 10915 29464 10924 29504
rect 10964 29464 13708 29504
rect 13748 29464 13757 29504
rect 14275 29464 14284 29504
rect 14324 29464 15436 29504
rect 15476 29464 15485 29504
rect 20039 29464 20048 29504
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20416 29464 20425 29504
rect 20707 29464 20716 29504
rect 20756 29464 21504 29504
rect 6604 29420 6644 29464
rect 21424 29444 21504 29464
rect 1132 29380 2572 29420
rect 2612 29380 2621 29420
rect 3052 29380 6644 29420
rect 6787 29420 6845 29421
rect 6787 29380 6796 29420
rect 6836 29380 6988 29420
rect 7028 29380 7037 29420
rect 14083 29380 14092 29420
rect 14132 29380 15532 29420
rect 15572 29380 15581 29420
rect 18211 29380 18220 29420
rect 18260 29380 19276 29420
rect 19316 29380 19325 29420
rect 0 29336 80 29356
rect 1132 29336 1172 29380
rect 0 29296 1172 29336
rect 2467 29336 2525 29337
rect 3052 29336 3092 29380
rect 6787 29379 6845 29380
rect 6691 29336 6749 29337
rect 13795 29336 13853 29337
rect 14275 29336 14333 29337
rect 14947 29336 15005 29337
rect 2467 29296 2476 29336
rect 2516 29296 3092 29336
rect 3139 29296 3148 29336
rect 3188 29296 3532 29336
rect 3572 29296 3581 29336
rect 6606 29296 6700 29336
rect 6740 29296 7276 29336
rect 7316 29296 7325 29336
rect 8995 29296 9004 29336
rect 9044 29296 9292 29336
rect 9332 29296 9341 29336
rect 11299 29296 11308 29336
rect 11348 29296 13652 29336
rect 13710 29296 13804 29336
rect 13844 29296 13853 29336
rect 14190 29296 14284 29336
rect 14324 29296 14333 29336
rect 14851 29296 14860 29336
rect 14900 29296 14956 29336
rect 14996 29296 15005 29336
rect 0 29276 80 29296
rect 2467 29295 2525 29296
rect 6691 29295 6749 29296
rect 1123 29252 1181 29253
rect 13612 29252 13652 29296
rect 13795 29295 13853 29296
rect 14275 29295 14333 29296
rect 14947 29295 15005 29296
rect 1123 29212 1132 29252
rect 1172 29212 12652 29252
rect 12692 29212 12701 29252
rect 13612 29212 14956 29252
rect 14996 29212 15005 29252
rect 17635 29212 17644 29252
rect 17684 29212 18796 29252
rect 18836 29212 18988 29252
rect 19028 29212 19037 29252
rect 1123 29211 1181 29212
rect 5347 29168 5405 29169
rect 5827 29168 5885 29169
rect 9379 29168 9437 29169
rect 9859 29168 9917 29169
rect 21424 29168 21504 29188
rect 2563 29128 2572 29168
rect 2612 29128 5356 29168
rect 5396 29128 5836 29168
rect 5876 29128 5885 29168
rect 6019 29128 6028 29168
rect 6068 29128 7852 29168
rect 7892 29128 7901 29168
rect 9294 29128 9388 29168
rect 9428 29128 9437 29168
rect 9774 29128 9868 29168
rect 9908 29128 9917 29168
rect 11395 29128 11404 29168
rect 11444 29128 11453 29168
rect 12355 29128 12364 29168
rect 12404 29128 13132 29168
rect 13172 29128 13181 29168
rect 15811 29128 15820 29168
rect 15860 29128 17932 29168
rect 17972 29128 17981 29168
rect 20707 29128 20716 29168
rect 20756 29128 21504 29168
rect 5347 29127 5405 29128
rect 5827 29127 5885 29128
rect 9379 29127 9437 29128
rect 9859 29127 9917 29128
rect 7843 29084 7901 29085
rect 11404 29084 11444 29128
rect 21424 29108 21504 29128
rect 14275 29084 14333 29085
rect 76 29044 2860 29084
rect 2900 29044 2909 29084
rect 3139 29044 3148 29084
rect 3188 29044 3436 29084
rect 3476 29044 3485 29084
rect 6124 29044 6412 29084
rect 6452 29044 6461 29084
rect 6979 29044 6988 29084
rect 7028 29044 7037 29084
rect 7747 29044 7756 29084
rect 7796 29044 7852 29084
rect 7892 29044 7901 29084
rect 76 29020 116 29044
rect 0 28960 116 29020
rect 6124 29000 6164 29044
rect 6988 29000 7028 29044
rect 7843 29043 7901 29044
rect 9292 29044 10924 29084
rect 10964 29044 10973 29084
rect 11404 29044 11788 29084
rect 11828 29044 12404 29084
rect 12451 29044 12460 29084
rect 12500 29044 13420 29084
rect 13460 29044 13469 29084
rect 13708 29044 13804 29084
rect 13844 29044 13853 29084
rect 13900 29044 14284 29084
rect 14324 29044 14333 29084
rect 9292 29000 9332 29044
rect 5731 28960 5740 29000
rect 5780 28960 6164 29000
rect 6499 28960 6508 29000
rect 6548 28960 7028 29000
rect 9252 28960 9292 29000
rect 9332 28960 9341 29000
rect 0 28940 80 28960
rect 12364 28916 12404 29044
rect 13507 29000 13565 29001
rect 13708 29000 13748 29044
rect 13900 29000 13940 29044
rect 14275 29043 14333 29044
rect 14467 29084 14525 29085
rect 14467 29044 14476 29084
rect 14516 29044 14610 29084
rect 16867 29044 16876 29084
rect 16916 29044 17548 29084
rect 17588 29044 17597 29084
rect 17731 29044 17740 29084
rect 17780 29044 18412 29084
rect 18452 29044 18461 29084
rect 14467 29043 14525 29044
rect 14947 29000 15005 29001
rect 12643 28960 12652 29000
rect 12692 28960 13516 29000
rect 13556 28960 13748 29000
rect 13860 28960 13900 29000
rect 13940 28960 13949 29000
rect 14862 28960 14956 29000
rect 14996 28960 15005 29000
rect 13507 28959 13565 28960
rect 14947 28959 15005 28960
rect 13795 28916 13853 28917
rect 14851 28916 14909 28917
rect 739 28876 748 28916
rect 788 28876 8840 28916
rect 12364 28876 13036 28916
rect 13076 28876 13085 28916
rect 13710 28876 13804 28916
rect 13844 28876 13853 28916
rect 8800 28832 8840 28876
rect 13795 28875 13853 28876
rect 14572 28876 14804 28916
rect 14572 28832 14612 28876
rect 8800 28792 14612 28832
rect 14764 28832 14804 28876
rect 14851 28876 14860 28916
rect 14900 28876 15244 28916
rect 15284 28876 15293 28916
rect 17251 28876 17260 28916
rect 17300 28876 18028 28916
rect 18068 28876 18077 28916
rect 14851 28875 14909 28876
rect 21424 28832 21504 28852
rect 14764 28792 20180 28832
rect 20227 28792 20236 28832
rect 20276 28792 21504 28832
rect 6307 28748 6365 28749
rect 14755 28748 14813 28749
rect 20140 28748 20180 28792
rect 21424 28772 21504 28792
rect 3679 28708 3688 28748
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 4056 28708 4065 28748
rect 6211 28708 6220 28748
rect 6260 28708 6316 28748
rect 6356 28708 6365 28748
rect 7075 28708 7084 28748
rect 7124 28708 7564 28748
rect 7604 28708 7613 28748
rect 9868 28708 11116 28748
rect 11156 28708 11165 28748
rect 12835 28708 12844 28748
rect 12884 28708 14572 28748
rect 14612 28708 14621 28748
rect 14755 28708 14764 28748
rect 14804 28708 14860 28748
rect 14900 28708 15724 28748
rect 15764 28708 15916 28748
rect 15956 28708 15965 28748
rect 18799 28708 18808 28748
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 19176 28708 19185 28748
rect 20140 28708 20908 28748
rect 20948 28708 20957 28748
rect 6307 28707 6365 28708
rect 0 28664 80 28684
rect 5635 28664 5693 28665
rect 9868 28664 9908 28708
rect 14755 28707 14813 28708
rect 0 28624 4684 28664
rect 4724 28624 4733 28664
rect 5635 28624 5644 28664
rect 5684 28624 9908 28664
rect 9955 28664 10013 28665
rect 9955 28624 9964 28664
rect 10004 28624 13516 28664
rect 13556 28624 13565 28664
rect 13699 28624 13708 28664
rect 13748 28624 14375 28664
rect 14415 28624 14424 28664
rect 14467 28624 14476 28664
rect 14516 28624 15148 28664
rect 15188 28624 15197 28664
rect 17923 28624 17932 28664
rect 17972 28624 18508 28664
rect 18548 28624 18557 28664
rect 0 28604 80 28624
rect 5635 28623 5693 28624
rect 9955 28623 10013 28624
rect 6403 28580 6461 28581
rect 5731 28540 5740 28580
rect 5780 28540 6124 28580
rect 6164 28540 6173 28580
rect 6403 28540 6412 28580
rect 6452 28540 21100 28580
rect 21140 28540 21149 28580
rect 6403 28539 6461 28540
rect 3139 28496 3197 28497
rect 21424 28496 21504 28516
rect 3054 28456 3148 28496
rect 3188 28456 3197 28496
rect 4003 28456 4012 28496
rect 4052 28456 4492 28496
rect 4532 28456 4541 28496
rect 6019 28456 6028 28496
rect 6068 28456 7372 28496
rect 7412 28456 7421 28496
rect 11011 28456 11020 28496
rect 11060 28456 21504 28496
rect 3139 28455 3197 28456
rect 21424 28436 21504 28456
rect 5827 28412 5885 28413
rect 11491 28412 11549 28413
rect 5742 28372 5836 28412
rect 5876 28372 5885 28412
rect 6595 28372 6604 28412
rect 6644 28372 7756 28412
rect 7796 28372 7805 28412
rect 11491 28372 11500 28412
rect 11540 28372 13708 28412
rect 13748 28372 13757 28412
rect 14083 28372 14092 28412
rect 14132 28372 14668 28412
rect 14708 28372 14717 28412
rect 5827 28371 5885 28372
rect 11491 28371 11549 28372
rect 0 28328 80 28348
rect 7363 28328 7421 28329
rect 12739 28328 12797 28329
rect 0 28288 2540 28328
rect 2659 28288 2668 28328
rect 2708 28288 3148 28328
rect 3188 28288 3197 28328
rect 4099 28288 4108 28328
rect 4148 28288 5644 28328
rect 5684 28288 6412 28328
rect 6452 28288 6461 28328
rect 6691 28288 6700 28328
rect 6740 28288 7372 28328
rect 7412 28288 7421 28328
rect 7843 28288 7852 28328
rect 7892 28288 10348 28328
rect 10388 28288 10397 28328
rect 12654 28288 12748 28328
rect 12788 28288 12797 28328
rect 0 28268 80 28288
rect 2500 28160 2540 28288
rect 7363 28287 7421 28288
rect 12739 28287 12797 28288
rect 13708 28244 13748 28372
rect 14851 28328 14909 28329
rect 15619 28328 15677 28329
rect 16675 28328 16733 28329
rect 19267 28328 19325 28329
rect 14851 28288 14860 28328
rect 14900 28288 15052 28328
rect 15092 28288 15101 28328
rect 15619 28288 15628 28328
rect 15668 28288 16684 28328
rect 16724 28288 16780 28328
rect 16820 28288 16829 28328
rect 17827 28288 17836 28328
rect 17876 28288 18604 28328
rect 18644 28288 18653 28328
rect 18979 28288 18988 28328
rect 19028 28288 19276 28328
rect 19316 28288 19325 28328
rect 20035 28288 20044 28328
rect 20084 28288 20524 28328
rect 20564 28288 20573 28328
rect 14851 28287 14909 28288
rect 15619 28287 15677 28288
rect 16675 28287 16733 28288
rect 19267 28287 19325 28288
rect 16291 28244 16349 28245
rect 3907 28204 3916 28244
rect 3956 28204 5548 28244
rect 5588 28204 5597 28244
rect 5740 28204 8812 28244
rect 8852 28204 8861 28244
rect 13708 28204 16244 28244
rect 5740 28160 5780 28204
rect 6787 28160 6845 28161
rect 14755 28160 14813 28161
rect 16204 28160 16244 28204
rect 16291 28204 16300 28244
rect 16340 28204 19564 28244
rect 19604 28204 19613 28244
rect 16291 28203 16349 28204
rect 21424 28160 21504 28180
rect 2500 28120 5780 28160
rect 5827 28120 5836 28160
rect 5876 28120 6028 28160
rect 6068 28120 6077 28160
rect 6403 28120 6412 28160
rect 6452 28120 6796 28160
rect 6836 28120 6845 28160
rect 12643 28120 12652 28160
rect 12692 28120 13708 28160
rect 13748 28120 13757 28160
rect 14371 28120 14380 28160
rect 14420 28120 14764 28160
rect 14804 28120 14813 28160
rect 14947 28120 14956 28160
rect 14996 28120 15572 28160
rect 16204 28120 16396 28160
rect 16436 28120 16445 28160
rect 16579 28120 16588 28160
rect 16628 28120 21504 28160
rect 6787 28119 6845 28120
rect 14755 28119 14813 28120
rect 5731 28076 5789 28077
rect 6499 28076 6557 28077
rect 15532 28076 15572 28120
rect 21424 28100 21504 28120
rect 4675 28036 4684 28076
rect 4724 28036 5396 28076
rect 0 27992 80 28012
rect 2947 27992 3005 27993
rect 5356 27992 5396 28036
rect 5731 28036 5740 28076
rect 5780 28036 5932 28076
rect 5972 28036 5981 28076
rect 6414 28036 6508 28076
rect 6548 28036 6557 28076
rect 5731 28035 5789 28036
rect 6499 28035 6557 28036
rect 6604 28036 11500 28076
rect 11540 28036 15436 28076
rect 15476 28036 15485 28076
rect 15532 28036 17932 28076
rect 17972 28036 17981 28076
rect 6604 27992 6644 28036
rect 7363 27992 7421 27993
rect 0 27952 2324 27992
rect 2862 27952 2956 27992
rect 2996 27952 3005 27992
rect 4919 27952 4928 27992
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 5296 27952 5305 27992
rect 5356 27952 6644 27992
rect 7267 27952 7276 27992
rect 7316 27952 7372 27992
rect 7412 27952 7421 27992
rect 0 27932 80 27952
rect 2284 27824 2324 27952
rect 2947 27951 3005 27952
rect 7363 27951 7421 27952
rect 7747 27992 7805 27993
rect 19459 27992 19517 27993
rect 7747 27952 7756 27992
rect 7796 27952 13132 27992
rect 13172 27952 13181 27992
rect 13507 27952 13516 27992
rect 13556 27952 15916 27992
rect 15956 27952 19084 27992
rect 19124 27952 19468 27992
rect 19508 27952 19517 27992
rect 20039 27952 20048 27992
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20416 27952 20425 27992
rect 7747 27951 7805 27952
rect 19459 27951 19517 27952
rect 12259 27908 12317 27909
rect 12547 27908 12605 27909
rect 14371 27908 14429 27909
rect 2371 27868 2380 27908
rect 2420 27868 7756 27908
rect 7796 27868 7805 27908
rect 11395 27868 11404 27908
rect 11444 27868 12076 27908
rect 12116 27868 12125 27908
rect 12259 27868 12268 27908
rect 12308 27868 12402 27908
rect 12547 27868 12556 27908
rect 12596 27868 12690 27908
rect 12844 27868 13460 27908
rect 12259 27867 12317 27868
rect 12547 27867 12605 27868
rect 12844 27824 12884 27868
rect 13420 27824 13460 27868
rect 14371 27868 14380 27908
rect 14420 27868 17836 27908
rect 17876 27868 17885 27908
rect 14371 27867 14429 27868
rect 21424 27824 21504 27844
rect 2284 27784 12884 27824
rect 12931 27784 12940 27824
rect 12980 27784 13324 27824
rect 13364 27784 13373 27824
rect 13420 27784 16204 27824
rect 16244 27784 16628 27824
rect 19267 27784 19276 27824
rect 19316 27784 21504 27824
rect 4579 27740 4637 27741
rect 8803 27740 8861 27741
rect 13219 27740 13277 27741
rect 14851 27740 14909 27741
rect 16291 27740 16349 27741
rect 1219 27700 1228 27740
rect 1268 27700 3340 27740
rect 3380 27700 3389 27740
rect 4494 27700 4588 27740
rect 4628 27700 4637 27740
rect 5347 27700 5356 27740
rect 5396 27700 5548 27740
rect 5588 27700 5972 27740
rect 6019 27700 6028 27740
rect 6068 27700 7372 27740
rect 7412 27700 7421 27740
rect 8803 27700 8812 27740
rect 8852 27700 10924 27740
rect 10964 27700 10973 27740
rect 13134 27700 13228 27740
rect 13268 27700 13277 27740
rect 4579 27699 4637 27700
rect 0 27656 80 27676
rect 2467 27656 2525 27657
rect 5635 27656 5693 27657
rect 0 27616 2476 27656
rect 2516 27616 2525 27656
rect 2947 27616 2956 27656
rect 2996 27616 3244 27656
rect 3284 27616 3293 27656
rect 4867 27616 4876 27656
rect 4916 27616 5644 27656
rect 5684 27616 5693 27656
rect 5932 27656 5972 27700
rect 8803 27699 8861 27700
rect 13219 27699 13277 27700
rect 13324 27700 14860 27740
rect 14900 27700 14909 27740
rect 15811 27700 15820 27740
rect 15860 27700 16300 27740
rect 16340 27700 16349 27740
rect 9763 27656 9821 27657
rect 13324 27656 13364 27700
rect 14851 27699 14909 27700
rect 16291 27699 16349 27700
rect 14467 27656 14525 27657
rect 16588 27656 16628 27784
rect 21424 27764 21504 27784
rect 17923 27700 17932 27740
rect 17972 27700 18796 27740
rect 18836 27700 18845 27740
rect 5932 27616 6124 27656
rect 6164 27616 6173 27656
rect 6979 27616 6988 27656
rect 7028 27616 8044 27656
rect 8084 27616 8093 27656
rect 8707 27616 8716 27656
rect 8756 27616 9484 27656
rect 9524 27616 9533 27656
rect 9678 27616 9772 27656
rect 9812 27616 9821 27656
rect 11587 27616 11596 27656
rect 11636 27616 11980 27656
rect 12020 27616 12029 27656
rect 12259 27616 12268 27656
rect 12308 27616 12844 27656
rect 12884 27616 12893 27656
rect 13315 27616 13324 27656
rect 13364 27616 13373 27656
rect 14275 27616 14284 27656
rect 14324 27616 14476 27656
rect 14516 27616 14525 27656
rect 14851 27616 14860 27656
rect 14900 27616 15436 27656
rect 15476 27616 15485 27656
rect 16579 27616 16588 27656
rect 16628 27616 16637 27656
rect 18019 27616 18028 27656
rect 18068 27616 20044 27656
rect 20084 27616 20093 27656
rect 0 27596 80 27616
rect 2467 27615 2525 27616
rect 5635 27615 5693 27616
rect 9763 27615 9821 27616
rect 14467 27615 14525 27616
rect 15235 27572 15293 27573
rect 7459 27532 7468 27572
rect 7508 27532 8524 27572
rect 8564 27532 8573 27572
rect 9667 27532 9676 27572
rect 9716 27532 15244 27572
rect 15284 27532 15293 27572
rect 15235 27531 15293 27532
rect 16579 27572 16637 27573
rect 16579 27532 16588 27572
rect 16628 27532 16780 27572
rect 16820 27532 17068 27572
rect 17108 27532 17117 27572
rect 16579 27531 16637 27532
rect 7555 27488 7613 27489
rect 10243 27488 10301 27489
rect 3907 27448 3916 27488
rect 3956 27448 7316 27488
rect 4195 27404 4253 27405
rect 7171 27404 7229 27405
rect 3619 27364 3628 27404
rect 3668 27364 3708 27404
rect 4195 27364 4204 27404
rect 4244 27364 5548 27404
rect 5588 27364 5597 27404
rect 7086 27364 7180 27404
rect 7220 27364 7229 27404
rect 7276 27404 7316 27448
rect 7555 27448 7564 27488
rect 7604 27448 9868 27488
rect 9908 27448 9917 27488
rect 10156 27448 10252 27488
rect 10292 27448 10301 27488
rect 7555 27447 7613 27448
rect 8995 27404 9053 27405
rect 10156 27404 10196 27448
rect 10243 27447 10301 27448
rect 11491 27488 11549 27489
rect 15811 27488 15869 27489
rect 21424 27488 21504 27508
rect 11491 27448 11500 27488
rect 11540 27448 11634 27488
rect 11813 27448 11822 27488
rect 11862 27448 12172 27488
rect 12212 27448 12596 27488
rect 12643 27448 12652 27488
rect 12692 27448 13228 27488
rect 13268 27448 15820 27488
rect 15860 27448 15869 27488
rect 17347 27448 17356 27488
rect 17396 27448 18124 27488
rect 18164 27448 18173 27488
rect 20899 27448 20908 27488
rect 20948 27448 21504 27488
rect 11491 27447 11549 27448
rect 12556 27404 12596 27448
rect 15811 27447 15869 27448
rect 21424 27428 21504 27448
rect 15907 27404 15965 27405
rect 7276 27364 9004 27404
rect 9044 27364 10196 27404
rect 10243 27364 10252 27404
rect 10292 27364 12364 27404
rect 12404 27364 12413 27404
rect 12547 27364 12556 27404
rect 12596 27364 12605 27404
rect 13507 27364 13516 27404
rect 13556 27364 15916 27404
rect 15956 27364 15965 27404
rect 0 27320 80 27340
rect 1123 27320 1181 27321
rect 3628 27320 3668 27364
rect 4195 27363 4253 27364
rect 7171 27363 7229 27364
rect 8995 27363 9053 27364
rect 15907 27363 15965 27364
rect 12547 27320 12605 27321
rect 0 27280 1132 27320
rect 1172 27280 1181 27320
rect 2947 27280 2956 27320
rect 2996 27280 4244 27320
rect 5731 27280 5740 27320
rect 5780 27280 11828 27320
rect 11875 27280 11884 27320
rect 11924 27280 12556 27320
rect 12596 27280 12605 27320
rect 13699 27280 13708 27320
rect 13748 27280 14956 27320
rect 14996 27280 15005 27320
rect 0 27260 80 27280
rect 1123 27279 1181 27280
rect 2851 27236 2909 27237
rect 4204 27236 4244 27280
rect 2755 27196 2764 27236
rect 2804 27196 2860 27236
rect 2900 27196 2909 27236
rect 3679 27196 3688 27236
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 4056 27196 4065 27236
rect 4204 27196 9676 27236
rect 9716 27196 9725 27236
rect 2851 27195 2909 27196
rect 11491 27152 11549 27153
rect 3331 27112 3340 27152
rect 3380 27112 11500 27152
rect 11540 27112 11549 27152
rect 11491 27111 11549 27112
rect 643 27068 701 27069
rect 11395 27068 11453 27069
rect 11788 27068 11828 27280
rect 12547 27279 12605 27280
rect 15139 27236 15197 27237
rect 14179 27196 14188 27236
rect 14228 27196 15148 27236
rect 15188 27196 15197 27236
rect 18799 27196 18808 27236
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 19176 27196 19185 27236
rect 15139 27195 15197 27196
rect 15043 27152 15101 27153
rect 21424 27152 21504 27172
rect 13315 27112 13324 27152
rect 13364 27112 15052 27152
rect 15092 27112 15148 27152
rect 15188 27112 15197 27152
rect 21091 27112 21100 27152
rect 21140 27112 21504 27152
rect 15043 27111 15101 27112
rect 21424 27092 21504 27112
rect 12355 27068 12413 27069
rect 14275 27068 14333 27069
rect 643 27028 652 27068
rect 692 27028 844 27068
rect 884 27028 893 27068
rect 3427 27028 3436 27068
rect 3476 27028 3628 27068
rect 3668 27028 3677 27068
rect 6211 27028 6220 27068
rect 6260 27028 6892 27068
rect 6932 27028 6941 27068
rect 11395 27028 11404 27068
rect 11444 27028 11692 27068
rect 11732 27028 11741 27068
rect 11788 27028 12364 27068
rect 12404 27028 14284 27068
rect 14324 27028 14333 27068
rect 14755 27028 14764 27068
rect 14804 27028 14956 27068
rect 14996 27028 15005 27068
rect 643 27027 701 27028
rect 11395 27027 11453 27028
rect 12355 27027 12413 27028
rect 14275 27027 14333 27028
rect 0 26984 80 27004
rect 3139 26984 3197 26985
rect 6499 26984 6557 26985
rect 0 26944 1652 26984
rect 0 26924 80 26944
rect 1612 26900 1652 26944
rect 3139 26944 3148 26984
rect 3188 26944 3340 26984
rect 3380 26944 3389 26984
rect 6499 26944 6508 26984
rect 6548 26944 6604 26984
rect 6644 26944 6653 26984
rect 7267 26944 7276 26984
rect 7316 26944 7468 26984
rect 7508 26944 7517 26984
rect 8515 26944 8524 26984
rect 8564 26944 13172 26984
rect 14563 26944 14572 26984
rect 14612 26944 15724 26984
rect 15764 26944 15773 26984
rect 16963 26944 16972 26984
rect 17012 26944 17260 26984
rect 17300 26944 17309 26984
rect 3139 26943 3197 26944
rect 6499 26943 6557 26944
rect 6211 26900 6269 26901
rect 1612 26860 6220 26900
rect 6260 26860 6269 26900
rect 6211 26859 6269 26860
rect 6403 26900 6461 26901
rect 9667 26900 9725 26901
rect 13132 26900 13172 26944
rect 14851 26900 14909 26901
rect 17827 26900 17885 26901
rect 6403 26860 6412 26900
rect 6452 26860 6892 26900
rect 6932 26860 6941 26900
rect 8995 26860 9004 26900
rect 9044 26860 9676 26900
rect 9716 26860 9725 26900
rect 6403 26859 6461 26860
rect 9667 26859 9725 26860
rect 11320 26860 11980 26900
rect 12020 26860 12029 26900
rect 13132 26860 14860 26900
rect 14900 26860 14909 26900
rect 17731 26860 17740 26900
rect 17780 26860 17836 26900
rect 17876 26860 17885 26900
rect 2851 26816 2909 26817
rect 1795 26776 1804 26816
rect 1844 26776 2476 26816
rect 2516 26776 2525 26816
rect 2766 26776 2860 26816
rect 2900 26776 2909 26816
rect 2851 26775 2909 26776
rect 3235 26816 3293 26817
rect 4483 26816 4541 26817
rect 11320 26816 11360 26860
rect 14851 26859 14909 26860
rect 17827 26859 17885 26860
rect 12547 26816 12605 26817
rect 15811 26816 15869 26817
rect 17059 26816 17117 26817
rect 21424 26816 21504 26836
rect 3235 26776 3244 26816
rect 3284 26776 3436 26816
rect 3476 26776 3485 26816
rect 4195 26776 4204 26816
rect 4244 26776 4492 26816
rect 4532 26776 4541 26816
rect 6307 26776 6316 26816
rect 6356 26776 6700 26816
rect 6740 26776 6749 26816
rect 6979 26776 6988 26816
rect 7028 26776 7468 26816
rect 7508 26776 7517 26816
rect 9475 26776 9484 26816
rect 9524 26776 10252 26816
rect 10292 26776 11360 26816
rect 12067 26776 12076 26816
rect 12116 26776 12268 26816
rect 12308 26776 12317 26816
rect 12462 26776 12556 26816
rect 12596 26776 12605 26816
rect 15235 26776 15244 26816
rect 15284 26776 15820 26816
rect 15860 26776 15869 26816
rect 16387 26776 16396 26816
rect 16436 26776 16780 26816
rect 16820 26776 16829 26816
rect 17059 26776 17068 26816
rect 17108 26776 21504 26816
rect 3235 26775 3293 26776
rect 4483 26775 4541 26776
rect 12547 26775 12605 26776
rect 15811 26775 15869 26776
rect 17059 26775 17117 26776
rect 21424 26756 21504 26776
rect 19267 26732 19325 26733
rect 1996 26692 19276 26732
rect 19316 26692 19325 26732
rect 0 26648 80 26668
rect 1996 26648 2036 26692
rect 19267 26691 19325 26692
rect 6307 26648 6365 26649
rect 11299 26648 11357 26649
rect 16675 26648 16733 26649
rect 0 26608 2036 26648
rect 4099 26608 4108 26648
rect 4148 26608 6316 26648
rect 6356 26608 6365 26648
rect 6787 26608 6796 26648
rect 6836 26608 7180 26648
rect 7220 26608 7229 26648
rect 7555 26608 7564 26648
rect 7604 26608 8564 26648
rect 8611 26608 8620 26648
rect 8660 26608 10252 26648
rect 10292 26608 10301 26648
rect 11299 26608 11308 26648
rect 11348 26608 11884 26648
rect 11924 26608 14572 26648
rect 14612 26608 14860 26648
rect 14900 26608 14909 26648
rect 16675 26608 16684 26648
rect 16724 26608 16972 26648
rect 17012 26608 17021 26648
rect 18307 26608 18316 26648
rect 18356 26608 18365 26648
rect 0 26588 80 26608
rect 6307 26607 6365 26608
rect 6883 26564 6941 26565
rect 8524 26564 8564 26608
rect 11299 26607 11357 26608
rect 16675 26607 16733 26608
rect 11491 26564 11549 26565
rect 1315 26524 1324 26564
rect 1364 26524 5740 26564
rect 5780 26524 5789 26564
rect 6307 26524 6316 26564
rect 6356 26524 6604 26564
rect 6644 26524 6653 26564
rect 6883 26524 6892 26564
rect 6932 26524 7084 26564
rect 7124 26524 7133 26564
rect 7651 26524 7660 26564
rect 7700 26524 8044 26564
rect 8084 26524 8093 26564
rect 8515 26524 8524 26564
rect 8564 26524 8573 26564
rect 11491 26524 11500 26564
rect 11540 26524 12844 26564
rect 12884 26524 12893 26564
rect 6883 26523 6941 26524
rect 11491 26523 11549 26524
rect 3139 26480 3197 26481
rect 5635 26480 5693 26481
rect 10339 26480 10397 26481
rect 15619 26480 15677 26481
rect 16099 26480 16157 26481
rect 16579 26480 16637 26481
rect 2467 26440 2476 26480
rect 2516 26440 2900 26480
rect 3054 26440 3148 26480
rect 3188 26440 3197 26480
rect 2860 26396 2900 26440
rect 3139 26439 3197 26440
rect 3724 26440 4492 26480
rect 4532 26440 4541 26480
rect 4919 26440 4928 26480
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 5296 26440 5305 26480
rect 5635 26440 5644 26480
rect 5684 26440 9292 26480
rect 9332 26440 9341 26480
rect 10254 26440 10348 26480
rect 10388 26440 10397 26480
rect 10627 26440 10636 26480
rect 10676 26440 11020 26480
rect 11060 26440 11069 26480
rect 14467 26440 14476 26480
rect 14516 26440 15052 26480
rect 15092 26440 15101 26480
rect 15619 26440 15628 26480
rect 15668 26440 15820 26480
rect 15860 26440 15869 26480
rect 16014 26440 16108 26480
rect 16148 26440 16157 26480
rect 16494 26440 16588 26480
rect 16628 26440 16637 26480
rect 18316 26480 18356 26608
rect 20611 26480 20669 26481
rect 21424 26480 21504 26500
rect 18316 26440 19276 26480
rect 19316 26440 19325 26480
rect 20039 26440 20048 26480
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20416 26440 20425 26480
rect 20611 26440 20620 26480
rect 20660 26440 21504 26480
rect 2947 26396 3005 26397
rect 3331 26396 3389 26397
rect 3724 26396 3764 26440
rect 5635 26439 5693 26440
rect 10339 26439 10397 26440
rect 15619 26439 15677 26440
rect 16099 26439 16157 26440
rect 16579 26439 16637 26440
rect 20611 26439 20669 26440
rect 21424 26420 21504 26440
rect 6787 26396 6845 26397
rect 10627 26396 10685 26397
rect 2860 26356 2956 26396
rect 2996 26356 3340 26396
rect 3380 26356 3764 26396
rect 6499 26356 6508 26396
rect 6548 26356 6796 26396
rect 6836 26356 6845 26396
rect 7843 26356 7852 26396
rect 7892 26356 10636 26396
rect 10676 26356 10685 26396
rect 2947 26355 3005 26356
rect 3331 26355 3389 26356
rect 6787 26355 6845 26356
rect 10627 26355 10685 26356
rect 14755 26396 14813 26397
rect 14755 26356 14764 26396
rect 14804 26356 17740 26396
rect 17780 26356 18508 26396
rect 18548 26356 18557 26396
rect 14755 26355 14813 26356
rect 0 26312 80 26332
rect 1699 26312 1757 26313
rect 7939 26312 7997 26313
rect 20707 26312 20765 26313
rect 0 26272 1708 26312
rect 1748 26272 1757 26312
rect 1987 26272 1996 26312
rect 2036 26272 2668 26312
rect 2708 26272 2717 26312
rect 7939 26272 7948 26312
rect 7988 26272 16492 26312
rect 16532 26272 16541 26312
rect 17923 26272 17932 26312
rect 17972 26272 18700 26312
rect 18740 26272 18749 26312
rect 20707 26272 20716 26312
rect 20756 26272 21428 26312
rect 0 26252 80 26272
rect 1699 26271 1757 26272
rect 7939 26271 7997 26272
rect 20707 26271 20765 26272
rect 3235 26188 3244 26228
rect 3284 26188 7372 26228
rect 7412 26188 7948 26228
rect 7988 26188 7997 26228
rect 8323 26188 8332 26228
rect 8372 26188 8620 26228
rect 8660 26188 8669 26228
rect 9283 26188 9292 26228
rect 9332 26188 9772 26228
rect 9812 26188 10156 26228
rect 10196 26188 10205 26228
rect 10435 26188 10444 26228
rect 10484 26188 20180 26228
rect 2371 26144 2429 26145
rect 3427 26144 3485 26145
rect 4675 26144 4733 26145
rect 10627 26144 10685 26145
rect 12259 26144 12317 26145
rect 14947 26144 15005 26145
rect 1219 26104 1228 26144
rect 1268 26104 2380 26144
rect 2420 26104 2429 26144
rect 3043 26104 3052 26144
rect 3092 26104 3436 26144
rect 3476 26104 3485 26144
rect 3811 26104 3820 26144
rect 3860 26104 4300 26144
rect 4340 26104 4349 26144
rect 4590 26104 4684 26144
rect 4724 26104 4733 26144
rect 6019 26104 6028 26144
rect 6068 26104 6412 26144
rect 6452 26104 6461 26144
rect 7075 26104 7084 26144
rect 7124 26104 7276 26144
rect 7316 26104 7325 26144
rect 7651 26104 7660 26144
rect 7700 26104 8524 26144
rect 8564 26104 8812 26144
rect 8852 26104 9580 26144
rect 9620 26104 9629 26144
rect 9955 26104 9964 26144
rect 10004 26104 10348 26144
rect 10388 26104 10397 26144
rect 10542 26104 10636 26144
rect 10676 26104 10685 26144
rect 12163 26104 12172 26144
rect 12212 26104 12268 26144
rect 12308 26104 12317 26144
rect 13123 26104 13132 26144
rect 13172 26104 13612 26144
rect 13652 26104 13661 26144
rect 14851 26104 14860 26144
rect 14900 26104 14956 26144
rect 14996 26104 15005 26144
rect 16195 26104 16204 26144
rect 16244 26104 16876 26144
rect 16916 26104 16925 26144
rect 17347 26104 17356 26144
rect 17396 26104 18316 26144
rect 18356 26104 18365 26144
rect 18499 26104 18508 26144
rect 18548 26104 18796 26144
rect 18836 26104 18845 26144
rect 2371 26103 2429 26104
rect 3427 26103 3485 26104
rect 3820 26060 3860 26104
rect 4675 26103 4733 26104
rect 6412 26060 6452 26104
rect 10627 26103 10685 26104
rect 12259 26103 12317 26104
rect 14947 26103 15005 26104
rect 7747 26060 7805 26061
rect 16483 26060 16541 26061
rect 2947 26020 2956 26060
rect 2996 26020 3860 26060
rect 6115 26020 6124 26060
rect 6164 26020 6356 26060
rect 6412 26020 7468 26060
rect 7508 26020 7517 26060
rect 7747 26020 7756 26060
rect 7796 26020 7852 26060
rect 7892 26020 7901 26060
rect 9187 26020 9196 26060
rect 9236 26020 11500 26060
rect 11540 26020 11549 26060
rect 15331 26020 15340 26060
rect 15380 26020 16492 26060
rect 16532 26020 16541 26060
rect 0 25976 80 25996
rect 4483 25976 4541 25977
rect 0 25936 4492 25976
rect 4532 25936 4541 25976
rect 0 25916 80 25936
rect 4483 25935 4541 25936
rect 6316 25892 6356 26020
rect 7747 26019 7805 26020
rect 16483 26019 16541 26020
rect 6403 25976 6461 25977
rect 16195 25976 16253 25977
rect 6403 25936 6412 25976
rect 6452 25936 15436 25976
rect 15476 25936 15485 25976
rect 16110 25936 16204 25976
rect 16244 25936 16253 25976
rect 16387 25936 16396 25976
rect 16436 25936 17740 25976
rect 17780 25936 17789 25976
rect 6403 25935 6461 25936
rect 16195 25935 16253 25936
rect 5923 25852 5932 25892
rect 5972 25852 6124 25892
rect 6164 25852 6173 25892
rect 6316 25852 6604 25892
rect 6644 25852 6653 25892
rect 18691 25852 18700 25892
rect 18740 25852 19276 25892
rect 19316 25852 19325 25892
rect 8611 25808 8669 25809
rect 8995 25808 9053 25809
rect 3523 25768 3532 25808
rect 3572 25768 5780 25808
rect 5827 25768 5836 25808
rect 5876 25768 6316 25808
rect 6356 25768 6365 25808
rect 6499 25768 6508 25808
rect 6548 25768 6892 25808
rect 6932 25768 6941 25808
rect 7468 25768 8620 25808
rect 8660 25768 8716 25808
rect 8756 25768 8765 25808
rect 8910 25768 9004 25808
rect 9044 25768 9053 25808
rect 20140 25808 20180 26188
rect 21388 26164 21428 26272
rect 21388 26104 21504 26164
rect 21424 26084 21504 26104
rect 21424 25808 21504 25828
rect 20140 25768 21504 25808
rect 5740 25724 5780 25768
rect 7468 25724 7508 25768
rect 8611 25767 8669 25768
rect 8995 25767 9053 25768
rect 21424 25748 21504 25768
rect 931 25684 940 25724
rect 980 25684 3244 25724
rect 3284 25684 3293 25724
rect 3679 25684 3688 25724
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 4056 25684 4065 25724
rect 5740 25684 7508 25724
rect 7555 25684 7564 25724
rect 7604 25684 8236 25724
rect 8276 25684 8285 25724
rect 9859 25684 9868 25724
rect 9908 25684 10156 25724
rect 10196 25684 15628 25724
rect 15668 25684 16684 25724
rect 16724 25684 16733 25724
rect 18799 25684 18808 25724
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 19176 25684 19185 25724
rect 0 25640 80 25660
rect 17827 25640 17885 25641
rect 0 25600 17836 25640
rect 17876 25600 18604 25640
rect 18644 25600 18653 25640
rect 0 25580 80 25600
rect 17827 25599 17885 25600
rect 16291 25556 16349 25557
rect 2371 25516 2380 25556
rect 2420 25516 2860 25556
rect 2900 25516 2909 25556
rect 5548 25516 7124 25556
rect 16099 25516 16108 25556
rect 16148 25516 16300 25556
rect 16340 25516 16349 25556
rect 3427 25472 3485 25473
rect 2467 25432 2476 25472
rect 2516 25432 3052 25472
rect 3092 25432 3101 25472
rect 3427 25432 3436 25472
rect 3476 25432 4300 25472
rect 4340 25432 4349 25472
rect 3427 25431 3485 25432
rect 2947 25388 3005 25389
rect 1699 25348 1708 25388
rect 1748 25348 2540 25388
rect 0 25304 80 25324
rect 1315 25304 1373 25305
rect 0 25264 556 25304
rect 596 25264 605 25304
rect 1219 25264 1228 25304
rect 1268 25264 1324 25304
rect 1364 25264 1373 25304
rect 2500 25304 2540 25348
rect 2947 25348 2956 25388
rect 2996 25348 5452 25388
rect 5492 25348 5501 25388
rect 2947 25347 3005 25348
rect 4387 25304 4445 25305
rect 2500 25264 4340 25304
rect 0 25244 80 25264
rect 1315 25263 1373 25264
rect 1324 25136 1364 25263
rect 4300 25220 4340 25264
rect 4387 25264 4396 25304
rect 4436 25264 4492 25304
rect 4532 25264 4541 25304
rect 4387 25263 4445 25264
rect 5548 25220 5588 25516
rect 7084 25472 7124 25516
rect 16291 25515 16349 25516
rect 21424 25472 21504 25492
rect 6115 25432 6124 25472
rect 6164 25432 6173 25472
rect 7075 25432 7084 25472
rect 7124 25432 11020 25472
rect 11060 25432 11069 25472
rect 16771 25432 16780 25472
rect 16820 25432 21504 25472
rect 6124 25304 6164 25432
rect 21424 25412 21504 25432
rect 6403 25388 6461 25389
rect 7939 25388 7997 25389
rect 6403 25348 6412 25388
rect 6452 25348 7948 25388
rect 7988 25348 7997 25388
rect 6403 25347 6461 25348
rect 7939 25347 7997 25348
rect 8515 25388 8573 25389
rect 8515 25348 8524 25388
rect 8564 25348 13036 25388
rect 13076 25348 13085 25388
rect 16099 25348 16108 25388
rect 16148 25348 18700 25388
rect 18740 25348 18749 25388
rect 8515 25347 8573 25348
rect 12643 25304 12701 25305
rect 5731 25264 5740 25304
rect 5780 25264 8332 25304
rect 8372 25264 9196 25304
rect 9236 25264 9245 25304
rect 9763 25264 9772 25304
rect 9812 25264 10156 25304
rect 10196 25264 10205 25304
rect 12558 25264 12652 25304
rect 12692 25264 12701 25304
rect 13123 25264 13132 25304
rect 13172 25264 13900 25304
rect 13940 25264 13949 25304
rect 15139 25264 15148 25304
rect 15188 25264 16012 25304
rect 16052 25264 16061 25304
rect 16291 25264 16300 25304
rect 16340 25264 16492 25304
rect 16532 25264 16541 25304
rect 16963 25264 16972 25304
rect 17012 25264 18316 25304
rect 18356 25264 18365 25304
rect 12643 25263 12701 25264
rect 2467 25180 2476 25220
rect 2516 25180 2956 25220
rect 2996 25180 3005 25220
rect 4300 25180 5588 25220
rect 5635 25220 5693 25221
rect 5827 25220 5885 25221
rect 8227 25220 8285 25221
rect 8515 25220 8573 25221
rect 5635 25180 5644 25220
rect 5684 25180 5778 25220
rect 5827 25180 5836 25220
rect 5876 25180 8236 25220
rect 8276 25180 8285 25220
rect 8419 25180 8428 25220
rect 8468 25180 8524 25220
rect 8564 25180 8573 25220
rect 8707 25180 8716 25220
rect 8756 25180 9388 25220
rect 9428 25180 9437 25220
rect 15235 25180 15244 25220
rect 15284 25180 15532 25220
rect 15572 25180 15581 25220
rect 16579 25180 16588 25220
rect 16628 25180 18124 25220
rect 18164 25180 18173 25220
rect 5635 25179 5693 25180
rect 5827 25179 5885 25180
rect 8227 25179 8285 25180
rect 8515 25179 8573 25180
rect 6499 25136 6557 25137
rect 21424 25136 21504 25156
rect 1324 25096 6316 25136
rect 6356 25096 6365 25136
rect 6499 25096 6508 25136
rect 6548 25096 6700 25136
rect 6740 25096 6749 25136
rect 6883 25096 6892 25136
rect 6932 25096 21504 25136
rect 6499 25095 6557 25096
rect 21424 25076 21504 25096
rect 12259 25052 12317 25053
rect 1411 25012 1420 25052
rect 1460 25012 3532 25052
rect 3572 25012 3581 25052
rect 4780 25012 5932 25052
rect 5972 25012 5981 25052
rect 8515 25012 8524 25052
rect 8564 25012 9292 25052
rect 9332 25012 9341 25052
rect 11683 25012 11692 25052
rect 11732 25012 12268 25052
rect 12308 25012 12317 25052
rect 0 24968 80 24988
rect 4780 24968 4820 25012
rect 12259 25011 12317 25012
rect 6403 24968 6461 24969
rect 14467 24968 14525 24969
rect 16195 24968 16253 24969
rect 0 24928 2540 24968
rect 3427 24928 3436 24968
rect 3476 24928 4820 24968
rect 4919 24928 4928 24968
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 5296 24928 5305 24968
rect 6115 24928 6124 24968
rect 6164 24928 6412 24968
rect 6452 24928 6461 24968
rect 7363 24928 7372 24968
rect 7412 24928 8908 24968
rect 8948 24928 9484 24968
rect 9524 24928 9533 24968
rect 11875 24928 11884 24968
rect 11924 24928 12268 24968
rect 12308 24928 12317 24968
rect 14275 24928 14284 24968
rect 14324 24928 14476 24968
rect 14516 24928 14525 24968
rect 16110 24928 16204 24968
rect 16244 24928 16253 24968
rect 20039 24928 20048 24968
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20416 24928 20425 24968
rect 0 24908 80 24928
rect 2500 24884 2540 24928
rect 6403 24927 6461 24928
rect 14467 24927 14525 24928
rect 16195 24927 16253 24928
rect 7459 24884 7517 24885
rect 16387 24884 16445 24885
rect 2500 24844 7468 24884
rect 7508 24844 7517 24884
rect 16302 24844 16396 24884
rect 16436 24844 16445 24884
rect 7459 24843 7517 24844
rect 16387 24843 16445 24844
rect 5539 24800 5597 24801
rect 6403 24800 6461 24801
rect 10243 24800 10301 24801
rect 21424 24800 21504 24820
rect 2092 24760 2540 24800
rect 3907 24760 3916 24800
rect 3956 24760 5548 24800
rect 5588 24760 5597 24800
rect 6211 24760 6220 24800
rect 6260 24760 6412 24800
rect 6452 24760 6461 24800
rect 7075 24760 7084 24800
rect 7124 24760 7756 24800
rect 7796 24760 7805 24800
rect 10243 24760 10252 24800
rect 10292 24760 21504 24800
rect 0 24632 80 24652
rect 2092 24632 2132 24760
rect 2500 24716 2540 24760
rect 5539 24759 5597 24760
rect 6403 24759 6461 24760
rect 10243 24759 10301 24760
rect 21424 24740 21504 24760
rect 8707 24716 8765 24717
rect 10819 24716 10877 24717
rect 2500 24676 8716 24716
rect 8756 24676 8765 24716
rect 9571 24676 9580 24716
rect 9620 24676 10828 24716
rect 10868 24676 10877 24716
rect 8707 24675 8765 24676
rect 10819 24675 10877 24676
rect 12268 24676 18988 24716
rect 19028 24676 19372 24716
rect 19412 24676 19421 24716
rect 20227 24676 20236 24716
rect 20276 24676 20716 24716
rect 20756 24676 20765 24716
rect 2755 24632 2813 24633
rect 8611 24632 8669 24633
rect 11683 24632 11741 24633
rect 0 24592 2132 24632
rect 2179 24592 2188 24632
rect 2228 24592 2540 24632
rect 2670 24592 2764 24632
rect 2804 24592 2813 24632
rect 3235 24592 3244 24632
rect 3284 24592 3532 24632
rect 3572 24592 3581 24632
rect 5155 24592 5164 24632
rect 5204 24592 5548 24632
rect 5588 24592 5740 24632
rect 5780 24592 5789 24632
rect 8419 24592 8428 24632
rect 8468 24592 8620 24632
rect 8660 24592 8669 24632
rect 10243 24592 10252 24632
rect 10292 24592 10732 24632
rect 10772 24592 10781 24632
rect 11491 24592 11500 24632
rect 11540 24592 11692 24632
rect 11732 24592 11741 24632
rect 0 24572 80 24592
rect 2500 24548 2540 24592
rect 2755 24591 2813 24592
rect 8611 24591 8669 24592
rect 11683 24591 11741 24592
rect 6211 24548 6269 24549
rect 12268 24548 12308 24676
rect 16291 24632 16349 24633
rect 12355 24592 12364 24632
rect 12404 24592 15340 24632
rect 15380 24592 15389 24632
rect 16206 24592 16300 24632
rect 16340 24592 16349 24632
rect 16291 24591 16349 24592
rect 2500 24508 3052 24548
rect 3092 24508 3101 24548
rect 5251 24508 5260 24548
rect 5300 24508 6028 24548
rect 6068 24508 6077 24548
rect 6211 24508 6220 24548
rect 6260 24508 12308 24548
rect 13987 24508 13996 24548
rect 14036 24508 15244 24548
rect 15284 24508 15916 24548
rect 15956 24508 15965 24548
rect 16099 24508 16108 24548
rect 16148 24508 17740 24548
rect 17780 24508 17789 24548
rect 6211 24507 6269 24508
rect 21424 24464 21504 24484
rect 4291 24424 4300 24464
rect 4340 24424 9484 24464
rect 9524 24424 12748 24464
rect 12788 24424 12797 24464
rect 13228 24424 21504 24464
rect 4291 24380 4349 24381
rect 13228 24380 13268 24424
rect 21424 24404 21504 24424
rect 16675 24380 16733 24381
rect 2947 24340 2956 24380
rect 2996 24340 3724 24380
rect 3764 24340 3773 24380
rect 4195 24340 4204 24380
rect 4244 24340 4300 24380
rect 4340 24340 10828 24380
rect 10868 24340 10877 24380
rect 12163 24340 12172 24380
rect 12212 24340 13268 24380
rect 15715 24340 15724 24380
rect 15764 24340 16108 24380
rect 16148 24340 16684 24380
rect 16724 24340 16733 24380
rect 4291 24339 4349 24340
rect 16675 24339 16733 24340
rect 0 24296 80 24316
rect 0 24256 18604 24296
rect 18644 24256 18653 24296
rect 0 24236 80 24256
rect 10531 24212 10589 24213
rect 16771 24212 16829 24213
rect 3679 24172 3688 24212
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 4056 24172 4065 24212
rect 6307 24172 6316 24212
rect 6356 24172 6796 24212
rect 6836 24172 6845 24212
rect 10446 24172 10540 24212
rect 10580 24172 10589 24212
rect 11107 24172 11116 24212
rect 11156 24172 12364 24212
rect 12404 24172 12413 24212
rect 14476 24172 14668 24212
rect 14708 24172 15092 24212
rect 10531 24171 10589 24172
rect 2755 24128 2813 24129
rect 14371 24128 14429 24129
rect 2755 24088 2764 24128
rect 2804 24088 14380 24128
rect 14420 24088 14429 24128
rect 2755 24087 2813 24088
rect 14371 24087 14429 24088
rect 3523 24004 3532 24044
rect 3572 24004 11116 24044
rect 11156 24004 11165 24044
rect 0 23960 80 23980
rect 355 23960 413 23961
rect 3235 23960 3293 23961
rect 14476 23960 14516 24172
rect 0 23920 364 23960
rect 404 23920 413 23960
rect 2179 23920 2188 23960
rect 2228 23920 2764 23960
rect 2804 23920 2813 23960
rect 3235 23920 3244 23960
rect 3284 23920 8180 23960
rect 8419 23920 8428 23960
rect 8468 23920 9964 23960
rect 10004 23920 10013 23960
rect 10723 23920 10732 23960
rect 10772 23920 11500 23960
rect 11540 23920 12460 23960
rect 12500 23920 12509 23960
rect 12835 23920 12844 23960
rect 12884 23920 13228 23960
rect 13268 23920 13277 23960
rect 14083 23920 14092 23960
rect 14132 23920 14516 23960
rect 15052 23960 15092 24172
rect 16771 24172 16780 24212
rect 16820 24172 17068 24212
rect 17108 24172 17117 24212
rect 18799 24172 18808 24212
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 19176 24172 19185 24212
rect 16771 24171 16829 24172
rect 21424 24129 21504 24148
rect 17443 24128 17501 24129
rect 21379 24128 21504 24129
rect 16483 24088 16492 24128
rect 16532 24088 16972 24128
rect 17012 24088 17021 24128
rect 17443 24088 17452 24128
rect 17492 24088 17548 24128
rect 17588 24088 17597 24128
rect 21379 24088 21388 24128
rect 21428 24088 21504 24128
rect 17443 24087 17501 24088
rect 21379 24087 21504 24088
rect 21424 24068 21504 24087
rect 16675 24004 16684 24044
rect 16724 24004 16733 24044
rect 16684 23960 16724 24004
rect 17155 23960 17213 23961
rect 15052 23920 16724 23960
rect 17070 23920 17164 23960
rect 17204 23920 17213 23960
rect 18595 23920 18604 23960
rect 18644 23920 20044 23960
rect 20084 23920 20093 23960
rect 0 23900 80 23920
rect 355 23919 413 23920
rect 3235 23919 3293 23920
rect 8140 23876 8180 23920
rect 17155 23919 17213 23920
rect 9379 23876 9437 23877
rect 14371 23876 14429 23877
rect 1987 23836 1996 23876
rect 2036 23836 5644 23876
rect 5684 23836 5932 23876
rect 5972 23836 5981 23876
rect 6499 23836 6508 23876
rect 6548 23836 7852 23876
rect 7892 23836 8044 23876
rect 8084 23836 8093 23876
rect 8140 23836 9388 23876
rect 9428 23836 9437 23876
rect 14286 23836 14380 23876
rect 14420 23836 14429 23876
rect 9379 23835 9437 23836
rect 14371 23835 14429 23836
rect 14668 23836 14764 23876
rect 14804 23836 14813 23876
rect 15427 23836 15436 23876
rect 15476 23836 15724 23876
rect 15764 23836 15773 23876
rect 16291 23836 16300 23876
rect 16340 23836 17644 23876
rect 17684 23836 18124 23876
rect 18164 23836 18173 23876
rect 3235 23792 3293 23793
rect 5539 23792 5597 23793
rect 172 23752 3244 23792
rect 3284 23752 3293 23792
rect 5155 23752 5164 23792
rect 5204 23752 5452 23792
rect 5492 23752 5548 23792
rect 5588 23752 5616 23792
rect 5827 23752 5836 23792
rect 5876 23752 6124 23792
rect 6164 23752 6173 23792
rect 7363 23752 7372 23792
rect 7412 23752 7756 23792
rect 7796 23752 7805 23792
rect 8803 23752 8812 23792
rect 8852 23752 10636 23792
rect 10676 23752 10685 23792
rect 10915 23752 10924 23792
rect 10964 23752 11596 23792
rect 11636 23752 11884 23792
rect 11924 23752 11933 23792
rect 12835 23752 12844 23792
rect 12884 23752 13132 23792
rect 13172 23752 13181 23792
rect 0 23624 80 23644
rect 0 23564 116 23624
rect 76 23540 116 23564
rect 172 23540 212 23752
rect 3235 23751 3293 23752
rect 5539 23751 5597 23752
rect 4579 23708 4637 23709
rect 8995 23708 9053 23709
rect 10051 23708 10109 23709
rect 14563 23708 14621 23709
rect 355 23668 364 23708
rect 404 23668 2860 23708
rect 2900 23668 4436 23708
rect 4291 23624 4349 23625
rect 3331 23584 3340 23624
rect 3380 23584 3532 23624
rect 3572 23584 3581 23624
rect 4003 23584 4012 23624
rect 4052 23584 4300 23624
rect 4340 23584 4349 23624
rect 4396 23624 4436 23668
rect 4579 23668 4588 23708
rect 4628 23668 5260 23708
rect 5300 23668 5309 23708
rect 7939 23668 7948 23708
rect 7988 23668 8332 23708
rect 8372 23668 8381 23708
rect 8899 23668 8908 23708
rect 8948 23668 9004 23708
rect 9044 23668 9053 23708
rect 9966 23668 10060 23708
rect 10100 23668 10109 23708
rect 14371 23668 14380 23708
rect 14420 23668 14572 23708
rect 14612 23668 14621 23708
rect 4579 23667 4637 23668
rect 8995 23667 9053 23668
rect 10051 23667 10109 23668
rect 14563 23667 14621 23668
rect 14668 23624 14708 23836
rect 20131 23792 20189 23793
rect 21424 23792 21504 23812
rect 15139 23752 15148 23792
rect 15188 23752 16684 23792
rect 16724 23752 17260 23792
rect 17300 23752 17309 23792
rect 18019 23752 18028 23792
rect 18068 23752 18412 23792
rect 18452 23752 19852 23792
rect 19892 23752 20084 23792
rect 20044 23708 20084 23752
rect 20131 23752 20140 23792
rect 20180 23752 21504 23792
rect 20131 23751 20189 23752
rect 21424 23732 21504 23752
rect 15523 23668 15532 23708
rect 15572 23668 17356 23708
rect 17396 23668 17405 23708
rect 20035 23668 20044 23708
rect 20084 23668 20093 23708
rect 4396 23584 10156 23624
rect 10196 23584 10205 23624
rect 14563 23584 14572 23624
rect 14612 23584 14708 23624
rect 14851 23584 14860 23624
rect 14900 23584 17644 23624
rect 17684 23584 17693 23624
rect 4291 23583 4349 23584
rect 11683 23540 11741 23541
rect 17827 23540 17885 23541
rect 76 23500 212 23540
rect 7555 23500 7564 23540
rect 7604 23500 8236 23540
rect 8276 23500 8285 23540
rect 11299 23500 11308 23540
rect 11348 23500 11692 23540
rect 11732 23500 11741 23540
rect 12739 23500 12748 23540
rect 12788 23500 15724 23540
rect 15764 23500 15773 23540
rect 17827 23500 17836 23540
rect 17876 23500 20564 23540
rect 11683 23499 11741 23500
rect 17827 23499 17885 23500
rect 20524 23456 20564 23500
rect 21424 23456 21504 23476
rect 4919 23416 4928 23456
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 5296 23416 5305 23456
rect 8803 23416 8812 23456
rect 8852 23416 9676 23456
rect 9716 23416 9725 23456
rect 11683 23416 11692 23456
rect 11732 23416 11884 23456
rect 11924 23416 11933 23456
rect 12835 23416 12844 23456
rect 12884 23416 17260 23456
rect 17300 23416 19468 23456
rect 19508 23416 19517 23456
rect 20039 23416 20048 23456
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20416 23416 20425 23456
rect 20524 23416 21504 23456
rect 21424 23396 21504 23416
rect 2083 23372 2141 23373
rect 268 23332 2092 23372
rect 2132 23332 2141 23372
rect 0 23288 80 23308
rect 268 23288 308 23332
rect 2083 23331 2141 23332
rect 4972 23332 5356 23372
rect 5396 23332 5405 23372
rect 8035 23332 8044 23372
rect 8084 23332 13324 23372
rect 13364 23332 13373 23372
rect 15619 23332 15628 23372
rect 15668 23332 17452 23372
rect 17492 23332 17501 23372
rect 4972 23288 5012 23332
rect 10243 23288 10301 23289
rect 14179 23288 14237 23289
rect 0 23248 308 23288
rect 2083 23248 2092 23288
rect 2132 23248 2668 23288
rect 2708 23248 2717 23288
rect 4963 23248 4972 23288
rect 5012 23248 5021 23288
rect 5443 23248 5452 23288
rect 5492 23248 5932 23288
rect 5972 23248 5981 23288
rect 6115 23248 6124 23288
rect 6164 23248 10252 23288
rect 10292 23248 10301 23288
rect 13987 23248 13996 23288
rect 14036 23248 14188 23288
rect 14228 23248 14237 23288
rect 14755 23248 14764 23288
rect 14804 23248 15052 23288
rect 15092 23248 17356 23288
rect 17396 23248 17932 23288
rect 17972 23248 17981 23288
rect 0 23228 80 23248
rect 10243 23247 10301 23248
rect 14179 23247 14237 23248
rect 163 23164 172 23204
rect 212 23164 3724 23204
rect 3764 23164 3773 23204
rect 9283 23164 9292 23204
rect 9332 23164 16204 23204
rect 16244 23164 16253 23204
rect 16867 23164 16876 23204
rect 16916 23164 18028 23204
rect 18068 23164 18077 23204
rect 10051 23120 10109 23121
rect 17443 23120 17501 23121
rect 21424 23120 21504 23140
rect 1891 23080 1900 23120
rect 1940 23080 5356 23120
rect 5396 23080 5405 23120
rect 6307 23080 6316 23120
rect 6356 23080 6796 23120
rect 6836 23080 8044 23120
rect 8084 23080 8093 23120
rect 9475 23080 9484 23120
rect 9524 23080 9868 23120
rect 9908 23080 9917 23120
rect 10051 23080 10060 23120
rect 10100 23080 10194 23120
rect 10531 23080 10540 23120
rect 10580 23080 11884 23120
rect 11924 23080 11933 23120
rect 12259 23080 12268 23120
rect 12308 23080 13996 23120
rect 14036 23080 14188 23120
rect 14228 23080 14237 23120
rect 14755 23080 14764 23120
rect 14804 23080 15148 23120
rect 15188 23080 15197 23120
rect 15811 23080 15820 23120
rect 15860 23080 16972 23120
rect 17012 23080 17021 23120
rect 17358 23080 17452 23120
rect 17492 23080 17501 23120
rect 18211 23080 18220 23120
rect 18260 23080 18700 23120
rect 18740 23080 18749 23120
rect 20995 23080 21004 23120
rect 21044 23080 21504 23120
rect 10051 23079 10109 23080
rect 17443 23079 17501 23080
rect 21424 23060 21504 23080
rect 16483 23036 16541 23037
rect 17155 23036 17213 23037
rect 3715 22996 3724 23036
rect 3764 22996 12556 23036
rect 12596 22996 12605 23036
rect 13219 22996 13228 23036
rect 13268 22996 16340 23036
rect 0 22952 80 22972
rect 16300 22952 16340 22996
rect 16483 22996 16492 23036
rect 16532 22996 17164 23036
rect 17204 22996 18796 23036
rect 18836 22996 18845 23036
rect 16483 22995 16541 22996
rect 17155 22995 17213 22996
rect 19267 22952 19325 22953
rect 0 22912 15532 22952
rect 15572 22912 15581 22952
rect 16300 22912 19276 22952
rect 19316 22912 19325 22952
rect 0 22892 80 22912
rect 19267 22911 19325 22912
rect 4579 22868 4637 22869
rect 5539 22868 5597 22869
rect 1219 22828 1228 22868
rect 1268 22828 4588 22868
rect 4628 22828 4637 22868
rect 5454 22828 5548 22868
rect 5588 22828 5597 22868
rect 4579 22827 4637 22828
rect 5539 22827 5597 22828
rect 8323 22868 8381 22869
rect 15043 22868 15101 22869
rect 16675 22868 16733 22869
rect 8323 22828 8332 22868
rect 8372 22828 15052 22868
rect 15092 22828 15101 22868
rect 16590 22828 16684 22868
rect 16724 22828 16733 22868
rect 8323 22827 8381 22828
rect 15043 22827 15101 22828
rect 16675 22827 16733 22828
rect 14947 22784 15005 22785
rect 19747 22784 19805 22785
rect 21424 22784 21504 22804
rect 4963 22744 4972 22784
rect 5012 22744 5644 22784
rect 5684 22744 5693 22784
rect 10627 22744 10636 22784
rect 10676 22744 11308 22784
rect 11348 22744 11357 22784
rect 13123 22744 13132 22784
rect 13172 22744 14572 22784
rect 14612 22744 14621 22784
rect 14947 22744 14956 22784
rect 14996 22744 15052 22784
rect 15092 22744 15101 22784
rect 15715 22744 15724 22784
rect 15764 22744 18316 22784
rect 18356 22744 18365 22784
rect 19747 22744 19756 22784
rect 19796 22744 21504 22784
rect 14947 22743 15005 22744
rect 19747 22743 19805 22744
rect 21424 22724 21504 22744
rect 8323 22700 8381 22701
rect 3679 22660 3688 22700
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 4056 22660 4065 22700
rect 7843 22660 7852 22700
rect 7892 22660 8332 22700
rect 8372 22660 8381 22700
rect 8323 22659 8381 22660
rect 12547 22700 12605 22701
rect 12547 22660 12556 22700
rect 12596 22660 12652 22700
rect 12692 22660 12701 22700
rect 14083 22660 14092 22700
rect 14132 22660 14284 22700
rect 14324 22660 16780 22700
rect 16820 22660 16829 22700
rect 17923 22660 17932 22700
rect 17972 22660 18412 22700
rect 18452 22660 18461 22700
rect 18799 22660 18808 22700
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 19176 22660 19185 22700
rect 12547 22659 12605 22660
rect 0 22616 80 22636
rect 0 22576 2188 22616
rect 2228 22576 2237 22616
rect 4771 22576 4780 22616
rect 4820 22576 5164 22616
rect 5204 22576 5213 22616
rect 11875 22576 11884 22616
rect 11924 22576 12556 22616
rect 12596 22576 13364 22616
rect 16387 22576 16396 22616
rect 16436 22576 19276 22616
rect 19316 22576 19564 22616
rect 19604 22576 19613 22616
rect 0 22556 80 22576
rect 3331 22532 3389 22533
rect 13324 22532 13364 22576
rect 19267 22532 19325 22533
rect 19459 22532 19517 22533
rect 1699 22492 1708 22532
rect 1748 22492 2380 22532
rect 2420 22492 2429 22532
rect 3331 22492 3340 22532
rect 3380 22492 4012 22532
rect 4052 22492 7372 22532
rect 7412 22492 9100 22532
rect 9140 22492 9580 22532
rect 9620 22492 9629 22532
rect 10243 22492 10252 22532
rect 10292 22492 13228 22532
rect 13268 22492 13277 22532
rect 13324 22492 16588 22532
rect 16628 22492 16637 22532
rect 19075 22492 19084 22532
rect 19124 22492 19276 22532
rect 19316 22492 19468 22532
rect 19508 22492 19517 22532
rect 3331 22491 3389 22492
rect 19267 22491 19325 22492
rect 19459 22491 19517 22492
rect 6019 22448 6077 22449
rect 14755 22448 14813 22449
rect 20131 22448 20189 22449
rect 21424 22448 21504 22468
rect 1603 22408 1612 22448
rect 1652 22408 5260 22448
rect 5300 22408 5309 22448
rect 6019 22408 6028 22448
rect 6068 22408 8332 22448
rect 8372 22408 8381 22448
rect 12355 22408 12364 22448
rect 12404 22408 12748 22448
rect 12788 22408 12797 22448
rect 14371 22408 14380 22448
rect 14420 22408 14764 22448
rect 14804 22408 14813 22448
rect 18211 22408 18220 22448
rect 18260 22408 18508 22448
rect 18548 22408 18557 22448
rect 18979 22408 18988 22448
rect 19028 22408 19372 22448
rect 19412 22408 19421 22448
rect 20131 22408 20140 22448
rect 20180 22408 21504 22448
rect 6019 22407 6077 22408
rect 14755 22407 14813 22408
rect 20131 22407 20189 22408
rect 21424 22388 21504 22408
rect 4675 22364 4733 22365
rect 6691 22364 6749 22365
rect 4675 22324 4684 22364
rect 4724 22324 4876 22364
rect 4916 22324 6700 22364
rect 6740 22324 6749 22364
rect 4675 22323 4733 22324
rect 6691 22323 6749 22324
rect 7363 22364 7421 22365
rect 7363 22324 7372 22364
rect 7412 22324 20180 22364
rect 7363 22323 7421 22324
rect 0 22280 80 22300
rect 2851 22280 2909 22281
rect 18595 22280 18653 22281
rect 0 22240 2860 22280
rect 2900 22240 2909 22280
rect 5827 22240 5836 22280
rect 5876 22240 6700 22280
rect 6740 22240 6749 22280
rect 10147 22240 10156 22280
rect 10196 22240 12748 22280
rect 12788 22240 13132 22280
rect 13172 22240 13181 22280
rect 13315 22240 13324 22280
rect 13364 22240 13516 22280
rect 13556 22240 15724 22280
rect 15764 22240 15773 22280
rect 18510 22240 18604 22280
rect 18644 22240 18892 22280
rect 18932 22240 18941 22280
rect 0 22220 80 22240
rect 2851 22239 2909 22240
rect 18595 22239 18653 22240
rect 5347 22196 5405 22197
rect 2851 22156 2860 22196
rect 2900 22156 4684 22196
rect 4724 22156 5356 22196
rect 5396 22156 5405 22196
rect 5347 22155 5405 22156
rect 6499 22112 6557 22113
rect 4291 22072 4300 22112
rect 4340 22072 5836 22112
rect 5876 22072 5885 22112
rect 6414 22072 6508 22112
rect 6548 22072 6557 22112
rect 6499 22071 6557 22072
rect 8995 22112 9053 22113
rect 20140 22112 20180 22324
rect 21424 22112 21504 22132
rect 8995 22072 9004 22112
rect 9044 22072 9484 22112
rect 9524 22072 9533 22112
rect 20140 22072 21504 22112
rect 8995 22071 9053 22072
rect 21424 22052 21504 22072
rect 3523 22028 3581 22029
rect 1123 21988 1132 22028
rect 1172 21988 3532 22028
rect 3572 21988 3581 22028
rect 14462 21988 14471 22028
rect 14511 21988 15916 22028
rect 15956 21988 15965 22028
rect 3523 21987 3581 21988
rect 0 21944 80 21964
rect 1891 21944 1949 21945
rect 0 21904 1900 21944
rect 1940 21904 1949 21944
rect 4919 21904 4928 21944
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 5296 21904 5305 21944
rect 7651 21904 7660 21944
rect 7700 21904 7852 21944
rect 7892 21904 12364 21944
rect 12404 21904 12413 21944
rect 20039 21904 20048 21944
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20416 21904 20425 21944
rect 0 21884 80 21904
rect 1891 21903 1949 21904
rect 13891 21820 13900 21860
rect 13940 21820 14476 21860
rect 14516 21820 14525 21860
rect 3427 21776 3485 21777
rect 20131 21776 20189 21777
rect 21424 21776 21504 21796
rect 3427 21736 3436 21776
rect 3476 21736 13652 21776
rect 14947 21736 14956 21776
rect 14996 21736 15340 21776
rect 15380 21736 15820 21776
rect 15860 21736 15869 21776
rect 20131 21736 20140 21776
rect 20180 21736 21504 21776
rect 3427 21735 3485 21736
rect 3148 21652 4012 21692
rect 4052 21652 4061 21692
rect 11320 21652 11596 21692
rect 11636 21652 11980 21692
rect 12020 21652 12029 21692
rect 0 21608 80 21628
rect 0 21568 1420 21608
rect 1460 21568 1469 21608
rect 0 21548 80 21568
rect 3148 21524 3188 21652
rect 7843 21608 7901 21609
rect 11320 21608 11360 21652
rect 3235 21568 3244 21608
rect 3284 21568 4204 21608
rect 4244 21568 4253 21608
rect 5731 21568 5740 21608
rect 5780 21568 6028 21608
rect 6068 21568 6077 21608
rect 7758 21568 7852 21608
rect 7892 21568 7901 21608
rect 9091 21568 9100 21608
rect 9140 21568 10388 21608
rect 10723 21568 10732 21608
rect 10772 21568 11360 21608
rect 13612 21608 13652 21736
rect 20131 21735 20189 21736
rect 21424 21716 21504 21736
rect 15523 21692 15581 21693
rect 15523 21652 15532 21692
rect 15572 21652 15668 21692
rect 18115 21652 18124 21692
rect 18164 21652 18412 21692
rect 18452 21652 18461 21692
rect 15523 21651 15581 21652
rect 14275 21608 14333 21609
rect 14467 21608 14525 21609
rect 15628 21608 15668 21652
rect 19267 21608 19325 21609
rect 13612 21568 13708 21608
rect 13748 21568 13757 21608
rect 13891 21568 13900 21608
rect 13940 21568 14284 21608
rect 14324 21568 14476 21608
rect 14516 21568 14525 21608
rect 14755 21568 14764 21608
rect 14804 21568 15532 21608
rect 15572 21568 15581 21608
rect 15628 21568 18644 21608
rect 18979 21568 18988 21608
rect 19028 21568 19276 21608
rect 19316 21568 19325 21608
rect 7843 21567 7901 21568
rect 3523 21524 3581 21525
rect 10243 21524 10301 21525
rect 2275 21484 2284 21524
rect 2324 21484 3188 21524
rect 3504 21484 3532 21524
rect 3572 21484 3628 21524
rect 3668 21484 10252 21524
rect 10292 21484 10301 21524
rect 10348 21524 10388 21568
rect 14275 21567 14333 21568
rect 14467 21567 14525 21568
rect 10348 21484 11788 21524
rect 11828 21484 13516 21524
rect 13556 21484 15244 21524
rect 15284 21484 15293 21524
rect 15715 21484 15724 21524
rect 15764 21484 17068 21524
rect 17108 21484 18548 21524
rect 3523 21483 3581 21484
rect 10243 21483 10301 21484
rect 14179 21440 14237 21441
rect 1315 21400 1324 21440
rect 1364 21400 5492 21440
rect 5539 21400 5548 21440
rect 5588 21400 6028 21440
rect 6068 21400 6077 21440
rect 6124 21400 8840 21440
rect 12259 21400 12268 21440
rect 12308 21400 14188 21440
rect 14228 21400 14764 21440
rect 14804 21400 14813 21440
rect 14947 21400 14956 21440
rect 14996 21400 15148 21440
rect 15188 21400 15340 21440
rect 15380 21400 16017 21440
rect 16057 21400 16066 21440
rect 5452 21356 5492 21400
rect 6124 21356 6164 21400
rect 8800 21356 8840 21400
rect 14179 21399 14237 21400
rect 10531 21356 10589 21357
rect 14659 21356 14717 21357
rect 18508 21356 18548 21484
rect 18604 21440 18644 21568
rect 19267 21567 19325 21568
rect 21424 21440 21504 21460
rect 18604 21400 21504 21440
rect 21424 21380 21504 21400
rect 5452 21316 6164 21356
rect 6211 21316 6220 21356
rect 6260 21316 7084 21356
rect 7124 21316 7133 21356
rect 8800 21316 10540 21356
rect 10580 21316 12844 21356
rect 12884 21316 12893 21356
rect 14659 21316 14668 21356
rect 14708 21316 16300 21356
rect 16340 21316 16349 21356
rect 17923 21316 17932 21356
rect 17972 21316 18316 21356
rect 18356 21316 18365 21356
rect 18499 21316 18508 21356
rect 18548 21316 18557 21356
rect 10531 21315 10589 21316
rect 14659 21315 14717 21316
rect 0 21272 80 21292
rect 13891 21272 13949 21273
rect 15619 21272 15677 21273
rect 0 21232 8236 21272
rect 8276 21232 8285 21272
rect 10732 21232 11212 21272
rect 11252 21232 11261 21272
rect 13891 21232 13900 21272
rect 13940 21232 15628 21272
rect 15668 21232 15677 21272
rect 0 21212 80 21232
rect 10732 21188 10772 21232
rect 13891 21231 13949 21232
rect 15619 21231 15677 21232
rect 3679 21148 3688 21188
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 4056 21148 4065 21188
rect 5731 21148 5740 21188
rect 5780 21148 6124 21188
rect 6164 21148 6173 21188
rect 10723 21148 10732 21188
rect 10772 21148 10781 21188
rect 18799 21148 18808 21188
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 19176 21148 19185 21188
rect 14179 21104 14237 21105
rect 13987 21064 13996 21104
rect 14036 21064 14188 21104
rect 14228 21064 14237 21104
rect 14179 21063 14237 21064
rect 16387 21104 16445 21105
rect 21424 21104 21504 21124
rect 16387 21064 16396 21104
rect 16436 21064 21504 21104
rect 16387 21063 16445 21064
rect 21424 21044 21504 21064
rect 9475 20980 9484 21020
rect 9524 20980 15724 21020
rect 15764 20980 15773 21020
rect 0 20936 80 20956
rect 16099 20936 16157 20937
rect 0 20896 6316 20936
rect 6356 20896 7276 20936
rect 7316 20896 7325 20936
rect 16099 20896 16108 20936
rect 16148 20896 21428 20936
rect 0 20876 80 20896
rect 16099 20895 16157 20896
rect 8323 20852 8381 20853
rect 9091 20852 9149 20853
rect 4003 20812 4012 20852
rect 4052 20812 8332 20852
rect 8372 20812 8381 20852
rect 9006 20812 9100 20852
rect 9140 20812 9292 20852
rect 9332 20812 9341 20852
rect 9955 20812 9964 20852
rect 10004 20812 11116 20852
rect 11156 20812 11165 20852
rect 8323 20811 8381 20812
rect 9091 20811 9149 20812
rect 21388 20788 21428 20896
rect 9571 20768 9629 20769
rect 15427 20768 15485 20769
rect 3139 20728 3148 20768
rect 3188 20728 6796 20768
rect 6836 20728 6845 20768
rect 9486 20728 9580 20768
rect 9620 20728 9772 20768
rect 9812 20728 9821 20768
rect 11011 20728 11020 20768
rect 11060 20728 11308 20768
rect 11348 20728 11357 20768
rect 13987 20728 13996 20768
rect 14036 20728 14956 20768
rect 14996 20728 15005 20768
rect 15342 20728 15436 20768
rect 15476 20728 15485 20768
rect 16099 20728 16108 20768
rect 16148 20728 16396 20768
rect 16436 20728 16445 20768
rect 16867 20728 16876 20768
rect 16916 20728 17644 20768
rect 17684 20728 17693 20768
rect 21388 20728 21504 20788
rect 9571 20727 9629 20728
rect 15427 20727 15485 20728
rect 21424 20708 21504 20728
rect 10339 20684 10397 20685
rect 16675 20684 16733 20685
rect 6307 20644 6316 20684
rect 6356 20644 7180 20684
rect 7220 20644 7229 20684
rect 10243 20644 10252 20684
rect 10292 20644 10348 20684
rect 10388 20644 10397 20684
rect 16590 20644 16684 20684
rect 16724 20644 16733 20684
rect 10339 20643 10397 20644
rect 16675 20643 16733 20644
rect 0 20600 80 20620
rect 0 20560 5164 20600
rect 5204 20560 5213 20600
rect 15331 20560 15340 20600
rect 15380 20560 16972 20600
rect 17012 20560 17021 20600
rect 17251 20560 17260 20600
rect 17300 20560 17548 20600
rect 17588 20560 17597 20600
rect 0 20540 80 20560
rect 10243 20476 10252 20516
rect 10292 20476 10636 20516
rect 10676 20476 10685 20516
rect 13219 20476 13228 20516
rect 13268 20476 20564 20516
rect 4919 20392 4928 20432
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 5296 20392 5305 20432
rect 10636 20348 10676 20476
rect 20524 20432 20564 20476
rect 21424 20432 21504 20452
rect 16579 20392 16588 20432
rect 16628 20392 17932 20432
rect 17972 20392 17981 20432
rect 20039 20392 20048 20432
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20416 20392 20425 20432
rect 20524 20392 21504 20432
rect 21424 20372 21504 20392
rect 12643 20348 12701 20349
rect 4771 20308 4780 20348
rect 4820 20308 7564 20348
rect 7604 20308 7613 20348
rect 10636 20308 12652 20348
rect 12692 20308 16876 20348
rect 16916 20308 16925 20348
rect 17059 20308 17068 20348
rect 17108 20308 17356 20348
rect 17396 20308 17405 20348
rect 12643 20307 12701 20308
rect 0 20264 80 20284
rect 15139 20264 15197 20265
rect 17827 20264 17885 20265
rect 0 20224 11020 20264
rect 11060 20224 11069 20264
rect 15139 20224 15148 20264
rect 15188 20224 15244 20264
rect 15284 20224 15293 20264
rect 17443 20224 17452 20264
rect 17492 20224 17836 20264
rect 17876 20224 17885 20264
rect 0 20204 80 20224
rect 15139 20223 15197 20224
rect 17827 20223 17885 20224
rect 16579 20180 16637 20181
rect 18595 20180 18653 20181
rect 20995 20180 21053 20181
rect 1987 20140 1996 20180
rect 2036 20140 2540 20180
rect 7524 20140 7564 20180
rect 7604 20140 7613 20180
rect 11212 20140 11596 20180
rect 11636 20140 11645 20180
rect 16579 20140 16588 20180
rect 16628 20140 16972 20180
rect 17012 20140 17021 20180
rect 18019 20140 18028 20180
rect 18068 20140 18220 20180
rect 18260 20140 18269 20180
rect 18595 20140 18604 20180
rect 18644 20140 18988 20180
rect 19028 20140 19037 20180
rect 20227 20140 20236 20180
rect 20276 20140 21004 20180
rect 21044 20140 21053 20180
rect 2500 20096 2540 20140
rect 3139 20096 3197 20097
rect 7564 20096 7604 20140
rect 11212 20096 11252 20140
rect 16579 20139 16637 20140
rect 18595 20139 18653 20140
rect 20995 20139 21053 20140
rect 15139 20096 15197 20097
rect 21424 20096 21504 20116
rect 2500 20056 2668 20096
rect 2708 20056 2717 20096
rect 3139 20056 3148 20096
rect 3188 20056 6988 20096
rect 7028 20056 7037 20096
rect 7564 20056 7852 20096
rect 7892 20056 7901 20096
rect 8707 20056 8716 20096
rect 8756 20056 8765 20096
rect 9379 20056 9388 20096
rect 9428 20056 11252 20096
rect 11320 20056 14284 20096
rect 14324 20056 14333 20096
rect 15139 20056 15148 20096
rect 15188 20056 15916 20096
rect 15956 20056 15965 20096
rect 16108 20056 21504 20096
rect 3139 20055 3197 20056
rect 8716 20012 8756 20056
rect 11320 20012 11360 20056
rect 15139 20055 15197 20056
rect 12931 20012 12989 20013
rect 3715 19972 3724 20012
rect 3764 19972 4492 20012
rect 4532 19972 8756 20012
rect 10819 19972 10828 20012
rect 10868 19972 11360 20012
rect 12835 19972 12844 20012
rect 12884 19972 12940 20012
rect 12980 19972 12989 20012
rect 0 19928 80 19948
rect 0 19888 1708 19928
rect 1748 19888 1757 19928
rect 0 19868 80 19888
rect 3724 19760 3764 19972
rect 12931 19971 12989 19972
rect 15331 20012 15389 20013
rect 16108 20012 16148 20056
rect 21424 20036 21504 20056
rect 19267 20012 19325 20013
rect 15331 19972 15340 20012
rect 15380 19972 16148 20012
rect 18604 19972 18796 20012
rect 18836 19972 18845 20012
rect 19075 19972 19084 20012
rect 19124 19972 19276 20012
rect 19316 19972 19468 20012
rect 19508 19972 19517 20012
rect 15331 19971 15389 19972
rect 16675 19928 16733 19929
rect 18604 19928 18644 19972
rect 19267 19971 19325 19972
rect 5347 19888 5356 19928
rect 5396 19888 8332 19928
rect 8372 19888 8381 19928
rect 11299 19888 11308 19928
rect 11348 19888 16684 19928
rect 16724 19888 16972 19928
rect 17012 19888 17021 19928
rect 17251 19888 17260 19928
rect 17300 19888 17740 19928
rect 17780 19888 17789 19928
rect 18595 19888 18604 19928
rect 18644 19888 18653 19928
rect 16675 19887 16733 19888
rect 5731 19844 5789 19845
rect 10051 19844 10109 19845
rect 4483 19804 4492 19844
rect 4532 19804 5164 19844
rect 5204 19804 5213 19844
rect 5731 19804 5740 19844
rect 5780 19804 10060 19844
rect 10100 19804 10109 19844
rect 15043 19804 15052 19844
rect 15092 19804 17452 19844
rect 17492 19804 17501 19844
rect 5731 19803 5789 19804
rect 10051 19803 10109 19804
rect 20611 19760 20669 19761
rect 21424 19760 21504 19780
rect 1987 19720 1996 19760
rect 2036 19720 3764 19760
rect 5443 19720 5452 19760
rect 5492 19720 6124 19760
rect 6164 19720 6604 19760
rect 6644 19720 11980 19760
rect 12020 19720 15436 19760
rect 15476 19720 16108 19760
rect 16148 19720 16157 19760
rect 20611 19720 20620 19760
rect 20660 19720 21504 19760
rect 20611 19719 20669 19720
rect 21424 19700 21504 19720
rect 3679 19636 3688 19676
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 4056 19636 4065 19676
rect 12067 19636 12076 19676
rect 12116 19636 14092 19676
rect 14132 19636 14141 19676
rect 18799 19636 18808 19676
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 19176 19636 19185 19676
rect 20035 19636 20044 19676
rect 20084 19636 20524 19676
rect 20564 19636 20573 19676
rect 0 19592 80 19612
rect 1987 19592 2045 19593
rect 10051 19592 10109 19593
rect 14755 19592 14813 19593
rect 0 19552 1804 19592
rect 1844 19552 1853 19592
rect 1987 19552 1996 19592
rect 2036 19552 2092 19592
rect 2132 19552 5356 19592
rect 5396 19552 5405 19592
rect 10051 19552 10060 19592
rect 10100 19552 10828 19592
rect 10868 19552 11404 19592
rect 11444 19552 11453 19592
rect 14755 19552 14764 19592
rect 14804 19552 14860 19592
rect 14900 19552 14909 19592
rect 16003 19552 16012 19592
rect 16052 19552 18220 19592
rect 18260 19552 19756 19592
rect 19796 19552 19805 19592
rect 0 19532 80 19552
rect 1987 19551 2045 19552
rect 10051 19551 10109 19552
rect 14755 19551 14813 19552
rect 16291 19508 16349 19509
rect 3427 19468 3436 19508
rect 3476 19468 3628 19508
rect 3668 19468 3677 19508
rect 8323 19468 8332 19508
rect 8372 19468 16300 19508
rect 16340 19468 16349 19508
rect 16291 19467 16349 19468
rect 5731 19424 5789 19425
rect 15523 19424 15581 19425
rect 19363 19424 19421 19425
rect 1315 19384 1324 19424
rect 1364 19384 5740 19424
rect 5780 19384 5789 19424
rect 9187 19384 9196 19424
rect 9236 19384 10060 19424
rect 10100 19384 10109 19424
rect 13891 19384 13900 19424
rect 13940 19384 14188 19424
rect 14228 19384 14237 19424
rect 15523 19384 15532 19424
rect 15572 19384 15724 19424
rect 15764 19384 15773 19424
rect 16483 19384 16492 19424
rect 16532 19384 19372 19424
rect 19412 19384 19421 19424
rect 5731 19383 5789 19384
rect 15523 19383 15581 19384
rect 19363 19383 19421 19384
rect 20803 19424 20861 19425
rect 21424 19424 21504 19444
rect 20803 19384 20812 19424
rect 20852 19384 21504 19424
rect 20803 19383 20861 19384
rect 21424 19364 21504 19384
rect 2371 19340 2429 19341
rect 2371 19300 2380 19340
rect 2420 19300 4396 19340
rect 4436 19300 6988 19340
rect 7028 19300 11308 19340
rect 11348 19300 11357 19340
rect 16387 19300 16396 19340
rect 16436 19300 17164 19340
rect 17204 19300 17213 19340
rect 2371 19299 2429 19300
rect 0 19256 80 19276
rect 13603 19256 13661 19257
rect 0 19216 76 19256
rect 116 19216 125 19256
rect 2755 19216 2764 19256
rect 2804 19216 3244 19256
rect 3284 19216 3293 19256
rect 4003 19216 4012 19256
rect 4052 19216 4300 19256
rect 4340 19216 4349 19256
rect 10243 19216 10252 19256
rect 10292 19216 10540 19256
rect 10580 19216 10589 19256
rect 13518 19216 13612 19256
rect 13652 19216 13804 19256
rect 13844 19216 13853 19256
rect 15619 19216 15628 19256
rect 15668 19216 18028 19256
rect 18068 19216 18077 19256
rect 18307 19216 18316 19256
rect 18356 19216 19852 19256
rect 19892 19216 19901 19256
rect 0 19196 80 19216
rect 13603 19215 13661 19216
rect 4387 19172 4445 19173
rect 1315 19132 1324 19172
rect 1364 19132 4396 19172
rect 4436 19132 4445 19172
rect 6691 19132 6700 19172
rect 6740 19132 11360 19172
rect 11587 19132 11596 19172
rect 11636 19132 14668 19172
rect 14708 19132 14717 19172
rect 14851 19132 14860 19172
rect 14900 19132 15820 19172
rect 15860 19132 15869 19172
rect 16099 19132 16108 19172
rect 16148 19132 16300 19172
rect 16340 19132 16684 19172
rect 16724 19132 16733 19172
rect 4387 19131 4445 19132
rect 3523 19048 3532 19088
rect 3572 19048 6316 19088
rect 6356 19048 10484 19088
rect 3139 19004 3197 19005
rect 10444 19004 10484 19048
rect 11320 19004 11360 19132
rect 14371 19088 14429 19089
rect 21424 19088 21504 19108
rect 14083 19048 14092 19088
rect 14132 19048 14380 19088
rect 14420 19048 14429 19088
rect 14755 19048 14764 19088
rect 14804 19048 17164 19088
rect 17204 19048 17213 19088
rect 20140 19048 21504 19088
rect 14371 19047 14429 19048
rect 15715 19004 15773 19005
rect 20140 19004 20180 19048
rect 21424 19028 21504 19048
rect 1219 18964 1228 19004
rect 1268 18964 3148 19004
rect 3188 18964 3197 19004
rect 8227 18964 8236 19004
rect 8276 18964 9964 19004
rect 10004 18964 10252 19004
rect 10292 18964 10301 19004
rect 10435 18964 10444 19004
rect 10484 18964 10493 19004
rect 11320 18964 13420 19004
rect 13460 18964 14284 19004
rect 14324 18964 14333 19004
rect 14467 18964 14476 19004
rect 14516 18964 14525 19004
rect 15139 18964 15148 19004
rect 15188 18964 15532 19004
rect 15572 18964 15581 19004
rect 15715 18964 15724 19004
rect 15764 18964 20180 19004
rect 3139 18963 3197 18964
rect 0 18920 80 18940
rect 2275 18920 2333 18921
rect 14476 18920 14516 18964
rect 15715 18963 15773 18964
rect 15907 18920 15965 18921
rect 16579 18920 16637 18921
rect 0 18880 940 18920
rect 980 18880 989 18920
rect 2275 18880 2284 18920
rect 2324 18880 4684 18920
rect 4724 18880 4733 18920
rect 4919 18880 4928 18920
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 5296 18880 5305 18920
rect 5347 18880 5356 18920
rect 5396 18880 7084 18920
rect 7124 18880 10732 18920
rect 10772 18880 10781 18920
rect 11971 18880 11980 18920
rect 12020 18880 12364 18920
rect 12404 18880 12413 18920
rect 14476 18880 14612 18920
rect 14659 18880 14668 18920
rect 14708 18880 15628 18920
rect 15668 18880 15677 18920
rect 15907 18880 15916 18920
rect 15956 18880 16588 18920
rect 16628 18880 16637 18920
rect 18595 18880 18604 18920
rect 18644 18880 18796 18920
rect 18836 18880 18845 18920
rect 20039 18880 20048 18920
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20416 18880 20425 18920
rect 0 18860 80 18880
rect 2275 18879 2333 18880
rect 14572 18836 14612 18880
rect 15907 18879 15965 18880
rect 16579 18879 16637 18880
rect 3139 18796 3148 18836
rect 3188 18796 4012 18836
rect 4052 18796 4061 18836
rect 5443 18796 5452 18836
rect 5492 18796 6028 18836
rect 6068 18796 6604 18836
rect 6644 18796 6653 18836
rect 10243 18796 10252 18836
rect 10292 18796 12076 18836
rect 12116 18796 12268 18836
rect 12308 18796 12317 18836
rect 14572 18796 16780 18836
rect 16820 18796 16829 18836
rect 14755 18752 14813 18753
rect 10339 18712 10348 18752
rect 10388 18712 10828 18752
rect 10868 18712 10877 18752
rect 14179 18712 14188 18752
rect 14228 18712 14572 18752
rect 14612 18712 14621 18752
rect 14670 18712 14764 18752
rect 14804 18712 14813 18752
rect 14755 18711 14813 18712
rect 16867 18752 16925 18753
rect 21424 18752 21504 18772
rect 16867 18712 16876 18752
rect 16916 18712 21504 18752
rect 16867 18711 16925 18712
rect 21424 18692 21504 18712
rect 1411 18628 1420 18668
rect 1460 18628 2476 18668
rect 2516 18628 2525 18668
rect 9571 18628 9580 18668
rect 9620 18628 13516 18668
rect 13556 18628 14476 18668
rect 14516 18628 14525 18668
rect 16099 18628 16108 18668
rect 16148 18628 18508 18668
rect 18548 18628 19660 18668
rect 19700 18628 19709 18668
rect 0 18584 80 18604
rect 6019 18584 6077 18585
rect 14851 18584 14909 18585
rect 19267 18584 19325 18585
rect 0 18544 6028 18584
rect 6068 18544 6077 18584
rect 12259 18544 12268 18584
rect 12308 18544 14668 18584
rect 14708 18544 14717 18584
rect 14851 18544 14860 18584
rect 14900 18544 15052 18584
rect 15092 18544 15101 18584
rect 15427 18544 15436 18584
rect 15476 18544 16300 18584
rect 16340 18544 16349 18584
rect 16579 18544 16588 18584
rect 16628 18544 16876 18584
rect 16916 18544 17644 18584
rect 17684 18544 17693 18584
rect 19182 18544 19276 18584
rect 19316 18544 19325 18584
rect 0 18524 80 18544
rect 6019 18543 6077 18544
rect 14851 18543 14909 18544
rect 19267 18543 19325 18544
rect 3331 18460 3340 18500
rect 3380 18460 3628 18500
rect 3668 18460 6700 18500
rect 6740 18460 6749 18500
rect 9091 18460 9100 18500
rect 9140 18460 9868 18500
rect 9908 18460 18796 18500
rect 18836 18460 18845 18500
rect 6787 18416 6845 18417
rect 17827 18416 17885 18417
rect 6115 18376 6124 18416
rect 6164 18376 6796 18416
rect 6836 18376 6845 18416
rect 17443 18376 17452 18416
rect 17492 18376 17836 18416
rect 17876 18376 17885 18416
rect 6787 18375 6845 18376
rect 17827 18375 17885 18376
rect 18211 18416 18269 18417
rect 21424 18416 21504 18436
rect 18211 18376 18220 18416
rect 18260 18376 21504 18416
rect 18211 18375 18269 18376
rect 21424 18356 21504 18376
rect 6403 18332 6461 18333
rect 6211 18292 6220 18332
rect 6260 18292 6412 18332
rect 6452 18292 6461 18332
rect 17539 18292 17548 18332
rect 17588 18292 18316 18332
rect 18356 18292 18365 18332
rect 6403 18291 6461 18292
rect 0 18248 80 18268
rect 0 18208 6028 18248
rect 6068 18208 6077 18248
rect 7555 18208 7564 18248
rect 7604 18208 7756 18248
rect 7796 18208 7805 18248
rect 8995 18208 9004 18248
rect 9044 18208 14476 18248
rect 14516 18208 18412 18248
rect 18452 18208 18461 18248
rect 0 18188 80 18208
rect 2755 18164 2813 18165
rect 2659 18124 2668 18164
rect 2708 18124 2764 18164
rect 2804 18124 2813 18164
rect 3679 18124 3688 18164
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 4056 18124 4065 18164
rect 18799 18124 18808 18164
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 19176 18124 19185 18164
rect 2755 18123 2813 18124
rect 21424 18080 21504 18100
rect 7747 18040 7756 18080
rect 7796 18040 21504 18080
rect 21424 18020 21504 18040
rect 14275 17956 14284 17996
rect 14324 17956 14860 17996
rect 14900 17956 14909 17996
rect 16291 17956 16300 17996
rect 16340 17956 16684 17996
rect 16724 17956 16733 17996
rect 17635 17956 17644 17996
rect 17684 17956 18604 17996
rect 18644 17956 19564 17996
rect 19604 17956 19613 17996
rect 0 17912 80 17932
rect 13219 17912 13277 17913
rect 17347 17912 17405 17913
rect 0 17872 1612 17912
rect 1652 17872 1661 17912
rect 13219 17872 13228 17912
rect 13268 17872 17356 17912
rect 17396 17872 17405 17912
rect 0 17852 80 17872
rect 13219 17871 13277 17872
rect 17347 17871 17405 17872
rect 9379 17828 9437 17829
rect 9091 17788 9100 17828
rect 9140 17788 9388 17828
rect 9428 17788 9437 17828
rect 9379 17787 9437 17788
rect 10627 17828 10685 17829
rect 10627 17788 10636 17828
rect 10676 17788 12460 17828
rect 12500 17788 12509 17828
rect 15427 17788 15436 17828
rect 15476 17788 16204 17828
rect 16244 17788 16253 17828
rect 16675 17788 16684 17828
rect 16724 17788 18604 17828
rect 18644 17788 19180 17828
rect 19220 17788 19229 17828
rect 10627 17787 10685 17788
rect 21424 17744 21504 17764
rect 2467 17704 2476 17744
rect 2516 17704 5452 17744
rect 5492 17704 5644 17744
rect 5684 17704 5693 17744
rect 6019 17704 6028 17744
rect 6068 17704 21504 17744
rect 2755 17660 2813 17661
rect 6028 17660 6068 17704
rect 21424 17684 21504 17704
rect 12451 17660 12509 17661
rect 2659 17620 2668 17660
rect 2708 17620 2764 17660
rect 2804 17620 2813 17660
rect 3427 17620 3436 17660
rect 3476 17620 6068 17660
rect 12366 17620 12460 17660
rect 12500 17620 12509 17660
rect 15235 17620 15244 17660
rect 15284 17620 16780 17660
rect 16820 17620 16829 17660
rect 2755 17619 2813 17620
rect 12451 17619 12509 17620
rect 0 17576 80 17596
rect 12460 17576 12500 17619
rect 0 17536 11116 17576
rect 11156 17536 11165 17576
rect 12460 17536 13420 17576
rect 13460 17536 13469 17576
rect 17923 17536 17932 17576
rect 17972 17536 19852 17576
rect 19892 17536 19901 17576
rect 0 17516 80 17536
rect 18691 17452 18700 17492
rect 18740 17452 19372 17492
rect 19412 17452 19421 17492
rect 6883 17408 6941 17409
rect 20611 17408 20669 17409
rect 21424 17408 21504 17428
rect 3139 17368 3148 17408
rect 3188 17368 3340 17408
rect 3380 17368 3389 17408
rect 4919 17368 4928 17408
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 5296 17368 5305 17408
rect 6691 17368 6700 17408
rect 6740 17368 6892 17408
rect 6932 17368 6941 17408
rect 11107 17368 11116 17408
rect 11156 17368 11308 17408
rect 11348 17368 11357 17408
rect 20039 17368 20048 17408
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20416 17368 20425 17408
rect 20611 17368 20620 17408
rect 20660 17368 21504 17408
rect 6883 17367 6941 17368
rect 20611 17367 20669 17368
rect 21424 17348 21504 17368
rect 2500 17284 10156 17324
rect 10196 17284 10205 17324
rect 0 17240 80 17260
rect 2500 17240 2540 17284
rect 15715 17240 15773 17241
rect 0 17200 2540 17240
rect 3235 17200 3244 17240
rect 3284 17200 3860 17240
rect 7363 17200 7372 17240
rect 7412 17200 8332 17240
rect 8372 17200 10444 17240
rect 10484 17200 12556 17240
rect 12596 17200 13996 17240
rect 14036 17200 14572 17240
rect 14612 17200 14621 17240
rect 15630 17200 15724 17240
rect 15764 17200 15773 17240
rect 17731 17200 17740 17240
rect 17780 17200 18316 17240
rect 18356 17200 18796 17240
rect 18836 17200 19084 17240
rect 19124 17200 20044 17240
rect 20084 17200 20093 17240
rect 0 17180 80 17200
rect 3820 17072 3860 17200
rect 15715 17199 15773 17200
rect 16483 17156 16541 17157
rect 9187 17116 9196 17156
rect 9236 17116 9484 17156
rect 9524 17116 9533 17156
rect 13324 17116 16492 17156
rect 16532 17116 16541 17156
rect 19267 17116 19276 17156
rect 19316 17116 20140 17156
rect 20180 17116 20189 17156
rect 13324 17072 13364 17116
rect 16483 17115 16541 17116
rect 21424 17073 21504 17092
rect 13891 17072 13949 17073
rect 19459 17072 19517 17073
rect 21379 17072 21504 17073
rect 3811 17032 3820 17072
rect 3860 17032 4684 17072
rect 4724 17032 5356 17072
rect 5396 17032 5548 17072
rect 5588 17032 5597 17072
rect 5644 17032 6316 17072
rect 6356 17032 6365 17072
rect 8611 17032 8620 17072
rect 8660 17032 10156 17072
rect 10196 17032 10732 17072
rect 10772 17032 10781 17072
rect 11299 17032 11308 17072
rect 11348 17032 11596 17072
rect 11636 17032 11884 17072
rect 11924 17032 11933 17072
rect 13315 17032 13324 17072
rect 13364 17032 13373 17072
rect 13891 17032 13900 17072
rect 13940 17032 15148 17072
rect 15188 17032 15724 17072
rect 15764 17032 15773 17072
rect 16387 17032 16396 17072
rect 16436 17032 17356 17072
rect 17396 17032 17405 17072
rect 19459 17032 19468 17072
rect 19508 17032 19948 17072
rect 19988 17032 19997 17072
rect 21379 17032 21388 17072
rect 21428 17032 21504 17072
rect 3331 16988 3389 16989
rect 5644 16988 5684 17032
rect 3246 16948 3340 16988
rect 3380 16948 5684 16988
rect 5827 16948 5836 16988
rect 5876 16948 6124 16988
rect 6164 16948 9964 16988
rect 10004 16948 10013 16988
rect 3331 16947 3389 16948
rect 0 16904 80 16924
rect 4675 16904 4733 16905
rect 13324 16904 13364 17032
rect 13891 17031 13949 17032
rect 19459 17031 19517 17032
rect 21379 17031 21504 17032
rect 21424 17012 21504 17031
rect 14563 16948 14572 16988
rect 14612 16948 15244 16988
rect 15284 16948 15293 16988
rect 0 16864 4684 16904
rect 4724 16864 4733 16904
rect 7843 16864 7852 16904
rect 7892 16864 8140 16904
rect 8180 16864 13364 16904
rect 0 16844 80 16864
rect 4675 16863 4733 16864
rect 2659 16780 2668 16820
rect 2708 16780 3436 16820
rect 3476 16780 3485 16820
rect 6499 16780 6508 16820
rect 6548 16780 7180 16820
rect 7220 16780 7229 16820
rect 14275 16780 14284 16820
rect 14324 16780 14764 16820
rect 14804 16780 14813 16820
rect 9379 16736 9437 16737
rect 2500 16696 5932 16736
rect 5972 16696 5981 16736
rect 9294 16696 9388 16736
rect 9428 16696 9437 16736
rect 0 16568 80 16588
rect 2500 16568 2540 16696
rect 9379 16695 9437 16696
rect 16387 16736 16445 16737
rect 21424 16736 21504 16756
rect 16387 16696 16396 16736
rect 16436 16696 21504 16736
rect 16387 16695 16445 16696
rect 21424 16676 21504 16696
rect 6691 16652 6749 16653
rect 2851 16612 2860 16652
rect 2900 16612 3340 16652
rect 3380 16612 3389 16652
rect 3679 16612 3688 16652
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 4056 16612 4065 16652
rect 6606 16612 6700 16652
rect 6740 16612 6749 16652
rect 9283 16612 9292 16652
rect 9332 16612 9868 16652
rect 9908 16612 9917 16652
rect 18799 16612 18808 16652
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 19176 16612 19185 16652
rect 6691 16611 6749 16612
rect 6595 16568 6653 16569
rect 7843 16568 7901 16569
rect 0 16528 2540 16568
rect 5731 16528 5740 16568
rect 5780 16528 5789 16568
rect 6595 16528 6604 16568
rect 6644 16528 7852 16568
rect 7892 16528 7901 16568
rect 0 16508 80 16528
rect 5740 16484 5780 16528
rect 6595 16527 6653 16528
rect 7843 16527 7901 16528
rect 19267 16484 19325 16485
rect 3043 16444 3052 16484
rect 3092 16444 3532 16484
rect 3572 16444 11360 16484
rect 18307 16444 18316 16484
rect 18356 16444 18892 16484
rect 18932 16444 18941 16484
rect 19267 16444 19276 16484
rect 19316 16444 19372 16484
rect 19412 16444 19421 16484
rect 4483 16400 4541 16401
rect 11320 16400 11360 16444
rect 19267 16443 19325 16444
rect 21424 16400 21504 16420
rect 3139 16360 3148 16400
rect 3188 16360 3724 16400
rect 3764 16360 3773 16400
rect 4387 16360 4396 16400
rect 4436 16360 4492 16400
rect 4532 16360 6164 16400
rect 6403 16360 6412 16400
rect 6452 16360 6700 16400
rect 6740 16360 6749 16400
rect 9676 16360 10252 16400
rect 10292 16360 10301 16400
rect 11320 16360 21504 16400
rect 4483 16359 4541 16360
rect 6124 16316 6164 16360
rect 3523 16276 3532 16316
rect 3572 16276 6028 16316
rect 6068 16276 6077 16316
rect 6124 16276 9484 16316
rect 9524 16276 9533 16316
rect 0 16232 80 16252
rect 0 16192 7660 16232
rect 7700 16192 7709 16232
rect 8707 16192 8716 16232
rect 8756 16192 9100 16232
rect 9140 16192 9149 16232
rect 0 16172 80 16192
rect 7363 16064 7421 16065
rect 67 16024 76 16064
rect 116 16024 1228 16064
rect 1268 16024 1277 16064
rect 7278 16024 7372 16064
rect 7412 16024 7421 16064
rect 7363 16023 7421 16024
rect 9676 15980 9716 16360
rect 21424 16340 21504 16360
rect 19939 16316 19997 16317
rect 9955 16276 9964 16316
rect 10004 16276 10828 16316
rect 10868 16276 10877 16316
rect 17251 16276 17260 16316
rect 17300 16276 17644 16316
rect 17684 16276 17693 16316
rect 18508 16276 19948 16316
rect 19988 16276 20044 16316
rect 20084 16276 20093 16316
rect 15523 16232 15581 16233
rect 10723 16192 10732 16232
rect 10772 16192 13804 16232
rect 13844 16192 13853 16232
rect 15523 16192 15532 16232
rect 15572 16192 15724 16232
rect 15764 16192 16588 16232
rect 16628 16192 16637 16232
rect 18019 16192 18028 16232
rect 18068 16192 18077 16232
rect 15523 16191 15581 16192
rect 15907 16148 15965 16149
rect 10531 16108 10540 16148
rect 10580 16108 11308 16148
rect 11348 16108 11357 16148
rect 15822 16108 15916 16148
rect 15956 16108 15965 16148
rect 15907 16107 15965 16108
rect 11491 16064 11549 16065
rect 11491 16024 11500 16064
rect 11540 16024 12172 16064
rect 12212 16024 12221 16064
rect 14083 16024 14092 16064
rect 14132 16024 14476 16064
rect 14516 16024 14525 16064
rect 15523 16024 15532 16064
rect 15572 16024 15724 16064
rect 15764 16024 15773 16064
rect 16003 16024 16012 16064
rect 16052 16024 16300 16064
rect 16340 16024 16349 16064
rect 16483 16024 16492 16064
rect 16532 16024 17164 16064
rect 17204 16024 17213 16064
rect 11491 16023 11549 16024
rect 16300 15980 16340 16024
rect 2755 15940 2764 15980
rect 2804 15940 3244 15980
rect 3284 15940 4492 15980
rect 4532 15940 5740 15980
rect 5780 15940 8908 15980
rect 8948 15940 8957 15980
rect 9667 15940 9676 15980
rect 9716 15940 9725 15980
rect 10147 15940 10156 15980
rect 10196 15940 16204 15980
rect 16244 15940 16253 15980
rect 16300 15940 17588 15980
rect 0 15896 80 15916
rect 0 15856 2540 15896
rect 4919 15856 4928 15896
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 5296 15856 5305 15896
rect 6211 15856 6220 15896
rect 6260 15856 10540 15896
rect 10580 15856 10589 15896
rect 10723 15856 10732 15896
rect 10772 15856 11116 15896
rect 11156 15856 11165 15896
rect 11320 15856 17452 15896
rect 17492 15856 17501 15896
rect 0 15836 80 15856
rect 2500 15812 2540 15856
rect 11320 15812 11360 15856
rect 2500 15772 11360 15812
rect 15331 15812 15389 15813
rect 17548 15812 17588 15940
rect 18028 15896 18068 16192
rect 18508 16148 18548 16276
rect 19939 16275 19997 16276
rect 18595 16192 18604 16232
rect 18644 16192 19852 16232
rect 19892 16192 19901 16232
rect 18499 16108 18508 16148
rect 18548 16108 18557 16148
rect 18691 16108 18700 16148
rect 18740 16108 19756 16148
rect 19796 16108 19805 16148
rect 21424 16064 21504 16084
rect 18403 16024 18412 16064
rect 18452 16024 19084 16064
rect 19124 16024 19133 16064
rect 19363 16024 19372 16064
rect 19412 16024 20044 16064
rect 20084 16024 20093 16064
rect 20524 16024 21504 16064
rect 20524 15980 20564 16024
rect 21424 16004 21504 16024
rect 19171 15940 19180 15980
rect 19220 15940 20564 15980
rect 17933 15856 18028 15896
rect 18068 15856 19276 15896
rect 19316 15856 19325 15896
rect 20039 15856 20048 15896
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20416 15856 20425 15896
rect 19267 15812 19325 15813
rect 15331 15772 15340 15812
rect 15380 15772 16108 15812
rect 16148 15772 16157 15812
rect 16492 15772 16972 15812
rect 17012 15772 17021 15812
rect 17548 15772 19276 15812
rect 19316 15772 19325 15812
rect 15331 15771 15389 15772
rect 1219 15688 1228 15728
rect 1268 15688 1996 15728
rect 2036 15688 2045 15728
rect 15715 15688 15724 15728
rect 15764 15688 16012 15728
rect 16052 15688 16061 15728
rect 2755 15644 2813 15645
rect 16099 15644 16157 15645
rect 16492 15644 16532 15772
rect 19267 15771 19325 15772
rect 21424 15728 21504 15748
rect 16579 15688 16588 15728
rect 16628 15688 21504 15728
rect 21424 15668 21504 15688
rect 2083 15604 2092 15644
rect 2132 15604 2764 15644
rect 2804 15604 3724 15644
rect 3764 15604 3773 15644
rect 11683 15604 11692 15644
rect 11732 15604 13132 15644
rect 13172 15604 13181 15644
rect 16099 15604 16108 15644
rect 16148 15604 16492 15644
rect 16532 15604 16541 15644
rect 16867 15604 16876 15644
rect 16916 15604 17452 15644
rect 17492 15604 17501 15644
rect 19555 15604 19564 15644
rect 19604 15604 20044 15644
rect 20084 15604 20093 15644
rect 2755 15603 2813 15604
rect 16099 15603 16157 15604
rect 0 15560 80 15580
rect 15139 15560 15197 15561
rect 17635 15560 17693 15561
rect 18595 15560 18653 15561
rect 0 15520 2860 15560
rect 2900 15520 2909 15560
rect 4963 15520 4972 15560
rect 5012 15520 6604 15560
rect 6644 15520 10060 15560
rect 10100 15520 10109 15560
rect 10339 15520 10348 15560
rect 10388 15520 11116 15560
rect 11156 15520 13228 15560
rect 13268 15520 13277 15560
rect 14659 15520 14668 15560
rect 14708 15520 15148 15560
rect 15188 15520 15436 15560
rect 15476 15520 15485 15560
rect 15619 15520 15628 15560
rect 15668 15520 16300 15560
rect 16340 15520 16349 15560
rect 17635 15520 17644 15560
rect 17684 15520 17740 15560
rect 17780 15520 18604 15560
rect 18644 15520 18653 15560
rect 18883 15520 18892 15560
rect 18932 15520 19372 15560
rect 19412 15520 19421 15560
rect 0 15500 80 15520
rect 15139 15519 15197 15520
rect 17635 15519 17693 15520
rect 18595 15519 18653 15520
rect 4483 15476 4541 15477
rect 7459 15476 7517 15477
rect 18211 15476 18269 15477
rect 19939 15476 19997 15477
rect 1603 15436 1612 15476
rect 1652 15436 4492 15476
rect 4532 15436 5260 15476
rect 5300 15436 5309 15476
rect 7374 15436 7468 15476
rect 7508 15436 7517 15476
rect 8227 15436 8236 15476
rect 8276 15436 9676 15476
rect 9716 15436 9725 15476
rect 11683 15436 11692 15476
rect 11732 15436 13324 15476
rect 13364 15436 13373 15476
rect 15331 15436 15340 15476
rect 15380 15436 18220 15476
rect 18260 15436 18269 15476
rect 19854 15436 19948 15476
rect 19988 15436 19997 15476
rect 4483 15435 4541 15436
rect 7459 15435 7517 15436
rect 18211 15435 18269 15436
rect 19939 15435 19997 15436
rect 21424 15392 21504 15412
rect 1507 15352 1516 15392
rect 1556 15352 2476 15392
rect 2516 15352 2525 15392
rect 3811 15352 3820 15392
rect 3860 15352 4820 15392
rect 8611 15352 8620 15392
rect 8660 15352 8812 15392
rect 8852 15352 9772 15392
rect 9812 15352 9821 15392
rect 10051 15352 10060 15392
rect 10100 15352 11500 15392
rect 11540 15352 11788 15392
rect 11828 15352 11837 15392
rect 16195 15352 16204 15392
rect 16244 15352 16492 15392
rect 16532 15352 17780 15392
rect 17827 15352 17836 15392
rect 17876 15352 20044 15392
rect 20084 15352 20093 15392
rect 20140 15352 21504 15392
rect 4780 15308 4820 15352
rect 16099 15308 16157 15309
rect 17740 15308 17780 15352
rect 1891 15268 1900 15308
rect 1940 15268 1949 15308
rect 3139 15268 3148 15308
rect 3188 15268 4012 15308
rect 4052 15268 4061 15308
rect 4771 15268 4780 15308
rect 4820 15268 6412 15308
rect 6452 15268 7180 15308
rect 7220 15268 7229 15308
rect 11011 15268 11020 15308
rect 11060 15268 12940 15308
rect 12980 15268 13228 15308
rect 13268 15268 13277 15308
rect 16003 15268 16012 15308
rect 16052 15268 16108 15308
rect 16148 15268 16157 15308
rect 16291 15268 16300 15308
rect 16340 15268 16684 15308
rect 16724 15268 16733 15308
rect 16963 15268 16972 15308
rect 17012 15268 17548 15308
rect 17588 15268 17597 15308
rect 17740 15268 18124 15308
rect 18164 15268 18173 15308
rect 19171 15268 19180 15308
rect 19220 15268 19564 15308
rect 19604 15268 19613 15308
rect 0 15224 80 15244
rect 1900 15224 1940 15268
rect 16099 15267 16157 15268
rect 20140 15224 20180 15352
rect 21424 15332 21504 15352
rect 0 15184 1940 15224
rect 3043 15184 3052 15224
rect 3092 15184 7948 15224
rect 7988 15184 7997 15224
rect 11320 15184 12268 15224
rect 12308 15184 20180 15224
rect 0 15164 80 15184
rect 11320 15140 11360 15184
rect 3052 15100 3244 15140
rect 3284 15100 3293 15140
rect 3679 15100 3688 15140
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 4056 15100 4065 15140
rect 4387 15100 4396 15140
rect 4436 15100 5356 15140
rect 5396 15100 5405 15140
rect 5539 15100 5548 15140
rect 5588 15100 11360 15140
rect 14947 15100 14956 15140
rect 14996 15100 15532 15140
rect 15572 15100 15581 15140
rect 15715 15100 15724 15140
rect 15764 15100 18028 15140
rect 18068 15100 18077 15140
rect 18799 15100 18808 15140
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 19176 15100 19185 15140
rect 3052 15056 3092 15100
rect 12067 15056 12125 15057
rect 15235 15056 15293 15057
rect 3043 15016 3052 15056
rect 3092 15016 3101 15056
rect 4675 15016 4684 15056
rect 4724 15016 9772 15056
rect 9812 15016 12076 15056
rect 12116 15016 12125 15056
rect 15150 15016 15244 15056
rect 15284 15016 15293 15056
rect 12067 15015 12125 15016
rect 15235 15015 15293 15016
rect 16099 15056 16157 15057
rect 21424 15056 21504 15076
rect 16099 15016 16108 15056
rect 16148 15016 21504 15056
rect 16099 15015 16157 15016
rect 21424 14996 21504 15016
rect 4579 14972 4637 14973
rect 4579 14932 4588 14972
rect 4628 14932 6028 14972
rect 6068 14932 8428 14972
rect 8468 14932 8477 14972
rect 9955 14932 9964 14972
rect 10004 14932 13612 14972
rect 13652 14932 16204 14972
rect 16244 14932 16253 14972
rect 18307 14932 18316 14972
rect 18356 14932 19180 14972
rect 19220 14932 19229 14972
rect 4579 14931 4637 14932
rect 0 14888 80 14908
rect 2179 14888 2237 14889
rect 0 14848 2188 14888
rect 2228 14848 2237 14888
rect 4195 14848 4204 14888
rect 4244 14848 6988 14888
rect 7028 14848 8620 14888
rect 8660 14848 8669 14888
rect 14764 14848 18796 14888
rect 18836 14848 18845 14888
rect 0 14828 80 14848
rect 2179 14847 2237 14848
rect 14764 14804 14804 14848
rect 3811 14764 3820 14804
rect 3860 14764 7084 14804
rect 7124 14764 7133 14804
rect 7363 14764 7372 14804
rect 7412 14764 10636 14804
rect 10676 14764 11360 14804
rect 14371 14764 14380 14804
rect 14420 14764 14764 14804
rect 14804 14764 14813 14804
rect 15235 14764 15244 14804
rect 15284 14764 16588 14804
rect 16628 14764 16637 14804
rect 16867 14764 16876 14804
rect 16916 14764 17260 14804
rect 17300 14764 17309 14804
rect 11320 14720 11360 14764
rect 21424 14720 21504 14740
rect 3235 14680 3244 14720
rect 3284 14680 5452 14720
rect 5492 14680 7276 14720
rect 7316 14680 7325 14720
rect 8419 14680 8428 14720
rect 8468 14680 10540 14720
rect 10580 14680 10589 14720
rect 11320 14680 17548 14720
rect 17588 14680 17597 14720
rect 19363 14680 19372 14720
rect 19412 14680 19660 14720
rect 19700 14680 19709 14720
rect 19843 14680 19852 14720
rect 19892 14680 21504 14720
rect 3244 14636 3284 14680
rect 21424 14660 21504 14680
rect 15907 14636 15965 14637
rect 2467 14596 2476 14636
rect 2516 14596 3284 14636
rect 15619 14596 15628 14636
rect 15668 14596 15916 14636
rect 15956 14596 15965 14636
rect 15907 14595 15965 14596
rect 0 14552 80 14572
rect 1219 14552 1277 14553
rect 5539 14552 5597 14553
rect 8803 14552 8861 14553
rect 0 14512 1228 14552
rect 1268 14512 1277 14552
rect 2275 14512 2284 14552
rect 2324 14512 4684 14552
rect 4724 14512 4733 14552
rect 5539 14512 5548 14552
rect 5588 14512 8756 14552
rect 0 14492 80 14512
rect 1219 14511 1277 14512
rect 5539 14511 5597 14512
rect 8611 14468 8669 14469
rect 1699 14428 1708 14468
rect 1748 14428 8620 14468
rect 8660 14428 8669 14468
rect 8716 14468 8756 14512
rect 8803 14512 8812 14552
rect 8852 14512 17068 14552
rect 17108 14512 17117 14552
rect 18403 14512 18412 14552
rect 18452 14512 18988 14552
rect 19028 14512 19037 14552
rect 8803 14511 8861 14512
rect 14659 14468 14717 14469
rect 8716 14428 11308 14468
rect 11348 14428 12844 14468
rect 12884 14428 12893 14468
rect 14659 14428 14668 14468
rect 14708 14428 14956 14468
rect 14996 14428 20564 14468
rect 8611 14427 8669 14428
rect 14659 14427 14717 14428
rect 20524 14384 20564 14428
rect 21424 14384 21504 14404
rect 4919 14344 4928 14384
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 5296 14344 5305 14384
rect 6979 14344 6988 14384
rect 7028 14344 14188 14384
rect 14228 14344 14237 14384
rect 20039 14344 20048 14384
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20416 14344 20425 14384
rect 20524 14344 21504 14384
rect 21424 14324 21504 14344
rect 6307 14260 6316 14300
rect 6356 14260 19660 14300
rect 19700 14260 20180 14300
rect 0 14216 80 14236
rect 6691 14216 6749 14217
rect 15715 14216 15773 14217
rect 0 14176 1804 14216
rect 1844 14176 1853 14216
rect 2659 14176 2668 14216
rect 2708 14176 4108 14216
rect 4148 14176 4157 14216
rect 6606 14176 6700 14216
rect 6740 14176 6749 14216
rect 8035 14176 8044 14216
rect 8084 14176 8428 14216
rect 8468 14176 8477 14216
rect 13027 14176 13036 14216
rect 13076 14176 13228 14216
rect 13268 14176 13277 14216
rect 13795 14176 13804 14216
rect 13844 14176 15724 14216
rect 15764 14176 20044 14216
rect 20084 14176 20093 14216
rect 0 14156 80 14176
rect 6691 14175 6749 14176
rect 15715 14175 15773 14176
rect 4579 14132 4637 14133
rect 20140 14132 20180 14260
rect 3235 14092 3244 14132
rect 3284 14092 4588 14132
rect 4628 14092 4637 14132
rect 9091 14092 9100 14132
rect 9140 14092 11828 14132
rect 11875 14092 11884 14132
rect 11924 14092 12940 14132
rect 12980 14092 12989 14132
rect 20140 14092 20276 14132
rect 4579 14091 4637 14092
rect 3523 14048 3581 14049
rect 11788 14048 11828 14092
rect 17251 14048 17309 14049
rect 20236 14048 20276 14092
rect 21424 14048 21504 14068
rect 3438 14008 3532 14048
rect 3572 14008 3581 14048
rect 6403 14008 6412 14048
rect 6452 14008 6796 14048
rect 6836 14008 6845 14048
rect 8323 14008 8332 14048
rect 8372 14008 8524 14048
rect 8564 14008 8716 14048
rect 8756 14008 8765 14048
rect 10915 14008 10924 14048
rect 10964 14008 11212 14048
rect 11252 14008 11261 14048
rect 11788 14008 13324 14048
rect 13364 14008 13373 14048
rect 15331 14008 15340 14048
rect 15380 14008 16012 14048
rect 16052 14008 16061 14048
rect 16579 14008 16588 14048
rect 16628 14008 16972 14048
rect 17012 14008 17021 14048
rect 17251 14008 17260 14048
rect 17300 14008 18700 14048
rect 18740 14008 18988 14048
rect 19028 14008 19037 14048
rect 20236 14008 21504 14048
rect 3523 14007 3581 14008
rect 17251 14007 17309 14008
rect 21424 13988 21504 14008
rect 3331 13964 3389 13965
rect 2851 13924 2860 13964
rect 2900 13924 3340 13964
rect 3380 13924 4012 13964
rect 4052 13924 4061 13964
rect 18595 13924 18604 13964
rect 18644 13924 18796 13964
rect 18836 13924 20084 13964
rect 3331 13923 3389 13924
rect 0 13880 80 13900
rect 0 13840 3628 13880
rect 3668 13840 3677 13880
rect 0 13820 80 13840
rect 4012 13796 4052 13924
rect 5731 13880 5789 13881
rect 14659 13880 14717 13881
rect 5731 13840 5740 13880
rect 5780 13840 6508 13880
rect 6548 13840 6557 13880
rect 6796 13840 7372 13880
rect 7412 13840 7421 13880
rect 11683 13840 11692 13880
rect 11732 13840 14668 13880
rect 14708 13840 14717 13880
rect 5731 13839 5789 13840
rect 5347 13796 5405 13797
rect 5635 13796 5693 13797
rect 6796 13796 6836 13840
rect 14659 13839 14717 13840
rect 15619 13880 15677 13881
rect 20044 13880 20084 13924
rect 15619 13840 15628 13880
rect 15668 13840 16492 13880
rect 16532 13840 16541 13880
rect 18883 13840 18892 13880
rect 18932 13840 19276 13880
rect 19316 13840 19325 13880
rect 20035 13840 20044 13880
rect 20084 13840 20093 13880
rect 15619 13839 15677 13840
rect 4012 13756 5300 13796
rect 5260 13712 5300 13756
rect 5347 13756 5356 13796
rect 5396 13756 5644 13796
rect 5684 13756 5693 13796
rect 6787 13756 6796 13796
rect 6836 13756 6845 13796
rect 11299 13756 11308 13796
rect 11348 13756 12076 13796
rect 12116 13756 12125 13796
rect 13219 13756 13228 13796
rect 13268 13756 13804 13796
rect 13844 13756 13853 13796
rect 5347 13755 5405 13756
rect 5635 13755 5693 13756
rect 21424 13712 21504 13732
rect 1027 13672 1036 13712
rect 1076 13672 4396 13712
rect 4436 13672 4445 13712
rect 5260 13672 6508 13712
rect 6548 13672 6557 13712
rect 8899 13672 8908 13712
rect 8948 13672 18412 13712
rect 18452 13672 21504 13712
rect 21424 13652 21504 13672
rect 2083 13588 2092 13628
rect 2132 13588 2380 13628
rect 2420 13588 2429 13628
rect 3679 13588 3688 13628
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 4056 13588 4065 13628
rect 8611 13588 8620 13628
rect 8660 13588 8812 13628
rect 8852 13588 8861 13628
rect 18799 13588 18808 13628
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 19176 13588 19185 13628
rect 0 13544 80 13564
rect 15331 13544 15389 13545
rect 0 13504 12172 13544
rect 12212 13504 12221 13544
rect 15139 13504 15148 13544
rect 15188 13504 15340 13544
rect 15380 13504 15389 13544
rect 0 13484 80 13504
rect 15331 13503 15389 13504
rect 2179 13460 2237 13461
rect 15523 13460 15581 13461
rect 2179 13420 2188 13460
rect 2228 13420 13996 13460
rect 14036 13420 14045 13460
rect 15438 13420 15532 13460
rect 15572 13420 15581 13460
rect 15715 13420 15724 13460
rect 15764 13420 16204 13460
rect 16244 13420 16588 13460
rect 16628 13420 16637 13460
rect 2179 13419 2237 13420
rect 15523 13419 15581 13420
rect 21424 13376 21504 13396
rect 2755 13336 2764 13376
rect 2804 13336 3436 13376
rect 3476 13336 3485 13376
rect 5923 13336 5932 13376
rect 5972 13336 6700 13376
rect 6740 13336 6749 13376
rect 9091 13336 9100 13376
rect 9140 13336 9484 13376
rect 9524 13336 9533 13376
rect 12652 13336 13324 13376
rect 13364 13336 21504 13376
rect 12652 13292 12692 13336
rect 21424 13316 21504 13336
rect 15235 13292 15293 13293
rect 16771 13292 16829 13293
rect 1603 13252 1612 13292
rect 1652 13252 10348 13292
rect 10388 13252 10397 13292
rect 12643 13252 12652 13292
rect 12692 13252 12701 13292
rect 15235 13252 15244 13292
rect 15284 13252 15724 13292
rect 15764 13252 15773 13292
rect 16483 13252 16492 13292
rect 16532 13252 16780 13292
rect 16820 13252 16829 13292
rect 17731 13252 17740 13292
rect 17780 13252 18124 13292
rect 18164 13252 18173 13292
rect 15235 13251 15293 13252
rect 16771 13251 16829 13252
rect 0 13208 80 13228
rect 5635 13208 5693 13209
rect 16099 13208 16157 13209
rect 0 13168 788 13208
rect 835 13168 844 13208
rect 884 13168 1420 13208
rect 1460 13168 1469 13208
rect 5635 13168 5644 13208
rect 5684 13168 7468 13208
rect 7508 13168 7517 13208
rect 7747 13168 7756 13208
rect 7796 13168 8236 13208
rect 8276 13168 8285 13208
rect 10723 13168 10732 13208
rect 10772 13168 12364 13208
rect 12404 13168 12413 13208
rect 12739 13168 12748 13208
rect 12788 13168 14380 13208
rect 14420 13168 15244 13208
rect 15284 13168 15820 13208
rect 15860 13168 15869 13208
rect 16014 13168 16108 13208
rect 16148 13168 16157 13208
rect 0 13148 80 13168
rect 748 12956 788 13168
rect 5635 13167 5693 13168
rect 16099 13167 16157 13168
rect 1987 13084 1996 13124
rect 2036 13084 7180 13124
rect 7220 13084 7229 13124
rect 17059 13084 17068 13124
rect 17108 13084 18124 13124
rect 18164 13084 18316 13124
rect 18356 13084 18365 13124
rect 1411 13040 1469 13041
rect 1326 13000 1420 13040
rect 1460 13000 1469 13040
rect 1411 12999 1469 13000
rect 2500 13000 17932 13040
rect 17972 13000 17981 13040
rect 2500 12956 2540 13000
rect 3331 12956 3389 12957
rect 748 12916 2540 12956
rect 2947 12916 2956 12956
rect 2996 12916 3340 12956
rect 3380 12916 3389 12956
rect 4195 12916 4204 12956
rect 4244 12916 7276 12956
rect 7316 12916 7325 12956
rect 10627 12916 10636 12956
rect 10676 12916 11116 12956
rect 11156 12916 11165 12956
rect 18019 12916 18028 12956
rect 18068 12916 18412 12956
rect 18452 12916 18461 12956
rect 3331 12915 3389 12916
rect 0 12872 80 12892
rect 0 12832 2036 12872
rect 2755 12832 2764 12872
rect 2804 12832 3244 12872
rect 3284 12832 3293 12872
rect 4003 12832 4012 12872
rect 4052 12832 4820 12872
rect 4919 12832 4928 12872
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 5296 12832 5305 12872
rect 5731 12832 5740 12872
rect 5780 12832 6124 12872
rect 6164 12832 9100 12872
rect 9140 12832 9149 12872
rect 14275 12832 14284 12872
rect 14324 12832 14764 12872
rect 14804 12832 18796 12872
rect 18836 12832 18845 12872
rect 20039 12832 20048 12872
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20416 12832 20425 12872
rect 0 12812 80 12832
rect 1996 12704 2036 12832
rect 2083 12788 2141 12789
rect 4780 12788 4820 12832
rect 6019 12788 6077 12789
rect 2083 12748 2092 12788
rect 2132 12748 4684 12788
rect 4724 12748 4733 12788
rect 4780 12748 6028 12788
rect 6068 12748 6077 12788
rect 7939 12748 7948 12788
rect 7988 12748 9580 12788
rect 9620 12748 14092 12788
rect 14132 12748 14141 12788
rect 2083 12747 2141 12748
rect 6019 12747 6077 12748
rect 1996 12664 10444 12704
rect 10484 12664 10493 12704
rect 15811 12664 15820 12704
rect 15860 12664 17548 12704
rect 17588 12664 17597 12704
rect 2467 12620 2525 12621
rect 16099 12620 16157 12621
rect 2382 12580 2476 12620
rect 2516 12580 2525 12620
rect 5251 12580 5260 12620
rect 5300 12580 5932 12620
rect 5972 12580 8044 12620
rect 8084 12580 8093 12620
rect 8707 12580 8716 12620
rect 8756 12580 10060 12620
rect 10100 12580 10732 12620
rect 10772 12580 10781 12620
rect 16099 12580 16108 12620
rect 16148 12580 18796 12620
rect 18836 12580 19276 12620
rect 19316 12580 19325 12620
rect 2467 12579 2525 12580
rect 16099 12579 16157 12580
rect 0 12536 80 12556
rect 15043 12536 15101 12537
rect 16291 12536 16349 12537
rect 19363 12536 19421 12537
rect 19939 12536 19997 12537
rect 0 12496 11116 12536
rect 11156 12496 11165 12536
rect 11491 12496 11500 12536
rect 11540 12496 12844 12536
rect 12884 12496 12893 12536
rect 14563 12496 14572 12536
rect 14612 12496 15052 12536
rect 15092 12496 15101 12536
rect 16206 12496 16300 12536
rect 16340 12496 16349 12536
rect 16963 12496 16972 12536
rect 17012 12496 17452 12536
rect 17492 12496 17501 12536
rect 19363 12496 19372 12536
rect 19412 12496 19948 12536
rect 19988 12496 20044 12536
rect 20084 12496 20093 12536
rect 0 12476 80 12496
rect 15043 12495 15101 12496
rect 16291 12495 16349 12496
rect 19363 12495 19421 12496
rect 19939 12495 19997 12496
rect 1699 12412 1708 12452
rect 1748 12412 1757 12452
rect 2083 12412 2092 12452
rect 2132 12412 16340 12452
rect 1708 12368 1748 12412
rect 16300 12368 16340 12412
rect 1708 12328 8908 12368
rect 8948 12328 8957 12368
rect 10540 12328 11596 12368
rect 11636 12328 11645 12368
rect 11779 12328 11788 12368
rect 11828 12328 12748 12368
rect 12788 12328 12797 12368
rect 16291 12328 16300 12368
rect 16340 12328 16349 12368
rect 2275 12284 2333 12285
rect 10540 12284 10580 12328
rect 1795 12244 1804 12284
rect 1844 12244 2284 12284
rect 2324 12244 2333 12284
rect 3331 12244 3340 12284
rect 3380 12244 3820 12284
rect 3860 12244 3869 12284
rect 4003 12244 4012 12284
rect 4052 12244 4492 12284
rect 4532 12244 8716 12284
rect 8756 12244 8765 12284
rect 10531 12244 10540 12284
rect 10580 12244 10589 12284
rect 2275 12243 2333 12244
rect 0 12200 80 12220
rect 0 12160 11596 12200
rect 11636 12160 11645 12200
rect 0 12140 80 12160
rect 2083 12116 2141 12117
rect 4675 12116 4733 12117
rect 1998 12076 2092 12116
rect 2132 12076 2141 12116
rect 2755 12076 2764 12116
rect 2804 12076 3148 12116
rect 3188 12076 3197 12116
rect 3679 12076 3688 12116
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 4056 12076 4065 12116
rect 4590 12076 4684 12116
rect 4724 12076 14764 12116
rect 14804 12076 14813 12116
rect 18799 12076 18808 12116
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 19176 12076 19185 12116
rect 2083 12075 2141 12076
rect 4675 12075 4733 12076
rect 8323 12032 8381 12033
rect 2179 11992 2188 12032
rect 2228 11992 2476 12032
rect 2516 11992 2525 12032
rect 8323 11992 8332 12032
rect 8372 11992 14572 12032
rect 14612 11992 14621 12032
rect 18307 11992 18316 12032
rect 18356 11992 18700 12032
rect 18740 11992 18749 12032
rect 8323 11991 8381 11992
rect 3139 11948 3197 11949
rect 3139 11908 3148 11948
rect 3188 11908 9484 11948
rect 9524 11908 9533 11948
rect 10435 11908 10444 11948
rect 10484 11908 19564 11948
rect 19604 11908 19613 11948
rect 3139 11907 3197 11908
rect 0 11864 80 11884
rect 6211 11864 6269 11865
rect 6883 11864 6941 11865
rect 14947 11864 15005 11865
rect 0 11824 1900 11864
rect 1940 11824 1949 11864
rect 2467 11824 2476 11864
rect 2516 11824 4204 11864
rect 4244 11824 4253 11864
rect 6211 11824 6220 11864
rect 6260 11824 6892 11864
rect 6932 11824 6941 11864
rect 8131 11824 8140 11864
rect 8180 11824 8716 11864
rect 8756 11824 8765 11864
rect 14947 11824 14956 11864
rect 14996 11824 15052 11864
rect 15092 11824 15101 11864
rect 0 11804 80 11824
rect 6211 11823 6269 11824
rect 6883 11823 6941 11824
rect 14947 11823 15005 11824
rect 3043 11740 3052 11780
rect 3092 11740 7564 11780
rect 7604 11740 7613 11780
rect 11011 11740 11020 11780
rect 11060 11740 11212 11780
rect 11252 11740 15244 11780
rect 15284 11740 15628 11780
rect 15668 11740 15677 11780
rect 4099 11696 4157 11697
rect 2956 11656 3244 11696
rect 3284 11656 3293 11696
rect 4014 11656 4108 11696
rect 4148 11656 4157 11696
rect 5923 11656 5932 11696
rect 5972 11656 6124 11696
rect 6164 11656 6173 11696
rect 6307 11656 6316 11696
rect 6356 11656 7852 11696
rect 7892 11656 7901 11696
rect 8131 11656 8140 11696
rect 8180 11656 8620 11696
rect 8660 11656 8669 11696
rect 9187 11656 9196 11696
rect 9236 11656 10540 11696
rect 10580 11656 10589 11696
rect 11320 11656 17260 11696
rect 17300 11656 17309 11696
rect 17923 11656 17932 11696
rect 17972 11656 18508 11696
rect 18548 11656 19468 11696
rect 19508 11656 19852 11696
rect 19892 11656 19901 11696
rect 2179 11612 2237 11613
rect 2179 11572 2188 11612
rect 2228 11572 2572 11612
rect 2612 11572 2621 11612
rect 2179 11571 2237 11572
rect 0 11528 80 11548
rect 0 11488 2860 11528
rect 2900 11488 2909 11528
rect 0 11468 80 11488
rect 2467 11444 2525 11445
rect 2956 11444 2996 11656
rect 4099 11655 4157 11656
rect 3043 11612 3101 11613
rect 11320 11612 11360 11656
rect 12931 11612 12989 11613
rect 3043 11572 3052 11612
rect 3092 11572 3668 11612
rect 7747 11572 7756 11612
rect 7796 11572 11360 11612
rect 12643 11572 12652 11612
rect 12692 11572 12940 11612
rect 12980 11572 12989 11612
rect 3043 11571 3101 11572
rect 3628 11528 3668 11572
rect 12931 11571 12989 11572
rect 3619 11488 3628 11528
rect 3668 11488 3677 11528
rect 14275 11488 14284 11528
rect 14324 11488 14476 11528
rect 14516 11488 14525 11528
rect 2382 11404 2476 11444
rect 2516 11404 2525 11444
rect 2467 11403 2525 11404
rect 2572 11404 2996 11444
rect 6883 11404 6892 11444
rect 6932 11404 8044 11444
rect 8084 11404 9868 11444
rect 9908 11404 11788 11444
rect 11828 11404 11837 11444
rect 13699 11404 13708 11444
rect 13748 11404 17164 11444
rect 17204 11404 17300 11444
rect 835 11276 893 11277
rect 2572 11276 2612 11404
rect 4919 11320 4928 11360
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 5296 11320 5305 11360
rect 16387 11276 16445 11277
rect 17260 11276 17300 11404
rect 20039 11320 20048 11360
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20416 11320 20425 11360
rect 835 11236 844 11276
rect 884 11236 2612 11276
rect 5923 11236 5932 11276
rect 5972 11236 16396 11276
rect 16436 11236 16445 11276
rect 17155 11236 17164 11276
rect 17204 11236 17300 11276
rect 835 11235 893 11236
rect 16387 11235 16445 11236
rect 0 11192 80 11212
rect 6019 11192 6077 11193
rect 0 11152 1900 11192
rect 1940 11152 1949 11192
rect 2179 11152 2188 11192
rect 2228 11152 4012 11192
rect 4052 11152 4061 11192
rect 5635 11152 5644 11192
rect 5684 11152 6028 11192
rect 6068 11152 6077 11192
rect 11971 11152 11980 11192
rect 12020 11152 12364 11192
rect 12404 11152 12413 11192
rect 14467 11152 14476 11192
rect 14516 11152 14668 11192
rect 14708 11152 14717 11192
rect 16291 11152 16300 11192
rect 16340 11152 18604 11192
rect 18644 11152 18653 11192
rect 0 11132 80 11152
rect 6019 11151 6077 11152
rect 1699 11068 1708 11108
rect 1748 11068 7180 11108
rect 7220 11068 7229 11108
rect 4195 11024 4253 11025
rect 15811 11024 15869 11025
rect 16771 11024 16829 11025
rect 2563 10984 2572 11024
rect 2612 10984 2956 11024
rect 2996 10984 3005 11024
rect 3811 10984 3820 11024
rect 3860 10984 4204 11024
rect 4244 10984 4253 11024
rect 4302 10984 4311 11024
rect 4351 10984 5204 11024
rect 5251 10984 5260 11024
rect 5300 10984 5548 11024
rect 5588 10984 5597 11024
rect 8035 10984 8044 11024
rect 8084 10984 8524 11024
rect 8564 10984 8573 11024
rect 15726 10984 15820 11024
rect 15860 10984 15869 11024
rect 16686 10984 16780 11024
rect 16820 10984 19276 11024
rect 19316 10984 19325 11024
rect 4195 10983 4253 10984
rect 4867 10940 4925 10941
rect 4195 10900 4204 10940
rect 4244 10900 4492 10940
rect 4532 10900 4541 10940
rect 4782 10900 4876 10940
rect 4916 10900 4925 10940
rect 5164 10940 5204 10984
rect 15811 10983 15869 10984
rect 16771 10983 16829 10984
rect 16099 10940 16157 10941
rect 5164 10900 7468 10940
rect 7508 10900 7517 10940
rect 10531 10900 10540 10940
rect 10580 10900 10828 10940
rect 10868 10900 10877 10940
rect 16099 10900 16108 10940
rect 16148 10900 16204 10940
rect 16244 10900 16253 10940
rect 4867 10899 4925 10900
rect 16099 10899 16157 10900
rect 0 10856 80 10876
rect 0 10816 14476 10856
rect 14516 10816 14525 10856
rect 0 10796 80 10816
rect 3523 10772 3581 10773
rect 15619 10772 15677 10773
rect 3523 10732 3532 10772
rect 3572 10732 4492 10772
rect 4532 10732 4541 10772
rect 4675 10732 4684 10772
rect 4724 10732 15628 10772
rect 15668 10732 15677 10772
rect 3523 10731 3581 10732
rect 15619 10731 15677 10732
rect 163 10648 172 10688
rect 212 10648 5164 10688
rect 5204 10648 5213 10688
rect 6499 10648 6508 10688
rect 6548 10648 8428 10688
rect 8468 10648 8477 10688
rect 13027 10648 13036 10688
rect 13076 10648 13228 10688
rect 13268 10648 20180 10688
rect 3235 10604 3293 10605
rect 4195 10604 4253 10605
rect 3043 10564 3052 10604
rect 3092 10564 3244 10604
rect 3284 10564 3293 10604
rect 3679 10564 3688 10604
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 4056 10564 4065 10604
rect 4195 10564 4204 10604
rect 4244 10564 4396 10604
rect 4436 10564 4445 10604
rect 8515 10564 8524 10604
rect 8564 10564 18700 10604
rect 18740 10564 18749 10604
rect 18799 10564 18808 10604
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 19176 10564 19185 10604
rect 3235 10563 3293 10564
rect 4195 10563 4253 10564
rect 0 10520 80 10540
rect 5347 10520 5405 10521
rect 20140 10520 20180 10648
rect 20611 10520 20669 10521
rect 0 10480 2188 10520
rect 2228 10480 2237 10520
rect 4579 10480 4588 10520
rect 4628 10480 4972 10520
rect 5012 10480 5021 10520
rect 5347 10480 5356 10520
rect 5396 10480 5644 10520
rect 5684 10480 6220 10520
rect 6260 10480 6269 10520
rect 15907 10480 15916 10520
rect 15956 10480 17452 10520
rect 17492 10480 17501 10520
rect 18595 10480 18604 10520
rect 18644 10480 18836 10520
rect 20140 10480 20620 10520
rect 20660 10480 20669 10520
rect 0 10460 80 10480
rect 5347 10479 5405 10480
rect 18796 10436 18836 10480
rect 20611 10479 20669 10480
rect 1987 10396 1996 10436
rect 2036 10396 2668 10436
rect 2708 10396 2717 10436
rect 3523 10396 3532 10436
rect 3572 10396 3820 10436
rect 3860 10396 6508 10436
rect 6548 10396 6557 10436
rect 12547 10396 12556 10436
rect 12596 10396 12748 10436
rect 12788 10396 12797 10436
rect 17251 10396 17260 10436
rect 17300 10396 17836 10436
rect 17876 10396 17885 10436
rect 18211 10396 18220 10436
rect 18260 10396 18412 10436
rect 18452 10396 18461 10436
rect 18787 10396 18796 10436
rect 18836 10396 18845 10436
rect 1315 10352 1373 10353
rect 1315 10312 1324 10352
rect 1364 10312 2860 10352
rect 2900 10312 2909 10352
rect 3427 10312 3436 10352
rect 3476 10312 6316 10352
rect 6356 10312 6365 10352
rect 10531 10312 10540 10352
rect 10580 10312 17164 10352
rect 17204 10312 17213 10352
rect 18019 10312 18028 10352
rect 18068 10312 18604 10352
rect 18644 10312 18653 10352
rect 1315 10311 1373 10312
rect 14467 10268 14525 10269
rect 16099 10268 16157 10269
rect 3043 10228 3052 10268
rect 3092 10228 13420 10268
rect 13460 10228 13469 10268
rect 13891 10228 13900 10268
rect 13940 10228 14284 10268
rect 14324 10228 14333 10268
rect 14467 10228 14476 10268
rect 14516 10228 14764 10268
rect 14804 10228 14813 10268
rect 16099 10228 16108 10268
rect 16148 10228 18700 10268
rect 18740 10228 18749 10268
rect 14467 10227 14525 10228
rect 16099 10227 16157 10228
rect 0 10184 80 10204
rect 3139 10184 3197 10185
rect 0 10144 1516 10184
rect 1556 10144 1565 10184
rect 2500 10144 3148 10184
rect 3188 10144 3572 10184
rect 3715 10144 3724 10184
rect 3764 10144 6164 10184
rect 6211 10144 6220 10184
rect 6260 10144 16396 10184
rect 16436 10144 16972 10184
rect 17012 10144 17021 10184
rect 17068 10144 18316 10184
rect 18356 10144 18365 10184
rect 0 10124 80 10144
rect 2500 10100 2540 10144
rect 3139 10143 3197 10144
rect 3532 10100 3572 10144
rect 4291 10100 4349 10101
rect 6124 10100 6164 10144
rect 15811 10100 15869 10101
rect 17068 10100 17108 10144
rect 1516 10060 2540 10100
rect 3523 10060 3532 10100
rect 3572 10060 3581 10100
rect 4291 10060 4300 10100
rect 4340 10060 4684 10100
rect 4724 10060 4733 10100
rect 6115 10060 6124 10100
rect 6164 10060 7468 10100
rect 7508 10060 7517 10100
rect 11587 10060 11596 10100
rect 11636 10060 13516 10100
rect 13556 10060 13565 10100
rect 14275 10060 14284 10100
rect 14324 10060 15764 10100
rect 1516 10016 1556 10060
rect 4291 10059 4349 10060
rect 3331 10016 3389 10017
rect 14947 10016 15005 10017
rect 1507 9976 1516 10016
rect 1556 9976 1565 10016
rect 3331 9976 3340 10016
rect 3380 9976 3436 10016
rect 3476 9976 3485 10016
rect 4291 9976 4300 10016
rect 4340 9976 4780 10016
rect 4820 9976 4829 10016
rect 5059 9976 5068 10016
rect 5108 9976 6220 10016
rect 6260 9976 6269 10016
rect 6403 9976 6412 10016
rect 6452 9976 7276 10016
rect 7316 9976 7325 10016
rect 8803 9976 8812 10016
rect 8852 9976 9100 10016
rect 9140 9976 9149 10016
rect 11395 9976 11404 10016
rect 11444 9976 11788 10016
rect 11828 9976 11837 10016
rect 11971 9976 11980 10016
rect 12020 9976 12652 10016
rect 12692 9976 12701 10016
rect 14862 9976 14956 10016
rect 14996 9976 15005 10016
rect 15724 10016 15764 10060
rect 15811 10060 15820 10100
rect 15860 10060 17108 10100
rect 17155 10060 17164 10100
rect 17204 10060 19948 10100
rect 19988 10060 19997 10100
rect 15811 10059 15869 10060
rect 15724 9976 16012 10016
rect 16052 9976 16204 10016
rect 16244 9976 16253 10016
rect 3331 9975 3389 9976
rect 14947 9975 15005 9976
rect 2755 9932 2813 9933
rect 16195 9932 16253 9933
rect 1315 9892 1324 9932
rect 1364 9892 2764 9932
rect 2804 9892 2813 9932
rect 8899 9892 8908 9932
rect 8948 9892 16204 9932
rect 16244 9892 16253 9932
rect 17731 9892 17740 9932
rect 17780 9892 17932 9932
rect 17972 9892 17981 9932
rect 2755 9891 2813 9892
rect 16195 9891 16253 9892
rect 0 9848 80 9868
rect 12451 9848 12509 9849
rect 0 9808 1420 9848
rect 1460 9808 1469 9848
rect 2563 9808 2572 9848
rect 2612 9808 2764 9848
rect 2804 9808 2813 9848
rect 4919 9808 4928 9848
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 5296 9808 5305 9848
rect 12451 9808 12460 9848
rect 12500 9808 12556 9848
rect 12596 9808 12605 9848
rect 20039 9808 20048 9848
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20416 9808 20425 9848
rect 0 9788 80 9808
rect 12451 9807 12509 9808
rect 3139 9764 3197 9765
rect 4099 9764 4157 9765
rect 3139 9724 3148 9764
rect 3188 9724 4108 9764
rect 4148 9724 11360 9764
rect 19363 9724 19372 9764
rect 19412 9724 19948 9764
rect 19988 9724 19997 9764
rect 3139 9723 3197 9724
rect 4099 9723 4157 9724
rect 2275 9680 2333 9681
rect 11320 9680 11360 9724
rect 2190 9640 2284 9680
rect 2324 9640 2333 9680
rect 2755 9640 2764 9680
rect 2804 9640 3724 9680
rect 3764 9640 3773 9680
rect 7075 9640 7084 9680
rect 7124 9640 7372 9680
rect 7412 9640 7421 9680
rect 10147 9640 10156 9680
rect 10196 9640 11020 9680
rect 11060 9640 11069 9680
rect 11320 9640 14380 9680
rect 14420 9640 16492 9680
rect 16532 9640 16541 9680
rect 17923 9640 17932 9680
rect 17972 9640 18220 9680
rect 18260 9640 18269 9680
rect 2275 9639 2333 9640
rect 3235 9596 3293 9597
rect 3139 9556 3148 9596
rect 3188 9556 3244 9596
rect 3284 9556 5932 9596
rect 5972 9556 5981 9596
rect 11491 9556 11500 9596
rect 11540 9556 11884 9596
rect 11924 9556 11933 9596
rect 3235 9555 3293 9556
rect 0 9512 80 9532
rect 3331 9512 3389 9513
rect 5635 9512 5693 9513
rect 12067 9512 12125 9513
rect 0 9472 3052 9512
rect 3092 9472 3101 9512
rect 3331 9472 3340 9512
rect 3380 9472 3724 9512
rect 3764 9472 3773 9512
rect 4195 9472 4204 9512
rect 4244 9472 4396 9512
rect 4436 9472 4445 9512
rect 5550 9472 5644 9512
rect 5684 9472 6124 9512
rect 6164 9472 6173 9512
rect 6883 9472 6892 9512
rect 6932 9472 7084 9512
rect 7124 9472 7133 9512
rect 11982 9472 12076 9512
rect 12116 9472 12268 9512
rect 12308 9472 12317 9512
rect 12835 9472 12844 9512
rect 12884 9472 13324 9512
rect 13364 9472 13373 9512
rect 15619 9472 15628 9512
rect 15668 9472 17836 9512
rect 17876 9472 17885 9512
rect 19267 9472 19276 9512
rect 19316 9472 19660 9512
rect 19700 9472 19709 9512
rect 0 9452 80 9472
rect 3331 9471 3389 9472
rect 5635 9471 5693 9472
rect 12067 9471 12125 9472
rect 1603 9388 1612 9428
rect 1652 9388 1804 9428
rect 1844 9388 1853 9428
rect 1987 9388 1996 9428
rect 2036 9388 9908 9428
rect 2179 9344 2237 9345
rect 9868 9344 9908 9388
rect 2179 9304 2188 9344
rect 2228 9304 2764 9344
rect 2804 9304 2813 9344
rect 6883 9304 6892 9344
rect 6932 9304 7276 9344
rect 7316 9304 7756 9344
rect 7796 9304 7805 9344
rect 9859 9304 9868 9344
rect 9908 9304 9917 9344
rect 2179 9303 2237 9304
rect 4099 9260 4157 9261
rect 4099 9220 4108 9260
rect 4148 9220 4972 9260
rect 5012 9220 5021 9260
rect 8515 9220 8524 9260
rect 8564 9220 10060 9260
rect 10100 9220 10348 9260
rect 10388 9220 11500 9260
rect 11540 9220 19276 9260
rect 19316 9220 19325 9260
rect 4099 9219 4157 9220
rect 0 9176 80 9196
rect 2851 9176 2909 9177
rect 0 9136 1900 9176
rect 1940 9136 1949 9176
rect 2851 9136 2860 9176
rect 2900 9136 6796 9176
rect 6836 9136 6845 9176
rect 9091 9136 9100 9176
rect 9140 9136 11360 9176
rect 14851 9136 14860 9176
rect 14900 9136 18028 9176
rect 18068 9136 18077 9176
rect 0 9116 80 9136
rect 2851 9135 2909 9136
rect 11320 9092 11360 9136
rect 2659 9052 2668 9092
rect 2708 9052 3532 9092
rect 3572 9052 3581 9092
rect 3679 9052 3688 9092
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 4056 9052 4065 9092
rect 6211 9052 6220 9092
rect 6260 9052 8812 9092
rect 8852 9052 8861 9092
rect 11320 9052 16492 9092
rect 16532 9052 16541 9092
rect 18799 9052 18808 9092
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 19176 9052 19185 9092
rect 2371 8968 2380 9008
rect 2420 8968 16396 9008
rect 16436 8968 16445 9008
rect 3331 8924 3389 8925
rect 4579 8924 4637 8925
rect 15427 8924 15485 8925
rect 3331 8884 3340 8924
rect 3380 8884 3628 8924
rect 3668 8884 3677 8924
rect 4494 8884 4588 8924
rect 4628 8884 4637 8924
rect 5155 8884 5164 8924
rect 5204 8884 10348 8924
rect 10388 8884 10397 8924
rect 15427 8884 15436 8924
rect 15476 8884 18508 8924
rect 18548 8884 18557 8924
rect 3331 8883 3389 8884
rect 4579 8883 4637 8884
rect 15427 8883 15485 8884
rect 0 8840 80 8860
rect 17644 8841 17684 8884
rect 6211 8840 6269 8841
rect 17635 8840 17693 8841
rect 18403 8840 18461 8841
rect 0 8800 3244 8840
rect 3284 8800 3293 8840
rect 4099 8800 4108 8840
rect 4148 8800 4157 8840
rect 4291 8800 4300 8840
rect 4340 8800 5452 8840
rect 5492 8800 5501 8840
rect 6126 8800 6220 8840
rect 6260 8800 6269 8840
rect 7075 8800 7084 8840
rect 7124 8800 8620 8840
rect 8660 8800 8840 8840
rect 12643 8800 12652 8840
rect 12692 8800 17356 8840
rect 17396 8800 17405 8840
rect 17635 8800 17644 8840
rect 17684 8800 17724 8840
rect 18318 8800 18412 8840
rect 18452 8800 18461 8840
rect 0 8780 80 8800
rect 4108 8756 4148 8800
rect 6211 8799 6269 8800
rect 4195 8756 4253 8757
rect 8800 8756 8840 8800
rect 1123 8716 1132 8756
rect 1172 8716 3820 8756
rect 3860 8716 3869 8756
rect 4108 8716 4204 8756
rect 4244 8716 4253 8756
rect 4579 8716 4588 8756
rect 4628 8716 4876 8756
rect 4916 8716 4925 8756
rect 5635 8716 5644 8756
rect 5684 8716 5932 8756
rect 5972 8716 5981 8756
rect 8800 8716 9620 8756
rect 10915 8716 10924 8756
rect 10964 8716 12940 8756
rect 12980 8716 12989 8756
rect 4195 8715 4253 8716
rect 2851 8672 2909 8673
rect 3235 8672 3293 8673
rect 2766 8632 2860 8672
rect 2900 8632 2909 8672
rect 3043 8632 3052 8672
rect 3092 8632 3244 8672
rect 3284 8632 3293 8672
rect 2851 8631 2909 8632
rect 3235 8631 3293 8632
rect 4387 8672 4445 8673
rect 9580 8672 9620 8716
rect 12067 8672 12125 8673
rect 12835 8672 12893 8673
rect 13420 8672 13460 8800
rect 17635 8799 17693 8800
rect 18403 8799 18461 8800
rect 18595 8840 18653 8841
rect 18595 8800 18604 8840
rect 18644 8800 18738 8840
rect 18595 8799 18653 8800
rect 15427 8756 15485 8757
rect 21379 8756 21437 8757
rect 15342 8716 15436 8756
rect 15476 8716 15485 8756
rect 16099 8716 16108 8756
rect 16148 8716 21388 8756
rect 21428 8716 21437 8756
rect 15427 8715 15485 8716
rect 21379 8715 21437 8716
rect 4387 8632 4396 8672
rect 4436 8632 7564 8672
rect 7604 8632 9100 8672
rect 9140 8632 9149 8672
rect 9571 8632 9580 8672
rect 9620 8632 11884 8672
rect 11924 8632 12076 8672
rect 12116 8632 12125 8672
rect 12750 8632 12844 8672
rect 12884 8632 12893 8672
rect 13411 8632 13420 8672
rect 13460 8632 13469 8672
rect 14755 8632 14764 8672
rect 14804 8632 16876 8672
rect 16916 8632 16925 8672
rect 19459 8632 19468 8672
rect 19508 8632 19756 8672
rect 19796 8632 19948 8672
rect 19988 8632 19997 8672
rect 4387 8631 4445 8632
rect 12067 8631 12125 8632
rect 12835 8631 12893 8632
rect 15523 8588 15581 8589
rect 2371 8548 2380 8588
rect 2420 8548 4108 8588
rect 4148 8548 4588 8588
rect 4628 8548 4637 8588
rect 5923 8548 5932 8588
rect 5972 8548 12460 8588
rect 12500 8548 12509 8588
rect 13699 8548 13708 8588
rect 13748 8548 14092 8588
rect 14132 8548 14141 8588
rect 15235 8548 15244 8588
rect 15284 8548 15532 8588
rect 15572 8548 15581 8588
rect 0 8504 80 8524
rect 3235 8504 3293 8505
rect 4483 8504 4541 8505
rect 12460 8504 12500 8548
rect 15523 8547 15581 8548
rect 0 8464 1420 8504
rect 1460 8464 1469 8504
rect 2860 8464 3244 8504
rect 3284 8464 3293 8504
rect 3619 8464 3628 8504
rect 3668 8464 4492 8504
rect 4532 8464 4541 8504
rect 4867 8464 4876 8504
rect 4916 8464 9580 8504
rect 9620 8464 9629 8504
rect 12460 8464 18412 8504
rect 18452 8464 18461 8504
rect 0 8444 80 8464
rect 2860 8420 2900 8464
rect 3235 8463 3293 8464
rect 4483 8463 4541 8464
rect 19939 8420 19997 8421
rect 2851 8380 2860 8420
rect 2900 8380 2909 8420
rect 3139 8380 3148 8420
rect 3188 8380 11692 8420
rect 11732 8380 11741 8420
rect 12931 8380 12940 8420
rect 12980 8380 19948 8420
rect 19988 8380 19997 8420
rect 19939 8379 19997 8380
rect 2467 8296 2476 8336
rect 2516 8296 4204 8336
rect 4244 8296 4253 8336
rect 4919 8296 4928 8336
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 5296 8296 5305 8336
rect 5356 8296 8332 8336
rect 8372 8296 8381 8336
rect 15331 8296 15340 8336
rect 15380 8296 15820 8336
rect 15860 8296 15869 8336
rect 20039 8296 20048 8336
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20416 8296 20425 8336
rect 5356 8252 5396 8296
rect 14947 8252 15005 8253
rect 15235 8252 15293 8253
rect 2500 8212 5396 8252
rect 8227 8212 8236 8252
rect 8276 8212 13036 8252
rect 13076 8212 13085 8252
rect 14179 8212 14188 8252
rect 14228 8212 14956 8252
rect 14996 8212 15005 8252
rect 15150 8212 15244 8252
rect 15284 8212 15293 8252
rect 15523 8212 15532 8252
rect 15572 8212 16588 8252
rect 16628 8212 16637 8252
rect 0 8168 80 8188
rect 0 8128 1804 8168
rect 1844 8128 1853 8168
rect 0 8108 80 8128
rect 2500 8084 2540 8212
rect 14947 8211 15005 8212
rect 15235 8211 15293 8212
rect 2755 8168 2813 8169
rect 7939 8168 7997 8169
rect 14275 8168 14333 8169
rect 2755 8128 2764 8168
rect 2804 8128 3532 8168
rect 3572 8128 3581 8168
rect 5251 8128 5260 8168
rect 5300 8128 5452 8168
rect 5492 8128 5501 8168
rect 5548 8128 6412 8168
rect 6452 8128 6461 8168
rect 6979 8128 6988 8168
rect 7028 8128 7276 8168
rect 7316 8128 7325 8168
rect 7939 8128 7948 8168
rect 7988 8128 8044 8168
rect 8084 8128 8093 8168
rect 14190 8128 14284 8168
rect 14324 8128 14333 8168
rect 15043 8128 15052 8168
rect 15092 8128 15724 8168
rect 15764 8128 15773 8168
rect 16003 8128 16012 8168
rect 16052 8128 19660 8168
rect 19700 8128 19709 8168
rect 2755 8127 2813 8128
rect 4291 8084 4349 8085
rect 5548 8084 5588 8128
rect 7939 8127 7997 8128
rect 14275 8127 14333 8128
rect 8515 8084 8573 8085
rect 1987 8044 1996 8084
rect 2036 8044 2540 8084
rect 2668 8044 3436 8084
rect 3476 8044 3485 8084
rect 4291 8044 4300 8084
rect 4340 8044 5588 8084
rect 6115 8044 6124 8084
rect 6164 8044 8524 8084
rect 8564 8044 18700 8084
rect 18740 8044 18749 8084
rect 2467 8000 2525 8001
rect 2668 8000 2708 8044
rect 4291 8043 4349 8044
rect 8515 8043 8573 8044
rect 4387 8000 4445 8001
rect 1219 7960 1228 8000
rect 1268 7960 2092 8000
rect 2132 7960 2141 8000
rect 2382 7960 2476 8000
rect 2516 7960 2525 8000
rect 2659 7960 2668 8000
rect 2708 7960 2717 8000
rect 4195 7960 4204 8000
rect 4244 7960 4396 8000
rect 4436 7960 4445 8000
rect 2467 7959 2525 7960
rect 4387 7959 4445 7960
rect 4675 8000 4733 8001
rect 10051 8000 10109 8001
rect 12067 8000 12125 8001
rect 4675 7960 4684 8000
rect 4724 7960 5740 8000
rect 5780 7960 5789 8000
rect 10051 7960 10060 8000
rect 10100 7960 10194 8000
rect 10435 7960 10444 8000
rect 10484 7960 10732 8000
rect 10772 7960 10781 8000
rect 12067 7960 12076 8000
rect 12116 7960 13708 8000
rect 13748 7960 14036 8000
rect 14083 7960 14092 8000
rect 14132 7960 17068 8000
rect 17108 7960 17117 8000
rect 18115 7960 18124 8000
rect 18164 7960 19852 8000
rect 19892 7960 19901 8000
rect 4675 7959 4733 7960
rect 10051 7959 10109 7960
rect 12067 7959 12125 7960
rect 2851 7916 2909 7917
rect 8611 7916 8669 7917
rect 13996 7916 14036 7960
rect 15235 7916 15293 7917
rect 1315 7876 1324 7916
rect 1364 7876 2860 7916
rect 2900 7876 2909 7916
rect 3427 7876 3436 7916
rect 3476 7876 6892 7916
rect 6932 7876 6941 7916
rect 7075 7876 7084 7916
rect 7124 7876 7133 7916
rect 8611 7876 8620 7916
rect 8660 7876 13804 7916
rect 13844 7876 13853 7916
rect 13996 7876 15244 7916
rect 15284 7876 15916 7916
rect 15956 7876 16204 7916
rect 16244 7876 16253 7916
rect 2851 7875 2909 7876
rect 0 7832 80 7852
rect 7084 7832 7124 7876
rect 8611 7875 8669 7876
rect 15235 7875 15293 7876
rect 19267 7832 19325 7833
rect 0 7792 1132 7832
rect 1172 7792 1181 7832
rect 4003 7792 4012 7832
rect 4052 7792 4061 7832
rect 6412 7792 7124 7832
rect 12835 7792 12844 7832
rect 12884 7792 18988 7832
rect 19028 7792 19276 7832
rect 19316 7792 19325 7832
rect 0 7772 80 7792
rect 2179 7708 2188 7748
rect 2228 7708 2476 7748
rect 2516 7708 2525 7748
rect 4012 7664 4052 7792
rect 6412 7749 6452 7792
rect 19267 7791 19325 7792
rect 6403 7748 6461 7749
rect 4579 7708 4588 7748
rect 4628 7708 5452 7748
rect 5492 7708 6412 7748
rect 6452 7708 6461 7748
rect 6403 7707 6461 7708
rect 6595 7748 6653 7749
rect 6595 7708 6604 7748
rect 6644 7708 6738 7748
rect 7075 7708 7084 7748
rect 7124 7708 7468 7748
rect 7508 7708 7517 7748
rect 8035 7708 8044 7748
rect 8084 7708 19372 7748
rect 19412 7708 19421 7748
rect 6595 7707 6653 7708
rect 15523 7664 15581 7665
rect 4012 7624 10060 7664
rect 10100 7624 10109 7664
rect 15235 7624 15244 7664
rect 15284 7624 15532 7664
rect 15572 7624 15581 7664
rect 15523 7623 15581 7624
rect 17923 7664 17981 7665
rect 17923 7624 17932 7664
rect 17972 7624 18028 7664
rect 18068 7624 18077 7664
rect 17923 7623 17981 7624
rect 12163 7580 12221 7581
rect 12643 7580 12701 7581
rect 15139 7580 15197 7581
rect 3679 7540 3688 7580
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 4056 7540 4065 7580
rect 6019 7540 6028 7580
rect 6068 7540 6796 7580
rect 6836 7540 6845 7580
rect 12163 7540 12172 7580
rect 12212 7540 12652 7580
rect 12692 7540 12701 7580
rect 14179 7540 14188 7580
rect 14228 7540 14860 7580
rect 14900 7540 14909 7580
rect 15139 7540 15148 7580
rect 15188 7540 15340 7580
rect 15380 7540 15389 7580
rect 17155 7540 17164 7580
rect 17204 7540 18508 7580
rect 18548 7540 18557 7580
rect 18799 7540 18808 7580
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 19176 7540 19185 7580
rect 12163 7539 12221 7540
rect 12643 7539 12701 7540
rect 15139 7539 15197 7540
rect 0 7496 80 7516
rect 0 7456 1612 7496
rect 1652 7456 1661 7496
rect 2956 7456 3340 7496
rect 3380 7456 3389 7496
rect 5155 7456 5164 7496
rect 5204 7456 8716 7496
rect 8756 7456 10252 7496
rect 10292 7456 10301 7496
rect 10531 7456 10540 7496
rect 10580 7456 12460 7496
rect 12500 7456 13612 7496
rect 13652 7456 13661 7496
rect 14659 7456 14668 7496
rect 14708 7456 16492 7496
rect 16532 7456 19372 7496
rect 19412 7456 19421 7496
rect 0 7436 80 7456
rect 2956 7412 2996 7456
rect 9571 7412 9629 7413
rect 2947 7372 2956 7412
rect 2996 7372 3005 7412
rect 3811 7372 3820 7412
rect 3860 7372 5836 7412
rect 5876 7372 6220 7412
rect 6260 7372 6269 7412
rect 9486 7372 9580 7412
rect 9620 7372 9629 7412
rect 9571 7371 9629 7372
rect 10051 7412 10109 7413
rect 10051 7372 10060 7412
rect 10100 7372 11692 7412
rect 11732 7372 11741 7412
rect 14755 7372 14764 7412
rect 14804 7372 14813 7412
rect 10051 7371 10109 7372
rect 8419 7328 8477 7329
rect 3715 7288 3724 7328
rect 3764 7288 7948 7328
rect 7988 7288 7997 7328
rect 8419 7288 8428 7328
rect 8468 7288 10828 7328
rect 10868 7288 10877 7328
rect 8419 7287 8477 7288
rect 8803 7244 8861 7245
rect 3628 7204 5260 7244
rect 5300 7204 5309 7244
rect 8718 7204 8812 7244
rect 8852 7204 8861 7244
rect 0 7160 80 7180
rect 3628 7160 3668 7204
rect 8803 7203 8861 7204
rect 12067 7160 12125 7161
rect 0 7120 1036 7160
rect 1076 7120 1085 7160
rect 2563 7120 2572 7160
rect 2612 7120 2764 7160
rect 2804 7120 2813 7160
rect 3331 7120 3340 7160
rect 3380 7120 3628 7160
rect 3668 7120 3677 7160
rect 4003 7120 4012 7160
rect 4052 7120 4300 7160
rect 4340 7120 4349 7160
rect 4588 7120 6412 7160
rect 6452 7120 7276 7160
rect 7316 7120 7325 7160
rect 7459 7120 7468 7160
rect 7508 7120 7660 7160
rect 7700 7120 7709 7160
rect 7939 7120 7948 7160
rect 7988 7120 8332 7160
rect 8372 7120 10540 7160
rect 10580 7120 10589 7160
rect 10723 7120 10732 7160
rect 10772 7120 11500 7160
rect 11540 7120 12076 7160
rect 12116 7120 12125 7160
rect 0 7100 80 7120
rect 2764 7076 2804 7120
rect 4588 7076 4628 7120
rect 12067 7119 12125 7120
rect 2764 7036 4628 7076
rect 4675 7076 4733 7077
rect 14764 7076 14804 7372
rect 16579 7288 16588 7328
rect 16628 7288 18604 7328
rect 18644 7288 18653 7328
rect 17827 7120 17836 7160
rect 17876 7120 19756 7160
rect 19796 7120 19805 7160
rect 15043 7076 15101 7077
rect 4675 7036 4684 7076
rect 4724 7036 7852 7076
rect 7892 7036 7901 7076
rect 8035 7036 8044 7076
rect 8084 7036 12556 7076
rect 12596 7036 12605 7076
rect 14275 7036 14284 7076
rect 14324 7036 14572 7076
rect 14612 7036 14621 7076
rect 14764 7036 14860 7076
rect 14900 7036 14909 7076
rect 15043 7036 15052 7076
rect 15092 7036 15186 7076
rect 4675 7035 4733 7036
rect 15043 7035 15101 7036
rect 2179 6952 2188 6992
rect 2228 6952 2540 6992
rect 6307 6952 6316 6992
rect 6356 6952 6796 6992
rect 6836 6952 6845 6992
rect 8515 6952 8524 6992
rect 8564 6952 9388 6992
rect 9428 6952 9437 6992
rect 11107 6952 11116 6992
rect 11156 6952 16300 6992
rect 16340 6952 16349 6992
rect 2500 6908 2540 6952
rect 2500 6868 11360 6908
rect 12835 6868 12844 6908
rect 12884 6868 13132 6908
rect 13172 6868 16588 6908
rect 16628 6868 16637 6908
rect 0 6824 80 6844
rect 11320 6824 11360 6868
rect 15811 6824 15869 6825
rect 0 6784 844 6824
rect 884 6784 893 6824
rect 3139 6784 3148 6824
rect 3188 6784 3628 6824
rect 3668 6784 3677 6824
rect 4771 6784 4780 6824
rect 4820 6784 4829 6824
rect 4919 6784 4928 6824
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 5296 6784 5305 6824
rect 6115 6784 6124 6824
rect 6164 6784 8140 6824
rect 8180 6784 8189 6824
rect 11320 6784 15820 6824
rect 15860 6784 15869 6824
rect 20039 6784 20048 6824
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20416 6784 20425 6824
rect 0 6764 80 6784
rect 4780 6740 4820 6784
rect 15811 6783 15869 6784
rect 3427 6700 3436 6740
rect 3476 6700 4820 6740
rect 5164 6700 5740 6740
rect 5780 6700 5789 6740
rect 6595 6700 6604 6740
rect 6644 6700 6988 6740
rect 7028 6700 7037 6740
rect 7651 6700 7660 6740
rect 7700 6700 7852 6740
rect 7892 6700 7901 6740
rect 5164 6656 5204 6700
rect 6307 6656 6365 6657
rect 2275 6616 2284 6656
rect 2324 6616 5204 6656
rect 5251 6616 5260 6656
rect 5300 6616 6316 6656
rect 6356 6616 6365 6656
rect 7267 6616 7276 6656
rect 7316 6616 8908 6656
rect 8948 6616 8957 6656
rect 10723 6616 10732 6656
rect 10772 6616 11596 6656
rect 11636 6616 11645 6656
rect 19459 6616 19468 6656
rect 19508 6616 19948 6656
rect 19988 6616 19997 6656
rect 6307 6615 6365 6616
rect 5155 6532 5164 6572
rect 5204 6532 5548 6572
rect 5588 6532 5597 6572
rect 5731 6532 5740 6572
rect 5780 6532 8812 6572
rect 8852 6532 8861 6572
rect 14851 6532 14860 6572
rect 14900 6532 18508 6572
rect 18548 6532 18557 6572
rect 0 6488 80 6508
rect 2371 6488 2429 6489
rect 16291 6488 16349 6489
rect 0 6428 116 6488
rect 1219 6448 1228 6488
rect 1268 6448 2380 6488
rect 2420 6448 2429 6488
rect 3043 6448 3052 6488
rect 3092 6448 11360 6488
rect 12547 6448 12556 6488
rect 12596 6448 13228 6488
rect 13268 6448 13277 6488
rect 13507 6448 13516 6488
rect 13556 6448 14092 6488
rect 14132 6448 16108 6488
rect 16148 6448 16157 6488
rect 16291 6448 16300 6488
rect 16340 6448 16492 6488
rect 16532 6448 16541 6488
rect 2371 6447 2429 6448
rect 76 6404 116 6428
rect 11320 6404 11360 6448
rect 16291 6447 16349 6448
rect 16300 6404 16340 6447
rect 76 6364 10964 6404
rect 11320 6364 12364 6404
rect 12404 6364 12413 6404
rect 14371 6364 14380 6404
rect 14420 6364 16340 6404
rect 18211 6364 18220 6404
rect 18260 6364 18269 6404
rect 6595 6320 6653 6321
rect 7939 6320 7997 6321
rect 10723 6320 10781 6321
rect 10924 6320 10964 6364
rect 18220 6320 18260 6364
rect 2659 6280 2668 6320
rect 2708 6280 4972 6320
rect 5012 6280 5021 6320
rect 5068 6280 6604 6320
rect 6644 6280 6653 6320
rect 7651 6280 7660 6320
rect 7700 6280 7948 6320
rect 7988 6280 7997 6320
rect 8227 6280 8236 6320
rect 8276 6280 10732 6320
rect 10772 6280 10781 6320
rect 10915 6280 10924 6320
rect 10964 6280 10973 6320
rect 11395 6280 11404 6320
rect 11444 6280 13132 6320
rect 13172 6280 15628 6320
rect 15668 6280 16204 6320
rect 16244 6280 16253 6320
rect 16483 6280 16492 6320
rect 16532 6280 16780 6320
rect 16820 6280 16829 6320
rect 18220 6280 18508 6320
rect 18548 6280 18557 6320
rect 5068 6236 5108 6280
rect 6595 6279 6653 6280
rect 7939 6279 7997 6280
rect 10723 6279 10781 6280
rect 1699 6196 1708 6236
rect 1748 6196 5108 6236
rect 6403 6236 6461 6237
rect 6403 6196 6412 6236
rect 6452 6196 6546 6236
rect 8707 6196 8716 6236
rect 8756 6196 9100 6236
rect 9140 6196 9149 6236
rect 15427 6196 15436 6236
rect 15476 6196 19276 6236
rect 19316 6196 19325 6236
rect 6403 6195 6461 6196
rect 0 6152 80 6172
rect 0 6112 212 6152
rect 5539 6112 5548 6152
rect 5588 6112 9292 6152
rect 9332 6112 9484 6152
rect 9524 6112 9533 6152
rect 12643 6112 12652 6152
rect 12692 6112 13324 6152
rect 13364 6112 13373 6152
rect 0 6092 80 6112
rect 172 5984 212 6112
rect 6499 6068 6557 6069
rect 3679 6028 3688 6068
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 4056 6028 4065 6068
rect 6499 6028 6508 6068
rect 6548 6028 7660 6068
rect 7700 6028 7709 6068
rect 8995 6028 9004 6068
rect 9044 6028 11116 6068
rect 11156 6028 11165 6068
rect 18799 6028 18808 6068
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 19176 6028 19185 6068
rect 6499 6027 6557 6028
rect 11683 5984 11741 5985
rect 172 5944 4396 5984
rect 4436 5944 4445 5984
rect 6211 5944 6220 5984
rect 6260 5944 10156 5984
rect 10196 5944 10205 5984
rect 11683 5944 11692 5984
rect 11732 5944 11788 5984
rect 11828 5944 11837 5984
rect 11683 5943 11741 5944
rect 4195 5900 4253 5901
rect 9283 5900 9341 5901
rect 12259 5900 12317 5901
rect 3811 5860 3820 5900
rect 3860 5860 4204 5900
rect 4244 5860 4253 5900
rect 7363 5860 7372 5900
rect 7412 5860 8332 5900
rect 8372 5860 8381 5900
rect 9198 5860 9292 5900
rect 9332 5860 9772 5900
rect 9812 5860 9821 5900
rect 11587 5860 11596 5900
rect 11636 5860 12268 5900
rect 12308 5860 12317 5900
rect 17251 5860 17260 5900
rect 17300 5860 18220 5900
rect 18260 5860 18412 5900
rect 18452 5860 18461 5900
rect 4195 5859 4253 5860
rect 9283 5859 9341 5860
rect 12259 5859 12317 5860
rect 0 5816 80 5836
rect 10243 5816 10301 5817
rect 17635 5816 17693 5817
rect 0 5776 2540 5816
rect 9187 5776 9196 5816
rect 9236 5776 9245 5816
rect 10243 5776 10252 5816
rect 10292 5776 11692 5816
rect 11732 5776 11741 5816
rect 14467 5776 14476 5816
rect 14516 5776 14764 5816
rect 14804 5776 14813 5816
rect 17347 5776 17356 5816
rect 17396 5776 17644 5816
rect 17684 5776 17693 5816
rect 17923 5776 17932 5816
rect 17972 5776 18316 5816
rect 18356 5776 18365 5816
rect 0 5756 80 5776
rect 2500 5732 2540 5776
rect 6115 5732 6173 5733
rect 8899 5732 8957 5733
rect 2500 5692 2668 5732
rect 2708 5692 2717 5732
rect 3043 5692 3052 5732
rect 3092 5692 4876 5732
rect 4916 5692 6124 5732
rect 6164 5692 6173 5732
rect 7267 5692 7276 5732
rect 7316 5692 8044 5732
rect 8084 5692 8093 5732
rect 8814 5692 8908 5732
rect 8948 5692 8957 5732
rect 6115 5691 6173 5692
rect 8899 5691 8957 5692
rect 643 5648 701 5649
rect 5347 5648 5405 5649
rect 643 5608 652 5648
rect 692 5608 4204 5648
rect 4244 5608 4253 5648
rect 5059 5608 5068 5648
rect 5108 5608 5356 5648
rect 5396 5608 5644 5648
rect 5684 5608 5693 5648
rect 6883 5608 6892 5648
rect 6932 5608 8428 5648
rect 8468 5608 8477 5648
rect 643 5607 701 5608
rect 5347 5607 5405 5608
rect 5539 5564 5597 5565
rect 1987 5524 1996 5564
rect 2036 5524 5548 5564
rect 5588 5524 5597 5564
rect 5731 5524 5740 5564
rect 5780 5524 5932 5564
rect 5972 5524 5981 5564
rect 5539 5523 5597 5524
rect 0 5480 80 5500
rect 9196 5480 9236 5776
rect 10243 5775 10301 5776
rect 17635 5775 17693 5776
rect 9475 5732 9533 5733
rect 9475 5692 9484 5732
rect 9524 5692 10252 5732
rect 10292 5692 10301 5732
rect 14563 5692 14572 5732
rect 14612 5692 18508 5732
rect 18548 5692 18557 5732
rect 9475 5691 9533 5692
rect 10723 5648 10781 5649
rect 14275 5648 14333 5649
rect 15043 5648 15101 5649
rect 19267 5648 19325 5649
rect 10638 5608 10732 5648
rect 10772 5608 10781 5648
rect 11587 5608 11596 5648
rect 11636 5608 12172 5648
rect 12212 5608 12221 5648
rect 14083 5608 14092 5648
rect 14132 5608 14284 5648
rect 14324 5608 14333 5648
rect 14958 5608 15052 5648
rect 15092 5608 15101 5648
rect 17827 5608 17836 5648
rect 17876 5608 18796 5648
rect 18836 5608 19276 5648
rect 19316 5608 19325 5648
rect 10723 5607 10781 5608
rect 14275 5607 14333 5608
rect 15043 5607 15101 5608
rect 19267 5607 19325 5608
rect 16675 5524 16684 5564
rect 16724 5524 17260 5564
rect 17300 5524 17309 5564
rect 0 5440 9236 5480
rect 9379 5480 9437 5481
rect 9379 5440 9388 5480
rect 9428 5440 9522 5480
rect 0 5420 80 5440
rect 9379 5439 9437 5440
rect 2083 5356 2092 5396
rect 2132 5356 14188 5396
rect 14228 5356 14237 5396
rect 16771 5356 16780 5396
rect 16820 5356 17356 5396
rect 17396 5356 17405 5396
rect 4483 5312 4541 5313
rect 2467 5272 2476 5312
rect 2516 5272 2764 5312
rect 2804 5272 3628 5312
rect 3668 5272 3677 5312
rect 4483 5272 4492 5312
rect 4532 5272 4780 5312
rect 4820 5272 4829 5312
rect 4919 5272 4928 5312
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 5296 5272 5305 5312
rect 6307 5272 6316 5312
rect 6356 5272 6365 5312
rect 7459 5272 7468 5312
rect 7508 5272 9772 5312
rect 9812 5272 11980 5312
rect 12020 5272 12029 5312
rect 14284 5272 18700 5312
rect 18740 5272 18749 5312
rect 20039 5272 20048 5312
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20416 5272 20425 5312
rect 4483 5271 4541 5272
rect 1411 5188 1420 5228
rect 1460 5188 6028 5228
rect 6068 5188 6077 5228
rect 0 5144 80 5164
rect 1315 5144 1373 5145
rect 0 5104 1324 5144
rect 1364 5104 1373 5144
rect 0 5084 80 5104
rect 1315 5103 1373 5104
rect 3427 5144 3485 5145
rect 6316 5144 6356 5272
rect 7267 5228 7325 5229
rect 12931 5228 12989 5229
rect 14284 5228 14324 5272
rect 7267 5188 7276 5228
rect 7316 5188 12940 5228
rect 12980 5188 14324 5228
rect 15619 5228 15677 5229
rect 15619 5188 15628 5228
rect 15668 5188 18316 5228
rect 18356 5188 18365 5228
rect 7267 5187 7325 5188
rect 12931 5187 12989 5188
rect 15619 5187 15677 5188
rect 7843 5144 7901 5145
rect 3427 5104 3436 5144
rect 3476 5104 4204 5144
rect 4244 5104 4253 5144
rect 4387 5104 4396 5144
rect 4436 5104 6356 5144
rect 7171 5104 7180 5144
rect 7220 5104 7852 5144
rect 7892 5104 7901 5144
rect 8995 5104 9004 5144
rect 9044 5104 9676 5144
rect 9716 5104 9725 5144
rect 12067 5104 12076 5144
rect 12116 5104 12308 5144
rect 3427 5103 3485 5104
rect 7843 5103 7901 5104
rect 12268 5060 12308 5104
rect 17635 5060 17693 5061
rect 7180 5020 7468 5060
rect 7508 5020 7517 5060
rect 9283 5020 9292 5060
rect 9332 5020 11404 5060
rect 11444 5020 11453 5060
rect 12259 5020 12268 5060
rect 12308 5020 12317 5060
rect 15724 5020 16204 5060
rect 16244 5020 16253 5060
rect 17635 5020 17644 5060
rect 17684 5020 18412 5060
rect 18452 5020 19468 5060
rect 19508 5020 19517 5060
rect 5443 4976 5501 4977
rect 7180 4976 7220 5020
rect 10435 4976 10493 4977
rect 15724 4976 15764 5020
rect 17635 5019 17693 5020
rect 5358 4936 5452 4976
rect 5492 4936 5501 4976
rect 7171 4936 7180 4976
rect 7220 4936 7229 4976
rect 7276 4936 8468 4976
rect 8803 4936 8812 4976
rect 8852 4936 10444 4976
rect 10484 4936 10493 4976
rect 12067 4936 12076 4976
rect 12116 4936 13516 4976
rect 13556 4936 13565 4976
rect 13795 4936 13804 4976
rect 13844 4936 15532 4976
rect 15572 4936 15581 4976
rect 15715 4936 15724 4976
rect 15764 4936 15773 4976
rect 16291 4936 16300 4976
rect 16340 4936 17164 4976
rect 17204 4936 17644 4976
rect 17684 4936 17693 4976
rect 18979 4936 18988 4976
rect 19028 4936 19372 4976
rect 19412 4936 19421 4976
rect 5443 4935 5501 4936
rect 2947 4852 2956 4892
rect 2996 4852 3244 4892
rect 3284 4852 3293 4892
rect 0 4808 80 4828
rect 4291 4808 4349 4809
rect 5452 4808 5492 4935
rect 7276 4892 7316 4936
rect 8428 4892 8468 4936
rect 10435 4935 10493 4936
rect 9091 4892 9149 4893
rect 17923 4892 17981 4893
rect 5923 4852 5932 4892
rect 5972 4852 7316 4892
rect 7363 4852 7372 4892
rect 7412 4852 8044 4892
rect 8084 4852 8093 4892
rect 8428 4852 9100 4892
rect 9140 4852 9149 4892
rect 9091 4851 9149 4852
rect 9964 4852 13228 4892
rect 13268 4852 13277 4892
rect 14947 4852 14956 4892
rect 14996 4852 15916 4892
rect 15956 4852 15965 4892
rect 17923 4852 17932 4892
rect 17972 4852 19948 4892
rect 19988 4852 19997 4892
rect 0 4768 4300 4808
rect 4340 4768 4349 4808
rect 4579 4768 4588 4808
rect 4628 4768 5492 4808
rect 6115 4808 6173 4809
rect 6787 4808 6845 4809
rect 9964 4808 10004 4852
rect 14956 4808 14996 4852
rect 17923 4851 17981 4852
rect 6115 4768 6124 4808
rect 6164 4768 6412 4808
rect 6452 4768 6461 4808
rect 6702 4768 6796 4808
rect 6836 4768 6845 4808
rect 7555 4768 7564 4808
rect 7604 4768 10004 4808
rect 10243 4768 10252 4808
rect 10292 4768 11596 4808
rect 11636 4768 11645 4808
rect 12547 4768 12556 4808
rect 12596 4768 14996 4808
rect 0 4748 80 4768
rect 4291 4767 4349 4768
rect 6115 4767 6173 4768
rect 6787 4767 6845 4768
rect 18403 4724 18461 4725
rect 4003 4684 4012 4724
rect 4052 4684 4204 4724
rect 4244 4684 4253 4724
rect 6979 4684 6988 4724
rect 7028 4684 12172 4724
rect 12212 4684 12221 4724
rect 18211 4684 18220 4724
rect 18260 4684 18412 4724
rect 18452 4684 18461 4724
rect 18403 4683 18461 4684
rect 8707 4640 8765 4641
rect 13027 4640 13085 4641
rect 2851 4600 2860 4640
rect 2900 4600 5876 4640
rect 5923 4600 5932 4640
rect 5972 4600 6220 4640
rect 6260 4600 6269 4640
rect 7180 4600 7948 4640
rect 7988 4600 7997 4640
rect 8707 4600 8716 4640
rect 8756 4600 13036 4640
rect 13076 4600 13085 4640
rect 4963 4556 5021 4557
rect 1891 4516 1900 4556
rect 1940 4516 2188 4556
rect 2228 4516 2237 4556
rect 3679 4516 3688 4556
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 4056 4516 4065 4556
rect 4878 4516 4972 4556
rect 5012 4516 5021 4556
rect 5836 4556 5876 4600
rect 7180 4556 7220 4600
rect 8707 4599 8765 4600
rect 13027 4599 13085 4600
rect 17923 4556 17981 4557
rect 5836 4516 7220 4556
rect 7267 4516 7276 4556
rect 7316 4516 10828 4556
rect 10868 4516 10877 4556
rect 12556 4516 16972 4556
rect 17012 4516 17932 4556
rect 17972 4516 17981 4556
rect 18799 4516 18808 4556
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 19176 4516 19185 4556
rect 4963 4515 5021 4516
rect 0 4472 80 4492
rect 9379 4472 9437 4473
rect 0 4432 76 4472
rect 116 4432 125 4472
rect 1699 4432 1708 4472
rect 1748 4432 9388 4472
rect 9428 4432 9437 4472
rect 10627 4432 10636 4472
rect 10676 4432 11212 4472
rect 11252 4432 11261 4472
rect 0 4412 80 4432
rect 9379 4431 9437 4432
rect 12556 4388 12596 4516
rect 17923 4515 17981 4516
rect 4579 4348 4588 4388
rect 4628 4348 5356 4388
rect 5396 4348 5405 4388
rect 6787 4348 6796 4388
rect 6836 4348 8620 4388
rect 8660 4348 8669 4388
rect 9004 4348 9196 4388
rect 9236 4348 9245 4388
rect 11320 4348 12596 4388
rect 12739 4348 12748 4388
rect 12788 4348 13132 4388
rect 13172 4348 13516 4388
rect 13556 4348 13565 4388
rect 2563 4304 2621 4305
rect 2563 4264 2572 4304
rect 2612 4264 2860 4304
rect 2900 4264 2909 4304
rect 2563 4263 2621 4264
rect 3139 4220 3197 4221
rect 8515 4220 8573 4221
rect 9004 4220 9044 4348
rect 11320 4304 11360 4348
rect 3054 4180 3148 4220
rect 3188 4180 3197 4220
rect 6307 4180 6316 4220
rect 6356 4180 8524 4220
rect 8564 4180 9044 4220
rect 9100 4264 11360 4304
rect 11875 4264 11884 4304
rect 11924 4264 14284 4304
rect 14324 4264 14333 4304
rect 3139 4179 3197 4180
rect 8515 4179 8573 4180
rect 0 4136 80 4156
rect 4099 4136 4157 4137
rect 9100 4136 9140 4264
rect 10819 4220 10877 4221
rect 9187 4180 9196 4220
rect 9236 4180 9868 4220
rect 9908 4180 9917 4220
rect 10734 4180 10828 4220
rect 10868 4180 10877 4220
rect 11203 4180 11212 4220
rect 11252 4180 13516 4220
rect 13556 4180 13565 4220
rect 0 4096 4108 4136
rect 4148 4096 4157 4136
rect 7555 4096 7564 4136
rect 7604 4096 8140 4136
rect 8180 4096 8189 4136
rect 8236 4096 9140 4136
rect 9868 4136 9908 4180
rect 10819 4179 10877 4180
rect 13891 4136 13949 4137
rect 16771 4136 16829 4137
rect 17923 4136 17981 4137
rect 9868 4096 11308 4136
rect 11348 4096 11357 4136
rect 13699 4096 13708 4136
rect 13748 4096 13900 4136
rect 13940 4096 13949 4136
rect 14947 4096 14956 4136
rect 14996 4096 15532 4136
rect 15572 4096 16588 4136
rect 16628 4096 16780 4136
rect 16820 4096 16829 4136
rect 17838 4096 17932 4136
rect 17972 4096 17981 4136
rect 0 4076 80 4096
rect 4099 4095 4157 4096
rect 8236 4052 8276 4096
rect 13891 4095 13949 4096
rect 16771 4095 16829 4096
rect 17923 4095 17981 4096
rect 2500 4012 8276 4052
rect 8899 4052 8957 4053
rect 8899 4012 8908 4052
rect 8948 4012 15820 4052
rect 15860 4012 15869 4052
rect 2500 3968 2540 4012
rect 8899 4011 8957 4012
rect 5731 3968 5789 3969
rect 9091 3968 9149 3969
rect 10147 3968 10205 3969
rect 1795 3928 1804 3968
rect 1844 3928 2540 3968
rect 4195 3928 4204 3968
rect 4244 3928 4492 3968
rect 4532 3928 4541 3968
rect 5155 3928 5164 3968
rect 5204 3928 5740 3968
rect 5780 3928 5789 3968
rect 7747 3928 7756 3968
rect 7796 3928 8620 3968
rect 8660 3928 8669 3968
rect 9091 3928 9100 3968
rect 9140 3928 10156 3968
rect 10196 3928 10205 3968
rect 5731 3927 5789 3928
rect 9091 3927 9149 3928
rect 10147 3927 10205 3928
rect 10339 3968 10397 3969
rect 10339 3928 10348 3968
rect 10388 3928 10482 3968
rect 11395 3928 11404 3968
rect 11444 3928 11980 3968
rect 12020 3928 12029 3968
rect 10339 3927 10397 3928
rect 2467 3884 2525 3885
rect 8323 3884 8381 3885
rect 2448 3844 2476 3884
rect 2516 3844 2572 3884
rect 2612 3844 4108 3884
rect 4148 3844 8236 3884
rect 8276 3844 8332 3884
rect 8372 3844 8381 3884
rect 2467 3843 2525 3844
rect 8323 3843 8381 3844
rect 10051 3884 10109 3885
rect 10051 3844 10060 3884
rect 10100 3844 12556 3884
rect 12596 3844 12605 3884
rect 15331 3844 15340 3884
rect 15380 3844 15820 3884
rect 15860 3844 15869 3884
rect 10051 3843 10109 3844
rect 0 3800 80 3820
rect 7459 3800 7517 3801
rect 0 3760 1900 3800
rect 1940 3760 1949 3800
rect 4919 3760 4928 3800
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 5296 3760 5305 3800
rect 7459 3760 7468 3800
rect 7508 3760 8140 3800
rect 8180 3760 8189 3800
rect 9283 3760 9292 3800
rect 9332 3760 9676 3800
rect 9716 3760 9725 3800
rect 20039 3760 20048 3800
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20416 3760 20425 3800
rect 0 3740 80 3760
rect 7459 3759 7517 3760
rect 11683 3716 11741 3717
rect 1411 3676 1420 3716
rect 1460 3676 3148 3716
rect 3188 3676 3197 3716
rect 7459 3676 7468 3716
rect 7508 3676 11692 3716
rect 11732 3676 12788 3716
rect 15619 3676 15628 3716
rect 15668 3676 16108 3716
rect 16148 3676 16157 3716
rect 18499 3676 18508 3716
rect 18548 3676 20180 3716
rect 11683 3675 11741 3676
rect 2083 3632 2141 3633
rect 2467 3632 2525 3633
rect 12748 3632 12788 3676
rect 16195 3632 16253 3633
rect 1998 3592 2092 3632
rect 2132 3592 2141 3632
rect 2382 3592 2476 3632
rect 2516 3592 3532 3632
rect 3572 3592 3581 3632
rect 5443 3592 5452 3632
rect 5492 3592 10156 3632
rect 10196 3592 10205 3632
rect 12748 3592 13132 3632
rect 13172 3592 13181 3632
rect 16110 3592 16204 3632
rect 16244 3592 16253 3632
rect 2083 3591 2141 3592
rect 2467 3591 2525 3592
rect 16195 3591 16253 3592
rect 16876 3592 19660 3632
rect 19700 3592 19709 3632
rect 2563 3548 2621 3549
rect 3331 3548 3389 3549
rect 5923 3548 5981 3549
rect 16876 3548 16916 3592
rect 1315 3508 1324 3548
rect 1364 3508 2572 3548
rect 2612 3508 2764 3548
rect 2804 3508 2813 3548
rect 3331 3508 3340 3548
rect 3380 3508 4204 3548
rect 4244 3508 5932 3548
rect 5972 3508 5981 3548
rect 8707 3508 8716 3548
rect 8756 3508 10252 3548
rect 10292 3508 10301 3548
rect 11875 3508 11884 3548
rect 11924 3508 14092 3548
rect 14132 3508 14141 3548
rect 15715 3508 15724 3548
rect 15764 3508 16012 3548
rect 16052 3508 16916 3548
rect 20140 3548 20180 3676
rect 20140 3508 20236 3548
rect 20276 3508 20285 3548
rect 2563 3507 2621 3508
rect 3331 3507 3389 3508
rect 5923 3507 5981 3508
rect 0 3464 80 3484
rect 0 3424 404 3464
rect 2275 3424 2284 3464
rect 2324 3424 5204 3464
rect 5251 3424 5260 3464
rect 5300 3424 7468 3464
rect 7508 3424 7517 3464
rect 7651 3424 7660 3464
rect 7700 3424 9292 3464
rect 9332 3424 9341 3464
rect 9580 3424 15052 3464
rect 15092 3424 15244 3464
rect 15284 3424 15293 3464
rect 0 3404 80 3424
rect 364 3380 404 3424
rect 4579 3380 4637 3381
rect 364 3340 4588 3380
rect 4628 3340 4637 3380
rect 5164 3380 5204 3424
rect 7747 3380 7805 3381
rect 9580 3380 9620 3424
rect 10051 3380 10109 3381
rect 10531 3380 10589 3381
rect 5164 3340 5548 3380
rect 5588 3340 5597 3380
rect 7662 3340 7756 3380
rect 7796 3340 7805 3380
rect 4579 3339 4637 3340
rect 7747 3339 7805 3340
rect 8716 3340 9196 3380
rect 9236 3340 9580 3380
rect 9620 3340 9629 3380
rect 9966 3340 10060 3380
rect 10100 3340 10109 3380
rect 10446 3340 10540 3380
rect 10580 3340 10589 3380
rect 931 3296 989 3297
rect 8716 3296 8756 3340
rect 10051 3339 10109 3340
rect 10531 3339 10589 3340
rect 11491 3380 11549 3381
rect 12355 3380 12413 3381
rect 16579 3380 16637 3381
rect 16963 3380 17021 3381
rect 11491 3340 11500 3380
rect 11540 3340 11634 3380
rect 12355 3340 12364 3380
rect 12404 3340 13708 3380
rect 13748 3340 13757 3380
rect 16494 3340 16588 3380
rect 16628 3340 16637 3380
rect 16878 3340 16972 3380
rect 17012 3340 17021 3380
rect 11491 3339 11549 3340
rect 12355 3339 12413 3340
rect 16579 3339 16637 3340
rect 16963 3339 17021 3340
rect 931 3256 940 3296
rect 980 3256 5164 3296
rect 5204 3256 5213 3296
rect 5347 3256 5356 3296
rect 5396 3256 8756 3296
rect 8803 3296 8861 3297
rect 8803 3256 8812 3296
rect 8852 3256 11020 3296
rect 11060 3256 11069 3296
rect 13123 3256 13132 3296
rect 13172 3256 18700 3296
rect 18740 3256 18749 3296
rect 931 3255 989 3256
rect 8803 3255 8861 3256
rect 4387 3172 4396 3212
rect 4436 3172 4684 3212
rect 4724 3172 4733 3212
rect 6019 3172 6028 3212
rect 6068 3172 6412 3212
rect 6452 3172 6461 3212
rect 7843 3172 7852 3212
rect 7892 3172 7901 3212
rect 8323 3172 8332 3212
rect 8372 3172 10540 3212
rect 10580 3172 10589 3212
rect 15043 3172 15052 3212
rect 15092 3172 16396 3212
rect 16436 3172 16445 3212
rect 0 3128 80 3148
rect 2275 3128 2333 3129
rect 7852 3128 7892 3172
rect 15043 3128 15101 3129
rect 0 3088 2284 3128
rect 2324 3088 2333 3128
rect 3043 3088 3052 3128
rect 3092 3088 7028 3128
rect 7075 3088 7084 3128
rect 7124 3088 7756 3128
rect 7796 3088 7805 3128
rect 7852 3088 8716 3128
rect 8756 3088 12844 3128
rect 12884 3088 15052 3128
rect 15092 3088 16204 3128
rect 16244 3088 16253 3128
rect 16579 3088 16588 3128
rect 16628 3088 17548 3128
rect 17588 3088 17597 3128
rect 0 3068 80 3088
rect 2275 3087 2333 3088
rect 6988 3044 7028 3088
rect 15043 3087 15101 3088
rect 8899 3044 8957 3045
rect 2755 3004 2764 3044
rect 2804 3004 3532 3044
rect 3572 3004 3581 3044
rect 3679 3004 3688 3044
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 4056 3004 4065 3044
rect 6988 3004 8908 3044
rect 8948 3004 8957 3044
rect 8899 3003 8957 3004
rect 11203 3044 11261 3045
rect 11203 3004 11212 3044
rect 11252 3004 18028 3044
rect 18068 3004 18077 3044
rect 18799 3004 18808 3044
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 19176 3004 19185 3044
rect 11203 3003 11261 3004
rect 4195 2920 4204 2960
rect 4244 2920 13612 2960
rect 13652 2920 13661 2960
rect 13708 2920 17068 2960
rect 17108 2920 17117 2960
rect 1795 2876 1853 2877
rect 13708 2876 13748 2920
rect 1795 2836 1804 2876
rect 1844 2836 3436 2876
rect 3476 2836 3485 2876
rect 9475 2836 9484 2876
rect 9524 2836 10828 2876
rect 10868 2836 10877 2876
rect 11107 2836 11116 2876
rect 11156 2836 12172 2876
rect 12212 2836 12221 2876
rect 13123 2836 13132 2876
rect 13172 2836 13748 2876
rect 14275 2836 14284 2876
rect 14324 2836 16780 2876
rect 16820 2836 16829 2876
rect 17827 2836 17836 2876
rect 17876 2836 18508 2876
rect 18548 2836 18557 2876
rect 1795 2835 1853 2836
rect 0 2792 80 2812
rect 835 2792 893 2793
rect 3619 2792 3677 2793
rect 4099 2792 4157 2793
rect 0 2752 844 2792
rect 884 2752 893 2792
rect 2851 2752 2860 2792
rect 2900 2752 2909 2792
rect 3534 2752 3628 2792
rect 3668 2752 3677 2792
rect 4003 2752 4012 2792
rect 4052 2752 4108 2792
rect 4148 2752 4157 2792
rect 6787 2752 6796 2792
rect 6836 2752 8524 2792
rect 8564 2752 8573 2792
rect 9859 2752 9868 2792
rect 9908 2752 11360 2792
rect 12259 2752 12268 2792
rect 12308 2752 15628 2792
rect 15668 2752 15677 2792
rect 0 2732 80 2752
rect 835 2751 893 2752
rect 2860 2708 2900 2752
rect 3619 2751 3677 2752
rect 4099 2751 4157 2752
rect 7555 2708 7613 2709
rect 8995 2708 9053 2709
rect 2860 2668 6988 2708
rect 7028 2668 7037 2708
rect 7470 2668 7564 2708
rect 7604 2668 7613 2708
rect 8899 2668 8908 2708
rect 8948 2668 9004 2708
rect 9044 2668 9053 2708
rect 7555 2667 7613 2668
rect 8995 2667 9053 2668
rect 9187 2708 9245 2709
rect 11320 2708 11360 2752
rect 11587 2708 11645 2709
rect 14179 2708 14237 2709
rect 14563 2708 14621 2709
rect 9187 2668 9196 2708
rect 9236 2668 9676 2708
rect 9716 2668 9725 2708
rect 11320 2668 11596 2708
rect 11636 2668 11645 2708
rect 14094 2668 14188 2708
rect 14228 2668 14237 2708
rect 14478 2668 14572 2708
rect 14612 2668 14621 2708
rect 9187 2667 9245 2668
rect 11587 2667 11645 2668
rect 14179 2667 14237 2668
rect 14563 2667 14621 2668
rect 6979 2624 7037 2625
rect 2668 2584 4876 2624
rect 4916 2584 6220 2624
rect 6260 2584 6269 2624
rect 6979 2584 6988 2624
rect 7028 2584 7084 2624
rect 7124 2584 7133 2624
rect 9091 2584 9100 2624
rect 9140 2584 10156 2624
rect 10196 2584 10205 2624
rect 10723 2584 10732 2624
rect 10772 2584 11360 2624
rect 2668 2540 2708 2584
rect 6979 2583 7037 2584
rect 3235 2540 3293 2541
rect 8035 2540 8093 2541
rect 8803 2540 8861 2541
rect 2659 2500 2668 2540
rect 2708 2500 2717 2540
rect 3150 2500 3244 2540
rect 3284 2500 3293 2540
rect 6403 2500 6412 2540
rect 6452 2500 6892 2540
rect 6932 2500 6941 2540
rect 7950 2500 8044 2540
rect 8084 2500 8093 2540
rect 8227 2500 8236 2540
rect 8276 2500 8620 2540
rect 8660 2500 8669 2540
rect 8772 2500 8812 2540
rect 8852 2500 8861 2540
rect 11320 2540 11360 2584
rect 11404 2584 11692 2624
rect 11732 2584 11741 2624
rect 12931 2584 12940 2624
rect 12980 2584 13364 2624
rect 14659 2584 14668 2624
rect 14708 2584 15244 2624
rect 15284 2584 15293 2624
rect 17731 2584 17740 2624
rect 17780 2584 18316 2624
rect 18356 2584 18365 2624
rect 19555 2584 19564 2624
rect 19604 2584 19948 2624
rect 19988 2584 19997 2624
rect 11404 2540 11444 2584
rect 11320 2500 11444 2540
rect 3235 2499 3293 2500
rect 8035 2499 8093 2500
rect 8800 2499 8861 2500
rect 0 2456 80 2476
rect 8800 2456 8840 2499
rect 13324 2456 13364 2584
rect 0 2416 8840 2456
rect 9859 2416 9868 2456
rect 9908 2416 13172 2456
rect 13315 2416 13324 2456
rect 13364 2416 13373 2456
rect 14179 2416 14188 2456
rect 14228 2416 14380 2456
rect 14420 2416 14429 2456
rect 0 2396 80 2416
rect 1219 2372 1277 2373
rect 1219 2332 1228 2372
rect 1268 2332 4396 2372
rect 4436 2332 4445 2372
rect 8227 2332 8236 2372
rect 8276 2332 9772 2372
rect 9812 2332 9821 2372
rect 11107 2332 11116 2372
rect 11156 2332 11308 2372
rect 11348 2332 12268 2372
rect 12308 2332 12317 2372
rect 13027 2332 13036 2372
rect 13076 2332 13085 2372
rect 1219 2331 1277 2332
rect 3043 2288 3101 2289
rect 556 2248 3052 2288
rect 3092 2248 3101 2288
rect 0 2120 80 2140
rect 556 2120 596 2248
rect 3043 2247 3101 2248
rect 3235 2288 3293 2289
rect 10243 2288 10301 2289
rect 3235 2248 3244 2288
rect 3284 2248 3378 2288
rect 4919 2248 4928 2288
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 5296 2248 5305 2288
rect 7075 2248 7084 2288
rect 7124 2248 10252 2288
rect 10292 2248 10301 2288
rect 3235 2247 3293 2248
rect 10243 2247 10301 2248
rect 11587 2204 11645 2205
rect 1123 2164 1132 2204
rect 1172 2164 2860 2204
rect 2900 2164 2909 2204
rect 3523 2164 3532 2204
rect 3572 2164 6316 2204
rect 6356 2164 6365 2204
rect 6979 2164 6988 2204
rect 7028 2164 8044 2204
rect 8084 2164 8093 2204
rect 8515 2164 8524 2204
rect 8564 2164 10060 2204
rect 10100 2164 11116 2204
rect 11156 2164 11165 2204
rect 11502 2164 11596 2204
rect 11636 2164 11645 2204
rect 11587 2163 11645 2164
rect 2755 2120 2813 2121
rect 13036 2120 13076 2332
rect 13132 2204 13172 2416
rect 20039 2248 20048 2288
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20416 2248 20425 2288
rect 13891 2204 13949 2205
rect 13132 2164 13900 2204
rect 13940 2164 16492 2204
rect 16532 2164 16541 2204
rect 13891 2163 13949 2164
rect 0 2080 596 2120
rect 2659 2080 2668 2120
rect 2708 2080 2764 2120
rect 2804 2080 2813 2120
rect 3331 2080 3340 2120
rect 3380 2080 6124 2120
rect 6164 2080 6173 2120
rect 6691 2080 6700 2120
rect 6740 2080 8428 2120
rect 8468 2080 8477 2120
rect 11299 2080 11308 2120
rect 11348 2080 11788 2120
rect 11828 2080 11837 2120
rect 12076 2080 15148 2120
rect 15188 2080 15197 2120
rect 0 2060 80 2080
rect 2755 2079 2813 2080
rect 5635 2036 5693 2037
rect 3340 1996 5644 2036
rect 5684 1996 5693 2036
rect 3340 1952 3380 1996
rect 5635 1995 5693 1996
rect 6979 2036 7037 2037
rect 6979 1996 6988 2036
rect 7028 1996 8812 2036
rect 8852 1996 8861 2036
rect 10339 1996 10348 2036
rect 10388 1996 10636 2036
rect 10676 1996 10685 2036
rect 6979 1995 7037 1996
rect 8419 1952 8477 1953
rect 3331 1912 3340 1952
rect 3380 1912 3389 1952
rect 5251 1912 5260 1952
rect 5300 1912 8372 1952
rect 7363 1868 7421 1869
rect 3139 1828 3148 1868
rect 3188 1828 7372 1868
rect 7412 1828 7421 1868
rect 7363 1827 7421 1828
rect 0 1784 80 1804
rect 7267 1784 7325 1785
rect 0 1744 172 1784
rect 212 1744 221 1784
rect 4291 1744 4300 1784
rect 4340 1744 4684 1784
rect 4724 1744 4733 1784
rect 7171 1744 7180 1784
rect 7220 1744 7276 1784
rect 7316 1744 7325 1784
rect 8332 1784 8372 1912
rect 8419 1912 8428 1952
rect 8468 1912 11980 1952
rect 12020 1912 12029 1952
rect 8419 1911 8477 1912
rect 9091 1868 9149 1869
rect 9475 1868 9533 1869
rect 12076 1868 12116 2080
rect 14380 1996 16052 2036
rect 14380 1952 14420 1996
rect 16012 1952 16052 1996
rect 12259 1912 12268 1952
rect 12308 1912 12748 1952
rect 12788 1912 14380 1952
rect 14420 1912 14429 1952
rect 14755 1912 14764 1952
rect 14804 1912 15244 1952
rect 15284 1912 15293 1952
rect 15811 1912 15820 1952
rect 15860 1912 15869 1952
rect 16003 1912 16012 1952
rect 16052 1912 16684 1952
rect 16724 1912 16733 1952
rect 9006 1828 9100 1868
rect 9140 1828 9149 1868
rect 9390 1828 9484 1868
rect 9524 1828 9533 1868
rect 9091 1827 9149 1828
rect 9475 1827 9533 1828
rect 11404 1828 12116 1868
rect 11404 1784 11444 1828
rect 15820 1784 15860 1912
rect 16003 1868 16061 1869
rect 16003 1828 16012 1868
rect 16052 1828 20236 1868
rect 20276 1828 20285 1868
rect 16003 1827 16061 1828
rect 8332 1744 11444 1784
rect 11491 1744 11500 1784
rect 11540 1744 18412 1784
rect 18452 1744 18461 1784
rect 0 1724 80 1744
rect 7267 1743 7325 1744
rect 15427 1700 15485 1701
rect 172 1660 6412 1700
rect 6452 1660 6461 1700
rect 9283 1660 9292 1700
rect 9332 1660 11980 1700
rect 12020 1660 12029 1700
rect 15427 1660 15436 1700
rect 15476 1660 16204 1700
rect 16244 1660 16253 1700
rect 0 1448 80 1468
rect 172 1448 212 1660
rect 15427 1659 15485 1660
rect 4867 1576 4876 1616
rect 4916 1576 15340 1616
rect 15380 1576 15389 1616
rect 3679 1492 3688 1532
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 4056 1492 4065 1532
rect 4675 1492 4684 1532
rect 4724 1492 6508 1532
rect 6548 1492 8428 1532
rect 8468 1492 8477 1532
rect 8899 1492 8908 1532
rect 8948 1492 9580 1532
rect 9620 1492 9629 1532
rect 15427 1492 15436 1532
rect 15476 1492 17164 1532
rect 17204 1492 17213 1532
rect 18799 1492 18808 1532
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 19176 1492 19185 1532
rect 10435 1448 10493 1449
rect 0 1408 212 1448
rect 1411 1408 1420 1448
rect 1460 1408 9772 1448
rect 9812 1408 9821 1448
rect 10435 1408 10444 1448
rect 10484 1408 10636 1448
rect 10676 1408 13460 1448
rect 0 1388 80 1408
rect 10435 1407 10493 1408
rect 2467 1364 2525 1365
rect 2467 1324 2476 1364
rect 2516 1324 4684 1364
rect 4724 1324 4733 1364
rect 4867 1324 4876 1364
rect 4916 1324 7468 1364
rect 7508 1324 7517 1364
rect 7852 1324 11500 1364
rect 11540 1324 11549 1364
rect 2467 1323 2525 1324
rect 2947 1280 3005 1281
rect 4675 1280 4733 1281
rect 7852 1280 7892 1324
rect 12739 1280 12797 1281
rect 2947 1240 2956 1280
rect 2996 1240 3724 1280
rect 3764 1240 3773 1280
rect 4675 1240 4684 1280
rect 4724 1240 4733 1280
rect 5251 1240 5260 1280
rect 5300 1240 7892 1280
rect 7939 1240 7948 1280
rect 7988 1240 8908 1280
rect 8948 1240 8957 1280
rect 9667 1240 9676 1280
rect 9716 1240 12364 1280
rect 12404 1240 12413 1280
rect 12654 1240 12748 1280
rect 12788 1240 12797 1280
rect 2947 1239 3005 1240
rect 4675 1239 4733 1240
rect 12739 1239 12797 1240
rect 13123 1280 13181 1281
rect 13420 1280 13460 1408
rect 13891 1324 13900 1364
rect 13940 1324 15140 1364
rect 15235 1324 15244 1364
rect 15284 1324 16780 1364
rect 16820 1324 18508 1364
rect 18548 1324 18557 1364
rect 15100 1280 15140 1324
rect 17731 1280 17789 1281
rect 18115 1280 18173 1281
rect 18691 1280 18749 1281
rect 13123 1240 13132 1280
rect 13172 1240 13324 1280
rect 13364 1240 13373 1280
rect 13420 1240 13940 1280
rect 15100 1240 17396 1280
rect 17646 1240 17740 1280
rect 17780 1240 17789 1280
rect 18030 1240 18124 1280
rect 18164 1240 18173 1280
rect 18606 1240 18700 1280
rect 18740 1240 18749 1280
rect 13123 1239 13181 1240
rect 4684 1196 4724 1239
rect 10339 1196 10397 1197
rect 13027 1196 13085 1197
rect 13900 1196 13940 1240
rect 17155 1196 17213 1197
rect 2380 1156 4724 1196
rect 6403 1156 6412 1196
rect 6452 1156 7660 1196
rect 7700 1156 7709 1196
rect 8611 1156 8620 1196
rect 8660 1156 10348 1196
rect 10388 1156 10397 1196
rect 11875 1156 11884 1196
rect 11924 1156 12652 1196
rect 12692 1156 12701 1196
rect 13027 1156 13036 1196
rect 13076 1156 13132 1196
rect 13172 1156 13181 1196
rect 13891 1156 13900 1196
rect 13940 1156 15572 1196
rect 17070 1156 17164 1196
rect 17204 1156 17213 1196
rect 0 1112 80 1132
rect 2380 1112 2420 1156
rect 10339 1155 10397 1156
rect 13027 1155 13085 1156
rect 0 1072 2420 1112
rect 2467 1112 2525 1113
rect 3331 1112 3389 1113
rect 6787 1112 6845 1113
rect 2467 1072 2476 1112
rect 2516 1072 2572 1112
rect 2612 1072 2621 1112
rect 2755 1072 2764 1112
rect 2804 1072 3340 1112
rect 3380 1072 3389 1112
rect 0 1052 80 1072
rect 2467 1071 2525 1072
rect 3331 1071 3389 1072
rect 4684 1072 5204 1112
rect 6702 1072 6796 1112
rect 6836 1072 6845 1112
rect 2659 1028 2717 1029
rect 4684 1028 4724 1072
rect 2659 988 2668 1028
rect 2708 988 3148 1028
rect 3188 988 3197 1028
rect 4483 988 4492 1028
rect 4532 988 4724 1028
rect 5164 1028 5204 1072
rect 6787 1071 6845 1072
rect 8323 1112 8381 1113
rect 15532 1112 15572 1156
rect 17155 1155 17213 1156
rect 8323 1072 8332 1112
rect 8372 1072 8428 1112
rect 8468 1072 8477 1112
rect 8707 1072 8716 1112
rect 8756 1072 13996 1112
rect 14036 1072 14045 1112
rect 15523 1072 15532 1112
rect 15572 1072 15820 1112
rect 15860 1072 16300 1112
rect 16340 1072 16349 1112
rect 8323 1071 8381 1072
rect 17356 1028 17396 1240
rect 17731 1239 17789 1240
rect 18115 1239 18173 1240
rect 18691 1239 18749 1240
rect 17539 1196 17597 1197
rect 17454 1156 17548 1196
rect 17588 1156 17597 1196
rect 17539 1155 17597 1156
rect 18019 1196 18077 1197
rect 18019 1156 18028 1196
rect 18068 1156 18316 1196
rect 18356 1156 18365 1196
rect 18019 1155 18077 1156
rect 17635 1072 17644 1112
rect 17684 1072 19660 1112
rect 19700 1072 19709 1112
rect 18307 1028 18365 1029
rect 5164 988 7564 1028
rect 7604 988 7613 1028
rect 9379 988 9388 1028
rect 9428 988 11212 1028
rect 11252 988 11261 1028
rect 17356 988 17588 1028
rect 2659 987 2717 988
rect 4771 944 4829 945
rect 11779 944 11837 945
rect 13315 944 13373 945
rect 13987 944 14045 945
rect 17548 944 17588 988
rect 18307 988 18316 1028
rect 18356 988 19084 1028
rect 19124 988 19133 1028
rect 18307 987 18365 988
rect 1027 904 1036 944
rect 1076 904 2956 944
rect 2996 904 3005 944
rect 4675 904 4684 944
rect 4724 904 4780 944
rect 4820 904 4829 944
rect 5539 904 5548 944
rect 5588 904 10444 944
rect 10484 904 10493 944
rect 11779 904 11788 944
rect 11828 904 12556 944
rect 12596 904 12605 944
rect 12931 904 12940 944
rect 12980 904 13324 944
rect 13364 904 13373 944
rect 13891 904 13900 944
rect 13940 904 13996 944
rect 14036 904 14045 944
rect 14275 904 14284 944
rect 14324 904 17356 944
rect 17396 904 17405 944
rect 17539 904 17548 944
rect 17588 904 17597 944
rect 4771 903 4829 904
rect 11779 903 11837 904
rect 13315 903 13373 904
rect 13987 903 14045 904
rect 739 860 797 861
rect 8227 860 8285 861
rect 14083 860 14141 861
rect 20515 860 20573 861
rect 739 820 748 860
rect 788 820 4492 860
rect 4532 820 4541 860
rect 5347 820 5356 860
rect 5396 820 8236 860
rect 8276 820 8285 860
rect 8803 820 8812 860
rect 8852 820 11884 860
rect 11924 820 11933 860
rect 13507 820 13516 860
rect 13556 820 14092 860
rect 14132 820 14141 860
rect 16003 820 16012 860
rect 16052 820 17644 860
rect 17684 820 17693 860
rect 18499 820 18508 860
rect 18548 820 20524 860
rect 20564 820 20573 860
rect 739 819 797 820
rect 8227 819 8285 820
rect 14083 819 14141 820
rect 20515 819 20573 820
rect 0 776 80 796
rect 1411 776 1469 777
rect 10435 776 10493 777
rect 13699 776 13757 777
rect 15619 776 15677 777
rect 16771 776 16829 777
rect 0 736 1420 776
rect 1460 736 1469 776
rect 4919 736 4928 776
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 5296 736 5305 776
rect 6499 736 6508 776
rect 6548 736 10444 776
rect 10484 736 10493 776
rect 13614 736 13708 776
rect 13748 736 13757 776
rect 15534 736 15628 776
rect 15668 736 15677 776
rect 16686 736 16780 776
rect 16820 736 16829 776
rect 20039 736 20048 776
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20416 736 20425 776
rect 0 716 80 736
rect 1411 735 1469 736
rect 10435 735 10493 736
rect 13699 735 13757 736
rect 15619 735 15677 736
rect 16771 735 16829 736
rect 11875 692 11933 693
rect 18883 692 18941 693
rect 3907 652 3916 692
rect 3956 652 6320 692
rect 6595 652 6604 692
rect 6644 652 11884 692
rect 11924 652 11933 692
rect 18798 652 18892 692
rect 18932 652 18941 692
rect 2947 608 3005 609
rect 6280 608 6320 652
rect 11875 651 11933 652
rect 18883 651 18941 652
rect 2862 568 2956 608
rect 2996 568 3005 608
rect 5059 568 5068 608
rect 5108 568 5932 608
rect 5972 568 5981 608
rect 6280 568 6892 608
rect 6932 568 6941 608
rect 10051 568 10060 608
rect 10100 568 10348 608
rect 10388 568 10397 608
rect 2947 567 3005 568
rect 6979 524 7037 525
rect 3331 484 3340 524
rect 3380 484 6988 524
rect 7028 484 7037 524
rect 8419 484 8428 524
rect 8468 484 8840 524
rect 9283 484 9292 524
rect 9332 484 14188 524
rect 14228 484 14237 524
rect 14851 484 14860 524
rect 14900 484 18028 524
rect 18068 484 18077 524
rect 6979 483 7037 484
rect 0 440 80 460
rect 8419 440 8477 441
rect 0 400 8428 440
rect 8468 400 8477 440
rect 8800 440 8840 484
rect 8800 400 17164 440
rect 17204 400 19564 440
rect 19604 400 19613 440
rect 0 380 80 400
rect 8419 399 8477 400
rect 6979 356 7037 357
rect 6894 316 6988 356
rect 7028 316 7037 356
rect 14659 316 14668 356
rect 14708 316 19948 356
rect 19988 316 19997 356
rect 6979 315 7037 316
rect 3523 272 3581 273
rect 11011 272 11069 273
rect 17347 272 17405 273
rect 172 232 3532 272
rect 3572 232 3581 272
rect 6115 232 6124 272
rect 6164 232 8524 272
rect 8564 232 8573 272
rect 10926 232 11020 272
rect 11060 232 11069 272
rect 15235 232 15244 272
rect 15284 232 16972 272
rect 17012 232 17021 272
rect 17347 232 17356 272
rect 17396 232 19276 272
rect 19316 232 19325 272
rect 0 104 80 124
rect 172 104 212 232
rect 3523 231 3581 232
rect 11011 231 11069 232
rect 17347 231 17405 232
rect 16099 188 16157 189
rect 19459 188 19517 189
rect 1891 148 1900 188
rect 1940 148 1949 188
rect 6211 148 6220 188
rect 6260 148 16108 188
rect 16148 148 16157 188
rect 16675 148 16684 188
rect 16724 148 17012 188
rect 19374 148 19468 188
rect 19508 148 19517 188
rect 0 64 212 104
rect 1900 104 1940 148
rect 16099 147 16157 148
rect 16972 104 17012 148
rect 19459 147 19517 148
rect 1900 64 7948 104
rect 7988 64 7997 104
rect 16963 64 16972 104
rect 17012 64 17021 104
rect 0 44 80 64
<< via3 >>
rect 7276 85660 7316 85700
rect 7756 85576 7796 85616
rect 940 85240 980 85280
rect 8524 84988 8564 85028
rect 3436 84904 3476 84944
rect 7660 84904 7700 84944
rect 12364 84904 12404 84944
rect 12844 84736 12884 84776
rect 2956 84652 2996 84692
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 4780 84652 4820 84692
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 11020 84484 11060 84524
rect 11980 84484 12020 84524
rect 6028 84400 6068 84440
rect 6412 84400 6452 84440
rect 6604 84400 6644 84440
rect 9676 84400 9716 84440
rect 9868 84400 9908 84440
rect 11212 84400 11252 84440
rect 12748 84400 12788 84440
rect 13900 84400 13940 84440
rect 1324 84316 1364 84356
rect 3532 84232 3572 84272
rect 16876 84400 16916 84440
rect 18028 84316 18068 84356
rect 19660 84316 19700 84356
rect 16588 84232 16628 84272
rect 12460 84064 12500 84104
rect 13228 84064 13268 84104
rect 17740 84064 17780 84104
rect 2572 83896 2612 83936
rect 4300 83896 4340 83936
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 10444 83644 10484 83684
rect 10060 83560 10100 83600
rect 1516 83476 1556 83516
rect 3340 83476 3380 83516
rect 10540 83476 10580 83516
rect 16972 83476 17012 83516
rect 8908 83392 8948 83432
rect 9292 83392 9332 83432
rect 12364 83308 12404 83348
rect 13612 83308 13652 83348
rect 14956 83308 14996 83348
rect 16012 83308 16052 83348
rect 6316 83224 6356 83264
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 13996 83140 14036 83180
rect 17452 83140 17492 83180
rect 3340 83056 3380 83096
rect 6316 82972 6356 83012
rect 10444 82972 10484 83012
rect 18412 83140 18452 83180
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 13804 82972 13844 83012
rect 5356 82888 5396 82928
rect 12652 82888 12692 82928
rect 5452 82804 5492 82844
rect 7468 82804 7508 82844
rect 5740 82720 5780 82760
rect 7372 82720 7412 82760
rect 14380 82720 14420 82760
rect 12172 82552 12212 82592
rect 12940 82552 12980 82592
rect 13132 82552 13172 82592
rect 14764 82552 14804 82592
rect 19564 82552 19604 82592
rect 2764 82384 2804 82424
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 11596 82384 11636 82424
rect 11884 82384 11924 82424
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 11980 82300 12020 82340
rect 19564 82300 19604 82340
rect 1324 82216 1364 82256
rect 4108 82132 4148 82172
rect 4780 82132 4820 82172
rect 5356 82132 5396 82172
rect 5836 82132 5876 82172
rect 6508 82132 6548 82172
rect 11788 82132 11828 82172
rect 1036 82048 1076 82088
rect 10348 82048 10388 82088
rect 3820 81964 3860 82004
rect 1804 81880 1844 81920
rect 4780 81880 4820 81920
rect 12652 81880 12692 81920
rect 14380 81880 14420 81920
rect 19276 81880 19316 81920
rect 11980 81796 12020 81836
rect 16396 81796 16436 81836
rect 3532 81712 3572 81752
rect 11596 81712 11636 81752
rect 14764 81712 14804 81752
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 1612 81460 1652 81500
rect 7852 81292 7892 81332
rect 3532 81208 3572 81248
rect 3916 81208 3956 81248
rect 18700 81208 18740 81248
rect 3628 81124 3668 81164
rect 10348 81124 10388 81164
rect 16396 81040 16436 81080
rect 16012 80956 16052 80996
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 17068 80872 17108 80912
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 1324 80788 1364 80828
rect 1900 80788 1940 80828
rect 14860 80620 14900 80660
rect 17932 80536 17972 80576
rect 4780 80452 4820 80492
rect 6988 80452 7028 80492
rect 7468 80452 7508 80492
rect 8044 80452 8084 80492
rect 14284 80452 14324 80492
rect 3148 80368 3188 80408
rect 18604 80368 18644 80408
rect 19948 80368 19988 80408
rect 15820 80284 15860 80324
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 7660 80116 7700 80156
rect 11404 80116 11444 80156
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 4492 80032 4532 80072
rect 5548 80032 5588 80072
rect 18508 80032 18548 80072
rect 19276 79948 19316 79988
rect 1420 79864 1460 79904
rect 5836 79780 5876 79820
rect 8044 79780 8084 79820
rect 17164 79780 17204 79820
rect 1324 79696 1364 79736
rect 1996 79696 2036 79736
rect 4684 79696 4724 79736
rect 6796 79696 6836 79736
rect 8620 79696 8660 79736
rect 18508 79696 18548 79736
rect 17068 79612 17108 79652
rect 18220 79612 18260 79652
rect 652 79528 692 79568
rect 2764 79528 2804 79568
rect 6124 79528 6164 79568
rect 1132 79444 1172 79484
rect 8236 79444 8276 79484
rect 2956 79360 2996 79400
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 6892 79360 6932 79400
rect 10444 79360 10484 79400
rect 10636 79360 10676 79400
rect 11980 79360 12020 79400
rect 17644 79360 17684 79400
rect 19564 79360 19604 79400
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 2284 79276 2324 79316
rect 12556 79276 12596 79316
rect 7180 79192 7220 79232
rect 7948 79192 7988 79232
rect 17356 79192 17396 79232
rect 1324 79108 1364 79148
rect 1612 79024 1652 79064
rect 18316 79108 18356 79148
rect 2476 78940 2516 78980
rect 7180 78940 7220 78980
rect 19276 78940 19316 78980
rect 3340 78856 3380 78896
rect 7084 78856 7124 78896
rect 8236 78856 8276 78896
rect 17260 78856 17300 78896
rect 17068 78688 17108 78728
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 3244 78520 3284 78560
rect 13036 78520 13076 78560
rect 14284 78520 14324 78560
rect 18316 78436 18356 78476
rect 1228 78352 1268 78392
rect 10828 78352 10868 78392
rect 18700 78352 18740 78392
rect 2284 78268 2324 78308
rect 11788 78268 11828 78308
rect 18028 78268 18068 78308
rect 8428 78184 8468 78224
rect 15724 78184 15764 78224
rect 4684 78100 4724 78140
rect 15532 78100 15572 78140
rect 1996 78016 2036 78056
rect 10444 77932 10484 77972
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 9580 77848 9620 77888
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 1996 77764 2036 77804
rect 1900 77680 1940 77720
rect 17356 77680 17396 77720
rect 18220 77680 18260 77720
rect 13324 77596 13364 77636
rect 1324 77512 1364 77552
rect 17068 77512 17108 77552
rect 3532 77428 3572 77468
rect 4204 77428 4244 77468
rect 10636 77428 10676 77468
rect 17164 77428 17204 77468
rect 1612 77344 1652 77384
rect 2380 77344 2420 77384
rect 18316 77344 18356 77384
rect 15052 77260 15092 77300
rect 2092 77176 2132 77216
rect 2860 77092 2900 77132
rect 3244 77092 3284 77132
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 10828 77092 10868 77132
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 3532 77008 3572 77048
rect 4108 76924 4148 76964
rect 17932 76924 17972 76964
rect 3436 76840 3476 76880
rect 8236 76840 8276 76880
rect 10444 76840 10484 76880
rect 17452 76840 17492 76880
rect 19276 76840 19316 76880
rect 5356 76756 5396 76796
rect 1420 76672 1460 76712
rect 2188 76672 2228 76712
rect 3244 76672 3284 76712
rect 10156 76672 10196 76712
rect 2092 76588 2132 76628
rect 2572 76504 2612 76544
rect 8332 76504 8372 76544
rect 16300 76504 16340 76544
rect 2380 76420 2420 76460
rect 2572 76336 2612 76376
rect 4780 76336 4820 76376
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 8428 76336 8468 76376
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 18028 76252 18068 76292
rect 19660 76252 19700 76292
rect 1804 76168 1844 76208
rect 6700 76168 6740 76208
rect 18412 76168 18452 76208
rect 1420 76084 1460 76124
rect 1324 76000 1364 76040
rect 1804 76000 1844 76040
rect 15532 76000 15572 76040
rect 19948 75748 19988 75788
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 1900 75496 1940 75536
rect 13420 75580 13460 75620
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 7564 75496 7604 75536
rect 4300 75412 4340 75452
rect 1420 75244 1460 75284
rect 3340 75244 3380 75284
rect 17260 75244 17300 75284
rect 2764 75160 2804 75200
rect 12556 75160 12596 75200
rect 15724 75160 15764 75200
rect 1228 74992 1268 75032
rect 4108 74992 4148 75032
rect 18700 74992 18740 75032
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 9196 74824 9236 74864
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 7756 74572 7796 74612
rect 15436 74572 15476 74612
rect 2764 74488 2804 74528
rect 3340 74404 3380 74444
rect 10732 74404 10772 74444
rect 17932 74404 17972 74444
rect 1708 74320 1748 74360
rect 3436 74236 3476 74276
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 16204 74068 16244 74108
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 14284 73984 14324 74024
rect 10444 73816 10484 73856
rect 8620 73648 8660 73688
rect 6892 73564 6932 73604
rect 7660 73480 7700 73520
rect 2956 73396 2996 73436
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 8236 73312 8276 73352
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 10444 73228 10484 73268
rect 652 73144 692 73184
rect 1132 73060 1172 73100
rect 12460 73144 12500 73184
rect 3148 73060 3188 73100
rect 10636 73060 10676 73100
rect 2380 72976 2420 73016
rect 13516 73144 13556 73184
rect 1324 72892 1364 72932
rect 13516 72808 13556 72848
rect 19660 72724 19700 72764
rect 3244 72640 3284 72680
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 9388 72388 9428 72428
rect 3436 72304 3476 72344
rect 460 72052 500 72092
rect 2668 71968 2708 72008
rect 11884 72220 11924 72260
rect 18412 72136 18452 72176
rect 19276 72052 19316 72092
rect 7948 71968 7988 72008
rect 17452 71968 17492 72008
rect 3532 71800 3572 71840
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 11212 71800 11252 71840
rect 12556 71800 12596 71840
rect 13228 71800 13268 71840
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 21388 71800 21428 71840
rect 10156 71716 10196 71756
rect 13804 71716 13844 71756
rect 13420 71632 13460 71672
rect 13324 71464 13364 71504
rect 14572 71464 14612 71504
rect 20812 71464 20852 71504
rect 1324 71296 1364 71336
rect 16204 71380 16244 71420
rect 4780 71296 4820 71336
rect 17644 71296 17684 71336
rect 9772 71212 9812 71252
rect 19852 71212 19892 71252
rect 1804 71128 1844 71168
rect 13228 71128 13268 71168
rect 13804 71128 13844 71168
rect 16780 71128 16820 71168
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 14380 71044 14420 71084
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 19564 71044 19604 71084
rect 3532 70876 3572 70916
rect 7852 70876 7892 70916
rect 8620 70876 8660 70916
rect 3340 70792 3380 70832
rect 5644 70792 5684 70832
rect 6988 70708 7028 70748
rect 15148 70792 15188 70832
rect 19660 70708 19700 70748
rect 7948 70624 7988 70664
rect 12556 70624 12596 70664
rect 4300 70540 4340 70580
rect 9004 70540 9044 70580
rect 15052 70540 15092 70580
rect 15532 70540 15572 70580
rect 20716 70456 20756 70496
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 18220 70288 18260 70328
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 11308 70204 11348 70244
rect 5356 70120 5396 70160
rect 7180 70120 7220 70160
rect 11212 70120 11252 70160
rect 14572 70120 14612 70160
rect 9484 70036 9524 70076
rect 4300 69952 4340 69992
rect 17836 70120 17876 70160
rect 19948 70036 19988 70076
rect 18508 69952 18548 69992
rect 11596 69868 11636 69908
rect 14572 69784 14612 69824
rect 19276 69784 19316 69824
rect 16108 69700 16148 69740
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 20620 69448 20660 69488
rect 2284 69364 2324 69404
rect 13612 69280 13652 69320
rect 17644 69196 17684 69236
rect 2092 69112 2132 69152
rect 2380 69112 2420 69152
rect 3148 69112 3188 69152
rect 19564 69028 19604 69068
rect 172 68944 212 68984
rect 6892 68944 6932 68984
rect 19276 68944 19316 68984
rect 3244 68860 3284 68900
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 2860 68692 2900 68732
rect 3340 68692 3380 68732
rect 13804 68692 13844 68732
rect 2860 68524 2900 68564
rect 11884 68524 11924 68564
rect 6316 68440 6356 68480
rect 6892 68440 6932 68480
rect 20908 68440 20948 68480
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 268 67936 308 67976
rect 13516 67936 13556 67976
rect 13996 67936 14036 67976
rect 5164 67768 5204 67808
rect 9100 67684 9140 67724
rect 11596 67684 11636 67724
rect 18220 67684 18260 67724
rect 76 67600 116 67640
rect 1036 67600 1076 67640
rect 5932 67600 5972 67640
rect 15916 67600 15956 67640
rect 6412 67516 6452 67556
rect 2668 67348 2708 67388
rect 17356 67348 17396 67388
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 11212 67264 11252 67304
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 1516 67096 1556 67136
rect 7660 67096 7700 67136
rect 16204 67012 16244 67052
rect 19660 67012 19700 67052
rect 16684 66928 16724 66968
rect 844 66760 884 66800
rect 7276 66760 7316 66800
rect 19756 66760 19796 66800
rect 1804 66676 1844 66716
rect 6700 66676 6740 66716
rect 8908 66676 8948 66716
rect 9100 66676 9140 66716
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 2284 66424 2324 66464
rect 7564 66424 7604 66464
rect 8332 66424 8372 66464
rect 7276 66340 7316 66380
rect 3340 66088 3380 66128
rect 6988 66004 7028 66044
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 14188 66424 14228 66464
rect 18508 66340 18548 66380
rect 17068 66004 17108 66044
rect 8332 65920 8372 65960
rect 7180 65836 7220 65876
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 7276 65752 7316 65792
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 1420 65668 1460 65708
rect 3148 65584 3188 65624
rect 3340 65416 3380 65456
rect 9388 65416 9428 65456
rect 11596 65416 11636 65456
rect 11980 65416 12020 65456
rect 15532 65416 15572 65456
rect 1708 65332 1748 65372
rect 16588 65248 16628 65288
rect 13228 65164 13268 65204
rect 17164 65164 17204 65204
rect 14476 65080 14516 65120
rect 21196 65080 21236 65120
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 14956 64912 14996 64952
rect 12556 64828 12596 64868
rect 20524 64828 20564 64868
rect 21004 64744 21044 64784
rect 2668 64660 2708 64700
rect 2188 64576 2228 64616
rect 15724 64660 15764 64700
rect 7564 64576 7604 64616
rect 19948 64576 19988 64616
rect 2476 64492 2516 64532
rect 6316 64408 6356 64448
rect 8140 64408 8180 64448
rect 11020 64408 11060 64448
rect 13228 64408 13268 64448
rect 19276 64408 19316 64448
rect 1036 64324 1076 64364
rect 6028 64324 6068 64364
rect 6892 64324 6932 64364
rect 16396 64324 16436 64364
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 8524 64240 8564 64280
rect 9100 64240 9140 64280
rect 11500 64240 11540 64280
rect 15820 64240 15860 64280
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 17260 64156 17300 64196
rect 17932 64072 17972 64112
rect 5836 63904 5876 63944
rect 17548 63904 17588 63944
rect 10540 63820 10580 63860
rect 14284 63736 14324 63776
rect 10828 63568 10868 63608
rect 18220 63568 18260 63608
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 8332 63484 8372 63524
rect 8524 63484 8564 63524
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 844 63400 884 63440
rect 19276 63400 19316 63440
rect 460 63232 500 63272
rect 1420 63232 1460 63272
rect 1996 63232 2036 63272
rect 9388 63232 9428 63272
rect 10348 63316 10388 63356
rect 10252 63232 10292 63272
rect 3436 63148 3476 63188
rect 8524 63148 8564 63188
rect 4396 63064 4436 63104
rect 6028 63064 6068 63104
rect 18508 63064 18548 63104
rect 16972 62980 17012 63020
rect 7756 62896 7796 62936
rect 460 62812 500 62852
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 5356 62728 5396 62768
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 4300 62644 4340 62684
rect 5836 62644 5876 62684
rect 9964 62644 10004 62684
rect 8620 62560 8660 62600
rect 14572 62560 14612 62600
rect 16876 62560 16916 62600
rect 1708 62476 1748 62516
rect 9964 62476 10004 62516
rect 15340 62308 15380 62348
rect 20236 62392 20276 62432
rect 3244 61972 3284 62012
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 3436 61888 3476 61928
rect 4396 61888 4436 61928
rect 11212 61888 11252 61928
rect 4588 61804 4628 61844
rect 17644 61804 17684 61844
rect 1132 61720 1172 61760
rect 4300 61720 4340 61760
rect 11500 61720 11540 61760
rect 11980 61720 12020 61760
rect 652 61636 692 61676
rect 4204 61636 4244 61676
rect 2764 61552 2804 61592
rect 3244 61552 3284 61592
rect 19468 61552 19508 61592
rect 15628 61468 15668 61508
rect 19852 61468 19892 61508
rect 10636 61384 10676 61424
rect 20716 61384 20756 61424
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 13228 61216 13268 61256
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 14860 61132 14900 61172
rect 6028 61048 6068 61088
rect 7564 61048 7604 61088
rect 9196 60964 9236 61004
rect 7564 60880 7604 60920
rect 8140 60880 8180 60920
rect 6988 60628 7028 60668
rect 7564 60544 7604 60584
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 13324 60460 13364 60500
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 14860 60376 14900 60416
rect 13228 60292 13268 60332
rect 6028 60208 6068 60248
rect 7756 60208 7796 60248
rect 3340 60124 3380 60164
rect 11020 60124 11060 60164
rect 11212 60124 11252 60164
rect 4108 60040 4148 60080
rect 12076 60040 12116 60080
rect 15916 60208 15956 60248
rect 4108 59872 4148 59912
rect 12460 59872 12500 59912
rect 12652 59872 12692 59912
rect 15820 59872 15860 59912
rect 11212 59788 11252 59828
rect 19948 59788 19988 59828
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 11980 59704 12020 59744
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 7276 59620 7316 59660
rect 11788 59452 11828 59492
rect 19564 59452 19604 59492
rect 4588 59368 4628 59408
rect 14668 59368 14708 59408
rect 19276 59368 19316 59408
rect 4204 59284 4244 59324
rect 4396 59284 4436 59324
rect 3148 59200 3188 59240
rect 6892 59200 6932 59240
rect 8524 59200 8564 59240
rect 9100 59200 9140 59240
rect 14860 59200 14900 59240
rect 12268 59032 12308 59072
rect 268 58948 308 58988
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 14092 58864 14132 58904
rect 10348 58696 10388 58736
rect 8332 58612 8372 58652
rect 8524 58612 8564 58652
rect 19276 58612 19316 58652
rect 15724 58528 15764 58568
rect 8140 58444 8180 58484
rect 8716 58444 8756 58484
rect 4108 58276 4148 58316
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 12364 58108 12404 58148
rect 19852 58024 19892 58064
rect 8236 57940 8276 57980
rect 16492 57940 16532 57980
rect 17644 57940 17684 57980
rect 1324 57856 1364 57896
rect 4204 57856 4244 57896
rect 8140 57856 8180 57896
rect 3244 57688 3284 57728
rect 4588 57688 4628 57728
rect 15340 57688 15380 57728
rect 11500 57520 11540 57560
rect 11788 57520 11828 57560
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 7660 57436 7700 57476
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 13996 57352 14036 57392
rect 20716 57352 20756 57392
rect 7276 57268 7316 57308
rect 3436 57184 3476 57224
rect 6988 57184 7028 57224
rect 7756 57184 7796 57224
rect 11788 56932 11828 56972
rect 13708 56764 13748 56804
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 7948 56680 7988 56720
rect 12364 56680 12404 56720
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 8716 56596 8756 56636
rect 14764 56596 14804 56636
rect 15724 56512 15764 56552
rect 16972 56260 17012 56300
rect 2764 56176 2804 56216
rect 14764 56176 14804 56216
rect 13996 56092 14036 56132
rect 14572 56092 14612 56132
rect 19948 56092 19988 56132
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 11500 55924 11540 55964
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 3244 55672 3284 55712
rect 8716 55672 8756 55712
rect 13420 55672 13460 55712
rect 12652 55588 12692 55628
rect 17644 55588 17684 55628
rect 7660 55504 7700 55544
rect 11596 55504 11636 55544
rect 14092 55504 14132 55544
rect 13420 55420 13460 55460
rect 8524 55252 8564 55292
rect 16972 55504 17012 55544
rect 13708 55252 13748 55292
rect 15340 55252 15380 55292
rect 16012 55252 16052 55292
rect 18124 55252 18164 55292
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 16396 55168 16436 55208
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 7756 54916 7796 54956
rect 14092 55084 14132 55124
rect 16012 55084 16052 55124
rect 19948 55000 19988 55040
rect 14092 54916 14132 54956
rect 1420 54832 1460 54872
rect 14476 54832 14516 54872
rect 11500 54748 11540 54788
rect 14668 54748 14708 54788
rect 15340 54748 15380 54788
rect 16396 54748 16436 54788
rect 8140 54664 8180 54704
rect 16588 54664 16628 54704
rect 3436 54580 3476 54620
rect 12460 54580 12500 54620
rect 1612 54496 1652 54536
rect 556 54412 596 54452
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 6028 54412 6068 54452
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 8140 54328 8180 54368
rect 13996 54160 14036 54200
rect 16108 54160 16148 54200
rect 19660 54160 19700 54200
rect 20524 54160 20564 54200
rect 2476 54076 2516 54116
rect 2764 54076 2804 54116
rect 11500 54076 11540 54116
rect 2380 53992 2420 54032
rect 7660 53992 7700 54032
rect 8332 53992 8372 54032
rect 10828 53992 10868 54032
rect 16972 53992 17012 54032
rect 17548 53740 17588 53780
rect 19372 53740 19412 53780
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 14284 53656 14324 53696
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 16396 53572 16436 53612
rect 3244 53488 3284 53528
rect 8716 53488 8756 53528
rect 12748 53488 12788 53528
rect 14956 53488 14996 53528
rect 4396 53320 4436 53360
rect 11500 53236 11540 53276
rect 13228 53236 13268 53276
rect 14284 53236 14324 53276
rect 11116 53152 11156 53192
rect 12460 53152 12500 53192
rect 14092 53152 14132 53192
rect 4588 52984 4628 53024
rect 12748 52984 12788 53024
rect 15052 52984 15092 53024
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 17740 52900 17780 52940
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 19852 52900 19892 52940
rect 13228 52816 13268 52856
rect 15628 52816 15668 52856
rect 19948 52816 19988 52856
rect 5068 52732 5108 52772
rect 19468 52732 19508 52772
rect 7852 52564 7892 52604
rect 6892 52480 6932 52520
rect 1612 52312 1652 52352
rect 16588 52312 16628 52352
rect 19468 52312 19508 52352
rect 11692 52228 11732 52268
rect 16108 52228 16148 52268
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 10540 52144 10580 52184
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 2380 52060 2420 52100
rect 2956 52060 2996 52100
rect 15724 52060 15764 52100
rect 16492 52060 16532 52100
rect 16588 51892 16628 51932
rect 20908 51892 20948 51932
rect 1900 51724 1940 51764
rect 6028 51724 6068 51764
rect 940 51640 980 51680
rect 8332 51724 8372 51764
rect 13420 51724 13460 51764
rect 16972 51724 17012 51764
rect 18508 51724 18548 51764
rect 19564 51472 19604 51512
rect 21004 51472 21044 51512
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 172 51304 212 51344
rect 15052 51304 15092 51344
rect 4396 51136 4436 51176
rect 4588 51136 4628 51176
rect 4108 50884 4148 50924
rect 10348 50884 10388 50924
rect 19276 50884 19316 50924
rect 4396 50716 4436 50756
rect 6028 50716 6068 50756
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 11692 50632 11732 50672
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 17740 50380 17780 50420
rect 19276 50296 19316 50336
rect 1708 50212 1748 50252
rect 76 49960 116 50000
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 20140 49876 20180 49916
rect 1900 49708 1940 49748
rect 15628 49708 15668 49748
rect 10444 49624 10484 49664
rect 20716 49624 20756 49664
rect 9676 49456 9716 49496
rect 18604 49288 18644 49328
rect 20524 49288 20564 49328
rect 13708 49204 13748 49244
rect 14476 49204 14516 49244
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 10444 49120 10484 49160
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 14668 48952 14708 48992
rect 15724 48952 15764 48992
rect 10348 48784 10388 48824
rect 13228 48784 13268 48824
rect 16588 48784 16628 48824
rect 15724 48700 15764 48740
rect 20908 48616 20948 48656
rect 1996 48448 2036 48488
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 19468 48196 19508 48236
rect 3148 48112 3188 48152
rect 8716 48028 8756 48068
rect 3148 47944 3188 47984
rect 18508 47860 18548 47900
rect 16300 47692 16340 47732
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 1900 47272 1940 47312
rect 4108 47272 4148 47312
rect 16588 47272 16628 47312
rect 20716 47272 20756 47312
rect 10828 47188 10868 47228
rect 8332 47104 8372 47144
rect 7852 47020 7892 47060
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 13420 46852 13460 46892
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 1132 46684 1172 46724
rect 940 46600 980 46640
rect 2764 46516 2804 46556
rect 6892 46432 6932 46472
rect 10540 46432 10580 46472
rect 11884 46432 11924 46472
rect 15724 46432 15764 46472
rect 7756 46348 7796 46388
rect 9772 46264 9812 46304
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 7852 45760 7892 45800
rect 12556 45508 12596 45548
rect 19948 45508 19988 45548
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 8140 45340 8180 45380
rect 11980 45340 12020 45380
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 17164 45256 17204 45296
rect 15916 45172 15956 45212
rect 10540 45088 10580 45128
rect 16108 45004 16148 45044
rect 7948 44920 7988 44960
rect 10636 44920 10676 44960
rect 18508 44920 18548 44960
rect 20140 44920 20180 44960
rect 8332 44836 8372 44876
rect 4108 44752 4148 44792
rect 10924 44668 10964 44708
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 13804 44500 13844 44540
rect 10156 44416 10196 44456
rect 8236 44164 8276 44204
rect 12460 44164 12500 44204
rect 15052 44164 15092 44204
rect 17356 44080 17396 44120
rect 19468 43996 19508 44036
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 2092 43744 2132 43784
rect 2476 43660 2516 43700
rect 6892 43660 6932 43700
rect 18412 43660 18452 43700
rect 19756 43660 19796 43700
rect 4780 43492 4820 43532
rect 2188 43324 2228 43364
rect 4108 43240 4148 43280
rect 12364 43240 12404 43280
rect 20908 43240 20948 43280
rect 7372 43156 7412 43196
rect 18604 43156 18644 43196
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 2380 42988 2420 43028
rect 6220 42988 6260 43028
rect 6508 42820 6548 42860
rect 14188 42820 14228 42860
rect 20044 42820 20084 42860
rect 21196 42820 21236 42860
rect 1324 42736 1364 42776
rect 2476 42736 2516 42776
rect 16588 42736 16628 42776
rect 21388 42736 21428 42776
rect 8524 42652 8564 42692
rect 10924 42652 10964 42692
rect 9676 42568 9716 42608
rect 15148 42568 15188 42608
rect 16780 42568 16820 42608
rect 17932 42568 17972 42608
rect 21004 42568 21044 42608
rect 17548 42484 17588 42524
rect 19948 42484 19988 42524
rect 11116 42400 11156 42440
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 17260 42316 17300 42356
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 4204 42148 4244 42188
rect 4492 42148 4532 42188
rect 7852 42148 7892 42188
rect 8524 42148 8564 42188
rect 15532 42148 15572 42188
rect 17836 42148 17876 42188
rect 19372 42148 19412 42188
rect 7756 41980 7796 42020
rect 10348 41980 10388 42020
rect 20812 42148 20852 42188
rect 3244 41896 3284 41936
rect 11020 41896 11060 41936
rect 13708 41896 13748 41936
rect 9772 41812 9812 41852
rect 10252 41812 10292 41852
rect 7180 41728 7220 41768
rect 7660 41728 7700 41768
rect 8716 41728 8756 41768
rect 17164 41728 17204 41768
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 8908 41560 8948 41600
rect 10444 41644 10484 41684
rect 16396 41560 16436 41600
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 4300 41476 4340 41516
rect 1996 41392 2036 41432
rect 6892 41392 6932 41432
rect 9772 41476 9812 41516
rect 17836 41476 17876 41516
rect 4108 41140 4148 41180
rect 4684 41056 4724 41096
rect 6892 41056 6932 41096
rect 8908 41056 8948 41096
rect 7660 40972 7700 41012
rect 9196 40972 9236 41012
rect 3436 40888 3476 40928
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 4204 40720 4244 40760
rect 8812 40888 8852 40928
rect 15052 41392 15092 41432
rect 20620 41392 20660 41432
rect 12652 41056 12692 41096
rect 14860 40972 14900 41012
rect 16108 40888 16148 40928
rect 8716 40720 8756 40760
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 6508 40636 6548 40676
rect 9196 40636 9236 40676
rect 10924 40636 10964 40676
rect 13516 40636 13556 40676
rect 7372 40552 7412 40592
rect 8236 40552 8276 40592
rect 13228 40552 13268 40592
rect 2956 40468 2996 40508
rect 3436 40468 3476 40508
rect 6892 40468 6932 40508
rect 20620 40552 20660 40592
rect 7180 40468 7220 40508
rect 11500 40468 11540 40508
rect 10348 40384 10388 40424
rect 3340 40300 3380 40340
rect 14092 40300 14132 40340
rect 14284 40300 14324 40340
rect 15052 40300 15092 40340
rect 19468 40300 19508 40340
rect 8908 40216 8948 40256
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 16108 40048 16148 40088
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 7852 39880 7892 39920
rect 8236 39880 8276 39920
rect 14188 39880 14228 39920
rect 4300 39712 4340 39752
rect 4684 39712 4724 39752
rect 8716 39712 8756 39752
rect 17932 39880 17972 39920
rect 8908 39544 8948 39584
rect 19372 39460 19412 39500
rect 1612 39376 1652 39416
rect 2092 39376 2132 39416
rect 6892 39376 6932 39416
rect 8812 39376 8852 39416
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 12556 39292 12596 39332
rect 13708 39292 13748 39332
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 9772 39208 9812 39248
rect 10252 39208 10292 39248
rect 20716 39208 20756 39248
rect 14188 39124 14228 39164
rect 18220 39124 18260 39164
rect 2380 39040 2420 39080
rect 6220 39040 6260 39080
rect 7180 39040 7220 39080
rect 10156 39040 10196 39080
rect 3052 38956 3092 38996
rect 4108 38956 4148 38996
rect 4780 38872 4820 38912
rect 18220 38872 18260 38912
rect 19468 38872 19508 38912
rect 4204 38788 4244 38828
rect 7468 38788 7508 38828
rect 13228 38788 13268 38828
rect 16300 38788 16340 38828
rect 19276 38788 19316 38828
rect 8716 38704 8756 38744
rect 4492 38620 4532 38660
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 1420 38452 1460 38492
rect 3340 38452 3380 38492
rect 19756 38452 19796 38492
rect 4684 38368 4724 38408
rect 5836 38368 5876 38408
rect 12556 38368 12596 38408
rect 19564 38368 19604 38408
rect 10252 38284 10292 38324
rect 12652 38284 12692 38324
rect 13420 38284 13460 38324
rect 20812 38284 20852 38324
rect 17836 38200 17876 38240
rect 19852 38200 19892 38240
rect 1996 38116 2036 38156
rect 2380 38116 2420 38156
rect 10252 38116 10292 38156
rect 2668 38032 2708 38072
rect 19948 38032 19988 38072
rect 9676 37864 9716 37904
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 1228 37696 1268 37736
rect 6028 37696 6068 37736
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 3820 37612 3860 37652
rect 20620 37612 20660 37652
rect 5356 37528 5396 37568
rect 6316 37444 6356 37484
rect 3244 37360 3284 37400
rect 4108 37276 4148 37316
rect 5644 37276 5684 37316
rect 9196 37276 9236 37316
rect 16204 37276 16244 37316
rect 7948 37108 7988 37148
rect 15724 37108 15764 37148
rect 17068 37108 17108 37148
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 11212 37024 11252 37064
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 6988 36856 7028 36896
rect 748 36772 788 36812
rect 5836 36688 5876 36728
rect 19372 36688 19412 36728
rect 12748 36604 12788 36644
rect 9100 36520 9140 36560
rect 16684 36520 16724 36560
rect 19276 36520 19316 36560
rect 2764 36352 2804 36392
rect 10444 36352 10484 36392
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 18412 36268 18452 36308
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 9868 36184 9908 36224
rect 9388 36016 9428 36056
rect 17068 36016 17108 36056
rect 7852 35848 7892 35888
rect 8620 35848 8660 35888
rect 17452 35848 17492 35888
rect 7468 35680 7508 35720
rect 11020 35680 11060 35720
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 5836 35512 5876 35552
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 8428 35344 8468 35384
rect 3532 35260 3572 35300
rect 8620 35260 8660 35300
rect 9676 35260 9716 35300
rect 19756 35260 19796 35300
rect 16876 35176 16916 35216
rect 12748 35092 12788 35132
rect 14764 34924 14804 34964
rect 11212 34840 11252 34880
rect 15628 34840 15668 34880
rect 18412 34840 18452 34880
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 16876 34756 16916 34796
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 2188 34672 2228 34712
rect 6892 34672 6932 34712
rect 20620 34672 20660 34712
rect 8812 34588 8852 34628
rect 20716 34588 20756 34628
rect 7756 34336 7796 34376
rect 12364 34336 12404 34376
rect 13420 34336 13460 34376
rect 21388 34336 21428 34376
rect 6700 34252 6740 34292
rect 7372 34252 7412 34292
rect 16780 34252 16820 34292
rect 10540 34168 10580 34208
rect 11308 34168 11348 34208
rect 1420 34084 1460 34124
rect 6028 34084 6068 34124
rect 4684 34000 4724 34040
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 8524 34000 8564 34040
rect 16780 34000 16820 34040
rect 17164 34000 17204 34040
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 14476 33916 14516 33956
rect 4012 33832 4052 33872
rect 8236 33832 8276 33872
rect 1996 33664 2036 33704
rect 2188 33664 2228 33704
rect 8428 33664 8468 33704
rect 11020 33664 11060 33704
rect 16588 33664 16628 33704
rect 6412 33580 6452 33620
rect 2764 33496 2804 33536
rect 8428 33496 8468 33536
rect 9100 33496 9140 33536
rect 18508 33496 18548 33536
rect 4684 33412 4724 33452
rect 8236 33412 8276 33452
rect 8812 33328 8852 33368
rect 9964 33328 10004 33368
rect 10156 33328 10196 33368
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 4684 32992 4724 33032
rect 8620 32992 8660 33032
rect 9388 32992 9428 33032
rect 13708 32992 13748 33032
rect 15244 32992 15284 33032
rect 18508 32908 18548 32948
rect 3244 32824 3284 32864
rect 17932 32824 17972 32864
rect 6892 32740 6932 32780
rect 8524 32740 8564 32780
rect 9388 32740 9428 32780
rect 14668 32740 14708 32780
rect 15532 32740 15572 32780
rect 5836 32656 5876 32696
rect 7468 32656 7508 32696
rect 10540 32656 10580 32696
rect 11500 32656 11540 32696
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 7756 32320 7796 32360
rect 15148 32320 15188 32360
rect 3532 32236 3572 32276
rect 8524 32236 8564 32276
rect 3052 32152 3092 32192
rect 1900 32068 1940 32108
rect 11020 32152 11060 32192
rect 15052 32152 15092 32192
rect 7564 32068 7604 32108
rect 5644 31900 5684 31940
rect 11308 31900 11348 31940
rect 1612 31816 1652 31856
rect 4588 31816 4628 31856
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 9868 31732 9908 31772
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 15244 31648 15284 31688
rect 14572 31480 14612 31520
rect 17548 31480 17588 31520
rect 20620 31480 20660 31520
rect 1612 31396 1652 31436
rect 14188 31396 14228 31436
rect 14668 31396 14708 31436
rect 18508 31396 18548 31436
rect 4204 31312 4244 31352
rect 11500 31312 11540 31352
rect 17644 31312 17684 31352
rect 5740 31228 5780 31268
rect 6508 31228 6548 31268
rect 8428 31228 8468 31268
rect 8716 31228 8756 31268
rect 7756 31144 7796 31184
rect 8908 31144 8948 31184
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 13516 30976 13556 31016
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 2764 30556 2804 30596
rect 9676 30724 9716 30764
rect 7852 30640 7892 30680
rect 11020 30640 11060 30680
rect 15148 30640 15188 30680
rect 18604 30640 18644 30680
rect 14572 30472 14612 30512
rect 2764 30388 2804 30428
rect 7756 30388 7796 30428
rect 14668 30304 14708 30344
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 5644 30220 5684 30260
rect 6508 30220 6548 30260
rect 14380 30220 14420 30260
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 2092 30136 2132 30176
rect 19756 30052 19796 30092
rect 13516 29968 13556 30008
rect 2956 29884 2996 29924
rect 6892 29884 6932 29924
rect 4300 29800 4340 29840
rect 6316 29800 6356 29840
rect 12748 29800 12788 29840
rect 9868 29716 9908 29756
rect 4108 29632 4148 29672
rect 14188 29632 14228 29672
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 6796 29380 6836 29420
rect 2476 29296 2516 29336
rect 6700 29296 6740 29336
rect 13804 29296 13844 29336
rect 14284 29296 14324 29336
rect 14956 29296 14996 29336
rect 1132 29212 1172 29252
rect 5356 29128 5396 29168
rect 5836 29128 5876 29168
rect 9388 29128 9428 29168
rect 9868 29128 9908 29168
rect 7852 29044 7892 29084
rect 14284 29044 14324 29084
rect 14476 29044 14516 29084
rect 13516 28960 13556 29000
rect 14956 28960 14996 29000
rect 13804 28876 13844 28916
rect 14860 28876 14900 28916
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 6316 28708 6356 28748
rect 14764 28708 14804 28748
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 5644 28624 5684 28664
rect 9964 28624 10004 28664
rect 6412 28540 6452 28580
rect 3148 28456 3188 28496
rect 5836 28372 5876 28412
rect 11500 28372 11540 28412
rect 7372 28288 7412 28328
rect 12748 28288 12788 28328
rect 14860 28288 14900 28328
rect 15628 28288 15668 28328
rect 16684 28288 16724 28328
rect 19276 28288 19316 28328
rect 16300 28204 16340 28244
rect 6796 28120 6836 28160
rect 14764 28120 14804 28160
rect 5740 28036 5780 28076
rect 6508 28036 6548 28076
rect 2956 27952 2996 27992
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 7372 27952 7412 27992
rect 7756 27952 7796 27992
rect 19468 27952 19508 27992
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 12268 27868 12308 27908
rect 12556 27868 12596 27908
rect 14380 27868 14420 27908
rect 4588 27700 4628 27740
rect 8812 27700 8852 27740
rect 13228 27700 13268 27740
rect 2476 27616 2516 27656
rect 5644 27616 5684 27656
rect 14860 27700 14900 27740
rect 16300 27700 16340 27740
rect 9772 27616 9812 27656
rect 14476 27616 14516 27656
rect 15244 27532 15284 27572
rect 16588 27532 16628 27572
rect 4204 27364 4244 27404
rect 7180 27364 7220 27404
rect 7564 27448 7604 27488
rect 10252 27448 10292 27488
rect 11500 27448 11540 27488
rect 15820 27448 15860 27488
rect 9004 27364 9044 27404
rect 15916 27364 15956 27404
rect 1132 27280 1172 27320
rect 12556 27280 12596 27320
rect 2860 27196 2900 27236
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 11500 27112 11540 27152
rect 15148 27196 15188 27236
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 15052 27112 15092 27152
rect 652 27028 692 27068
rect 11404 27028 11444 27068
rect 12364 27028 12404 27068
rect 14284 27028 14324 27068
rect 3148 26944 3188 26984
rect 6508 26944 6548 26984
rect 6220 26860 6260 26900
rect 6412 26860 6452 26900
rect 9676 26860 9716 26900
rect 14860 26860 14900 26900
rect 17836 26860 17876 26900
rect 2860 26776 2900 26816
rect 3244 26776 3284 26816
rect 4492 26776 4532 26816
rect 12556 26776 12596 26816
rect 15820 26776 15860 26816
rect 17068 26776 17108 26816
rect 19276 26692 19316 26732
rect 6316 26608 6356 26648
rect 11308 26608 11348 26648
rect 16684 26608 16724 26648
rect 6892 26524 6932 26564
rect 11500 26524 11540 26564
rect 3148 26440 3188 26480
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 5644 26440 5684 26480
rect 10348 26440 10388 26480
rect 15628 26440 15668 26480
rect 16108 26440 16148 26480
rect 16588 26440 16628 26480
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20620 26440 20660 26480
rect 2956 26356 2996 26396
rect 3340 26356 3380 26396
rect 6796 26356 6836 26396
rect 10636 26356 10676 26396
rect 14764 26356 14804 26396
rect 1708 26272 1748 26312
rect 7948 26272 7988 26312
rect 20716 26272 20756 26312
rect 2380 26104 2420 26144
rect 3436 26104 3476 26144
rect 4684 26104 4724 26144
rect 10636 26104 10676 26144
rect 12268 26104 12308 26144
rect 14956 26104 14996 26144
rect 7756 26020 7796 26060
rect 16492 26020 16532 26060
rect 4492 25936 4532 25976
rect 6412 25936 6452 25976
rect 16204 25936 16244 25976
rect 8620 25768 8660 25808
rect 9004 25768 9044 25808
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 17836 25600 17876 25640
rect 16300 25516 16340 25556
rect 3436 25432 3476 25472
rect 1324 25264 1364 25304
rect 2956 25348 2996 25388
rect 4396 25264 4436 25304
rect 6412 25348 6452 25388
rect 7948 25348 7988 25388
rect 8524 25348 8564 25388
rect 12652 25264 12692 25304
rect 5644 25180 5684 25220
rect 5836 25180 5876 25220
rect 8236 25180 8276 25220
rect 8524 25180 8564 25220
rect 6508 25096 6548 25136
rect 12268 25012 12308 25052
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 6412 24928 6452 24968
rect 14476 24928 14516 24968
rect 16204 24928 16244 24968
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 7468 24844 7508 24884
rect 16396 24844 16436 24884
rect 5548 24760 5588 24800
rect 6412 24760 6452 24800
rect 10252 24760 10292 24800
rect 8716 24676 8756 24716
rect 10828 24676 10868 24716
rect 2764 24592 2804 24632
rect 8620 24592 8660 24632
rect 11692 24592 11732 24632
rect 16300 24592 16340 24632
rect 6220 24508 6260 24548
rect 4300 24340 4340 24380
rect 16684 24340 16724 24380
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 10540 24172 10580 24212
rect 2764 24088 2804 24128
rect 14380 24088 14420 24128
rect 364 23920 404 23960
rect 3244 23920 3284 23960
rect 16780 24172 16820 24212
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 17452 24088 17492 24128
rect 21388 24088 21428 24128
rect 17164 23920 17204 23960
rect 9388 23836 9428 23876
rect 14380 23836 14420 23876
rect 3244 23752 3284 23792
rect 5548 23752 5588 23792
rect 4300 23584 4340 23624
rect 4588 23668 4628 23708
rect 9004 23668 9044 23708
rect 10060 23668 10100 23708
rect 14572 23668 14612 23708
rect 20140 23752 20180 23792
rect 11692 23500 11732 23540
rect 17836 23500 17876 23540
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 2092 23332 2132 23372
rect 10252 23248 10292 23288
rect 14188 23248 14228 23288
rect 10060 23080 10100 23120
rect 17452 23080 17492 23120
rect 16492 22996 16532 23036
rect 17164 22996 17204 23036
rect 19276 22912 19316 22952
rect 4588 22828 4628 22868
rect 5548 22828 5588 22868
rect 8332 22828 8372 22868
rect 15052 22828 15092 22868
rect 16684 22828 16724 22868
rect 14956 22744 14996 22784
rect 19756 22744 19796 22784
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 8332 22660 8372 22700
rect 12556 22660 12596 22700
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 3340 22492 3380 22532
rect 19276 22492 19316 22532
rect 19468 22492 19508 22532
rect 6028 22408 6068 22448
rect 14764 22408 14804 22448
rect 20140 22408 20180 22448
rect 4684 22324 4724 22364
rect 6700 22324 6740 22364
rect 7372 22324 7412 22364
rect 2860 22240 2900 22280
rect 18604 22240 18644 22280
rect 5356 22156 5396 22196
rect 6508 22072 6548 22112
rect 9004 22072 9044 22112
rect 3532 21988 3572 22028
rect 1900 21904 1940 21944
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 3436 21736 3476 21776
rect 20140 21736 20180 21776
rect 7852 21568 7892 21608
rect 15532 21652 15572 21692
rect 14284 21568 14324 21608
rect 14476 21568 14516 21608
rect 19276 21568 19316 21608
rect 3532 21484 3572 21524
rect 10252 21484 10292 21524
rect 14188 21400 14228 21440
rect 10540 21316 10580 21356
rect 14668 21316 14708 21356
rect 13900 21232 13940 21272
rect 15628 21232 15668 21272
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 14188 21064 14228 21104
rect 16396 21064 16436 21104
rect 16108 20896 16148 20936
rect 8332 20812 8372 20852
rect 9100 20812 9140 20852
rect 9580 20728 9620 20768
rect 15436 20728 15476 20768
rect 10348 20644 10388 20684
rect 16684 20644 16724 20684
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 12652 20308 12692 20348
rect 15148 20224 15188 20264
rect 17836 20224 17876 20264
rect 16588 20140 16628 20180
rect 18604 20140 18644 20180
rect 21004 20140 21044 20180
rect 3148 20056 3188 20096
rect 15148 20056 15188 20096
rect 12940 19972 12980 20012
rect 15340 19972 15380 20012
rect 19276 19972 19316 20012
rect 16684 19888 16724 19928
rect 5740 19804 5780 19844
rect 10060 19804 10100 19844
rect 20620 19720 20660 19760
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 1996 19552 2036 19592
rect 10060 19552 10100 19592
rect 14764 19552 14804 19592
rect 16300 19468 16340 19508
rect 5740 19384 5780 19424
rect 15532 19384 15572 19424
rect 19372 19384 19412 19424
rect 20812 19384 20852 19424
rect 2380 19300 2420 19340
rect 13612 19216 13652 19256
rect 4396 19132 4436 19172
rect 14380 19048 14420 19088
rect 3148 18964 3188 19004
rect 15724 18964 15764 19004
rect 2284 18880 2324 18920
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 15916 18880 15956 18920
rect 16588 18880 16628 18920
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 14764 18712 14804 18752
rect 16876 18712 16916 18752
rect 6028 18544 6068 18584
rect 14860 18544 14900 18584
rect 19276 18544 19316 18584
rect 6796 18376 6836 18416
rect 17836 18376 17876 18416
rect 18220 18376 18260 18416
rect 6412 18292 6452 18332
rect 2764 18124 2804 18164
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 13228 17872 13268 17912
rect 17356 17872 17396 17912
rect 9388 17788 9428 17828
rect 10636 17788 10676 17828
rect 2764 17620 2804 17660
rect 12460 17620 12500 17660
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 6892 17368 6932 17408
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20620 17368 20660 17408
rect 15724 17200 15764 17240
rect 16492 17116 16532 17156
rect 13900 17032 13940 17072
rect 19468 17032 19508 17072
rect 21388 17032 21428 17072
rect 3340 16948 3380 16988
rect 4684 16864 4724 16904
rect 9388 16696 9428 16736
rect 16396 16696 16436 16736
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 6700 16612 6740 16652
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 6604 16528 6644 16568
rect 7852 16528 7892 16568
rect 19276 16444 19316 16484
rect 4492 16360 4532 16400
rect 7372 16024 7412 16064
rect 19948 16276 19988 16316
rect 15532 16192 15572 16232
rect 15916 16108 15956 16148
rect 11500 16024 11540 16064
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 15340 15772 15380 15812
rect 19276 15772 19316 15812
rect 2764 15604 2804 15644
rect 16108 15604 16148 15644
rect 15148 15520 15188 15560
rect 17644 15520 17684 15560
rect 18604 15520 18644 15560
rect 4492 15436 4532 15476
rect 7468 15436 7508 15476
rect 18220 15436 18260 15476
rect 19948 15436 19988 15476
rect 16108 15268 16148 15308
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 12076 15016 12116 15056
rect 15244 15016 15284 15056
rect 16108 15016 16148 15056
rect 4588 14932 4628 14972
rect 2188 14848 2228 14888
rect 15916 14596 15956 14636
rect 1228 14512 1268 14552
rect 5548 14512 5588 14552
rect 8620 14428 8660 14468
rect 8812 14512 8852 14552
rect 14668 14428 14708 14468
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 6700 14176 6740 14216
rect 15724 14176 15764 14216
rect 4588 14092 4628 14132
rect 3532 14008 3572 14048
rect 17260 14008 17300 14048
rect 3340 13924 3380 13964
rect 5740 13840 5780 13880
rect 14668 13840 14708 13880
rect 15628 13840 15668 13880
rect 5356 13756 5396 13796
rect 5644 13756 5684 13796
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 15340 13504 15380 13544
rect 2188 13420 2228 13460
rect 15532 13420 15572 13460
rect 15244 13252 15284 13292
rect 16780 13252 16820 13292
rect 5644 13168 5684 13208
rect 16108 13168 16148 13208
rect 1420 13000 1460 13040
rect 3340 12916 3380 12956
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 2092 12748 2132 12788
rect 6028 12748 6068 12788
rect 2476 12580 2516 12620
rect 16108 12580 16148 12620
rect 15052 12496 15092 12536
rect 16300 12496 16340 12536
rect 19372 12496 19412 12536
rect 19948 12496 19988 12536
rect 2284 12244 2324 12284
rect 2092 12076 2132 12116
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 4684 12076 4724 12116
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 8332 11992 8372 12032
rect 3148 11908 3188 11948
rect 6220 11824 6260 11864
rect 6892 11824 6932 11864
rect 14956 11824 14996 11864
rect 4108 11656 4148 11696
rect 2188 11572 2228 11612
rect 3052 11572 3092 11612
rect 12940 11572 12980 11612
rect 2476 11404 2516 11444
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 844 11236 884 11276
rect 16396 11236 16436 11276
rect 6028 11152 6068 11192
rect 4204 10984 4244 11024
rect 15820 10984 15860 11024
rect 16780 10984 16820 11024
rect 4876 10900 4916 10940
rect 16108 10900 16148 10940
rect 3532 10732 3572 10772
rect 15628 10732 15668 10772
rect 3244 10564 3284 10604
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 4204 10564 4244 10604
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 5356 10480 5396 10520
rect 20620 10480 20660 10520
rect 1324 10312 1364 10352
rect 14476 10228 14516 10268
rect 16108 10228 16148 10268
rect 3148 10144 3188 10184
rect 4300 10060 4340 10100
rect 3340 9976 3380 10016
rect 14956 9976 14996 10016
rect 15820 10060 15860 10100
rect 2764 9892 2804 9932
rect 16204 9892 16244 9932
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 12460 9808 12500 9848
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 3148 9724 3188 9764
rect 4108 9724 4148 9764
rect 2284 9640 2324 9680
rect 3244 9556 3284 9596
rect 3340 9472 3380 9512
rect 5644 9472 5684 9512
rect 12076 9472 12116 9512
rect 2188 9304 2228 9344
rect 4108 9220 4148 9260
rect 2860 9136 2900 9176
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 3340 8884 3380 8924
rect 4588 8884 4628 8924
rect 15436 8884 15476 8924
rect 6220 8800 6260 8840
rect 17644 8800 17684 8840
rect 18412 8800 18452 8840
rect 4204 8716 4244 8756
rect 2860 8632 2900 8672
rect 3244 8632 3284 8672
rect 18604 8800 18644 8840
rect 15436 8716 15476 8756
rect 21388 8716 21428 8756
rect 4396 8632 4436 8672
rect 12076 8632 12116 8672
rect 12844 8632 12884 8672
rect 15532 8548 15572 8588
rect 3244 8464 3284 8504
rect 4492 8464 4532 8504
rect 19948 8380 19988 8420
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 14956 8212 14996 8252
rect 15244 8212 15284 8252
rect 2764 8128 2804 8168
rect 7948 8128 7988 8168
rect 14284 8128 14324 8168
rect 4300 8044 4340 8084
rect 8524 8044 8564 8084
rect 2476 7960 2516 8000
rect 4396 7960 4436 8000
rect 4684 7960 4724 8000
rect 10060 7960 10100 8000
rect 12076 7960 12116 8000
rect 2860 7876 2900 7916
rect 8620 7876 8660 7916
rect 15244 7876 15284 7916
rect 19276 7792 19316 7832
rect 6412 7708 6452 7748
rect 6604 7708 6644 7748
rect 15532 7624 15572 7664
rect 17932 7624 17972 7664
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 12172 7540 12212 7580
rect 12652 7540 12692 7580
rect 15148 7540 15188 7580
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 9580 7372 9620 7412
rect 10060 7372 10100 7412
rect 8428 7288 8468 7328
rect 8812 7204 8852 7244
rect 12076 7120 12116 7160
rect 4684 7036 4724 7076
rect 15052 7036 15092 7076
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 15820 6784 15860 6824
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 6316 6616 6356 6656
rect 2380 6448 2420 6488
rect 16300 6448 16340 6488
rect 6604 6280 6644 6320
rect 7948 6280 7988 6320
rect 10732 6280 10772 6320
rect 6412 6196 6452 6236
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 6508 6028 6548 6068
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 11692 5944 11732 5984
rect 4204 5860 4244 5900
rect 9292 5860 9332 5900
rect 12268 5860 12308 5900
rect 10252 5776 10292 5816
rect 17644 5776 17684 5816
rect 6124 5692 6164 5732
rect 8908 5692 8948 5732
rect 652 5608 692 5648
rect 5356 5608 5396 5648
rect 5548 5524 5588 5564
rect 9484 5692 9524 5732
rect 10732 5608 10772 5648
rect 14284 5608 14324 5648
rect 15052 5608 15092 5648
rect 19276 5608 19316 5648
rect 9388 5440 9428 5480
rect 4492 5272 4532 5312
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 1324 5104 1364 5144
rect 7276 5188 7316 5228
rect 12940 5188 12980 5228
rect 15628 5188 15668 5228
rect 3436 5104 3476 5144
rect 7852 5104 7892 5144
rect 17644 5020 17684 5060
rect 5452 4936 5492 4976
rect 10444 4936 10484 4976
rect 9100 4852 9140 4892
rect 17932 4852 17972 4892
rect 4300 4768 4340 4808
rect 6124 4768 6164 4808
rect 6796 4768 6836 4808
rect 18412 4684 18452 4724
rect 8716 4600 8756 4640
rect 13036 4600 13076 4640
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4972 4516 5012 4556
rect 17932 4516 17972 4556
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 9388 4432 9428 4472
rect 2572 4264 2612 4304
rect 3148 4180 3188 4220
rect 8524 4180 8564 4220
rect 10828 4180 10868 4220
rect 4108 4096 4148 4136
rect 13900 4096 13940 4136
rect 16780 4096 16820 4136
rect 17932 4096 17972 4136
rect 8908 4012 8948 4052
rect 5740 3928 5780 3968
rect 9100 3928 9140 3968
rect 10156 3928 10196 3968
rect 10348 3928 10388 3968
rect 2476 3844 2516 3884
rect 8332 3844 8372 3884
rect 10060 3844 10100 3884
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 7468 3760 7508 3800
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 11692 3676 11732 3716
rect 2092 3592 2132 3632
rect 2476 3592 2516 3632
rect 16204 3592 16244 3632
rect 2572 3508 2612 3548
rect 3340 3508 3380 3548
rect 5932 3508 5972 3548
rect 4588 3340 4628 3380
rect 7756 3340 7796 3380
rect 10060 3340 10100 3380
rect 10540 3340 10580 3380
rect 11500 3340 11540 3380
rect 12364 3340 12404 3380
rect 16588 3340 16628 3380
rect 16972 3340 17012 3380
rect 940 3256 980 3296
rect 8812 3256 8852 3296
rect 2284 3088 2324 3128
rect 15052 3088 15092 3128
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 8908 3004 8948 3044
rect 11212 3004 11252 3044
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 1804 2836 1844 2876
rect 844 2752 884 2792
rect 3628 2752 3668 2792
rect 4108 2752 4148 2792
rect 7564 2668 7604 2708
rect 9004 2668 9044 2708
rect 9196 2668 9236 2708
rect 11596 2668 11636 2708
rect 14188 2668 14228 2708
rect 14572 2668 14612 2708
rect 6988 2584 7028 2624
rect 3244 2500 3284 2540
rect 8044 2500 8084 2540
rect 8812 2500 8852 2540
rect 1228 2332 1268 2372
rect 3052 2248 3092 2288
rect 3244 2248 3284 2288
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 10252 2248 10292 2288
rect 11596 2164 11636 2204
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 13900 2164 13940 2204
rect 2764 2080 2804 2120
rect 5644 1996 5684 2036
rect 6988 1996 7028 2036
rect 7372 1828 7412 1868
rect 7276 1744 7316 1784
rect 8428 1912 8468 1952
rect 9100 1828 9140 1868
rect 9484 1828 9524 1868
rect 16012 1828 16052 1868
rect 15436 1660 15476 1700
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 10444 1408 10484 1448
rect 2476 1324 2516 1364
rect 2956 1240 2996 1280
rect 4684 1240 4724 1280
rect 12748 1240 12788 1280
rect 13132 1240 13172 1280
rect 17740 1240 17780 1280
rect 18124 1240 18164 1280
rect 18700 1240 18740 1280
rect 10348 1156 10388 1196
rect 13036 1156 13076 1196
rect 17164 1156 17204 1196
rect 2476 1072 2516 1112
rect 3340 1072 3380 1112
rect 6796 1072 6836 1112
rect 2668 988 2708 1028
rect 8332 1072 8372 1112
rect 17548 1156 17588 1196
rect 18028 1156 18068 1196
rect 18316 988 18356 1028
rect 4780 904 4820 944
rect 11788 904 11828 944
rect 13324 904 13364 944
rect 13996 904 14036 944
rect 748 820 788 860
rect 8236 820 8276 860
rect 14092 820 14132 860
rect 20524 820 20564 860
rect 1420 736 1460 776
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 10444 736 10484 776
rect 13708 736 13748 776
rect 15628 736 15668 776
rect 16780 736 16820 776
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 11884 652 11924 692
rect 18892 652 18932 692
rect 2956 568 2996 608
rect 6988 484 7028 524
rect 8428 400 8468 440
rect 6988 316 7028 356
rect 3532 232 3572 272
rect 11020 232 11060 272
rect 17356 232 17396 272
rect 16108 148 16148 188
rect 19468 148 19508 188
<< metal4 >>
rect 7276 85700 7316 85709
rect 940 85280 980 85289
rect 652 79568 692 79577
rect 555 75872 597 75881
rect 555 75832 556 75872
rect 596 75832 597 75872
rect 555 75823 597 75832
rect 556 73193 596 75823
rect 555 73184 597 73193
rect 555 73144 556 73184
rect 596 73144 597 73184
rect 555 73135 597 73144
rect 652 73184 692 79528
rect 652 73135 692 73144
rect 843 73100 885 73109
rect 843 73060 844 73100
rect 884 73060 885 73100
rect 843 73051 885 73060
rect 460 72092 500 72101
rect 172 68984 212 68993
rect 76 67640 116 67649
rect 76 50000 116 67600
rect 172 51344 212 68944
rect 268 67976 308 67985
rect 268 58988 308 67936
rect 460 63272 500 72052
rect 844 66800 884 73051
rect 844 66751 884 66760
rect 460 63223 500 63232
rect 844 63440 884 63449
rect 268 58939 308 58948
rect 460 62852 500 62861
rect 172 51295 212 51304
rect 76 49951 116 49960
rect 364 23960 404 23969
rect 364 23801 404 23920
rect 363 23792 405 23801
rect 363 23752 364 23792
rect 404 23752 405 23792
rect 363 23743 405 23752
rect 460 2885 500 62812
rect 652 61676 692 61685
rect 556 54452 596 54461
rect 556 23885 596 54412
rect 652 27749 692 61636
rect 748 36812 788 36821
rect 651 27740 693 27749
rect 651 27700 652 27740
rect 692 27700 693 27740
rect 651 27691 693 27700
rect 652 27068 692 27077
rect 555 23876 597 23885
rect 555 23836 556 23876
rect 596 23836 597 23876
rect 555 23827 597 23836
rect 652 5648 692 27028
rect 652 5599 692 5608
rect 459 2876 501 2885
rect 459 2836 460 2876
rect 500 2836 501 2876
rect 459 2827 501 2836
rect 748 860 788 36772
rect 844 26657 884 63400
rect 940 51680 980 85240
rect 3436 84944 3476 84953
rect 2956 84692 2996 84701
rect 1323 84356 1365 84365
rect 1323 84316 1324 84356
rect 1364 84316 1365 84356
rect 1323 84307 1365 84316
rect 1324 84222 1364 84307
rect 2572 83936 2612 83945
rect 1516 83516 1556 83525
rect 1324 82256 1364 82265
rect 1036 82088 1076 82097
rect 1036 67640 1076 82048
rect 1324 80828 1364 82216
rect 1324 80779 1364 80788
rect 1420 79904 1460 79913
rect 1324 79736 1364 79745
rect 1132 79484 1172 79493
rect 1132 74780 1172 79444
rect 1324 79148 1364 79696
rect 1324 79099 1364 79108
rect 1228 78392 1268 78401
rect 1228 75032 1268 78352
rect 1228 74983 1268 74992
rect 1324 77552 1364 77561
rect 1324 76040 1364 77512
rect 1420 76712 1460 79864
rect 1420 76124 1460 76672
rect 1420 76075 1460 76084
rect 1132 74740 1268 74780
rect 1036 67591 1076 67600
rect 1132 73100 1172 73109
rect 940 51631 980 51640
rect 1036 64364 1076 64373
rect 940 46640 980 46649
rect 843 26648 885 26657
rect 843 26608 844 26648
rect 884 26608 885 26648
rect 843 26599 885 26608
rect 844 11276 884 11285
rect 844 2792 884 11236
rect 940 3296 980 46600
rect 1036 10949 1076 64324
rect 1132 61760 1172 73060
rect 1132 61711 1172 61720
rect 1131 52772 1173 52781
rect 1131 52732 1132 52772
rect 1172 52732 1173 52772
rect 1131 52723 1173 52732
rect 1132 46724 1172 52723
rect 1132 46675 1172 46684
rect 1228 41600 1268 74740
rect 1324 73100 1364 76000
rect 1420 75284 1460 75293
rect 1420 75041 1460 75244
rect 1419 75032 1461 75041
rect 1419 74992 1420 75032
rect 1460 74992 1461 75032
rect 1419 74983 1461 74992
rect 1324 73060 1460 73100
rect 1324 72932 1364 72941
rect 1324 71336 1364 72892
rect 1324 71287 1364 71296
rect 1420 65708 1460 73060
rect 1516 67136 1556 83476
rect 1804 81920 1844 81929
rect 1612 81500 1652 81509
rect 1612 79064 1652 81460
rect 1612 77384 1652 79024
rect 1612 77335 1652 77344
rect 1804 76208 1844 81880
rect 1804 76159 1844 76168
rect 1900 80828 1940 80837
rect 1900 77720 1940 80788
rect 1804 76040 1844 76049
rect 1516 67087 1556 67096
rect 1708 74360 1748 74369
rect 1420 65659 1460 65668
rect 1708 65372 1748 74320
rect 1804 71168 1844 76000
rect 1900 75536 1940 77680
rect 1900 75487 1940 75496
rect 1996 79736 2036 79745
rect 1996 78056 2036 79696
rect 1996 77804 2036 78016
rect 1996 73100 2036 77764
rect 2284 79316 2324 79325
rect 2284 78308 2324 79276
rect 2092 77216 2132 77225
rect 2092 76628 2132 77176
rect 2092 76579 2132 76588
rect 2188 76712 2228 76721
rect 1996 73060 2132 73100
rect 1804 71119 1844 71128
rect 2092 69152 2132 73060
rect 2092 69103 2132 69112
rect 1708 65323 1748 65332
rect 1804 66716 1844 66725
rect 1420 63272 1460 63281
rect 1323 62180 1365 62189
rect 1323 62140 1324 62180
rect 1364 62140 1365 62180
rect 1323 62131 1365 62140
rect 1324 57896 1364 62131
rect 1324 57847 1364 57856
rect 1420 54872 1460 63232
rect 1420 54823 1460 54832
rect 1708 62516 1748 62525
rect 1612 54536 1652 54545
rect 1612 52352 1652 54496
rect 1612 52303 1652 52312
rect 1708 50252 1748 62476
rect 1708 50203 1748 50212
rect 1132 41560 1268 41600
rect 1324 42776 1364 42785
rect 1132 33452 1172 41560
rect 1228 37736 1268 37747
rect 1228 37661 1268 37696
rect 1227 37652 1269 37661
rect 1227 37612 1228 37652
rect 1268 37612 1269 37652
rect 1227 37603 1269 37612
rect 1132 33412 1268 33452
rect 1132 29252 1172 29261
rect 1132 27320 1172 29212
rect 1132 27271 1172 27280
rect 1228 15140 1268 33412
rect 1324 25304 1364 42736
rect 1612 39416 1652 39425
rect 1420 38492 1460 38501
rect 1420 34124 1460 38452
rect 1420 34075 1460 34084
rect 1612 31856 1652 39376
rect 1612 31436 1652 31816
rect 1612 31387 1652 31396
rect 1707 27488 1749 27497
rect 1707 27448 1708 27488
rect 1748 27448 1749 27488
rect 1707 27439 1749 27448
rect 1708 26312 1748 27439
rect 1708 26263 1748 26272
rect 1324 25255 1364 25264
rect 1132 15100 1268 15140
rect 1132 11360 1172 15100
rect 1227 14552 1269 14561
rect 1227 14512 1228 14552
rect 1268 14512 1269 14552
rect 1227 14503 1269 14512
rect 1228 14418 1268 14503
rect 1420 13040 1460 13049
rect 1132 11320 1268 11360
rect 1035 10940 1077 10949
rect 1035 10900 1036 10940
rect 1076 10900 1077 10940
rect 1035 10891 1077 10900
rect 940 3247 980 3256
rect 844 2743 884 2752
rect 1228 2372 1268 11320
rect 1324 10352 1364 10361
rect 1324 5144 1364 10312
rect 1324 5095 1364 5104
rect 1228 2323 1268 2332
rect 748 811 788 820
rect 1420 776 1460 13000
rect 1804 2876 1844 66676
rect 2188 64616 2228 76672
rect 2284 69404 2324 78268
rect 2476 78980 2516 78989
rect 2380 77384 2420 77393
rect 2380 76460 2420 77344
rect 2380 73016 2420 76420
rect 2380 72967 2420 72976
rect 2284 69355 2324 69364
rect 2380 69152 2420 69161
rect 2188 64567 2228 64576
rect 2284 66464 2324 66473
rect 1996 63272 2036 63281
rect 1900 51764 1940 51773
rect 1900 49748 1940 51724
rect 1900 47312 1940 49708
rect 1996 48488 2036 63232
rect 2284 53285 2324 66424
rect 2380 54032 2420 69112
rect 2476 64532 2516 78940
rect 2572 76544 2612 83896
rect 2764 82424 2804 82433
rect 2764 79568 2804 82384
rect 2764 79519 2804 79528
rect 2956 79400 2996 84652
rect 3340 83516 3380 83525
rect 3340 83096 3380 83476
rect 3340 83047 3380 83056
rect 3051 80660 3093 80669
rect 3051 80620 3052 80660
rect 3092 80620 3093 80660
rect 3051 80611 3093 80620
rect 2956 79351 2996 79360
rect 2572 76495 2612 76504
rect 2860 77132 2900 77141
rect 2476 64483 2516 64492
rect 2572 76376 2612 76385
rect 2475 59492 2517 59501
rect 2475 59452 2476 59492
rect 2516 59452 2517 59492
rect 2475 59443 2517 59452
rect 2476 54116 2516 59443
rect 2476 54067 2516 54076
rect 2380 53983 2420 53992
rect 2283 53276 2325 53285
rect 2283 53236 2284 53276
rect 2324 53236 2325 53276
rect 2283 53227 2325 53236
rect 1996 48439 2036 48448
rect 2380 52100 2420 52109
rect 1900 47263 1940 47272
rect 2092 43784 2132 43793
rect 1996 41432 2036 41441
rect 1996 38156 2036 41392
rect 2092 39416 2132 43744
rect 2092 39367 2132 39376
rect 2188 43364 2228 43373
rect 1996 38107 2036 38116
rect 2188 34712 2228 43324
rect 2380 43028 2420 52060
rect 2380 42979 2420 42988
rect 2476 43700 2516 43709
rect 2476 42776 2516 43660
rect 2476 42727 2516 42736
rect 2379 39080 2421 39089
rect 2379 39040 2380 39080
rect 2420 39040 2421 39080
rect 2379 39031 2421 39040
rect 2380 38946 2420 39031
rect 1996 33704 2036 33713
rect 1900 32108 1940 32117
rect 1900 21944 1940 32068
rect 1900 21895 1940 21904
rect 1996 19592 2036 33664
rect 2188 33704 2228 34672
rect 2188 33655 2228 33664
rect 2380 38156 2420 38165
rect 2092 30176 2132 30185
rect 2092 23372 2132 30136
rect 2380 26144 2420 38116
rect 2476 29336 2516 29345
rect 2476 27656 2516 29296
rect 2476 27607 2516 27616
rect 2380 26069 2420 26104
rect 2379 26060 2421 26069
rect 2379 26020 2380 26060
rect 2420 26020 2421 26060
rect 2379 26011 2421 26020
rect 2380 25980 2420 26011
rect 2092 23323 2132 23332
rect 1996 19543 2036 19552
rect 2380 19340 2420 19349
rect 2284 18920 2324 18929
rect 2188 14888 2228 14897
rect 2188 13460 2228 14848
rect 2188 13411 2228 13420
rect 2092 12788 2132 12797
rect 2092 12116 2132 12748
rect 2284 12284 2324 18880
rect 2284 12235 2324 12244
rect 2092 12067 2132 12076
rect 2188 11612 2228 11621
rect 2188 9344 2228 11572
rect 2188 9295 2228 9304
rect 2284 9680 2324 9689
rect 2091 3632 2133 3641
rect 2091 3592 2092 3632
rect 2132 3592 2133 3632
rect 2091 3583 2133 3592
rect 2092 3498 2132 3583
rect 2284 3128 2324 9640
rect 2380 6488 2420 19300
rect 2476 12620 2516 12629
rect 2476 11444 2516 12580
rect 2476 11395 2516 11404
rect 2380 6439 2420 6448
rect 2476 8000 2516 8009
rect 2476 3884 2516 7960
rect 2476 3835 2516 3844
rect 2572 4304 2612 76336
rect 2764 75200 2804 75209
rect 2764 74528 2804 75160
rect 2668 72008 2708 72017
rect 2668 67388 2708 71968
rect 2668 64700 2708 67348
rect 2668 64651 2708 64660
rect 2764 61592 2804 74488
rect 2860 68732 2900 77092
rect 2860 68683 2900 68692
rect 2956 73436 2996 73445
rect 2764 61543 2804 61552
rect 2860 68564 2900 68573
rect 2763 61088 2805 61097
rect 2763 61048 2764 61088
rect 2804 61048 2805 61088
rect 2763 61039 2805 61048
rect 2764 56216 2804 61039
rect 2764 56167 2804 56176
rect 2764 54116 2804 54125
rect 2764 46556 2804 54076
rect 2764 46507 2804 46516
rect 2284 3079 2324 3088
rect 2476 3632 2516 3641
rect 1804 2827 1844 2836
rect 2476 1364 2516 3592
rect 2572 3548 2612 4264
rect 2572 3499 2612 3508
rect 2668 38072 2708 38081
rect 2476 1112 2516 1324
rect 2476 1063 2516 1072
rect 2668 1028 2708 38032
rect 2860 37325 2900 68524
rect 2956 52100 2996 73396
rect 2956 52051 2996 52060
rect 2956 40508 2996 40517
rect 2859 37316 2901 37325
rect 2859 37276 2860 37316
rect 2900 37276 2901 37316
rect 2859 37267 2901 37276
rect 2764 36392 2804 36401
rect 2764 33536 2804 36352
rect 2764 30596 2804 33496
rect 2764 30547 2804 30556
rect 2764 30428 2804 30437
rect 2764 24632 2804 30388
rect 2956 29924 2996 40468
rect 3052 38996 3092 80611
rect 3148 80408 3188 80417
rect 3148 73100 3188 80368
rect 3340 78896 3380 78905
rect 3244 78560 3284 78569
rect 3244 77132 3284 78520
rect 3244 77083 3284 77092
rect 3148 73051 3188 73060
rect 3244 76712 3284 76721
rect 3244 72680 3284 76672
rect 3340 75284 3380 78856
rect 3436 76880 3476 84904
rect 3688 84692 4056 84701
rect 3728 84652 3770 84692
rect 3810 84652 3852 84692
rect 3892 84652 3934 84692
rect 3974 84652 4016 84692
rect 3688 84643 4056 84652
rect 4780 84692 4820 84701
rect 4683 84356 4725 84365
rect 4683 84316 4684 84356
rect 4724 84316 4725 84356
rect 4683 84307 4725 84316
rect 3532 84272 3572 84281
rect 3532 81752 3572 84232
rect 4300 83936 4340 83945
rect 3688 83180 4056 83189
rect 3728 83140 3770 83180
rect 3810 83140 3852 83180
rect 3892 83140 3934 83180
rect 3974 83140 4016 83180
rect 3688 83131 4056 83140
rect 4108 82172 4148 82181
rect 3820 82013 3860 82098
rect 3819 82004 3861 82013
rect 3819 81964 3820 82004
rect 3860 81964 3861 82004
rect 3819 81955 3861 81964
rect 3532 81500 3572 81712
rect 3688 81668 4056 81677
rect 3728 81628 3770 81668
rect 3810 81628 3852 81668
rect 3892 81628 3934 81668
rect 3974 81628 4016 81668
rect 3688 81619 4056 81628
rect 3532 81460 3668 81500
rect 3532 81248 3572 81257
rect 3532 77468 3572 81208
rect 3628 81164 3668 81460
rect 3628 81115 3668 81124
rect 3916 81248 3956 81257
rect 3916 80669 3956 81208
rect 3915 80660 3957 80669
rect 3915 80620 3916 80660
rect 3956 80620 3957 80660
rect 3915 80611 3957 80620
rect 3688 80156 4056 80165
rect 3728 80116 3770 80156
rect 3810 80116 3852 80156
rect 3892 80116 3934 80156
rect 3974 80116 4016 80156
rect 3688 80107 4056 80116
rect 3688 78644 4056 78653
rect 3728 78604 3770 78644
rect 3810 78604 3852 78644
rect 3892 78604 3934 78644
rect 3974 78604 4016 78644
rect 3688 78595 4056 78604
rect 3532 77419 3572 77428
rect 3688 77132 4056 77141
rect 3728 77092 3770 77132
rect 3810 77092 3852 77132
rect 3892 77092 3934 77132
rect 3974 77092 4016 77132
rect 3688 77083 4056 77092
rect 3436 76831 3476 76840
rect 3532 77048 3572 77057
rect 3340 75235 3380 75244
rect 3244 72631 3284 72640
rect 3340 74444 3380 74453
rect 3340 70832 3380 74404
rect 3436 74276 3476 74285
rect 3436 72344 3476 74236
rect 3436 72295 3476 72304
rect 3532 71840 3572 77008
rect 4108 76964 4148 82132
rect 4108 76915 4148 76924
rect 4204 77468 4244 77477
rect 3688 75620 4056 75629
rect 3728 75580 3770 75620
rect 3810 75580 3852 75620
rect 3892 75580 3934 75620
rect 3974 75580 4016 75620
rect 3688 75571 4056 75580
rect 4108 75032 4148 75041
rect 3688 74108 4056 74117
rect 3728 74068 3770 74108
rect 3810 74068 3852 74108
rect 3892 74068 3934 74108
rect 3974 74068 4016 74108
rect 3688 74059 4056 74068
rect 3688 72596 4056 72605
rect 3728 72556 3770 72596
rect 3810 72556 3852 72596
rect 3892 72556 3934 72596
rect 3974 72556 4016 72596
rect 3688 72547 4056 72556
rect 3532 71791 3572 71800
rect 3688 71084 4056 71093
rect 3728 71044 3770 71084
rect 3810 71044 3852 71084
rect 3892 71044 3934 71084
rect 3974 71044 4016 71084
rect 3688 71035 4056 71044
rect 3340 70783 3380 70792
rect 3532 70916 3572 70925
rect 3148 69152 3188 69161
rect 3148 65624 3188 69112
rect 3148 65575 3188 65584
rect 3244 68900 3284 68909
rect 3244 62012 3284 68860
rect 3340 68732 3380 68741
rect 3340 66128 3380 68692
rect 3340 66079 3380 66088
rect 3244 61963 3284 61972
rect 3340 65456 3380 65465
rect 3244 61592 3284 61601
rect 3148 59240 3188 59249
rect 3148 48152 3188 59200
rect 3244 57728 3284 61552
rect 3340 60164 3380 65416
rect 3340 60115 3380 60124
rect 3436 63188 3476 63197
rect 3436 61928 3476 63148
rect 3244 57679 3284 57688
rect 3436 57224 3476 61888
rect 3244 55712 3284 55721
rect 3244 53528 3284 55672
rect 3436 54620 3476 57184
rect 3436 54571 3476 54580
rect 3244 53479 3284 53488
rect 3148 48103 3188 48112
rect 3148 47984 3188 47993
rect 3148 41441 3188 47944
rect 3243 41936 3285 41945
rect 3243 41896 3244 41936
rect 3284 41896 3285 41936
rect 3243 41887 3285 41896
rect 3147 41432 3189 41441
rect 3147 41392 3148 41432
rect 3188 41392 3189 41432
rect 3147 41383 3189 41392
rect 3052 38947 3092 38956
rect 3244 37400 3284 41887
rect 3436 40928 3476 40937
rect 3436 40508 3476 40888
rect 3436 40459 3476 40468
rect 3244 37351 3284 37360
rect 3340 40340 3380 40349
rect 3340 38492 3380 40300
rect 3244 32864 3284 32873
rect 2956 29875 2996 29884
rect 3052 32192 3092 32201
rect 2956 27992 2996 28001
rect 2764 24583 2804 24592
rect 2860 27236 2900 27245
rect 2860 26816 2900 27196
rect 2764 24128 2804 24137
rect 2764 23801 2804 24088
rect 2763 23792 2805 23801
rect 2763 23752 2764 23792
rect 2804 23752 2805 23792
rect 2763 23743 2805 23752
rect 2860 22280 2900 26776
rect 2956 26396 2996 27952
rect 3052 26909 3092 32152
rect 3148 28496 3188 28505
rect 3148 26984 3188 28456
rect 3148 26935 3188 26944
rect 3051 26900 3093 26909
rect 3051 26860 3052 26900
rect 3092 26860 3093 26900
rect 3051 26851 3093 26860
rect 3244 26816 3284 32824
rect 3340 29000 3380 38452
rect 3532 35300 3572 70876
rect 3688 69572 4056 69581
rect 3728 69532 3770 69572
rect 3810 69532 3852 69572
rect 3892 69532 3934 69572
rect 3974 69532 4016 69572
rect 3688 69523 4056 69532
rect 3688 68060 4056 68069
rect 3728 68020 3770 68060
rect 3810 68020 3852 68060
rect 3892 68020 3934 68060
rect 3974 68020 4016 68060
rect 3688 68011 4056 68020
rect 3688 66548 4056 66557
rect 3728 66508 3770 66548
rect 3810 66508 3852 66548
rect 3892 66508 3934 66548
rect 3974 66508 4016 66548
rect 3688 66499 4056 66508
rect 3688 65036 4056 65045
rect 3728 64996 3770 65036
rect 3810 64996 3852 65036
rect 3892 64996 3934 65036
rect 3974 64996 4016 65036
rect 3688 64987 4056 64996
rect 3688 63524 4056 63533
rect 3728 63484 3770 63524
rect 3810 63484 3852 63524
rect 3892 63484 3934 63524
rect 3974 63484 4016 63524
rect 3688 63475 4056 63484
rect 3688 62012 4056 62021
rect 3728 61972 3770 62012
rect 3810 61972 3852 62012
rect 3892 61972 3934 62012
rect 3974 61972 4016 62012
rect 3688 61963 4056 61972
rect 3688 60500 4056 60509
rect 3728 60460 3770 60500
rect 3810 60460 3852 60500
rect 3892 60460 3934 60500
rect 3974 60460 4016 60500
rect 3688 60451 4056 60460
rect 4108 60080 4148 74992
rect 4204 61676 4244 77428
rect 4300 75452 4340 83896
rect 4684 81920 4724 84307
rect 4780 82172 4820 84652
rect 6028 84440 6068 84449
rect 4928 83936 5296 83945
rect 4968 83896 5010 83936
rect 5050 83896 5092 83936
rect 5132 83896 5174 83936
rect 5214 83896 5256 83936
rect 4928 83887 5296 83896
rect 5356 82928 5396 82937
rect 4928 82424 5296 82433
rect 4968 82384 5010 82424
rect 5050 82384 5092 82424
rect 5132 82384 5174 82424
rect 5214 82384 5256 82424
rect 4928 82375 5296 82384
rect 4780 82123 4820 82132
rect 5356 82172 5396 82888
rect 5451 82844 5493 82853
rect 5451 82804 5452 82844
rect 5492 82804 5493 82844
rect 5451 82795 5493 82804
rect 5452 82710 5492 82795
rect 5740 82760 5780 82769
rect 4780 81920 4820 81929
rect 4684 81880 4780 81920
rect 5356 81920 5396 82132
rect 5356 81880 5492 81920
rect 4300 75403 4340 75412
rect 4492 80072 4532 80081
rect 4300 70580 4340 70589
rect 4300 69992 4340 70540
rect 4300 62684 4340 69952
rect 4300 61760 4340 62644
rect 4396 63104 4436 63113
rect 4396 61928 4436 63064
rect 4396 61879 4436 61888
rect 4300 61711 4340 61720
rect 4204 61627 4244 61636
rect 4108 59912 4148 60040
rect 3688 58988 4056 58997
rect 3728 58948 3770 58988
rect 3810 58948 3852 58988
rect 3892 58948 3934 58988
rect 3974 58948 4016 58988
rect 3688 58939 4056 58948
rect 4108 58316 4148 59872
rect 4204 59324 4244 59335
rect 4204 59249 4244 59284
rect 4396 59324 4436 59333
rect 4203 59240 4245 59249
rect 4203 59200 4204 59240
rect 4244 59200 4245 59240
rect 4203 59191 4245 59200
rect 4108 58267 4148 58276
rect 4204 57896 4244 59191
rect 4204 57847 4244 57856
rect 3688 57476 4056 57485
rect 3728 57436 3770 57476
rect 3810 57436 3852 57476
rect 3892 57436 3934 57476
rect 3974 57436 4016 57476
rect 3688 57427 4056 57436
rect 3688 55964 4056 55973
rect 3728 55924 3770 55964
rect 3810 55924 3852 55964
rect 3892 55924 3934 55964
rect 3974 55924 4016 55964
rect 3688 55915 4056 55924
rect 3688 54452 4056 54461
rect 3728 54412 3770 54452
rect 3810 54412 3852 54452
rect 3892 54412 3934 54452
rect 3974 54412 4016 54452
rect 3688 54403 4056 54412
rect 4396 53360 4436 59284
rect 4396 53311 4436 53320
rect 3688 52940 4056 52949
rect 3728 52900 3770 52940
rect 3810 52900 3852 52940
rect 3892 52900 3934 52940
rect 3974 52900 4016 52940
rect 3688 52891 4056 52900
rect 3688 51428 4056 51437
rect 3728 51388 3770 51428
rect 3810 51388 3852 51428
rect 3892 51388 3934 51428
rect 3974 51388 4016 51428
rect 3688 51379 4056 51388
rect 4396 51176 4436 51185
rect 4108 50924 4148 50933
rect 3688 49916 4056 49925
rect 3728 49876 3770 49916
rect 3810 49876 3852 49916
rect 3892 49876 3934 49916
rect 3974 49876 4016 49916
rect 3688 49867 4056 49876
rect 3688 48404 4056 48413
rect 3728 48364 3770 48404
rect 3810 48364 3852 48404
rect 3892 48364 3934 48404
rect 3974 48364 4016 48404
rect 3688 48355 4056 48364
rect 4108 47312 4148 50884
rect 4396 50756 4436 51136
rect 4396 50707 4436 50716
rect 3688 46892 4056 46901
rect 3728 46852 3770 46892
rect 3810 46852 3852 46892
rect 3892 46852 3934 46892
rect 3974 46852 4016 46892
rect 3688 46843 4056 46852
rect 3688 45380 4056 45389
rect 3728 45340 3770 45380
rect 3810 45340 3852 45380
rect 3892 45340 3934 45380
rect 3974 45340 4016 45380
rect 3688 45331 4056 45340
rect 4108 44792 4148 47272
rect 4108 44743 4148 44752
rect 3688 43868 4056 43877
rect 3728 43828 3770 43868
rect 3810 43828 3852 43868
rect 3892 43828 3934 43868
rect 3974 43828 4016 43868
rect 3688 43819 4056 43828
rect 4108 43280 4148 43289
rect 3688 42356 4056 42365
rect 3728 42316 3770 42356
rect 3810 42316 3852 42356
rect 3892 42316 3934 42356
rect 3974 42316 4016 42356
rect 3688 42307 4056 42316
rect 4108 41180 4148 43240
rect 4108 41131 4148 41140
rect 4204 42188 4244 42197
rect 4204 41012 4244 42148
rect 4492 42188 4532 80032
rect 4684 79736 4724 81880
rect 4780 81871 4820 81880
rect 4928 80912 5296 80921
rect 4968 80872 5010 80912
rect 5050 80872 5092 80912
rect 5132 80872 5174 80912
rect 5214 80872 5256 80912
rect 4928 80863 5296 80872
rect 4684 79687 4724 79696
rect 4780 80492 4820 80501
rect 4684 78140 4724 78149
rect 4587 62180 4629 62189
rect 4587 62140 4588 62180
rect 4628 62140 4629 62180
rect 4587 62131 4629 62140
rect 4588 61844 4628 62131
rect 4588 61795 4628 61804
rect 4588 59408 4628 59417
rect 4588 57728 4628 59368
rect 4588 57679 4628 57688
rect 4588 53024 4628 53033
rect 4588 51176 4628 52984
rect 4588 51127 4628 51136
rect 4684 46640 4724 78100
rect 4780 76376 4820 80452
rect 4928 79400 5296 79409
rect 4968 79360 5010 79400
rect 5050 79360 5092 79400
rect 5132 79360 5174 79400
rect 5214 79360 5256 79400
rect 4928 79351 5296 79360
rect 4928 77888 5296 77897
rect 4968 77848 5010 77888
rect 5050 77848 5092 77888
rect 5132 77848 5174 77888
rect 5214 77848 5256 77888
rect 4928 77839 5296 77848
rect 5356 76796 5396 76805
rect 4780 76327 4820 76336
rect 4928 76376 5296 76385
rect 4968 76336 5010 76376
rect 5050 76336 5092 76376
rect 5132 76336 5174 76376
rect 5214 76336 5256 76376
rect 4928 76327 5296 76336
rect 4928 74864 5296 74873
rect 4968 74824 5010 74864
rect 5050 74824 5092 74864
rect 5132 74824 5174 74864
rect 5214 74824 5256 74864
rect 4928 74815 5296 74824
rect 4928 73352 5296 73361
rect 4968 73312 5010 73352
rect 5050 73312 5092 73352
rect 5132 73312 5174 73352
rect 5214 73312 5256 73352
rect 4928 73303 5296 73312
rect 4928 71840 5296 71849
rect 4968 71800 5010 71840
rect 5050 71800 5092 71840
rect 5132 71800 5174 71840
rect 5214 71800 5256 71840
rect 4928 71791 5296 71800
rect 4492 42139 4532 42148
rect 4588 46600 4724 46640
rect 4780 71336 4820 71345
rect 4108 40972 4244 41012
rect 4300 41516 4340 41525
rect 3688 40844 4056 40853
rect 3728 40804 3770 40844
rect 3810 40804 3852 40844
rect 3892 40804 3934 40844
rect 3974 40804 4016 40844
rect 3688 40795 4056 40804
rect 3688 39332 4056 39341
rect 3728 39292 3770 39332
rect 3810 39292 3852 39332
rect 3892 39292 3934 39332
rect 3974 39292 4016 39332
rect 3688 39283 4056 39292
rect 4108 38996 4148 40972
rect 4108 38947 4148 38956
rect 4204 40760 4244 40769
rect 4204 38828 4244 40720
rect 4300 39752 4340 41476
rect 4588 40676 4628 46600
rect 4780 43532 4820 71296
rect 4928 70328 5296 70337
rect 4968 70288 5010 70328
rect 5050 70288 5092 70328
rect 5132 70288 5174 70328
rect 5214 70288 5256 70328
rect 4928 70279 5296 70288
rect 5356 70160 5396 76756
rect 5356 70111 5396 70120
rect 4928 68816 5296 68825
rect 4968 68776 5010 68816
rect 5050 68776 5092 68816
rect 5132 68776 5174 68816
rect 5214 68776 5256 68816
rect 4928 68767 5296 68776
rect 5163 67808 5205 67817
rect 5163 67768 5164 67808
rect 5204 67768 5205 67808
rect 5163 67759 5205 67768
rect 5355 67808 5397 67817
rect 5355 67768 5356 67808
rect 5396 67768 5397 67808
rect 5355 67759 5397 67768
rect 5164 67674 5204 67759
rect 4928 67304 5296 67313
rect 4968 67264 5010 67304
rect 5050 67264 5092 67304
rect 5132 67264 5174 67304
rect 5214 67264 5256 67304
rect 4928 67255 5296 67264
rect 4928 65792 5296 65801
rect 4968 65752 5010 65792
rect 5050 65752 5092 65792
rect 5132 65752 5174 65792
rect 5214 65752 5256 65792
rect 4928 65743 5296 65752
rect 4928 64280 5296 64289
rect 4968 64240 5010 64280
rect 5050 64240 5092 64280
rect 5132 64240 5174 64280
rect 5214 64240 5256 64280
rect 4928 64231 5296 64240
rect 4928 62768 5296 62777
rect 4968 62728 5010 62768
rect 5050 62728 5092 62768
rect 5132 62728 5174 62768
rect 5214 62728 5256 62768
rect 4928 62719 5296 62728
rect 5356 62768 5396 67759
rect 5356 62719 5396 62728
rect 4928 61256 5296 61265
rect 4968 61216 5010 61256
rect 5050 61216 5092 61256
rect 5132 61216 5174 61256
rect 5214 61216 5256 61256
rect 4928 61207 5296 61216
rect 4928 59744 5296 59753
rect 4968 59704 5010 59744
rect 5050 59704 5092 59744
rect 5132 59704 5174 59744
rect 5214 59704 5256 59744
rect 4928 59695 5296 59704
rect 4928 58232 5296 58241
rect 4968 58192 5010 58232
rect 5050 58192 5092 58232
rect 5132 58192 5174 58232
rect 5214 58192 5256 58232
rect 4928 58183 5296 58192
rect 4928 56720 5296 56729
rect 4968 56680 5010 56720
rect 5050 56680 5092 56720
rect 5132 56680 5174 56720
rect 5214 56680 5256 56720
rect 4928 56671 5296 56680
rect 4928 55208 5296 55217
rect 4968 55168 5010 55208
rect 5050 55168 5092 55208
rect 5132 55168 5174 55208
rect 5214 55168 5256 55208
rect 4928 55159 5296 55168
rect 4928 53696 5296 53705
rect 4968 53656 5010 53696
rect 5050 53656 5092 53696
rect 5132 53656 5174 53696
rect 5214 53656 5256 53696
rect 4928 53647 5296 53656
rect 5067 52772 5109 52781
rect 5067 52732 5068 52772
rect 5108 52732 5109 52772
rect 5067 52723 5109 52732
rect 5068 52638 5108 52723
rect 4928 52184 5296 52193
rect 4968 52144 5010 52184
rect 5050 52144 5092 52184
rect 5132 52144 5174 52184
rect 5214 52144 5256 52184
rect 4928 52135 5296 52144
rect 4928 50672 5296 50681
rect 4968 50632 5010 50672
rect 5050 50632 5092 50672
rect 5132 50632 5174 50672
rect 5214 50632 5256 50672
rect 4928 50623 5296 50632
rect 4928 49160 5296 49169
rect 4968 49120 5010 49160
rect 5050 49120 5092 49160
rect 5132 49120 5174 49160
rect 5214 49120 5256 49160
rect 4928 49111 5296 49120
rect 4928 47648 5296 47657
rect 4968 47608 5010 47648
rect 5050 47608 5092 47648
rect 5132 47608 5174 47648
rect 5214 47608 5256 47648
rect 4928 47599 5296 47608
rect 4928 46136 5296 46145
rect 4968 46096 5010 46136
rect 5050 46096 5092 46136
rect 5132 46096 5174 46136
rect 5214 46096 5256 46136
rect 4928 46087 5296 46096
rect 4928 44624 5296 44633
rect 4968 44584 5010 44624
rect 5050 44584 5092 44624
rect 5132 44584 5174 44624
rect 5214 44584 5256 44624
rect 4928 44575 5296 44584
rect 4780 41945 4820 43492
rect 4928 43112 5296 43121
rect 4968 43072 5010 43112
rect 5050 43072 5092 43112
rect 5132 43072 5174 43112
rect 5214 43072 5256 43112
rect 4928 43063 5296 43072
rect 4779 41936 4821 41945
rect 4779 41896 4780 41936
rect 4820 41896 4821 41936
rect 4779 41887 4821 41896
rect 4928 41600 5296 41609
rect 4968 41560 5010 41600
rect 5050 41560 5092 41600
rect 5132 41560 5174 41600
rect 5214 41560 5256 41600
rect 4928 41551 5296 41560
rect 4300 39703 4340 39712
rect 4492 40636 4628 40676
rect 4684 41096 4724 41105
rect 4299 39080 4341 39089
rect 4299 39040 4300 39080
rect 4340 39040 4341 39080
rect 4299 39031 4341 39040
rect 4204 38779 4244 38788
rect 3688 37820 4056 37829
rect 3728 37780 3770 37820
rect 3810 37780 3852 37820
rect 3892 37780 3934 37820
rect 3974 37780 4016 37820
rect 3688 37771 4056 37780
rect 3820 37652 3860 37661
rect 3820 37493 3860 37612
rect 3819 37484 3861 37493
rect 3819 37444 3820 37484
rect 3860 37444 3861 37484
rect 3819 37435 3861 37444
rect 4107 37316 4149 37325
rect 4107 37276 4108 37316
rect 4148 37276 4149 37316
rect 4107 37267 4149 37276
rect 4108 36737 4148 37267
rect 4107 36728 4149 36737
rect 4107 36688 4108 36728
rect 4148 36688 4149 36728
rect 4107 36679 4149 36688
rect 3688 36308 4056 36317
rect 3728 36268 3770 36308
rect 3810 36268 3852 36308
rect 3892 36268 3934 36308
rect 3974 36268 4016 36308
rect 3688 36259 4056 36268
rect 3532 35251 3572 35260
rect 3688 34796 4056 34805
rect 3728 34756 3770 34796
rect 3810 34756 3852 34796
rect 3892 34756 3934 34796
rect 3974 34756 4016 34796
rect 3688 34747 4056 34756
rect 4011 33872 4053 33881
rect 4011 33832 4012 33872
rect 4052 33832 4053 33872
rect 4011 33823 4053 33832
rect 4012 33738 4052 33823
rect 3688 33284 4056 33293
rect 3728 33244 3770 33284
rect 3810 33244 3852 33284
rect 3892 33244 3934 33284
rect 3974 33244 4016 33284
rect 3688 33235 4056 33244
rect 3532 32276 3572 32285
rect 3340 28960 3476 29000
rect 3244 26767 3284 26776
rect 2956 26347 2996 26356
rect 3148 26480 3188 26489
rect 2860 22231 2900 22240
rect 2956 25388 2996 25397
rect 2764 18164 2804 18173
rect 2764 17660 2804 18124
rect 2764 17611 2804 17620
rect 2764 15644 2804 15653
rect 2764 9932 2804 15604
rect 2764 9883 2804 9892
rect 2860 9176 2900 9185
rect 2860 8672 2900 9136
rect 2764 8168 2804 8177
rect 2764 2120 2804 8128
rect 2860 7916 2900 8632
rect 2860 7867 2900 7876
rect 2764 2071 2804 2080
rect 2956 1280 2996 25348
rect 3148 20096 3188 26440
rect 3340 26396 3380 26405
rect 3244 23960 3284 23969
rect 3244 23792 3284 23920
rect 3244 23743 3284 23752
rect 3340 22532 3380 26356
rect 3340 22483 3380 22492
rect 3436 26144 3476 28960
rect 3436 25472 3476 26104
rect 3436 21776 3476 25432
rect 3532 22028 3572 32236
rect 3688 31772 4056 31781
rect 3728 31732 3770 31772
rect 3810 31732 3852 31772
rect 3892 31732 3934 31772
rect 3974 31732 4016 31772
rect 3688 31723 4056 31732
rect 4204 31352 4244 31361
rect 3688 30260 4056 30269
rect 3728 30220 3770 30260
rect 3810 30220 3852 30260
rect 3892 30220 3934 30260
rect 3974 30220 4016 30260
rect 3688 30211 4056 30220
rect 4107 29672 4149 29681
rect 4107 29632 4108 29672
rect 4148 29632 4149 29672
rect 4107 29623 4149 29632
rect 4108 29538 4148 29623
rect 3688 28748 4056 28757
rect 3728 28708 3770 28748
rect 3810 28708 3852 28748
rect 3892 28708 3934 28748
rect 3974 28708 4016 28748
rect 3688 28699 4056 28708
rect 4204 27404 4244 31312
rect 4204 27355 4244 27364
rect 4300 29840 4340 39031
rect 4492 38660 4532 40636
rect 4684 39752 4724 41056
rect 4928 40088 5296 40097
rect 4968 40048 5010 40088
rect 5050 40048 5092 40088
rect 5132 40048 5174 40088
rect 5214 40048 5256 40088
rect 4928 40039 5296 40048
rect 4684 39703 4724 39712
rect 4492 38611 4532 38620
rect 4780 38912 4820 38921
rect 4684 38408 4724 38417
rect 4684 35729 4724 38368
rect 4683 35720 4725 35729
rect 4683 35680 4684 35720
rect 4724 35680 4725 35720
rect 4683 35671 4725 35680
rect 4684 34040 4724 34049
rect 4684 33452 4724 34000
rect 3688 27236 4056 27245
rect 3728 27196 3770 27236
rect 3810 27196 3852 27236
rect 3892 27196 3934 27236
rect 3974 27196 4016 27236
rect 3688 27187 4056 27196
rect 3688 25724 4056 25733
rect 3728 25684 3770 25724
rect 3810 25684 3852 25724
rect 3892 25684 3934 25724
rect 3974 25684 4016 25724
rect 3688 25675 4056 25684
rect 4300 24380 4340 29800
rect 4492 33412 4684 33452
rect 4492 29000 4532 33412
rect 4684 33403 4724 33412
rect 4684 33032 4724 33041
rect 4300 24331 4340 24340
rect 4396 28960 4532 29000
rect 4588 31856 4628 31865
rect 4396 25304 4436 28960
rect 4588 27908 4628 31816
rect 4492 27868 4628 27908
rect 4492 26816 4532 27868
rect 4587 27740 4629 27749
rect 4587 27700 4588 27740
rect 4628 27700 4629 27740
rect 4587 27691 4629 27700
rect 4588 27606 4628 27691
rect 4492 26767 4532 26776
rect 4684 26144 4724 32992
rect 4684 26095 4724 26104
rect 4491 25976 4533 25985
rect 4491 25936 4492 25976
rect 4532 25936 4533 25976
rect 4491 25927 4533 25936
rect 4492 25842 4532 25927
rect 3688 24212 4056 24221
rect 3728 24172 3770 24212
rect 3810 24172 3852 24212
rect 3892 24172 3934 24212
rect 3974 24172 4016 24212
rect 3688 24163 4056 24172
rect 4300 23624 4340 23633
rect 3688 22700 4056 22709
rect 3728 22660 3770 22700
rect 3810 22660 3852 22700
rect 3892 22660 3934 22700
rect 3974 22660 4016 22700
rect 3688 22651 4056 22660
rect 3532 21979 3572 21988
rect 3436 21727 3476 21736
rect 3148 19004 3188 20056
rect 3148 18955 3188 18964
rect 3532 21524 3572 21533
rect 3340 16988 3380 16997
rect 3340 13964 3380 16948
rect 3532 14048 3572 21484
rect 3688 21188 4056 21197
rect 3728 21148 3770 21188
rect 3810 21148 3852 21188
rect 3892 21148 3934 21188
rect 3974 21148 4016 21188
rect 3688 21139 4056 21148
rect 3688 19676 4056 19685
rect 3728 19636 3770 19676
rect 3810 19636 3852 19676
rect 3892 19636 3934 19676
rect 3974 19636 4016 19676
rect 3688 19627 4056 19636
rect 3688 18164 4056 18173
rect 3728 18124 3770 18164
rect 3810 18124 3852 18164
rect 3892 18124 3934 18164
rect 3974 18124 4016 18164
rect 3688 18115 4056 18124
rect 3688 16652 4056 16661
rect 3728 16612 3770 16652
rect 3810 16612 3852 16652
rect 3892 16612 3934 16652
rect 3974 16612 4016 16652
rect 3688 16603 4056 16612
rect 3688 15140 4056 15149
rect 3728 15100 3770 15140
rect 3810 15100 3852 15140
rect 3892 15100 3934 15140
rect 3974 15100 4016 15140
rect 3688 15091 4056 15100
rect 3532 13999 3572 14008
rect 3340 13915 3380 13924
rect 3688 13628 4056 13637
rect 3728 13588 3770 13628
rect 3810 13588 3852 13628
rect 3892 13588 3934 13628
rect 3974 13588 4016 13628
rect 3688 13579 4056 13588
rect 3340 12956 3380 12965
rect 3148 11948 3188 11957
rect 3052 11612 3092 11621
rect 3052 2288 3092 11572
rect 3148 10184 3188 11908
rect 3148 10135 3188 10144
rect 3244 10604 3284 10613
rect 3148 9764 3188 9773
rect 3148 4220 3188 9724
rect 3244 9596 3284 10564
rect 3340 10016 3380 12916
rect 3688 12116 4056 12125
rect 3728 12076 3770 12116
rect 3810 12076 3852 12116
rect 3892 12076 3934 12116
rect 3974 12076 4016 12116
rect 3688 12067 4056 12076
rect 4108 11696 4148 11705
rect 3435 10940 3477 10949
rect 3435 10900 3436 10940
rect 3476 10900 3477 10940
rect 3435 10891 3477 10900
rect 3340 9967 3380 9976
rect 3244 9547 3284 9556
rect 3340 9512 3380 9521
rect 3340 8924 3380 9472
rect 3340 8875 3380 8884
rect 3244 8672 3284 8681
rect 3244 8504 3284 8632
rect 3244 8455 3284 8464
rect 3436 5144 3476 10891
rect 3436 5095 3476 5104
rect 3532 10772 3572 10781
rect 3148 4171 3188 4180
rect 3340 3548 3380 3557
rect 3052 2239 3092 2248
rect 3244 2540 3284 2549
rect 3244 2288 3284 2500
rect 3244 2239 3284 2248
rect 2956 1231 2996 1240
rect 3340 1112 3380 3508
rect 3340 1063 3380 1072
rect 2668 979 2708 988
rect 1420 727 1460 736
rect 2955 608 2997 617
rect 2955 568 2956 608
rect 2996 568 2997 608
rect 2955 559 2997 568
rect 2956 474 2996 559
rect 3532 272 3572 10732
rect 3688 10604 4056 10613
rect 3728 10564 3770 10604
rect 3810 10564 3852 10604
rect 3892 10564 3934 10604
rect 3974 10564 4016 10604
rect 3688 10555 4056 10564
rect 4108 9764 4148 11656
rect 4204 11024 4244 11033
rect 4204 10604 4244 10984
rect 4204 10555 4244 10564
rect 4300 10100 4340 23584
rect 4300 10051 4340 10060
rect 4396 19172 4436 25264
rect 4108 9715 4148 9724
rect 4108 9260 4148 9269
rect 3688 9092 4056 9101
rect 3728 9052 3770 9092
rect 3810 9052 3852 9092
rect 3892 9052 3934 9092
rect 3974 9052 4016 9092
rect 3688 9043 4056 9052
rect 3688 7580 4056 7589
rect 3728 7540 3770 7580
rect 3810 7540 3852 7580
rect 3892 7540 3934 7580
rect 3974 7540 4016 7580
rect 3688 7531 4056 7540
rect 3688 6068 4056 6077
rect 3728 6028 3770 6068
rect 3810 6028 3852 6068
rect 3892 6028 3934 6068
rect 3974 6028 4016 6068
rect 3688 6019 4056 6028
rect 3688 4556 4056 4565
rect 3728 4516 3770 4556
rect 3810 4516 3852 4556
rect 3892 4516 3934 4556
rect 3974 4516 4016 4556
rect 3688 4507 4056 4516
rect 4108 4136 4148 9220
rect 4204 8756 4244 8765
rect 4204 5900 4244 8716
rect 4396 8672 4436 19132
rect 4588 23708 4628 23717
rect 4588 22868 4628 23668
rect 4492 16400 4532 16409
rect 4492 15476 4532 16360
rect 4492 15427 4532 15436
rect 4588 14972 4628 22828
rect 4684 22364 4724 22373
rect 4684 16904 4724 22324
rect 4684 16855 4724 16864
rect 4588 14132 4628 14932
rect 4588 14083 4628 14092
rect 4684 12116 4724 12125
rect 4204 5851 4244 5860
rect 4300 8084 4340 8093
rect 4300 4808 4340 8044
rect 4396 8000 4436 8632
rect 4588 8924 4628 8933
rect 4396 7951 4436 7960
rect 4492 8504 4532 8513
rect 4492 5312 4532 8464
rect 4492 5263 4532 5272
rect 4300 4759 4340 4768
rect 4203 4556 4245 4565
rect 4203 4516 4204 4556
rect 4244 4516 4245 4556
rect 4203 4507 4245 4516
rect 4108 4087 4148 4096
rect 4204 3800 4244 4507
rect 4108 3760 4244 3800
rect 3688 3044 4056 3053
rect 3728 3004 3770 3044
rect 3810 3004 3852 3044
rect 3892 3004 3934 3044
rect 3974 3004 4016 3044
rect 3688 2995 4056 3004
rect 3627 2792 3669 2801
rect 3627 2752 3628 2792
rect 3668 2752 3669 2792
rect 3627 2743 3669 2752
rect 4108 2792 4148 3760
rect 4588 3380 4628 8884
rect 4684 8000 4724 12076
rect 4684 7951 4724 7960
rect 4588 3331 4628 3340
rect 4684 7076 4724 7085
rect 4108 2743 4148 2752
rect 3628 2658 3668 2743
rect 3688 1532 4056 1541
rect 3728 1492 3770 1532
rect 3810 1492 3852 1532
rect 3892 1492 3934 1532
rect 3974 1492 4016 1532
rect 3688 1483 4056 1492
rect 4684 1280 4724 7036
rect 4684 1231 4724 1240
rect 4780 944 4820 38872
rect 4928 38576 5296 38585
rect 4968 38536 5010 38576
rect 5050 38536 5092 38576
rect 5132 38536 5174 38576
rect 5214 38536 5256 38576
rect 4928 38527 5296 38536
rect 5356 37568 5396 37577
rect 4928 37064 5296 37073
rect 4968 37024 5010 37064
rect 5050 37024 5092 37064
rect 5132 37024 5174 37064
rect 5214 37024 5256 37064
rect 4928 37015 5296 37024
rect 4928 35552 5296 35561
rect 4968 35512 5010 35552
rect 5050 35512 5092 35552
rect 5132 35512 5174 35552
rect 5214 35512 5256 35552
rect 4928 35503 5296 35512
rect 4928 34040 5296 34049
rect 4968 34000 5010 34040
rect 5050 34000 5092 34040
rect 5132 34000 5174 34040
rect 5214 34000 5256 34040
rect 4928 33991 5296 34000
rect 4928 32528 5296 32537
rect 4968 32488 5010 32528
rect 5050 32488 5092 32528
rect 5132 32488 5174 32528
rect 5214 32488 5256 32528
rect 4928 32479 5296 32488
rect 4928 31016 5296 31025
rect 4968 30976 5010 31016
rect 5050 30976 5092 31016
rect 5132 30976 5174 31016
rect 5214 30976 5256 31016
rect 4928 30967 5296 30976
rect 4928 29504 5296 29513
rect 4968 29464 5010 29504
rect 5050 29464 5092 29504
rect 5132 29464 5174 29504
rect 5214 29464 5256 29504
rect 4928 29455 5296 29464
rect 5356 29168 5396 37528
rect 5356 29119 5396 29128
rect 4928 27992 5296 28001
rect 4968 27952 5010 27992
rect 5050 27952 5092 27992
rect 5132 27952 5174 27992
rect 5214 27952 5256 27992
rect 4928 27943 5296 27952
rect 4928 26480 5296 26489
rect 4968 26440 5010 26480
rect 5050 26440 5092 26480
rect 5132 26440 5174 26480
rect 5214 26440 5256 26480
rect 4928 26431 5296 26440
rect 4928 24968 5296 24977
rect 4968 24928 5010 24968
rect 5050 24928 5092 24968
rect 5132 24928 5174 24968
rect 5214 24928 5256 24968
rect 4928 24919 5296 24928
rect 4928 23456 5296 23465
rect 4968 23416 5010 23456
rect 5050 23416 5092 23456
rect 5132 23416 5174 23456
rect 5214 23416 5256 23456
rect 4928 23407 5296 23416
rect 5356 22196 5396 22205
rect 4928 21944 5296 21953
rect 4968 21904 5010 21944
rect 5050 21904 5092 21944
rect 5132 21904 5174 21944
rect 5214 21904 5256 21944
rect 4928 21895 5296 21904
rect 4928 20432 5296 20441
rect 4968 20392 5010 20432
rect 5050 20392 5092 20432
rect 5132 20392 5174 20432
rect 5214 20392 5256 20432
rect 4928 20383 5296 20392
rect 4928 18920 5296 18929
rect 4968 18880 5010 18920
rect 5050 18880 5092 18920
rect 5132 18880 5174 18920
rect 5214 18880 5256 18920
rect 4928 18871 5296 18880
rect 4928 17408 5296 17417
rect 4968 17368 5010 17408
rect 5050 17368 5092 17408
rect 5132 17368 5174 17408
rect 5214 17368 5256 17408
rect 4928 17359 5296 17368
rect 4928 15896 5296 15905
rect 4968 15856 5010 15896
rect 5050 15856 5092 15896
rect 5132 15856 5174 15896
rect 5214 15856 5256 15896
rect 4928 15847 5296 15856
rect 4928 14384 5296 14393
rect 4968 14344 5010 14384
rect 5050 14344 5092 14384
rect 5132 14344 5174 14384
rect 5214 14344 5256 14384
rect 4928 14335 5296 14344
rect 5356 13796 5396 22156
rect 5356 13747 5396 13756
rect 4928 12872 5296 12881
rect 4968 12832 5010 12872
rect 5050 12832 5092 12872
rect 5132 12832 5174 12872
rect 5214 12832 5256 12872
rect 4928 12823 5296 12832
rect 4928 11360 5296 11369
rect 4968 11320 5010 11360
rect 5050 11320 5092 11360
rect 5132 11320 5174 11360
rect 5214 11320 5256 11360
rect 4928 11311 5296 11320
rect 4875 10940 4917 10949
rect 4875 10900 4876 10940
rect 4916 10900 4917 10940
rect 4875 10891 4917 10900
rect 4876 10806 4916 10891
rect 5356 10520 5396 10529
rect 4928 9848 5296 9857
rect 4968 9808 5010 9848
rect 5050 9808 5092 9848
rect 5132 9808 5174 9848
rect 5214 9808 5256 9848
rect 4928 9799 5296 9808
rect 4928 8336 5296 8345
rect 4968 8296 5010 8336
rect 5050 8296 5092 8336
rect 5132 8296 5174 8336
rect 5214 8296 5256 8336
rect 4928 8287 5296 8296
rect 4928 6824 5296 6833
rect 4968 6784 5010 6824
rect 5050 6784 5092 6824
rect 5132 6784 5174 6824
rect 5214 6784 5256 6824
rect 4928 6775 5296 6784
rect 5356 5648 5396 10480
rect 5356 5599 5396 5608
rect 4928 5312 5296 5321
rect 4968 5272 5010 5312
rect 5050 5272 5092 5312
rect 5132 5272 5174 5312
rect 5214 5272 5256 5312
rect 4928 5263 5296 5272
rect 5452 4976 5492 81880
rect 5548 80072 5588 80081
rect 5548 75041 5588 80032
rect 5547 75032 5589 75041
rect 5547 74992 5548 75032
rect 5588 74992 5589 75032
rect 5547 74983 5589 74992
rect 5548 24800 5588 74983
rect 5644 70832 5684 70841
rect 5644 37316 5684 70792
rect 5644 36569 5684 37276
rect 5643 36560 5685 36569
rect 5643 36520 5644 36560
rect 5684 36520 5685 36560
rect 5643 36511 5685 36520
rect 5644 31940 5684 31949
rect 5644 30260 5684 31900
rect 5740 31268 5780 82720
rect 5836 82172 5876 82181
rect 5836 79820 5876 82132
rect 5836 79771 5876 79780
rect 5932 67640 5972 67649
rect 5836 63944 5876 63953
rect 5836 62684 5876 63904
rect 5836 62635 5876 62644
rect 5836 38408 5876 38417
rect 5836 36728 5876 38368
rect 5836 36679 5876 36688
rect 5835 35720 5877 35729
rect 5835 35680 5836 35720
rect 5876 35680 5877 35720
rect 5835 35671 5877 35680
rect 5836 35552 5876 35671
rect 5836 32696 5876 35512
rect 5836 32647 5876 32656
rect 5740 31219 5780 31228
rect 5644 30211 5684 30220
rect 5835 29168 5877 29177
rect 5835 29128 5836 29168
rect 5876 29128 5877 29168
rect 5835 29119 5877 29128
rect 5836 29034 5876 29119
rect 5644 28664 5684 28673
rect 5644 27656 5684 28624
rect 5836 28412 5876 28421
rect 5644 27607 5684 27616
rect 5740 28076 5780 28085
rect 5644 26480 5684 26489
rect 5644 25220 5684 26440
rect 5644 25171 5684 25180
rect 5548 24751 5588 24760
rect 5548 23792 5588 23801
rect 5548 22868 5588 23752
rect 5548 22819 5588 22828
rect 5740 19844 5780 28036
rect 5836 25220 5876 28372
rect 5836 25171 5876 25180
rect 5740 19424 5780 19804
rect 5740 19375 5780 19384
rect 5548 14552 5588 14561
rect 5548 5564 5588 14512
rect 5740 13880 5780 13889
rect 5644 13796 5684 13805
rect 5644 13208 5684 13756
rect 5644 9512 5684 13168
rect 5644 9463 5684 9472
rect 5740 5648 5780 13840
rect 5548 5515 5588 5524
rect 5644 5608 5780 5648
rect 5452 4927 5492 4936
rect 4971 4556 5013 4565
rect 4971 4516 4972 4556
rect 5012 4516 5013 4556
rect 4971 4507 5013 4516
rect 4972 4422 5012 4507
rect 4928 3800 5296 3809
rect 4968 3760 5010 3800
rect 5050 3760 5092 3800
rect 5132 3760 5174 3800
rect 5214 3760 5256 3800
rect 4928 3751 5296 3760
rect 4928 2288 5296 2297
rect 4968 2248 5010 2288
rect 5050 2248 5092 2288
rect 5132 2248 5174 2288
rect 5214 2248 5256 2288
rect 4928 2239 5296 2248
rect 5644 2036 5684 5608
rect 5644 1987 5684 1996
rect 5740 3968 5780 3977
rect 5740 1877 5780 3928
rect 5932 3548 5972 67600
rect 6028 64364 6068 84400
rect 6412 84440 6452 84449
rect 6316 83264 6356 83273
rect 6316 83012 6356 83224
rect 6028 64315 6068 64324
rect 6124 79568 6164 79577
rect 6028 63104 6068 63113
rect 6028 61088 6068 63064
rect 6028 61039 6068 61048
rect 6028 60248 6068 60257
rect 6028 54452 6068 60208
rect 6028 54403 6068 54412
rect 6028 51764 6068 51773
rect 6028 50756 6068 51724
rect 6028 50707 6068 50716
rect 6028 37736 6068 37745
rect 6028 34124 6068 37696
rect 6028 34075 6068 34084
rect 6027 30848 6069 30857
rect 6027 30808 6028 30848
rect 6068 30808 6069 30848
rect 6027 30799 6069 30808
rect 6028 22448 6068 30799
rect 6028 18584 6068 22408
rect 6028 18535 6068 18544
rect 6028 12788 6068 12797
rect 6028 11192 6068 12748
rect 6028 11143 6068 11152
rect 6124 5732 6164 79528
rect 6316 68480 6356 82972
rect 6412 76889 6452 84400
rect 6604 84440 6644 84449
rect 6508 82172 6548 82181
rect 6411 76880 6453 76889
rect 6411 76840 6412 76880
rect 6452 76840 6453 76880
rect 6411 76831 6453 76840
rect 6316 68431 6356 68440
rect 6412 67556 6452 67565
rect 6219 67472 6261 67481
rect 6219 67432 6220 67472
rect 6260 67432 6261 67472
rect 6219 67423 6261 67432
rect 6220 43028 6260 67423
rect 6220 42979 6260 42988
rect 6316 64448 6356 64457
rect 6220 39080 6260 39089
rect 6220 30857 6260 39040
rect 6316 37661 6356 64408
rect 6315 37652 6357 37661
rect 6315 37612 6316 37652
rect 6356 37612 6357 37652
rect 6315 37603 6357 37612
rect 6315 37484 6357 37493
rect 6315 37444 6316 37484
rect 6356 37444 6357 37484
rect 6315 37435 6357 37444
rect 6316 37350 6356 37435
rect 6412 33881 6452 67516
rect 6508 42860 6548 82132
rect 6508 42811 6548 42820
rect 6507 41684 6549 41693
rect 6507 41644 6508 41684
rect 6548 41644 6549 41684
rect 6507 41635 6549 41644
rect 6508 40676 6548 41635
rect 6508 40627 6548 40636
rect 6507 37652 6549 37661
rect 6507 37612 6508 37652
rect 6548 37612 6549 37652
rect 6507 37603 6549 37612
rect 6411 33872 6453 33881
rect 6411 33832 6412 33872
rect 6452 33832 6453 33872
rect 6411 33823 6453 33832
rect 6412 33620 6452 33629
rect 6219 30848 6261 30857
rect 6219 30808 6220 30848
rect 6260 30808 6261 30848
rect 6219 30799 6261 30808
rect 6316 29840 6356 29849
rect 6316 28748 6356 29800
rect 6316 28699 6356 28708
rect 6412 28580 6452 33580
rect 6508 31268 6548 37603
rect 6508 31219 6548 31228
rect 6412 28531 6452 28540
rect 6508 30260 6548 30269
rect 6508 28076 6548 30220
rect 6508 28027 6548 28036
rect 6508 26984 6548 26993
rect 6220 26900 6260 26909
rect 6220 24548 6260 26860
rect 6411 26900 6453 26909
rect 6411 26860 6412 26900
rect 6452 26860 6453 26900
rect 6411 26851 6453 26860
rect 6412 26766 6452 26851
rect 6220 24499 6260 24508
rect 6316 26648 6356 26657
rect 6220 11864 6260 11873
rect 6220 8840 6260 11824
rect 6220 8791 6260 8800
rect 6316 6656 6356 26608
rect 6411 25976 6453 25985
rect 6411 25936 6412 25976
rect 6452 25936 6453 25976
rect 6411 25927 6453 25936
rect 6412 25842 6452 25927
rect 6412 25388 6452 25397
rect 6412 24968 6452 25348
rect 6508 25136 6548 26944
rect 6508 25087 6548 25096
rect 6412 24919 6452 24928
rect 6412 24800 6452 24809
rect 6412 18332 6452 24760
rect 6412 18283 6452 18292
rect 6508 22112 6548 22121
rect 6316 6607 6356 6616
rect 6412 7748 6452 7757
rect 6412 6236 6452 7708
rect 6412 6187 6452 6196
rect 6508 6068 6548 22072
rect 6604 16568 6644 84400
rect 6987 80660 7029 80669
rect 6987 80620 6988 80660
rect 7028 80620 7029 80660
rect 6987 80611 7029 80620
rect 6988 80492 7028 80611
rect 6988 80443 7028 80452
rect 6796 79736 6836 79745
rect 6700 76208 6740 76217
rect 6700 75881 6740 76168
rect 6699 75872 6741 75881
rect 6699 75832 6700 75872
rect 6740 75832 6741 75872
rect 6699 75823 6741 75832
rect 6700 66716 6740 66725
rect 6700 34292 6740 66676
rect 6700 34243 6740 34252
rect 6796 29681 6836 79696
rect 6892 79400 6932 79409
rect 6892 73604 6932 79360
rect 7180 79232 7220 79241
rect 7180 78980 7220 79192
rect 7180 78931 7220 78940
rect 6892 73555 6932 73564
rect 7084 78896 7124 78905
rect 6988 70748 7028 70757
rect 6892 68984 6932 68993
rect 6892 68480 6932 68944
rect 6892 64364 6932 68440
rect 6988 66044 7028 70708
rect 6988 65995 7028 66004
rect 6892 64315 6932 64324
rect 6988 60668 7028 60677
rect 6891 59240 6933 59249
rect 6891 59200 6892 59240
rect 6932 59200 6933 59240
rect 6891 59191 6933 59200
rect 6892 59106 6932 59191
rect 6988 57224 7028 60628
rect 6988 57175 7028 57184
rect 6892 52520 6932 52529
rect 6892 46472 6932 52480
rect 6892 46423 6932 46432
rect 6892 43700 6932 43709
rect 6892 41693 6932 43660
rect 6891 41684 6933 41693
rect 6891 41644 6892 41684
rect 6932 41644 6933 41684
rect 6891 41635 6933 41644
rect 6987 41600 7029 41609
rect 6987 41560 6988 41600
rect 7028 41560 7029 41600
rect 6987 41551 7029 41560
rect 6892 41432 6932 41441
rect 6892 41096 6932 41392
rect 6892 41047 6932 41056
rect 6892 40508 6932 40517
rect 6892 39416 6932 40468
rect 6892 39367 6932 39376
rect 6988 36896 7028 41551
rect 6988 36847 7028 36856
rect 6987 36728 7029 36737
rect 6987 36688 6988 36728
rect 7028 36688 7029 36728
rect 6987 36679 7029 36688
rect 6892 34712 6932 34721
rect 6892 32780 6932 34672
rect 6892 32731 6932 32740
rect 6892 29924 6932 29933
rect 6795 29672 6837 29681
rect 6795 29632 6796 29672
rect 6836 29632 6837 29672
rect 6795 29623 6837 29632
rect 6796 29420 6836 29429
rect 6700 29336 6740 29345
rect 6700 22364 6740 29296
rect 6796 28160 6836 29380
rect 6796 28111 6836 28120
rect 6892 26564 6932 29884
rect 6892 26515 6932 26524
rect 6700 22315 6740 22324
rect 6796 26396 6836 26405
rect 6796 18416 6836 26356
rect 6796 18367 6836 18376
rect 6892 17408 6932 17417
rect 6604 16519 6644 16528
rect 6700 16652 6740 16661
rect 6700 14216 6740 16612
rect 6700 14167 6740 14176
rect 6892 11864 6932 17368
rect 6988 12629 7028 36679
rect 6987 12620 7029 12629
rect 6987 12580 6988 12620
rect 7028 12580 7029 12620
rect 6987 12571 7029 12580
rect 6892 11815 6932 11824
rect 7084 11360 7124 78856
rect 7180 70160 7220 70169
rect 7180 65876 7220 70120
rect 7276 66800 7316 85660
rect 7756 85616 7796 85625
rect 7660 84944 7700 84953
rect 7468 82844 7508 82853
rect 7276 66751 7316 66760
rect 7372 82760 7412 82769
rect 7180 65827 7220 65836
rect 7276 66380 7316 66389
rect 7276 65792 7316 66340
rect 7276 65743 7316 65752
rect 7276 59660 7316 59669
rect 7276 57308 7316 59620
rect 7276 57259 7316 57268
rect 7372 43196 7412 82720
rect 7468 80837 7508 82804
rect 7467 80828 7509 80837
rect 7467 80788 7468 80828
rect 7508 80788 7509 80828
rect 7467 80779 7509 80788
rect 7180 41768 7220 41777
rect 7180 40508 7220 41728
rect 7275 41432 7317 41441
rect 7275 41392 7276 41432
rect 7316 41392 7317 41432
rect 7275 41383 7317 41392
rect 7180 40459 7220 40468
rect 7179 39080 7221 39089
rect 7179 39040 7180 39080
rect 7220 39040 7221 39080
rect 7179 39031 7221 39040
rect 7180 38946 7220 39031
rect 7179 36560 7221 36569
rect 7179 36520 7180 36560
rect 7220 36520 7221 36560
rect 7179 36511 7221 36520
rect 7180 27572 7220 36511
rect 7276 27656 7316 41383
rect 7372 40592 7412 43156
rect 7372 40543 7412 40552
rect 7468 80492 7508 80501
rect 7468 38828 7508 80452
rect 7660 80156 7700 84904
rect 7660 80107 7700 80116
rect 7756 79493 7796 85576
rect 8524 85028 8564 85037
rect 8139 82844 8181 82853
rect 8139 82804 8140 82844
rect 8180 82804 8181 82844
rect 8139 82795 8181 82804
rect 7852 81332 7892 81341
rect 7755 79484 7797 79493
rect 7755 79444 7756 79484
rect 7796 79444 7797 79484
rect 7755 79435 7797 79444
rect 7564 75536 7604 75545
rect 7564 68396 7604 75496
rect 7756 74612 7796 74621
rect 7660 73520 7700 73529
rect 7660 73109 7700 73480
rect 7659 73100 7701 73109
rect 7659 73060 7660 73100
rect 7700 73060 7701 73100
rect 7659 73051 7701 73060
rect 7564 68356 7700 68396
rect 7660 67136 7700 68356
rect 7564 66464 7604 66473
rect 7564 64616 7604 66424
rect 7564 61853 7604 64576
rect 7563 61844 7605 61853
rect 7563 61804 7564 61844
rect 7604 61804 7605 61844
rect 7563 61795 7605 61804
rect 7564 61088 7604 61097
rect 7564 60920 7604 61048
rect 7564 60871 7604 60880
rect 7564 60584 7604 60593
rect 7564 41609 7604 60544
rect 7660 57476 7700 67096
rect 7756 62936 7796 74572
rect 7852 70916 7892 81292
rect 8044 80492 8084 80501
rect 8044 79820 8084 80452
rect 7948 79232 7988 79241
rect 7948 72008 7988 79192
rect 7948 71959 7988 71968
rect 7852 70867 7892 70876
rect 7756 62887 7796 62896
rect 7948 70664 7988 70673
rect 7851 61844 7893 61853
rect 7851 61804 7852 61844
rect 7892 61804 7893 61844
rect 7851 61795 7893 61804
rect 7660 57427 7700 57436
rect 7756 60248 7796 60257
rect 7756 57224 7796 60208
rect 7756 57175 7796 57184
rect 7660 55544 7700 55553
rect 7660 54032 7700 55504
rect 7660 53983 7700 53992
rect 7756 54956 7796 54965
rect 7756 46388 7796 54916
rect 7756 46339 7796 46348
rect 7852 52604 7892 61795
rect 7948 56720 7988 70624
rect 7948 56671 7988 56680
rect 7852 47060 7892 52564
rect 7852 45800 7892 47020
rect 7852 45751 7892 45760
rect 7948 44960 7988 44969
rect 7852 42188 7892 42197
rect 7756 42020 7796 42029
rect 7660 41768 7700 41777
rect 7563 41600 7605 41609
rect 7563 41560 7564 41600
rect 7604 41560 7605 41600
rect 7563 41551 7605 41560
rect 7660 41012 7700 41728
rect 7660 40963 7700 40972
rect 7468 38779 7508 38788
rect 7468 35720 7508 35729
rect 7372 34292 7412 34301
rect 7372 28328 7412 34252
rect 7468 32696 7508 35680
rect 7756 35300 7796 41980
rect 7852 39920 7892 42148
rect 7852 39871 7892 39880
rect 7851 37736 7893 37745
rect 7851 37696 7852 37736
rect 7892 37696 7893 37736
rect 7851 37687 7893 37696
rect 7468 32647 7508 32656
rect 7660 35260 7796 35300
rect 7852 35888 7892 37687
rect 7948 37148 7988 44920
rect 7948 37099 7988 37108
rect 7564 32108 7604 32117
rect 7564 28664 7604 32068
rect 7372 27992 7412 28288
rect 7372 27943 7412 27952
rect 7468 28624 7604 28664
rect 7276 27616 7412 27656
rect 7180 27532 7316 27572
rect 7179 27404 7221 27413
rect 7179 27364 7180 27404
rect 7220 27364 7221 27404
rect 7179 27355 7221 27364
rect 7180 27270 7220 27355
rect 7276 20180 7316 27532
rect 7372 22364 7412 27616
rect 7468 24884 7508 28624
rect 7563 27488 7605 27497
rect 7563 27448 7564 27488
rect 7604 27448 7605 27488
rect 7563 27439 7605 27448
rect 7564 27354 7604 27439
rect 7468 24835 7508 24844
rect 7372 22315 7412 22324
rect 6988 11320 7124 11360
rect 7180 20140 7316 20180
rect 6604 7748 6644 7757
rect 6604 6320 6644 7708
rect 6604 6271 6644 6280
rect 6508 6019 6548 6028
rect 6124 4808 6164 5692
rect 6124 4759 6164 4768
rect 6795 4808 6837 4817
rect 6795 4768 6796 4808
rect 6836 4768 6837 4808
rect 6795 4759 6837 4768
rect 6796 4674 6836 4759
rect 5932 3499 5972 3508
rect 6988 2624 7028 11320
rect 6988 2036 7028 2584
rect 7180 2540 7220 20140
rect 7372 16064 7412 16073
rect 7276 5228 7316 5237
rect 7276 2801 7316 5188
rect 7275 2792 7317 2801
rect 7275 2752 7276 2792
rect 7316 2752 7317 2792
rect 7275 2743 7317 2752
rect 5739 1868 5781 1877
rect 5739 1828 5740 1868
rect 5780 1828 5781 1868
rect 5739 1819 5781 1828
rect 6795 1112 6837 1121
rect 6795 1072 6796 1112
rect 6836 1072 6837 1112
rect 6795 1063 6837 1072
rect 6796 978 6836 1063
rect 4780 895 4820 904
rect 4928 776 5296 785
rect 4968 736 5010 776
rect 5050 736 5092 776
rect 5132 736 5174 776
rect 5214 736 5256 776
rect 4928 727 5296 736
rect 6988 524 7028 1996
rect 7084 2500 7220 2540
rect 7084 617 7124 2500
rect 7276 1784 7316 2743
rect 7372 1868 7412 16024
rect 7468 15476 7508 15485
rect 7468 3800 7508 15436
rect 7660 4565 7700 35260
rect 7756 34376 7796 34385
rect 7756 32360 7796 34336
rect 7756 31184 7796 32320
rect 7756 31135 7796 31144
rect 7852 30680 7892 35848
rect 7852 30631 7892 30640
rect 7756 30428 7796 30437
rect 7756 27992 7796 30388
rect 7852 29084 7892 29093
rect 7852 29000 7892 29044
rect 7852 28960 7988 29000
rect 7796 27952 7892 27992
rect 7756 27943 7796 27952
rect 7755 26060 7797 26069
rect 7755 26020 7756 26060
rect 7796 26020 7797 26060
rect 7755 26011 7797 26020
rect 7756 25926 7796 26011
rect 7755 23960 7797 23969
rect 7755 23920 7756 23960
rect 7796 23920 7797 23960
rect 7755 23911 7797 23920
rect 7659 4556 7701 4565
rect 7659 4516 7660 4556
rect 7700 4516 7701 4556
rect 7659 4507 7701 4516
rect 7468 3751 7508 3760
rect 7756 3380 7796 23911
rect 7852 21608 7892 27952
rect 7948 26312 7988 28960
rect 7948 25388 7988 26272
rect 7948 25339 7988 25348
rect 7852 21559 7892 21568
rect 7852 16568 7892 16577
rect 7852 5144 7892 16528
rect 7948 8168 7988 8177
rect 7948 6320 7988 8128
rect 7948 6271 7988 6280
rect 7852 5095 7892 5104
rect 7756 3331 7796 3340
rect 7563 2876 7605 2885
rect 7563 2836 7564 2876
rect 7604 2836 7605 2876
rect 7563 2827 7605 2836
rect 7564 2708 7604 2827
rect 7564 2659 7604 2668
rect 8044 2540 8084 79780
rect 8140 64448 8180 82795
rect 8236 79484 8276 79493
rect 8236 78896 8276 79444
rect 8236 78847 8276 78856
rect 8428 78224 8468 78233
rect 8236 76880 8276 76889
rect 8236 73352 8276 76840
rect 8236 73303 8276 73312
rect 8332 76544 8372 76553
rect 8332 66464 8372 76504
rect 8428 76376 8468 78184
rect 8428 76327 8468 76336
rect 8332 65960 8372 66424
rect 8332 65911 8372 65920
rect 8524 65885 8564 84988
rect 12364 84944 12404 84953
rect 11020 84524 11060 84533
rect 9676 84440 9716 84449
rect 8908 83432 8948 83441
rect 8620 79736 8660 79745
rect 8620 73688 8660 79696
rect 8620 70916 8660 73648
rect 8620 70867 8660 70876
rect 8908 66716 8948 83392
rect 9292 83432 9332 83441
rect 9196 74864 9236 74873
rect 8908 66667 8948 66676
rect 9004 70580 9044 70589
rect 8523 65876 8565 65885
rect 8523 65836 8524 65876
rect 8564 65836 8565 65876
rect 8523 65827 8565 65836
rect 8427 64868 8469 64877
rect 8427 64828 8428 64868
rect 8468 64828 8469 64868
rect 8427 64819 8469 64828
rect 8140 64399 8180 64408
rect 8332 63524 8372 63533
rect 8140 60920 8180 60929
rect 8140 58484 8180 60880
rect 8332 58652 8372 63484
rect 8332 58603 8372 58612
rect 8140 58435 8180 58444
rect 8236 57980 8276 57989
rect 8140 57896 8180 57905
rect 8140 54704 8180 57856
rect 8140 54368 8180 54664
rect 8140 54319 8180 54328
rect 8140 45380 8180 45389
rect 8140 22457 8180 45340
rect 8236 44204 8276 57940
rect 8332 54032 8372 54041
rect 8332 51764 8372 53992
rect 8332 47144 8372 51724
rect 8332 47095 8372 47104
rect 8236 44155 8276 44164
rect 8332 44876 8372 44885
rect 8236 40592 8276 40601
rect 8236 39920 8276 40552
rect 8236 39871 8276 39880
rect 8236 33872 8276 33881
rect 8236 33452 8276 33832
rect 8236 33403 8276 33412
rect 8236 25220 8276 25229
rect 8139 22448 8181 22457
rect 8139 22408 8140 22448
rect 8180 22408 8181 22448
rect 8139 22399 8181 22408
rect 8044 2491 8084 2500
rect 7372 1819 7412 1828
rect 7276 1735 7316 1744
rect 8236 860 8276 25180
rect 8332 22868 8372 44836
rect 8428 35384 8468 64819
rect 8524 64280 8564 64289
rect 8524 63524 8564 64240
rect 8524 63475 8564 63484
rect 8524 63188 8564 63197
rect 8524 59240 8564 63148
rect 8524 59191 8564 59200
rect 8620 62600 8660 62609
rect 8524 58652 8564 58661
rect 8524 55292 8564 58612
rect 8524 55243 8564 55252
rect 8523 49748 8565 49757
rect 8523 49708 8524 49748
rect 8564 49708 8565 49748
rect 8523 49699 8565 49708
rect 8524 42692 8564 49699
rect 8524 42643 8564 42652
rect 8524 42188 8564 42197
rect 8524 37745 8564 42148
rect 8523 37736 8565 37745
rect 8523 37696 8524 37736
rect 8564 37696 8565 37736
rect 8523 37687 8565 37696
rect 8620 35888 8660 62560
rect 8716 58484 8756 58493
rect 8716 56636 8756 58444
rect 8716 56587 8756 56596
rect 8716 55712 8756 55721
rect 8716 53528 8756 55672
rect 8716 53479 8756 53488
rect 8715 48068 8757 48077
rect 8715 48028 8716 48068
rect 8756 48028 8757 48068
rect 8715 48019 8757 48028
rect 8716 47934 8756 48019
rect 8716 41768 8756 41777
rect 8716 40760 8756 41728
rect 8908 41600 8948 41609
rect 8908 41096 8948 41560
rect 8908 41047 8948 41056
rect 8716 39752 8756 40720
rect 8716 39703 8756 39712
rect 8812 40928 8852 40937
rect 8812 39416 8852 40888
rect 8908 40256 8948 40265
rect 8908 39584 8948 40216
rect 8908 39535 8948 39544
rect 8812 39367 8852 39376
rect 8620 35839 8660 35848
rect 8716 38744 8756 38753
rect 8428 35335 8468 35344
rect 8620 35300 8660 35309
rect 8524 34040 8564 34049
rect 8428 33704 8468 33713
rect 8428 33536 8468 33664
rect 8428 33487 8468 33496
rect 8524 32780 8564 34000
rect 8620 33032 8660 35260
rect 8620 32983 8660 32992
rect 8524 32731 8564 32740
rect 8716 32612 8756 38704
rect 8812 34628 8852 34637
rect 8812 33368 8852 34588
rect 9004 33536 9044 70540
rect 9100 67724 9140 67733
rect 9100 66716 9140 67684
rect 9100 64280 9140 66676
rect 9100 64231 9140 64240
rect 9196 61004 9236 74824
rect 9196 60955 9236 60964
rect 9100 59240 9140 59249
rect 9100 36560 9140 59200
rect 9196 41012 9236 41021
rect 9196 40676 9236 40972
rect 9196 40627 9236 40636
rect 9100 36511 9140 36520
rect 9196 37316 9236 37325
rect 9100 33536 9140 33545
rect 9004 33496 9100 33536
rect 8812 33319 8852 33328
rect 8524 32572 8756 32612
rect 8524 32276 8564 32572
rect 8332 22819 8372 22828
rect 8428 31268 8468 31277
rect 8332 22700 8372 22709
rect 8332 20852 8372 22660
rect 8332 12032 8372 20812
rect 8332 11983 8372 11992
rect 8428 7328 8468 31228
rect 8524 25388 8564 32236
rect 8716 31268 8756 31277
rect 8524 25220 8564 25348
rect 8524 25171 8564 25180
rect 8620 25808 8660 25817
rect 8620 24632 8660 25768
rect 8716 24716 8756 31228
rect 8908 31184 8948 31193
rect 8716 24667 8756 24676
rect 8812 27740 8852 27749
rect 8620 24583 8660 24592
rect 8812 23969 8852 27700
rect 8811 23960 8853 23969
rect 8811 23920 8812 23960
rect 8852 23920 8853 23960
rect 8811 23911 8853 23920
rect 8811 14552 8853 14561
rect 8811 14512 8812 14552
rect 8852 14512 8853 14552
rect 8811 14503 8853 14512
rect 8620 14468 8660 14477
rect 8428 7279 8468 7288
rect 8524 8084 8564 8093
rect 8524 4220 8564 8044
rect 8620 7916 8660 14428
rect 8812 14418 8852 14503
rect 8811 12620 8853 12629
rect 8811 12580 8812 12620
rect 8852 12580 8853 12620
rect 8811 12571 8853 12580
rect 8620 7867 8660 7876
rect 8812 7244 8852 12571
rect 8812 7195 8852 7204
rect 8908 5732 8948 31144
rect 9004 27404 9044 27413
rect 9004 25808 9044 27364
rect 9004 25759 9044 25768
rect 9003 23708 9045 23717
rect 9003 23668 9004 23708
rect 9044 23668 9045 23708
rect 9003 23659 9045 23668
rect 9004 23574 9044 23659
rect 8908 5683 8948 5692
rect 9004 22112 9044 22121
rect 8524 4171 8564 4180
rect 8716 4640 8756 4649
rect 8332 3884 8372 3893
rect 8332 1112 8372 3844
rect 8332 1063 8372 1072
rect 8428 1952 8468 1961
rect 8236 811 8276 820
rect 7083 608 7125 617
rect 7083 568 7084 608
rect 7124 568 7125 608
rect 7083 559 7125 568
rect 6988 475 7028 484
rect 8428 440 8468 1912
rect 8428 391 8468 400
rect 8716 365 8756 4600
rect 8908 4052 8948 4061
rect 8812 3296 8852 3305
rect 8812 2540 8852 3256
rect 8908 3044 8948 4012
rect 8908 2995 8948 3004
rect 9004 2708 9044 22072
rect 9100 20852 9140 33496
rect 9100 20803 9140 20812
rect 9004 2659 9044 2668
rect 9100 4892 9140 4901
rect 9100 3968 9140 4852
rect 8812 2491 8852 2500
rect 9100 1868 9140 3928
rect 9196 2708 9236 37276
rect 9292 5900 9332 83392
rect 9580 77888 9620 77897
rect 9388 72428 9428 72437
rect 9388 65456 9428 72388
rect 9388 65407 9428 65416
rect 9484 70076 9524 70085
rect 9388 63272 9428 63281
rect 9388 36056 9428 63232
rect 9388 36007 9428 36016
rect 9388 33032 9428 33041
rect 9388 32780 9428 32992
rect 9388 32731 9428 32740
rect 9388 29168 9428 29177
rect 9388 23876 9428 29128
rect 9388 23827 9428 23836
rect 9388 17828 9428 17837
rect 9388 16736 9428 17788
rect 9388 16687 9428 16696
rect 9292 5851 9332 5860
rect 9484 5732 9524 70036
rect 9580 20768 9620 77848
rect 9676 67817 9716 84400
rect 9868 84440 9908 84449
rect 9868 73100 9908 84400
rect 10444 83684 10484 83693
rect 10060 83600 10100 83609
rect 9963 83180 10005 83189
rect 9963 83140 9964 83180
rect 10004 83140 10005 83180
rect 9963 83131 10005 83140
rect 9772 73060 9908 73100
rect 9772 71252 9812 73060
rect 9772 71203 9812 71212
rect 9771 68648 9813 68657
rect 9771 68608 9772 68648
rect 9812 68608 9813 68648
rect 9771 68599 9813 68608
rect 9675 67808 9717 67817
rect 9675 67768 9676 67808
rect 9716 67768 9717 67808
rect 9675 67759 9717 67768
rect 9675 49496 9717 49505
rect 9675 49456 9676 49496
rect 9716 49456 9717 49496
rect 9675 49447 9717 49456
rect 9676 49362 9716 49447
rect 9772 46304 9812 68599
rect 9867 64448 9909 64457
rect 9867 64408 9868 64448
rect 9908 64408 9909 64448
rect 9867 64399 9909 64408
rect 9772 46255 9812 46264
rect 9676 42608 9716 42617
rect 9676 37904 9716 42568
rect 9772 41852 9812 41861
rect 9772 41516 9812 41812
rect 9772 39248 9812 41476
rect 9772 39199 9812 39208
rect 9676 35300 9716 37864
rect 9868 36224 9908 64399
rect 9964 62684 10004 83131
rect 10060 82097 10100 83560
rect 10444 83012 10484 83644
rect 10539 83516 10581 83525
rect 10539 83476 10540 83516
rect 10580 83476 10581 83516
rect 10539 83467 10581 83476
rect 10540 83382 10580 83467
rect 10444 82963 10484 82972
rect 10059 82088 10101 82097
rect 10059 82048 10060 82088
rect 10100 82048 10101 82088
rect 10059 82039 10101 82048
rect 10348 82088 10388 82097
rect 9964 62635 10004 62644
rect 9868 36175 9908 36184
rect 9964 62516 10004 62525
rect 9676 30764 9716 35260
rect 9964 33368 10004 62476
rect 9964 33319 10004 33328
rect 9676 26900 9716 30724
rect 9868 31772 9908 31781
rect 9868 29756 9908 31732
rect 9868 29168 9908 29716
rect 9868 29119 9908 29128
rect 9963 29168 10005 29177
rect 9963 29128 9964 29168
rect 10004 29128 10005 29168
rect 9963 29119 10005 29128
rect 9964 28664 10004 29119
rect 9964 28615 10004 28624
rect 9771 27656 9813 27665
rect 9771 27616 9772 27656
rect 9812 27616 9813 27656
rect 9771 27607 9813 27616
rect 9772 27522 9812 27607
rect 9676 26851 9716 26860
rect 10060 23708 10100 82039
rect 10348 81164 10388 82048
rect 10348 81115 10388 81124
rect 10444 79400 10484 79409
rect 10444 77972 10484 79360
rect 10444 76880 10484 77932
rect 10636 79400 10676 79409
rect 10636 77468 10676 79360
rect 10636 77419 10676 77428
rect 10828 78392 10868 78401
rect 10828 77132 10868 78352
rect 10828 77083 10868 77092
rect 10444 76831 10484 76840
rect 10156 76712 10196 76721
rect 10156 71756 10196 76672
rect 10732 74444 10772 74453
rect 10444 73856 10484 73865
rect 10444 73268 10484 73816
rect 10444 73219 10484 73228
rect 10156 71707 10196 71716
rect 10636 73100 10676 73109
rect 10540 63860 10580 63869
rect 10348 63356 10388 63365
rect 10252 63272 10292 63283
rect 10252 63197 10292 63232
rect 10251 63188 10293 63197
rect 10251 63148 10252 63188
rect 10292 63148 10293 63188
rect 10251 63139 10293 63148
rect 10348 58736 10388 63316
rect 10348 58687 10388 58696
rect 10540 52184 10580 63820
rect 10636 61424 10676 73060
rect 10636 61375 10676 61384
rect 10348 50924 10388 50933
rect 10348 48824 10388 50884
rect 10444 49664 10484 49673
rect 10444 49160 10484 49624
rect 10444 49111 10484 49120
rect 10348 48775 10388 48784
rect 10540 46472 10580 52144
rect 10540 46423 10580 46432
rect 10540 45128 10580 45137
rect 10156 44456 10196 44465
rect 10156 39080 10196 44416
rect 10348 42020 10388 42029
rect 10252 41852 10292 41861
rect 10252 39248 10292 41812
rect 10348 40424 10388 41980
rect 10348 40375 10388 40384
rect 10444 41684 10484 41693
rect 10252 39199 10292 39208
rect 10156 39031 10196 39040
rect 10252 38324 10292 38333
rect 10252 38156 10292 38284
rect 10060 23659 10100 23668
rect 10156 33368 10196 33377
rect 9580 20719 9620 20728
rect 10060 23120 10100 23129
rect 10060 19844 10100 23080
rect 10060 19592 10100 19804
rect 10060 19543 10100 19552
rect 10060 8000 10100 8009
rect 9579 7412 9621 7421
rect 9579 7372 9580 7412
rect 9620 7372 9621 7412
rect 9579 7363 9621 7372
rect 10060 7412 10100 7960
rect 10060 7363 10100 7372
rect 9580 7278 9620 7363
rect 9388 5480 9428 5489
rect 9388 4472 9428 5440
rect 9388 4423 9428 4432
rect 9196 2659 9236 2668
rect 9100 1819 9140 1828
rect 9484 1868 9524 5692
rect 10156 3968 10196 33328
rect 10252 27488 10292 38116
rect 10444 36392 10484 41644
rect 10540 39929 10580 45088
rect 10636 44960 10676 44969
rect 10539 39920 10581 39929
rect 10539 39880 10540 39920
rect 10580 39880 10581 39920
rect 10539 39871 10581 39880
rect 10444 36343 10484 36352
rect 10540 34208 10580 34217
rect 10540 32696 10580 34168
rect 10540 32647 10580 32656
rect 10636 30941 10676 44920
rect 10635 30932 10677 30941
rect 10635 30892 10636 30932
rect 10676 30892 10677 30932
rect 10635 30883 10677 30892
rect 10252 27439 10292 27448
rect 10348 26480 10388 26489
rect 10252 24800 10292 24809
rect 10252 23288 10292 24760
rect 10252 23239 10292 23248
rect 10252 21524 10292 21552
rect 10348 21524 10388 26440
rect 10636 26396 10676 26405
rect 10636 26144 10676 26356
rect 10292 21484 10388 21524
rect 10252 21475 10292 21484
rect 10348 20684 10388 21484
rect 10540 24212 10580 24221
rect 10540 21356 10580 24172
rect 10540 21307 10580 21316
rect 10348 20635 10388 20644
rect 10636 17828 10676 26104
rect 10636 17779 10676 17788
rect 10732 6320 10772 74404
rect 11020 64448 11060 84484
rect 11980 84524 12020 84533
rect 11212 84440 11252 84449
rect 11115 78140 11157 78149
rect 11115 78100 11116 78140
rect 11156 78100 11157 78140
rect 11115 78091 11157 78100
rect 11020 64399 11060 64408
rect 10828 63608 10868 63617
rect 10828 55460 10868 63568
rect 11019 63188 11061 63197
rect 11019 63148 11020 63188
rect 11060 63148 11061 63188
rect 11019 63139 11061 63148
rect 10923 61424 10965 61433
rect 10923 61384 10924 61424
rect 10964 61384 10965 61424
rect 10923 61375 10965 61384
rect 10924 58400 10964 61375
rect 11020 60164 11060 63139
rect 11020 60115 11060 60124
rect 10924 58360 11060 58400
rect 10828 55420 10964 55460
rect 10827 54032 10869 54041
rect 10827 53992 10828 54032
rect 10868 53992 10869 54032
rect 10827 53983 10869 53992
rect 10828 53898 10868 53983
rect 10828 47228 10868 47237
rect 10828 24893 10868 47188
rect 10924 44708 10964 55420
rect 10924 44659 10964 44668
rect 10924 42692 10964 42701
rect 10924 40676 10964 42652
rect 11020 42533 11060 58360
rect 11116 53192 11156 78091
rect 11212 71840 11252 84400
rect 11596 82424 11636 82433
rect 11596 81752 11636 82384
rect 11884 82424 11924 82433
rect 11788 82172 11828 82200
rect 11884 82172 11924 82384
rect 11980 82340 12020 84484
rect 12364 83348 12404 84904
rect 12844 84776 12884 84785
rect 12748 84440 12788 84449
rect 12459 84104 12501 84113
rect 12459 84064 12460 84104
rect 12500 84064 12501 84104
rect 12459 84055 12501 84064
rect 12460 83970 12500 84055
rect 12364 83299 12404 83308
rect 12652 82928 12692 82937
rect 11980 82291 12020 82300
rect 12172 82592 12212 82601
rect 11828 82132 11924 82172
rect 11788 82123 11828 82132
rect 11596 81703 11636 81712
rect 11212 71791 11252 71800
rect 11404 80156 11444 80165
rect 11308 70244 11348 70253
rect 11212 70160 11252 70169
rect 11212 67304 11252 70120
rect 11212 67255 11252 67264
rect 11212 61928 11252 61937
rect 11212 60164 11252 61888
rect 11212 59828 11252 60124
rect 11212 59779 11252 59788
rect 11211 59408 11253 59417
rect 11211 59368 11212 59408
rect 11252 59368 11253 59408
rect 11211 59359 11253 59368
rect 11116 53143 11156 53152
rect 11019 42524 11061 42533
rect 11019 42484 11020 42524
rect 11060 42484 11061 42524
rect 11019 42475 11061 42484
rect 11116 42440 11156 42451
rect 11116 42365 11156 42400
rect 11115 42356 11157 42365
rect 11115 42316 11116 42356
rect 11156 42316 11157 42356
rect 11115 42307 11157 42316
rect 10924 40627 10964 40636
rect 11020 41936 11060 41945
rect 11020 35720 11060 41896
rect 11115 39920 11157 39929
rect 11115 39880 11116 39920
rect 11156 39880 11157 39920
rect 11115 39871 11157 39880
rect 11020 35671 11060 35680
rect 11019 33704 11061 33713
rect 11019 33664 11020 33704
rect 11060 33664 11061 33704
rect 11019 33655 11061 33664
rect 11020 33570 11060 33655
rect 11020 32192 11060 32201
rect 11020 30680 11060 32152
rect 11020 30631 11060 30640
rect 10827 24884 10869 24893
rect 10827 24844 10828 24884
rect 10868 24844 10869 24884
rect 10827 24835 10869 24844
rect 10732 6271 10772 6280
rect 10828 24716 10868 24725
rect 10156 3919 10196 3928
rect 10252 5816 10292 5825
rect 10060 3884 10100 3893
rect 10060 3380 10100 3844
rect 10060 3331 10100 3340
rect 10252 2288 10292 5776
rect 10731 5648 10773 5657
rect 10731 5608 10732 5648
rect 10772 5608 10773 5648
rect 10731 5599 10773 5608
rect 10732 5514 10772 5599
rect 10444 4976 10484 4985
rect 10252 2239 10292 2248
rect 10348 3968 10388 3977
rect 9484 1819 9524 1828
rect 10348 1196 10388 3928
rect 10348 1147 10388 1156
rect 10444 1448 10484 4936
rect 10828 4220 10868 24676
rect 11116 24557 11156 39871
rect 11212 37064 11252 59359
rect 11212 37015 11252 37024
rect 11212 34880 11252 34889
rect 11115 24548 11157 24557
rect 11115 24508 11116 24548
rect 11156 24508 11157 24548
rect 11115 24499 11157 24508
rect 10828 4171 10868 4180
rect 10540 3380 10580 3389
rect 10540 2885 10580 3340
rect 11212 3044 11252 34840
rect 11308 34208 11348 70204
rect 11308 34159 11348 34168
rect 11308 31940 11348 31949
rect 11308 26648 11348 31900
rect 11404 27068 11444 80116
rect 11788 78308 11828 78317
rect 11596 69908 11636 69917
rect 11596 67724 11636 69868
rect 11596 65456 11636 67684
rect 11500 64280 11540 64289
rect 11500 61760 11540 64240
rect 11500 61711 11540 61720
rect 11500 57560 11540 57569
rect 11500 55964 11540 57520
rect 11500 55915 11540 55924
rect 11596 55544 11636 65416
rect 11788 64280 11828 78268
rect 11884 72260 11924 82132
rect 11980 81836 12020 81845
rect 11980 79400 12020 81796
rect 11980 79351 12020 79360
rect 11884 68564 11924 72220
rect 11884 68515 11924 68524
rect 11980 65456 12020 65465
rect 11788 64240 11924 64280
rect 11787 59492 11829 59501
rect 11787 59452 11788 59492
rect 11828 59452 11829 59492
rect 11787 59443 11829 59452
rect 11788 59358 11828 59443
rect 11788 57560 11828 57569
rect 11788 56972 11828 57520
rect 11788 56923 11828 56932
rect 11500 54788 11540 54797
rect 11500 54116 11540 54748
rect 11500 53276 11540 54076
rect 11500 53227 11540 53236
rect 11500 40508 11540 40517
rect 11500 33713 11540 40468
rect 11499 33704 11541 33713
rect 11499 33664 11500 33704
rect 11540 33664 11541 33704
rect 11499 33655 11541 33664
rect 11500 32696 11540 33655
rect 11500 32647 11540 32656
rect 11500 31352 11540 31361
rect 11500 28412 11540 31312
rect 11500 27488 11540 28372
rect 11500 27439 11540 27448
rect 11404 27019 11444 27028
rect 11500 27152 11540 27161
rect 11308 26599 11348 26608
rect 11500 26564 11540 27112
rect 11500 26515 11540 26524
rect 11596 24044 11636 55504
rect 11692 52268 11732 52277
rect 11692 50672 11732 52228
rect 11692 50623 11732 50632
rect 11884 46640 11924 64240
rect 11980 61760 12020 65416
rect 11980 61711 12020 61720
rect 12076 60080 12116 60089
rect 11788 46600 11924 46640
rect 11980 59744 12020 59753
rect 11212 2995 11252 3004
rect 11308 24004 11636 24044
rect 11692 24632 11732 24641
rect 10539 2876 10581 2885
rect 10539 2836 10540 2876
rect 10580 2836 10581 2876
rect 10539 2827 10581 2836
rect 11019 1868 11061 1877
rect 11019 1828 11020 1868
rect 11060 1828 11061 1868
rect 11019 1819 11061 1828
rect 10444 776 10484 1408
rect 10444 727 10484 736
rect 6987 356 7029 365
rect 6987 316 6988 356
rect 7028 316 7029 356
rect 6987 307 7029 316
rect 8715 356 8757 365
rect 8715 316 8716 356
rect 8756 316 8757 356
rect 8715 307 8757 316
rect 3532 223 3572 232
rect 6988 222 7028 307
rect 11020 272 11060 1819
rect 11308 1121 11348 24004
rect 11692 23540 11732 24592
rect 11692 23491 11732 23500
rect 11500 16064 11540 16073
rect 11500 3380 11540 16024
rect 11692 5984 11732 5993
rect 11692 3716 11732 5944
rect 11692 3667 11732 3676
rect 11500 3331 11540 3340
rect 11596 2708 11636 2717
rect 11596 2204 11636 2668
rect 11596 2155 11636 2164
rect 11307 1112 11349 1121
rect 11307 1072 11308 1112
rect 11348 1072 11349 1112
rect 11307 1063 11349 1072
rect 11788 944 11828 46600
rect 11788 895 11828 904
rect 11884 46472 11924 46481
rect 11884 692 11924 46432
rect 11980 45380 12020 59704
rect 11980 45331 12020 45340
rect 12076 29000 12116 60040
rect 11980 28960 12116 29000
rect 11980 22709 12020 28960
rect 11979 22700 12021 22709
rect 11979 22660 11980 22700
rect 12020 22660 12021 22700
rect 11979 22651 12021 22660
rect 12075 15056 12117 15065
rect 12075 15016 12076 15056
rect 12116 15016 12117 15056
rect 12075 15007 12117 15016
rect 12076 14922 12116 15007
rect 12076 9512 12116 9521
rect 12076 8672 12116 9472
rect 12076 8000 12116 8632
rect 12076 7160 12116 7960
rect 12172 7580 12212 82552
rect 12652 81920 12692 82888
rect 12652 81871 12692 81880
rect 12556 79316 12596 79325
rect 12556 75200 12596 79276
rect 12556 75151 12596 75160
rect 12460 73184 12500 73193
rect 12363 63692 12405 63701
rect 12363 63652 12364 63692
rect 12404 63652 12405 63692
rect 12363 63643 12405 63652
rect 12268 59072 12308 59081
rect 12268 44969 12308 59032
rect 12364 58316 12404 63643
rect 12460 59912 12500 73144
rect 12556 71840 12596 71849
rect 12556 70664 12596 71800
rect 12556 70615 12596 70624
rect 12460 59863 12500 59872
rect 12556 64868 12596 64877
rect 12364 58276 12500 58316
rect 12364 58148 12404 58157
rect 12364 56720 12404 58108
rect 12364 56671 12404 56680
rect 12460 55460 12500 58276
rect 12364 55420 12500 55460
rect 12267 44960 12309 44969
rect 12267 44920 12268 44960
rect 12308 44920 12309 44960
rect 12267 44911 12309 44920
rect 12364 43280 12404 55420
rect 12459 54620 12501 54629
rect 12459 54580 12460 54620
rect 12500 54580 12501 54620
rect 12459 54571 12501 54580
rect 12460 53192 12500 54571
rect 12460 53143 12500 53152
rect 12556 45548 12596 64828
rect 12652 59912 12692 59921
rect 12652 55628 12692 59872
rect 12652 54629 12692 55588
rect 12651 54620 12693 54629
rect 12651 54580 12652 54620
rect 12692 54580 12693 54620
rect 12651 54571 12693 54580
rect 12748 53528 12788 84400
rect 12748 53024 12788 53488
rect 12748 52975 12788 52984
rect 12556 45499 12596 45508
rect 12364 43231 12404 43240
rect 12460 44204 12500 44213
rect 12364 34376 12404 34385
rect 12268 27908 12308 27917
rect 12268 26144 12308 27868
rect 12364 27068 12404 34336
rect 12364 27019 12404 27028
rect 12268 26095 12308 26104
rect 12363 25220 12405 25229
rect 12363 25180 12364 25220
rect 12404 25180 12405 25220
rect 12363 25171 12405 25180
rect 12172 7531 12212 7540
rect 12268 25052 12308 25061
rect 12076 7111 12116 7120
rect 12268 5900 12308 25012
rect 12268 5851 12308 5860
rect 12364 3380 12404 25171
rect 12460 24641 12500 44164
rect 12652 41096 12692 41105
rect 12556 39332 12596 39341
rect 12556 38408 12596 39292
rect 12556 38359 12596 38368
rect 12652 38324 12692 41056
rect 12652 38275 12692 38284
rect 12748 36644 12788 36653
rect 12748 35132 12788 36604
rect 12748 35083 12788 35092
rect 12748 29840 12788 29849
rect 12748 28328 12788 29800
rect 12748 28279 12788 28288
rect 12556 27908 12596 27917
rect 12556 27320 12596 27868
rect 12556 27271 12596 27280
rect 12556 26816 12596 26825
rect 12459 24632 12501 24641
rect 12459 24592 12460 24632
rect 12500 24592 12501 24632
rect 12459 24583 12501 24592
rect 12556 22700 12596 26776
rect 12556 22651 12596 22660
rect 12652 25304 12692 25313
rect 12652 20348 12692 25264
rect 12652 20299 12692 20308
rect 12460 17660 12500 17669
rect 12460 9848 12500 17620
rect 12460 9799 12500 9808
rect 12844 8672 12884 84736
rect 18808 84692 19176 84701
rect 18848 84652 18890 84692
rect 18930 84652 18972 84692
rect 19012 84652 19054 84692
rect 19094 84652 19136 84692
rect 18808 84643 19176 84652
rect 13900 84440 13940 84449
rect 13228 84104 13268 84113
rect 12940 82592 12980 82601
rect 12940 20273 12980 82552
rect 13132 82592 13172 82601
rect 13036 78560 13076 78569
rect 12939 20264 12981 20273
rect 12939 20224 12940 20264
rect 12980 20224 12981 20264
rect 12939 20215 12981 20224
rect 12844 8623 12884 8632
rect 12940 20012 12980 20021
rect 12940 11612 12980 19972
rect 12364 3331 12404 3340
rect 12652 7580 12692 7589
rect 11884 643 11924 652
rect 11020 223 11060 232
rect 12652 197 12692 7540
rect 12940 5228 12980 11572
rect 12940 5179 12980 5188
rect 13036 4640 13076 78520
rect 13036 4591 13076 4600
rect 13035 1868 13077 1877
rect 13035 1828 13036 1868
rect 13076 1828 13077 1868
rect 13035 1819 13077 1828
rect 12747 1280 12789 1289
rect 12747 1240 12748 1280
rect 12788 1240 12789 1280
rect 12747 1231 12789 1240
rect 12748 1146 12788 1231
rect 13036 1196 13076 1819
rect 13132 1280 13172 82552
rect 13228 71840 13268 84064
rect 13611 83348 13653 83357
rect 13611 83308 13612 83348
rect 13652 83308 13653 83348
rect 13611 83299 13653 83308
rect 13612 83214 13652 83299
rect 13804 83012 13844 83021
rect 13228 71791 13268 71800
rect 13324 77636 13364 77645
rect 13324 71504 13364 77596
rect 13420 75620 13460 75629
rect 13420 71672 13460 75580
rect 13516 73184 13556 73193
rect 13516 72848 13556 73144
rect 13516 72799 13556 72808
rect 13420 71623 13460 71632
rect 13804 71756 13844 82972
rect 13324 71455 13364 71464
rect 13228 71168 13268 71177
rect 13228 65204 13268 71128
rect 13804 71168 13844 71716
rect 13804 71119 13844 71128
rect 13612 69320 13652 69329
rect 13228 65155 13268 65164
rect 13516 67976 13556 67985
rect 13228 64448 13268 64457
rect 13228 61256 13268 64408
rect 13228 61207 13268 61216
rect 13324 60500 13364 60509
rect 13228 60332 13268 60341
rect 13228 54041 13268 60292
rect 13227 54032 13269 54041
rect 13227 53992 13228 54032
rect 13268 53992 13269 54032
rect 13227 53983 13269 53992
rect 13228 53276 13268 53983
rect 13228 53227 13268 53236
rect 13228 52856 13268 52865
rect 13228 48824 13268 52816
rect 13228 48775 13268 48784
rect 13228 40592 13268 40601
rect 13228 38828 13268 40552
rect 13228 38779 13268 38788
rect 13227 28916 13269 28925
rect 13227 28876 13228 28916
rect 13268 28876 13269 28916
rect 13227 28867 13269 28876
rect 13228 27740 13268 28867
rect 13228 27691 13268 27700
rect 13227 20096 13269 20105
rect 13227 20056 13228 20096
rect 13268 20056 13269 20096
rect 13227 20047 13269 20056
rect 13228 17912 13268 20047
rect 13228 17863 13268 17872
rect 13132 1231 13172 1240
rect 13036 1147 13076 1156
rect 13324 944 13364 60460
rect 13420 55712 13460 55721
rect 13420 55460 13460 55672
rect 13420 55411 13460 55420
rect 13420 51764 13460 51773
rect 13420 46892 13460 51724
rect 13420 46843 13460 46852
rect 13516 40676 13556 67936
rect 13516 40627 13556 40636
rect 13420 38324 13460 38333
rect 13420 34376 13460 38284
rect 13420 34327 13460 34336
rect 13516 31016 13556 31025
rect 13516 30008 13556 30976
rect 13516 29959 13556 29968
rect 13515 29672 13557 29681
rect 13515 29632 13516 29672
rect 13556 29632 13557 29672
rect 13515 29623 13557 29632
rect 13516 29000 13556 29623
rect 13516 28951 13556 28960
rect 13612 19256 13652 69280
rect 13804 68732 13844 68741
rect 13708 56804 13748 56813
rect 13708 55292 13748 56764
rect 13708 55243 13748 55252
rect 13707 55124 13749 55133
rect 13707 55084 13708 55124
rect 13748 55084 13749 55124
rect 13707 55075 13749 55084
rect 13708 49244 13748 55075
rect 13708 49195 13748 49204
rect 13804 44540 13844 68692
rect 13804 44491 13844 44500
rect 13708 41936 13748 41945
rect 13708 39332 13748 41896
rect 13708 39283 13748 39292
rect 13612 19207 13652 19216
rect 13708 33032 13748 33041
rect 13324 895 13364 904
rect 13708 776 13748 32992
rect 13804 29336 13844 29345
rect 13804 28916 13844 29296
rect 13804 28867 13844 28876
rect 13900 21272 13940 84400
rect 16876 84440 16916 84449
rect 16588 84272 16628 84281
rect 14956 83348 14996 83357
rect 13996 83180 14036 83189
rect 13996 67976 14036 83140
rect 14380 82760 14420 82769
rect 14380 81920 14420 82720
rect 14380 81871 14420 81880
rect 14764 82592 14804 82601
rect 14764 81752 14804 82552
rect 14764 81703 14804 81712
rect 14860 80660 14900 80669
rect 14284 80492 14324 80501
rect 14284 78560 14324 80452
rect 14284 78511 14324 78520
rect 13996 67927 14036 67936
rect 14284 74024 14324 74033
rect 14188 66464 14228 66473
rect 14092 58904 14132 58913
rect 13996 57392 14036 57401
rect 13996 56132 14036 57352
rect 13996 56083 14036 56092
rect 14092 55880 14132 58864
rect 13996 55840 14132 55880
rect 13996 55133 14036 55840
rect 14092 55544 14132 55553
rect 13995 55124 14037 55133
rect 13995 55084 13996 55124
rect 14036 55084 14037 55124
rect 13995 55075 14037 55084
rect 14092 55124 14132 55504
rect 14092 55075 14132 55084
rect 14092 54956 14132 54965
rect 13900 21223 13940 21232
rect 13996 54200 14036 54209
rect 13900 17072 13940 17081
rect 13900 4136 13940 17032
rect 13900 2204 13940 4096
rect 13900 2155 13940 2164
rect 13996 944 14036 54160
rect 14092 53192 14132 54916
rect 14092 53143 14132 53152
rect 14188 42860 14228 66424
rect 14284 64793 14324 73984
rect 14572 71504 14612 71513
rect 14380 71084 14420 71093
rect 14283 64784 14325 64793
rect 14283 64744 14284 64784
rect 14324 64744 14325 64784
rect 14283 64735 14325 64744
rect 14284 63776 14324 63785
rect 14284 63197 14324 63736
rect 14283 63188 14325 63197
rect 14283 63148 14284 63188
rect 14324 63148 14325 63188
rect 14283 63139 14325 63148
rect 14284 55460 14324 63139
rect 14380 59240 14420 71044
rect 14572 70160 14612 71464
rect 14572 70111 14612 70120
rect 14572 69824 14612 69833
rect 14475 69068 14517 69077
rect 14475 69028 14476 69068
rect 14516 69028 14517 69068
rect 14475 69019 14517 69028
rect 14476 65120 14516 69019
rect 14476 65071 14516 65080
rect 14572 65036 14612 69784
rect 14860 69077 14900 80620
rect 14859 69068 14901 69077
rect 14859 69028 14860 69068
rect 14900 69028 14901 69068
rect 14859 69019 14901 69028
rect 14956 68993 14996 83308
rect 16012 83348 16052 83357
rect 16012 83189 16052 83308
rect 16011 83180 16053 83189
rect 16011 83140 16012 83180
rect 16052 83140 16053 83180
rect 16011 83131 16053 83140
rect 16396 81836 16436 81845
rect 16396 81089 16436 81796
rect 16395 81080 16437 81089
rect 16395 81040 16396 81080
rect 16436 81040 16437 81080
rect 16395 81031 16437 81040
rect 16012 80996 16052 81005
rect 15820 80324 15860 80333
rect 15724 78224 15764 78233
rect 15532 78140 15572 78149
rect 15051 77300 15093 77309
rect 15051 77260 15052 77300
rect 15092 77260 15093 77300
rect 15051 77251 15093 77260
rect 15052 77166 15092 77251
rect 15532 76040 15572 78100
rect 15436 74612 15476 74621
rect 15148 70832 15188 70841
rect 15052 70580 15092 70589
rect 14763 68984 14805 68993
rect 14763 68944 14764 68984
rect 14804 68944 14805 68984
rect 14763 68935 14805 68944
rect 14955 68984 14997 68993
rect 14955 68944 14956 68984
rect 14996 68944 14997 68984
rect 14955 68935 14997 68944
rect 14572 64996 14708 65036
rect 14571 64784 14613 64793
rect 14571 64744 14572 64784
rect 14612 64744 14613 64784
rect 14571 64735 14613 64744
rect 14572 62600 14612 64735
rect 14572 62551 14612 62560
rect 14668 59408 14708 64996
rect 14668 59359 14708 59368
rect 14380 59200 14708 59240
rect 14572 56132 14612 56141
rect 14284 55420 14420 55460
rect 14284 53696 14324 53705
rect 14284 53285 14324 53656
rect 14283 53276 14325 53285
rect 14283 53236 14284 53276
rect 14324 53236 14325 53276
rect 14283 53227 14325 53236
rect 14284 53142 14324 53227
rect 14188 42811 14228 42820
rect 13996 895 14036 904
rect 14092 40340 14132 40349
rect 14092 860 14132 40300
rect 14284 40340 14324 40349
rect 14188 39920 14228 39929
rect 14188 39164 14228 39880
rect 14188 39115 14228 39124
rect 14284 37820 14324 40300
rect 14188 37780 14324 37820
rect 14188 31436 14228 37780
rect 14188 31387 14228 31396
rect 14380 30260 14420 55420
rect 14476 54872 14516 54881
rect 14476 49244 14516 54832
rect 14476 49195 14516 49204
rect 14380 30211 14420 30220
rect 14476 33956 14516 33965
rect 14187 29672 14229 29681
rect 14187 29632 14188 29672
rect 14228 29632 14229 29672
rect 14187 29623 14229 29632
rect 14188 29538 14228 29623
rect 14284 29336 14324 29345
rect 14284 29084 14324 29296
rect 14284 29035 14324 29044
rect 14476 29084 14516 33916
rect 14572 31520 14612 56092
rect 14668 54788 14708 59200
rect 14764 56636 14804 68935
rect 14956 64952 14996 64961
rect 14860 61172 14900 61181
rect 14860 60416 14900 61132
rect 14860 60367 14900 60376
rect 14764 56587 14804 56596
rect 14860 59240 14900 59249
rect 14860 56561 14900 59200
rect 14859 56552 14901 56561
rect 14859 56512 14860 56552
rect 14900 56512 14901 56552
rect 14859 56503 14901 56512
rect 14668 54739 14708 54748
rect 14764 56216 14804 56225
rect 14667 49496 14709 49505
rect 14667 49456 14668 49496
rect 14708 49456 14709 49496
rect 14667 49447 14709 49456
rect 14668 48992 14708 49447
rect 14668 48943 14708 48952
rect 14764 48152 14804 56176
rect 14956 55460 14996 64912
rect 15052 56729 15092 70540
rect 15051 56720 15093 56729
rect 15051 56680 15052 56720
rect 15092 56680 15093 56720
rect 15051 56671 15093 56680
rect 15051 56552 15093 56561
rect 15051 56512 15052 56552
rect 15092 56512 15093 56552
rect 15051 56503 15093 56512
rect 14668 48112 14804 48152
rect 14860 55420 14996 55460
rect 14668 32780 14708 48112
rect 14763 47984 14805 47993
rect 14763 47944 14764 47984
rect 14804 47944 14805 47984
rect 14763 47935 14805 47944
rect 14764 34964 14804 47935
rect 14860 41012 14900 55420
rect 14956 53528 14996 53537
rect 14956 47993 14996 53488
rect 15052 53024 15092 56503
rect 15052 52975 15092 52984
rect 15052 51344 15092 51353
rect 14955 47984 14997 47993
rect 14955 47944 14956 47984
rect 14996 47944 14997 47984
rect 14955 47935 14997 47944
rect 15052 44204 15092 51304
rect 15052 44155 15092 44164
rect 15148 42608 15188 70792
rect 15340 62348 15380 62357
rect 15340 57728 15380 62308
rect 15340 57679 15380 57688
rect 15148 42559 15188 42568
rect 15340 55292 15380 55301
rect 15340 54788 15380 55252
rect 14860 40963 14900 40972
rect 15052 41432 15092 41441
rect 15052 40340 15092 41392
rect 15052 40291 15092 40300
rect 14764 34915 14804 34924
rect 14668 32731 14708 32740
rect 15244 33032 15284 33041
rect 15148 32360 15188 32369
rect 14572 31471 14612 31480
rect 15052 32192 15092 32201
rect 14668 31436 14708 31445
rect 14380 27908 14420 27917
rect 14284 27068 14324 27077
rect 14188 23288 14228 23297
rect 14188 21440 14228 23248
rect 14284 21608 14324 27028
rect 14380 24128 14420 27868
rect 14476 27665 14516 29044
rect 14572 30512 14612 30521
rect 14475 27656 14517 27665
rect 14475 27616 14476 27656
rect 14516 27616 14517 27656
rect 14475 27607 14517 27616
rect 14476 27521 14516 27607
rect 14380 24079 14420 24088
rect 14476 24968 14516 24977
rect 14284 21559 14324 21568
rect 14380 23876 14420 23885
rect 14188 21391 14228 21400
rect 14188 21104 14228 21113
rect 14188 2708 14228 21064
rect 14380 19088 14420 23836
rect 14476 22616 14516 24928
rect 14572 23708 14612 30472
rect 14572 23659 14612 23668
rect 14668 30344 14708 31396
rect 14476 22576 14612 22616
rect 14380 19039 14420 19048
rect 14476 21608 14516 21617
rect 14476 10268 14516 21568
rect 14476 10219 14516 10228
rect 14284 8168 14324 8177
rect 14284 5648 14324 8128
rect 14284 5599 14324 5608
rect 14188 2659 14228 2668
rect 14572 2708 14612 22576
rect 14668 21356 14708 30304
rect 14956 29336 14996 29345
rect 14956 29000 14996 29296
rect 14956 28951 14996 28960
rect 14859 28916 14901 28925
rect 14859 28876 14860 28916
rect 14900 28876 14901 28916
rect 14859 28867 14901 28876
rect 14860 28782 14900 28867
rect 14764 28748 14804 28757
rect 14764 28160 14804 28708
rect 14764 28111 14804 28120
rect 14860 28328 14900 28337
rect 14860 27740 14900 28288
rect 14860 27691 14900 27700
rect 15052 27152 15092 32152
rect 15148 30680 15188 32320
rect 15148 27236 15188 30640
rect 15244 31688 15284 32992
rect 15244 27572 15284 31648
rect 15244 27523 15284 27532
rect 15148 27187 15188 27196
rect 15052 27103 15092 27112
rect 14860 26900 14900 26909
rect 14764 26396 14804 26405
rect 14764 23717 14804 26356
rect 14763 23708 14805 23717
rect 14763 23668 14764 23708
rect 14804 23668 14805 23708
rect 14763 23659 14805 23668
rect 14764 22448 14804 23659
rect 14764 22399 14804 22408
rect 14668 21307 14708 21316
rect 14764 19592 14804 19601
rect 14764 18752 14804 19552
rect 14764 18703 14804 18712
rect 14860 18584 14900 26860
rect 14956 26144 14996 26153
rect 14956 22784 14996 26104
rect 14956 22735 14996 22744
rect 15052 22868 15092 22877
rect 15052 21785 15092 22828
rect 15051 21776 15093 21785
rect 15051 21736 15052 21776
rect 15092 21736 15093 21776
rect 15051 21727 15093 21736
rect 15148 20264 15188 20273
rect 15148 20096 15188 20224
rect 15148 20047 15188 20056
rect 15340 20012 15380 54748
rect 15340 19963 15380 19972
rect 15436 20768 15476 74572
rect 15532 70580 15572 76000
rect 15724 75200 15764 78184
rect 15724 75151 15764 75160
rect 15532 70531 15572 70540
rect 15532 65456 15572 65465
rect 15532 42188 15572 65416
rect 15724 64700 15764 64709
rect 15628 61508 15668 61517
rect 15628 58568 15668 61468
rect 15724 60080 15764 64660
rect 15820 64280 15860 80284
rect 15820 64231 15860 64240
rect 15916 67640 15956 67649
rect 15916 60248 15956 67600
rect 15916 60199 15956 60208
rect 15724 60040 15956 60080
rect 15820 59912 15860 59921
rect 15724 58568 15764 58577
rect 15628 58528 15724 58568
rect 15724 56552 15764 58528
rect 15724 56503 15764 56512
rect 15628 52856 15668 52865
rect 15628 49748 15668 52816
rect 15628 49699 15668 49708
rect 15724 52100 15764 52109
rect 15724 48992 15764 52060
rect 15724 48943 15764 48952
rect 15724 48740 15764 48749
rect 15724 46472 15764 48700
rect 15724 46423 15764 46432
rect 15532 42139 15572 42148
rect 15724 37148 15764 37157
rect 15628 34880 15668 34889
rect 15532 32780 15572 32789
rect 15532 21692 15572 32740
rect 15628 28328 15668 34840
rect 15628 28279 15668 28288
rect 15532 21643 15572 21652
rect 15628 26480 15668 26489
rect 15628 21440 15668 26440
rect 14860 18535 14900 18544
rect 15340 15812 15380 15821
rect 15148 15560 15188 15569
rect 14668 14468 14708 14477
rect 14668 13880 14708 14428
rect 14668 13831 14708 13840
rect 15052 12536 15092 12545
rect 14956 11864 14996 11873
rect 14956 10016 14996 11824
rect 14956 9967 14996 9976
rect 14956 8252 14996 8261
rect 14956 5648 14996 8212
rect 15052 7076 15092 12496
rect 15148 7580 15188 15520
rect 15244 15056 15284 15065
rect 15244 13292 15284 15016
rect 15340 13544 15380 15772
rect 15340 13495 15380 13504
rect 15244 13243 15284 13252
rect 15436 8924 15476 20728
rect 15532 21400 15668 21440
rect 15532 19424 15572 21400
rect 15532 19375 15572 19384
rect 15628 21272 15668 21281
rect 15532 16232 15572 16241
rect 15532 13460 15572 16192
rect 15628 13880 15668 21232
rect 15724 19004 15764 37108
rect 15820 27488 15860 59872
rect 15916 45212 15956 60040
rect 16012 55292 16052 80956
rect 16396 80946 16436 81031
rect 16300 76544 16340 76553
rect 16204 74108 16244 74117
rect 16204 71420 16244 74068
rect 16204 71371 16244 71380
rect 16012 55243 16052 55252
rect 16108 69740 16148 69749
rect 15916 45163 15956 45172
rect 16012 55124 16052 55133
rect 15820 27439 15860 27448
rect 15916 27404 15956 27413
rect 15724 18955 15764 18964
rect 15820 26816 15860 26825
rect 15724 17240 15764 17249
rect 15724 14216 15764 17200
rect 15724 14167 15764 14176
rect 15628 13831 15668 13840
rect 15532 13411 15572 13420
rect 15820 11024 15860 26776
rect 15916 18920 15956 27364
rect 15916 18871 15956 18880
rect 15916 16148 15956 16157
rect 15916 14636 15956 16108
rect 15916 14587 15956 14596
rect 15436 8875 15476 8884
rect 15628 10772 15668 10781
rect 15436 8756 15476 8765
rect 15244 8252 15284 8261
rect 15244 7916 15284 8212
rect 15244 7867 15284 7876
rect 15148 7531 15188 7540
rect 15052 7027 15092 7036
rect 15052 5648 15092 5657
rect 14956 5608 15052 5648
rect 15052 3128 15092 5608
rect 15052 3079 15092 3088
rect 14572 2659 14612 2668
rect 15436 1700 15476 8716
rect 15532 8588 15572 8597
rect 15532 7664 15572 8548
rect 15532 7615 15572 7624
rect 15628 5228 15668 10732
rect 15820 10100 15860 10984
rect 15820 6824 15860 10060
rect 15820 6775 15860 6784
rect 15628 5179 15668 5188
rect 16012 1868 16052 55084
rect 16108 54200 16148 69700
rect 16108 54151 16148 54160
rect 16204 67052 16244 67061
rect 16108 52268 16148 52277
rect 16108 45044 16148 52228
rect 16108 44995 16148 45004
rect 16108 40928 16148 40937
rect 16108 40088 16148 40888
rect 16108 40039 16148 40048
rect 16204 37316 16244 67012
rect 16300 47732 16340 76504
rect 16588 65288 16628 84232
rect 16780 71168 16820 71177
rect 16683 66968 16725 66977
rect 16683 66928 16684 66968
rect 16724 66928 16725 66968
rect 16683 66919 16725 66928
rect 16684 66834 16724 66919
rect 16588 65239 16628 65248
rect 16396 64364 16436 64373
rect 16396 55208 16436 64324
rect 16396 54788 16436 55168
rect 16396 54739 16436 54748
rect 16492 57980 16532 57989
rect 16300 47683 16340 47692
rect 16396 53612 16436 53621
rect 16396 46640 16436 53572
rect 16492 52100 16532 57940
rect 16588 54704 16628 54713
rect 16588 52352 16628 54664
rect 16588 52303 16628 52312
rect 16492 52051 16532 52060
rect 16588 51932 16628 51941
rect 16588 48824 16628 51892
rect 16588 47312 16628 48784
rect 16588 47263 16628 47272
rect 16396 46600 16532 46640
rect 16396 41600 16436 41609
rect 16204 37267 16244 37276
rect 16300 38828 16340 38837
rect 16300 28244 16340 38788
rect 16300 27740 16340 28204
rect 16300 27691 16340 27700
rect 16108 26480 16148 26489
rect 16108 20936 16148 26440
rect 16204 25976 16244 25985
rect 16204 24968 16244 25936
rect 16204 24919 16244 24928
rect 16300 25556 16340 25565
rect 16300 24632 16340 25516
rect 16396 24884 16436 41560
rect 16396 24835 16436 24844
rect 16492 26060 16532 46600
rect 16588 42776 16628 42785
rect 16588 33704 16628 42736
rect 16780 42608 16820 71128
rect 16876 62600 16916 84400
rect 18028 84356 18068 84365
rect 17740 84104 17780 84113
rect 16972 83516 17012 83525
rect 16972 63020 17012 83476
rect 17452 83180 17492 83189
rect 17068 80912 17108 80921
rect 17068 79652 17108 80872
rect 17068 79603 17108 79612
rect 17164 79820 17204 79829
rect 17068 78728 17108 78737
rect 17068 77552 17108 78688
rect 17068 77503 17108 77512
rect 17164 77468 17204 79780
rect 17356 79232 17396 79241
rect 17164 77419 17204 77428
rect 17260 78896 17300 78905
rect 17260 75284 17300 78856
rect 17356 77720 17396 79192
rect 17356 77671 17396 77680
rect 17452 76880 17492 83140
rect 17452 76831 17492 76840
rect 17644 79400 17684 79409
rect 17260 75235 17300 75244
rect 17452 72008 17492 72017
rect 17356 67388 17396 67397
rect 16972 62971 17012 62980
rect 17068 66044 17108 66053
rect 16876 62551 16916 62560
rect 16972 56300 17012 56309
rect 16972 55544 17012 56260
rect 16972 54032 17012 55504
rect 16972 53983 17012 53992
rect 16780 42559 16820 42568
rect 16972 51764 17012 51773
rect 16588 33655 16628 33664
rect 16684 36560 16724 36569
rect 16684 28496 16724 36520
rect 16876 35216 16916 35225
rect 16876 34796 16916 35176
rect 16876 34747 16916 34756
rect 16588 28456 16724 28496
rect 16780 34292 16820 34301
rect 16780 34040 16820 34252
rect 16588 27572 16628 28456
rect 16588 27523 16628 27532
rect 16684 28328 16724 28337
rect 16684 26648 16724 28288
rect 16684 26599 16724 26608
rect 16300 24583 16340 24592
rect 16492 23465 16532 26020
rect 16588 26480 16628 26489
rect 16491 23456 16533 23465
rect 16491 23416 16492 23456
rect 16532 23416 16533 23456
rect 16491 23407 16533 23416
rect 16492 23036 16532 23045
rect 16395 22700 16437 22709
rect 16395 22660 16396 22700
rect 16436 22660 16437 22700
rect 16395 22651 16437 22660
rect 16396 21104 16436 22651
rect 16396 21055 16436 21064
rect 16108 20887 16148 20896
rect 16300 19508 16340 19517
rect 16108 15644 16148 15653
rect 16108 15308 16148 15604
rect 16108 15259 16148 15268
rect 16107 15056 16149 15065
rect 16107 15016 16108 15056
rect 16148 15016 16149 15056
rect 16107 15007 16149 15016
rect 16108 14922 16148 15007
rect 16012 1819 16052 1828
rect 16108 13208 16148 13217
rect 16108 12620 16148 13168
rect 16108 10940 16148 12580
rect 16108 10268 16148 10900
rect 15436 1651 15476 1660
rect 14092 811 14132 820
rect 13708 727 13748 736
rect 15627 776 15669 785
rect 15627 736 15628 776
rect 15668 736 15669 776
rect 15627 727 15669 736
rect 15628 642 15668 727
rect 12651 188 12693 197
rect 12651 148 12652 188
rect 12692 148 12693 188
rect 12651 139 12693 148
rect 16108 188 16148 10228
rect 16300 12536 16340 19468
rect 16492 17156 16532 22996
rect 16588 20180 16628 26440
rect 16684 24380 16724 24389
rect 16684 22868 16724 24340
rect 16780 24212 16820 34000
rect 16875 30932 16917 30941
rect 16875 30892 16876 30932
rect 16916 30892 16917 30932
rect 16875 30883 16917 30892
rect 16780 24163 16820 24172
rect 16684 22819 16724 22828
rect 16588 20131 16628 20140
rect 16684 20684 16724 20693
rect 16684 19928 16724 20644
rect 16684 19879 16724 19888
rect 16492 17107 16532 17116
rect 16588 18920 16628 18929
rect 16204 9932 16244 9941
rect 16204 3632 16244 9892
rect 16300 6488 16340 12496
rect 16396 16736 16436 16745
rect 16396 11276 16436 16696
rect 16396 11227 16436 11236
rect 16300 6439 16340 6448
rect 16204 3583 16244 3592
rect 16588 3380 16628 18880
rect 16876 18752 16916 30883
rect 16876 18703 16916 18712
rect 16780 13292 16820 13301
rect 16780 11024 16820 13252
rect 16780 10975 16820 10984
rect 16588 3331 16628 3340
rect 16780 4136 16820 4145
rect 16780 776 16820 4096
rect 16972 3380 17012 51724
rect 17068 37148 17108 66004
rect 17164 65204 17204 65213
rect 17164 45296 17204 65164
rect 17164 45247 17204 45256
rect 17260 64196 17300 64205
rect 17260 42356 17300 64156
rect 17356 44120 17396 67348
rect 17356 44071 17396 44080
rect 17260 42307 17300 42316
rect 17068 37099 17108 37108
rect 17164 41768 17204 41777
rect 17068 36056 17108 36065
rect 17068 26816 17108 36016
rect 17164 34040 17204 41728
rect 17452 35888 17492 71968
rect 17644 71336 17684 79360
rect 17644 71287 17684 71296
rect 17644 69236 17684 69245
rect 17548 63944 17588 63953
rect 17548 53780 17588 63904
rect 17644 61844 17684 69196
rect 17644 61795 17684 61804
rect 17644 57980 17684 57989
rect 17644 55628 17684 57940
rect 17644 55579 17684 55588
rect 17548 53731 17588 53740
rect 17740 52940 17780 84064
rect 17932 80576 17972 80585
rect 17932 76964 17972 80536
rect 18028 78308 18068 84316
rect 19660 84356 19700 84365
rect 18412 83180 18452 83189
rect 18028 78149 18068 78268
rect 18220 79652 18260 79661
rect 18027 78140 18069 78149
rect 18027 78100 18028 78140
rect 18068 78100 18069 78140
rect 18027 78091 18069 78100
rect 18220 77720 18260 79612
rect 18316 79148 18356 79157
rect 18316 78476 18356 79108
rect 18316 78427 18356 78436
rect 18220 77671 18260 77680
rect 17932 74444 17972 76924
rect 18316 77384 18356 77393
rect 17932 74395 17972 74404
rect 18028 76292 18068 76301
rect 17740 52891 17780 52900
rect 17836 70160 17876 70169
rect 17740 50420 17780 50429
rect 17548 42524 17588 42533
rect 17548 42365 17588 42484
rect 17547 42356 17589 42365
rect 17547 42316 17548 42356
rect 17588 42316 17589 42356
rect 17547 42307 17589 42316
rect 17452 35839 17492 35848
rect 17164 33991 17204 34000
rect 17548 31520 17588 31529
rect 17163 27404 17205 27413
rect 17163 27364 17164 27404
rect 17204 27364 17205 27404
rect 17163 27355 17205 27364
rect 17068 26767 17108 26776
rect 17164 26648 17204 27355
rect 17068 26608 17204 26648
rect 17068 20180 17108 26608
rect 17452 24128 17492 24137
rect 17164 23960 17204 23969
rect 17164 23036 17204 23920
rect 17259 23456 17301 23465
rect 17259 23416 17260 23456
rect 17300 23416 17301 23456
rect 17259 23407 17301 23416
rect 17164 22987 17204 22996
rect 17068 20140 17204 20180
rect 16972 3331 17012 3340
rect 17164 1196 17204 20140
rect 17260 14048 17300 23407
rect 17452 23120 17492 24088
rect 17452 23071 17492 23080
rect 17260 13999 17300 14008
rect 17356 17912 17396 17921
rect 17164 1147 17204 1156
rect 16780 727 16820 736
rect 17356 272 17396 17872
rect 17548 1196 17588 31480
rect 17644 31352 17684 31361
rect 17644 15560 17684 31312
rect 17644 15511 17684 15520
rect 17644 8840 17684 8849
rect 17644 5816 17684 8800
rect 17644 5060 17684 5776
rect 17644 5011 17684 5020
rect 17740 1280 17780 50380
rect 17836 42188 17876 70120
rect 17932 64112 17972 64121
rect 17932 42608 17972 64072
rect 17932 42559 17972 42568
rect 17836 42139 17876 42148
rect 17836 41516 17876 41525
rect 17836 38240 17876 41476
rect 17836 38191 17876 38200
rect 17932 39920 17972 39929
rect 17932 32864 17972 39880
rect 17932 32815 17972 32824
rect 17836 26900 17876 26909
rect 17836 25640 17876 26860
rect 17836 25591 17876 25600
rect 17835 24884 17877 24893
rect 17835 24844 17836 24884
rect 17876 24844 17877 24884
rect 17835 24835 17877 24844
rect 17836 23540 17876 24835
rect 17836 23491 17876 23500
rect 17836 20264 17876 20273
rect 17836 18416 17876 20224
rect 17836 18367 17876 18376
rect 17932 7664 17972 7673
rect 17932 4892 17972 7624
rect 17932 4556 17972 4852
rect 17932 4136 17972 4516
rect 17932 4087 17972 4096
rect 17740 1231 17780 1240
rect 17548 1147 17588 1156
rect 18028 1196 18068 76252
rect 18220 70328 18260 70337
rect 18220 67724 18260 70288
rect 18220 63608 18260 67684
rect 18220 63559 18260 63568
rect 18124 55292 18164 55301
rect 18124 1280 18164 55252
rect 18220 39164 18260 39173
rect 18220 38912 18260 39124
rect 18220 38863 18260 38872
rect 18220 18416 18260 18425
rect 18220 15476 18260 18376
rect 18220 15427 18260 15436
rect 18124 1231 18164 1240
rect 18028 1147 18068 1156
rect 18316 1028 18356 77344
rect 18412 76208 18452 83140
rect 18808 83180 19176 83189
rect 18848 83140 18890 83180
rect 18930 83140 18972 83180
rect 19012 83140 19054 83180
rect 19094 83140 19136 83180
rect 18808 83131 19176 83140
rect 19564 82592 19604 82601
rect 19564 82340 19604 82552
rect 19276 81920 19316 81929
rect 18808 81668 19176 81677
rect 18848 81628 18890 81668
rect 18930 81628 18972 81668
rect 19012 81628 19054 81668
rect 19094 81628 19136 81668
rect 18808 81619 19176 81628
rect 18700 81248 18740 81257
rect 18604 80408 18644 80417
rect 18412 76159 18452 76168
rect 18508 80072 18548 80081
rect 18508 79736 18548 80032
rect 18412 72176 18452 72185
rect 18412 43700 18452 72136
rect 18508 69992 18548 79696
rect 18508 69943 18548 69952
rect 18508 66380 18548 66389
rect 18508 63104 18548 66340
rect 18508 63055 18548 63064
rect 18508 51764 18548 51773
rect 18508 47900 18548 51724
rect 18604 49328 18644 80368
rect 18700 78392 18740 81208
rect 18808 80156 19176 80165
rect 18848 80116 18890 80156
rect 18930 80116 18972 80156
rect 19012 80116 19054 80156
rect 19094 80116 19136 80156
rect 18808 80107 19176 80116
rect 19276 79988 19316 81880
rect 19276 79939 19316 79948
rect 19564 79400 19604 82300
rect 19564 79351 19604 79360
rect 19276 78980 19316 78989
rect 18808 78644 19176 78653
rect 18848 78604 18890 78644
rect 18930 78604 18972 78644
rect 19012 78604 19054 78644
rect 19094 78604 19136 78644
rect 18808 78595 19176 78604
rect 18700 78343 18740 78352
rect 18808 77132 19176 77141
rect 18848 77092 18890 77132
rect 18930 77092 18972 77132
rect 19012 77092 19054 77132
rect 19094 77092 19136 77132
rect 18808 77083 19176 77092
rect 19276 76880 19316 78940
rect 19276 76831 19316 76840
rect 19660 76292 19700 84316
rect 20048 83936 20416 83945
rect 20088 83896 20130 83936
rect 20170 83896 20212 83936
rect 20252 83896 20294 83936
rect 20334 83896 20376 83936
rect 20048 83887 20416 83896
rect 20048 82424 20416 82433
rect 20088 82384 20130 82424
rect 20170 82384 20212 82424
rect 20252 82384 20294 82424
rect 20334 82384 20376 82424
rect 20048 82375 20416 82384
rect 20048 80912 20416 80921
rect 20088 80872 20130 80912
rect 20170 80872 20212 80912
rect 20252 80872 20294 80912
rect 20334 80872 20376 80912
rect 20048 80863 20416 80872
rect 19660 76243 19700 76252
rect 19948 80408 19988 80417
rect 19948 75788 19988 80368
rect 20048 79400 20416 79409
rect 20088 79360 20130 79400
rect 20170 79360 20212 79400
rect 20252 79360 20294 79400
rect 20334 79360 20376 79400
rect 20048 79351 20416 79360
rect 20048 77888 20416 77897
rect 20088 77848 20130 77888
rect 20170 77848 20212 77888
rect 20252 77848 20294 77888
rect 20334 77848 20376 77888
rect 20048 77839 20416 77848
rect 20048 76376 20416 76385
rect 20088 76336 20130 76376
rect 20170 76336 20212 76376
rect 20252 76336 20294 76376
rect 20334 76336 20376 76376
rect 20048 76327 20416 76336
rect 19948 75739 19988 75748
rect 18808 75620 19176 75629
rect 18848 75580 18890 75620
rect 18930 75580 18972 75620
rect 19012 75580 19054 75620
rect 19094 75580 19136 75620
rect 18808 75571 19176 75580
rect 18604 49279 18644 49288
rect 18700 75032 18740 75041
rect 18508 44960 18548 47860
rect 18508 44911 18548 44920
rect 18412 43651 18452 43660
rect 18604 43196 18644 43205
rect 18412 36308 18452 36317
rect 18412 34880 18452 36268
rect 18412 34831 18452 34840
rect 18508 33536 18548 33545
rect 18508 32948 18548 33496
rect 18508 31436 18548 32908
rect 18508 31387 18548 31396
rect 18604 30680 18644 43156
rect 18604 30631 18644 30640
rect 18604 22280 18644 22289
rect 18604 20180 18644 22240
rect 18604 20131 18644 20140
rect 18604 15560 18644 15569
rect 18412 8840 18452 8849
rect 18412 4724 18452 8800
rect 18604 8840 18644 15520
rect 18604 8791 18644 8800
rect 18412 4675 18452 4684
rect 18700 1280 18740 74992
rect 20048 74864 20416 74873
rect 20088 74824 20130 74864
rect 20170 74824 20212 74864
rect 20252 74824 20294 74864
rect 20334 74824 20376 74864
rect 20048 74815 20416 74824
rect 18808 74108 19176 74117
rect 18848 74068 18890 74108
rect 18930 74068 18972 74108
rect 19012 74068 19054 74108
rect 19094 74068 19136 74108
rect 18808 74059 19176 74068
rect 20048 73352 20416 73361
rect 20088 73312 20130 73352
rect 20170 73312 20212 73352
rect 20252 73312 20294 73352
rect 20334 73312 20376 73352
rect 20048 73303 20416 73312
rect 19660 72764 19700 72773
rect 18808 72596 19176 72605
rect 18848 72556 18890 72596
rect 18930 72556 18972 72596
rect 19012 72556 19054 72596
rect 19094 72556 19136 72596
rect 18808 72547 19176 72556
rect 19276 72092 19316 72101
rect 18808 71084 19176 71093
rect 18848 71044 18890 71084
rect 18930 71044 18972 71084
rect 19012 71044 19054 71084
rect 19094 71044 19136 71084
rect 18808 71035 19176 71044
rect 19276 69824 19316 72052
rect 19276 69775 19316 69784
rect 19564 71084 19604 71093
rect 18808 69572 19176 69581
rect 18848 69532 18890 69572
rect 18930 69532 18972 69572
rect 19012 69532 19054 69572
rect 19094 69532 19136 69572
rect 18808 69523 19176 69532
rect 19564 69068 19604 71044
rect 19660 70748 19700 72724
rect 20048 71840 20416 71849
rect 20088 71800 20130 71840
rect 20170 71800 20212 71840
rect 20252 71800 20294 71840
rect 20334 71800 20376 71840
rect 20048 71791 20416 71800
rect 21388 71840 21428 71849
rect 20812 71504 20852 71513
rect 19660 70699 19700 70708
rect 19852 71252 19892 71261
rect 19564 69019 19604 69028
rect 19276 68984 19316 68993
rect 18808 68060 19176 68069
rect 18848 68020 18890 68060
rect 18930 68020 18972 68060
rect 19012 68020 19054 68060
rect 19094 68020 19136 68060
rect 18808 68011 19176 68020
rect 18808 66548 19176 66557
rect 18848 66508 18890 66548
rect 18930 66508 18972 66548
rect 19012 66508 19054 66548
rect 19094 66508 19136 66548
rect 18808 66499 19176 66508
rect 18808 65036 19176 65045
rect 18848 64996 18890 65036
rect 18930 64996 18972 65036
rect 19012 64996 19054 65036
rect 19094 64996 19136 65036
rect 18808 64987 19176 64996
rect 19276 64877 19316 68944
rect 19660 67052 19700 67061
rect 19275 64868 19317 64877
rect 19275 64828 19276 64868
rect 19316 64828 19317 64868
rect 19275 64819 19317 64828
rect 19275 64448 19317 64457
rect 19275 64408 19276 64448
rect 19316 64408 19317 64448
rect 19275 64399 19317 64408
rect 19276 64314 19316 64399
rect 18808 63524 19176 63533
rect 18848 63484 18890 63524
rect 18930 63484 18972 63524
rect 19012 63484 19054 63524
rect 19094 63484 19136 63524
rect 18808 63475 19176 63484
rect 19276 63440 19316 63449
rect 18808 62012 19176 62021
rect 18848 61972 18890 62012
rect 18930 61972 18972 62012
rect 19012 61972 19054 62012
rect 19094 61972 19136 62012
rect 18808 61963 19176 61972
rect 18808 60500 19176 60509
rect 18848 60460 18890 60500
rect 18930 60460 18972 60500
rect 19012 60460 19054 60500
rect 19094 60460 19136 60500
rect 18808 60451 19176 60460
rect 19276 59408 19316 63400
rect 19276 59359 19316 59368
rect 19468 61592 19508 61601
rect 18808 58988 19176 58997
rect 18848 58948 18890 58988
rect 18930 58948 18972 58988
rect 19012 58948 19054 58988
rect 19094 58948 19136 58988
rect 18808 58939 19176 58948
rect 19276 58652 19316 58661
rect 18808 57476 19176 57485
rect 18848 57436 18890 57476
rect 18930 57436 18972 57476
rect 19012 57436 19054 57476
rect 19094 57436 19136 57476
rect 18808 57427 19176 57436
rect 18808 55964 19176 55973
rect 18848 55924 18890 55964
rect 18930 55924 18972 55964
rect 19012 55924 19054 55964
rect 19094 55924 19136 55964
rect 18808 55915 19176 55924
rect 18808 54452 19176 54461
rect 18848 54412 18890 54452
rect 18930 54412 18972 54452
rect 19012 54412 19054 54452
rect 19094 54412 19136 54452
rect 18808 54403 19176 54412
rect 18808 52940 19176 52949
rect 18848 52900 18890 52940
rect 18930 52900 18972 52940
rect 19012 52900 19054 52940
rect 19094 52900 19136 52940
rect 18808 52891 19176 52900
rect 18808 51428 19176 51437
rect 18848 51388 18890 51428
rect 18930 51388 18972 51428
rect 19012 51388 19054 51428
rect 19094 51388 19136 51428
rect 18808 51379 19176 51388
rect 19276 50924 19316 58612
rect 19276 50336 19316 50884
rect 19276 50287 19316 50296
rect 19372 53780 19412 53789
rect 18808 49916 19176 49925
rect 18848 49876 18890 49916
rect 18930 49876 18972 49916
rect 19012 49876 19054 49916
rect 19094 49876 19136 49916
rect 18808 49867 19176 49876
rect 18808 48404 19176 48413
rect 18848 48364 18890 48404
rect 18930 48364 18972 48404
rect 19012 48364 19054 48404
rect 19094 48364 19136 48404
rect 18808 48355 19176 48364
rect 18808 46892 19176 46901
rect 18848 46852 18890 46892
rect 18930 46852 18972 46892
rect 19012 46852 19054 46892
rect 19094 46852 19136 46892
rect 18808 46843 19176 46852
rect 18808 45380 19176 45389
rect 18848 45340 18890 45380
rect 18930 45340 18972 45380
rect 19012 45340 19054 45380
rect 19094 45340 19136 45380
rect 18808 45331 19176 45340
rect 18808 43868 19176 43877
rect 18848 43828 18890 43868
rect 18930 43828 18972 43868
rect 19012 43828 19054 43868
rect 19094 43828 19136 43868
rect 18808 43819 19176 43828
rect 18808 42356 19176 42365
rect 18848 42316 18890 42356
rect 18930 42316 18972 42356
rect 19012 42316 19054 42356
rect 19094 42316 19136 42356
rect 18808 42307 19176 42316
rect 19372 42188 19412 53740
rect 19468 52772 19508 61552
rect 19563 59492 19605 59501
rect 19563 59452 19564 59492
rect 19604 59452 19605 59492
rect 19563 59443 19605 59452
rect 19564 59358 19604 59443
rect 19660 54200 19700 67012
rect 19660 54151 19700 54160
rect 19756 66800 19796 66809
rect 19468 52723 19508 52732
rect 19468 52352 19508 52361
rect 19468 48236 19508 52312
rect 19468 48187 19508 48196
rect 19564 51512 19604 51521
rect 19372 42139 19412 42148
rect 19468 44036 19508 44045
rect 18808 40844 19176 40853
rect 18848 40804 18890 40844
rect 18930 40804 18972 40844
rect 19012 40804 19054 40844
rect 19094 40804 19136 40844
rect 18808 40795 19176 40804
rect 19468 40340 19508 43996
rect 19468 40291 19508 40300
rect 19372 39500 19412 39509
rect 18808 39332 19176 39341
rect 18848 39292 18890 39332
rect 18930 39292 18972 39332
rect 19012 39292 19054 39332
rect 19094 39292 19136 39332
rect 18808 39283 19176 39292
rect 19276 38828 19316 38837
rect 18808 37820 19176 37829
rect 18848 37780 18890 37820
rect 18930 37780 18972 37820
rect 19012 37780 19054 37820
rect 19094 37780 19136 37820
rect 18808 37771 19176 37780
rect 19276 36560 19316 38788
rect 18808 36308 19176 36317
rect 18848 36268 18890 36308
rect 18930 36268 18972 36308
rect 19012 36268 19054 36308
rect 19094 36268 19136 36308
rect 18808 36259 19176 36268
rect 18808 34796 19176 34805
rect 18848 34756 18890 34796
rect 18930 34756 18972 34796
rect 19012 34756 19054 34796
rect 19094 34756 19136 34796
rect 18808 34747 19176 34756
rect 18808 33284 19176 33293
rect 18848 33244 18890 33284
rect 18930 33244 18972 33284
rect 19012 33244 19054 33284
rect 19094 33244 19136 33284
rect 18808 33235 19176 33244
rect 18808 31772 19176 31781
rect 18848 31732 18890 31772
rect 18930 31732 18972 31772
rect 19012 31732 19054 31772
rect 19094 31732 19136 31772
rect 18808 31723 19176 31732
rect 18808 30260 19176 30269
rect 18848 30220 18890 30260
rect 18930 30220 18972 30260
rect 19012 30220 19054 30260
rect 19094 30220 19136 30260
rect 18808 30211 19176 30220
rect 18808 28748 19176 28757
rect 18848 28708 18890 28748
rect 18930 28708 18972 28748
rect 19012 28708 19054 28748
rect 19094 28708 19136 28748
rect 18808 28699 19176 28708
rect 19276 28328 19316 36520
rect 18808 27236 19176 27245
rect 18848 27196 18890 27236
rect 18930 27196 18972 27236
rect 19012 27196 19054 27236
rect 19094 27196 19136 27236
rect 18808 27187 19176 27196
rect 19276 26732 19316 28288
rect 19276 26683 19316 26692
rect 19372 36728 19412 39460
rect 18808 25724 19176 25733
rect 18848 25684 18890 25724
rect 18930 25684 18972 25724
rect 19012 25684 19054 25724
rect 19094 25684 19136 25724
rect 18808 25675 19176 25684
rect 18808 24212 19176 24221
rect 18848 24172 18890 24212
rect 18930 24172 18972 24212
rect 19012 24172 19054 24212
rect 19094 24172 19136 24212
rect 18808 24163 19176 24172
rect 19276 22952 19316 22961
rect 18808 22700 19176 22709
rect 18848 22660 18890 22700
rect 18930 22660 18972 22700
rect 19012 22660 19054 22700
rect 19094 22660 19136 22700
rect 18808 22651 19176 22660
rect 19276 22532 19316 22912
rect 19276 22483 19316 22492
rect 19276 21608 19316 21617
rect 18808 21188 19176 21197
rect 18848 21148 18890 21188
rect 18930 21148 18972 21188
rect 19012 21148 19054 21188
rect 19094 21148 19136 21188
rect 18808 21139 19176 21148
rect 19276 20012 19316 21568
rect 19276 19963 19316 19972
rect 18808 19676 19176 19685
rect 18848 19636 18890 19676
rect 18930 19636 18972 19676
rect 19012 19636 19054 19676
rect 19094 19636 19136 19676
rect 18808 19627 19176 19636
rect 19372 19424 19412 36688
rect 19468 38912 19508 38921
rect 19468 27992 19508 38872
rect 19564 38408 19604 51472
rect 19756 43700 19796 66760
rect 19852 64616 19892 71212
rect 20716 70496 20756 70505
rect 20048 70328 20416 70337
rect 20088 70288 20130 70328
rect 20170 70288 20212 70328
rect 20252 70288 20294 70328
rect 20334 70288 20376 70328
rect 20048 70279 20416 70288
rect 19948 70076 19988 70085
rect 19948 68657 19988 70036
rect 20620 69488 20660 69497
rect 20048 68816 20416 68825
rect 20088 68776 20130 68816
rect 20170 68776 20212 68816
rect 20252 68776 20294 68816
rect 20334 68776 20376 68816
rect 20048 68767 20416 68776
rect 19947 68648 19989 68657
rect 19947 68608 19948 68648
rect 19988 68608 19989 68648
rect 19947 68599 19989 68608
rect 20620 67481 20660 69448
rect 20619 67472 20661 67481
rect 20619 67432 20620 67472
rect 20660 67432 20661 67472
rect 20619 67423 20661 67432
rect 20048 67304 20416 67313
rect 20088 67264 20130 67304
rect 20170 67264 20212 67304
rect 20252 67264 20294 67304
rect 20334 67264 20376 67304
rect 20048 67255 20416 67264
rect 20048 65792 20416 65801
rect 20088 65752 20130 65792
rect 20170 65752 20212 65792
rect 20252 65752 20294 65792
rect 20334 65752 20376 65792
rect 20048 65743 20416 65752
rect 20524 64868 20564 64877
rect 19948 64616 19988 64625
rect 19852 64576 19948 64616
rect 19852 61508 19892 61517
rect 19852 58064 19892 61468
rect 19948 59828 19988 64576
rect 20048 64280 20416 64289
rect 20088 64240 20130 64280
rect 20170 64240 20212 64280
rect 20252 64240 20294 64280
rect 20334 64240 20376 64280
rect 20048 64231 20416 64240
rect 20048 62768 20416 62777
rect 20088 62728 20130 62768
rect 20170 62728 20212 62768
rect 20252 62728 20294 62768
rect 20334 62728 20376 62768
rect 20048 62719 20416 62728
rect 20236 62432 20276 62441
rect 20236 61433 20276 62392
rect 20235 61424 20277 61433
rect 20235 61384 20236 61424
rect 20276 61384 20277 61424
rect 20235 61375 20277 61384
rect 20048 61256 20416 61265
rect 20088 61216 20130 61256
rect 20170 61216 20212 61256
rect 20252 61216 20294 61256
rect 20334 61216 20376 61256
rect 20048 61207 20416 61216
rect 19948 59779 19988 59788
rect 20048 59744 20416 59753
rect 20088 59704 20130 59744
rect 20170 59704 20212 59744
rect 20252 59704 20294 59744
rect 20334 59704 20376 59744
rect 20048 59695 20416 59704
rect 20048 58232 20416 58241
rect 20088 58192 20130 58232
rect 20170 58192 20212 58232
rect 20252 58192 20294 58232
rect 20334 58192 20376 58232
rect 20048 58183 20416 58192
rect 19852 58015 19892 58024
rect 20048 56720 20416 56729
rect 20088 56680 20130 56720
rect 20170 56680 20212 56720
rect 20252 56680 20294 56720
rect 20334 56680 20376 56720
rect 20048 56671 20416 56680
rect 19948 56132 19988 56141
rect 19948 55040 19988 56092
rect 20048 55208 20416 55217
rect 20088 55168 20130 55208
rect 20170 55168 20212 55208
rect 20252 55168 20294 55208
rect 20334 55168 20376 55208
rect 20048 55159 20416 55168
rect 19948 54991 19988 55000
rect 20524 54200 20564 64828
rect 20716 62852 20756 70456
rect 20524 54151 20564 54160
rect 20620 62812 20756 62852
rect 20048 53696 20416 53705
rect 20088 53656 20130 53696
rect 20170 53656 20212 53696
rect 20252 53656 20294 53696
rect 20334 53656 20376 53696
rect 20048 53647 20416 53656
rect 19756 43651 19796 43660
rect 19852 52940 19892 52949
rect 19564 38359 19604 38368
rect 19756 38492 19796 38501
rect 19756 35300 19796 38452
rect 19852 38240 19892 52900
rect 19948 52856 19988 52865
rect 19948 45548 19988 52816
rect 20048 52184 20416 52193
rect 20088 52144 20130 52184
rect 20170 52144 20212 52184
rect 20252 52144 20294 52184
rect 20334 52144 20376 52184
rect 20048 52135 20416 52144
rect 20048 50672 20416 50681
rect 20088 50632 20130 50672
rect 20170 50632 20212 50672
rect 20252 50632 20294 50672
rect 20334 50632 20376 50672
rect 20048 50623 20416 50632
rect 20139 49916 20181 49925
rect 20139 49876 20140 49916
rect 20180 49876 20181 49916
rect 20139 49867 20181 49876
rect 20140 49782 20180 49867
rect 20524 49328 20564 49337
rect 20048 49160 20416 49169
rect 20088 49120 20130 49160
rect 20170 49120 20212 49160
rect 20252 49120 20294 49160
rect 20334 49120 20376 49160
rect 20048 49111 20416 49120
rect 20048 47648 20416 47657
rect 20088 47608 20130 47648
rect 20170 47608 20212 47648
rect 20252 47608 20294 47648
rect 20334 47608 20376 47648
rect 20048 47599 20416 47608
rect 20048 46136 20416 46145
rect 20088 46096 20130 46136
rect 20170 46096 20212 46136
rect 20252 46096 20294 46136
rect 20334 46096 20376 46136
rect 20048 46087 20416 46096
rect 19948 45499 19988 45508
rect 20139 44960 20181 44969
rect 20139 44920 20140 44960
rect 20180 44920 20181 44960
rect 20139 44911 20181 44920
rect 20140 44826 20180 44911
rect 20048 44624 20416 44633
rect 20088 44584 20130 44624
rect 20170 44584 20212 44624
rect 20252 44584 20294 44624
rect 20334 44584 20376 44624
rect 20048 44575 20416 44584
rect 20048 43112 20416 43121
rect 20088 43072 20130 43112
rect 20170 43072 20212 43112
rect 20252 43072 20294 43112
rect 20334 43072 20376 43112
rect 20048 43063 20416 43072
rect 20044 42860 20084 42869
rect 19947 42524 19989 42533
rect 19947 42484 19948 42524
rect 19988 42484 19989 42524
rect 19947 42475 19989 42484
rect 19948 42390 19988 42475
rect 20044 41768 20084 42820
rect 19852 38191 19892 38200
rect 19948 41728 20084 41768
rect 19948 38072 19988 41728
rect 20048 41600 20416 41609
rect 20088 41560 20130 41600
rect 20170 41560 20212 41600
rect 20252 41560 20294 41600
rect 20334 41560 20376 41600
rect 20048 41551 20416 41560
rect 20048 40088 20416 40097
rect 20088 40048 20130 40088
rect 20170 40048 20212 40088
rect 20252 40048 20294 40088
rect 20334 40048 20376 40088
rect 20048 40039 20416 40048
rect 20048 38576 20416 38585
rect 20088 38536 20130 38576
rect 20170 38536 20212 38576
rect 20252 38536 20294 38576
rect 20334 38536 20376 38576
rect 20048 38527 20416 38536
rect 19948 38023 19988 38032
rect 20048 37064 20416 37073
rect 20088 37024 20130 37064
rect 20170 37024 20212 37064
rect 20252 37024 20294 37064
rect 20334 37024 20376 37064
rect 20048 37015 20416 37024
rect 20048 35552 20416 35561
rect 20088 35512 20130 35552
rect 20170 35512 20212 35552
rect 20252 35512 20294 35552
rect 20334 35512 20376 35552
rect 20048 35503 20416 35512
rect 19756 35251 19796 35260
rect 20048 34040 20416 34049
rect 20088 34000 20130 34040
rect 20170 34000 20212 34040
rect 20252 34000 20294 34040
rect 20334 34000 20376 34040
rect 20048 33991 20416 34000
rect 20048 32528 20416 32537
rect 20088 32488 20130 32528
rect 20170 32488 20212 32528
rect 20252 32488 20294 32528
rect 20334 32488 20376 32528
rect 20048 32479 20416 32488
rect 20048 31016 20416 31025
rect 20088 30976 20130 31016
rect 20170 30976 20212 31016
rect 20252 30976 20294 31016
rect 20334 30976 20376 31016
rect 20048 30967 20416 30976
rect 19468 27943 19508 27952
rect 19756 30092 19796 30101
rect 19756 22784 19796 30052
rect 20048 29504 20416 29513
rect 20088 29464 20130 29504
rect 20170 29464 20212 29504
rect 20252 29464 20294 29504
rect 20334 29464 20376 29504
rect 20048 29455 20416 29464
rect 20048 27992 20416 28001
rect 20088 27952 20130 27992
rect 20170 27952 20212 27992
rect 20252 27952 20294 27992
rect 20334 27952 20376 27992
rect 20048 27943 20416 27952
rect 20048 26480 20416 26489
rect 20088 26440 20130 26480
rect 20170 26440 20212 26480
rect 20252 26440 20294 26480
rect 20334 26440 20376 26480
rect 20048 26431 20416 26440
rect 20048 24968 20416 24977
rect 20088 24928 20130 24968
rect 20170 24928 20212 24968
rect 20252 24928 20294 24968
rect 20334 24928 20376 24968
rect 20048 24919 20416 24928
rect 20139 23792 20181 23801
rect 20139 23752 20140 23792
rect 20180 23752 20181 23792
rect 20139 23743 20181 23752
rect 20140 23658 20180 23743
rect 20048 23456 20416 23465
rect 20088 23416 20130 23456
rect 20170 23416 20212 23456
rect 20252 23416 20294 23456
rect 20334 23416 20376 23456
rect 20048 23407 20416 23416
rect 19756 22735 19796 22744
rect 19276 18584 19316 18593
rect 18808 18164 19176 18173
rect 18848 18124 18890 18164
rect 18930 18124 18972 18164
rect 19012 18124 19054 18164
rect 19094 18124 19136 18164
rect 18808 18115 19176 18124
rect 18808 16652 19176 16661
rect 18848 16612 18890 16652
rect 18930 16612 18972 16652
rect 19012 16612 19054 16652
rect 19094 16612 19136 16652
rect 18808 16603 19176 16612
rect 19276 16484 19316 18544
rect 19276 15812 19316 16444
rect 19276 15763 19316 15772
rect 18808 15140 19176 15149
rect 18848 15100 18890 15140
rect 18930 15100 18972 15140
rect 19012 15100 19054 15140
rect 19094 15100 19136 15140
rect 18808 15091 19176 15100
rect 18808 13628 19176 13637
rect 18848 13588 18890 13628
rect 18930 13588 18972 13628
rect 19012 13588 19054 13628
rect 19094 13588 19136 13628
rect 18808 13579 19176 13588
rect 19372 12536 19412 19384
rect 19468 22532 19508 22541
rect 19468 17072 19508 22492
rect 20139 22448 20181 22457
rect 20139 22408 20140 22448
rect 20180 22408 20181 22448
rect 20139 22399 20181 22408
rect 20140 22314 20180 22399
rect 20048 21944 20416 21953
rect 20088 21904 20130 21944
rect 20170 21904 20212 21944
rect 20252 21904 20294 21944
rect 20334 21904 20376 21944
rect 20048 21895 20416 21904
rect 20139 21776 20181 21785
rect 20139 21736 20140 21776
rect 20180 21736 20181 21776
rect 20139 21727 20181 21736
rect 20140 21642 20180 21727
rect 20048 20432 20416 20441
rect 20088 20392 20130 20432
rect 20170 20392 20212 20432
rect 20252 20392 20294 20432
rect 20334 20392 20376 20432
rect 20048 20383 20416 20392
rect 20048 18920 20416 18929
rect 20088 18880 20130 18920
rect 20170 18880 20212 18920
rect 20252 18880 20294 18920
rect 20334 18880 20376 18920
rect 20048 18871 20416 18880
rect 20048 17408 20416 17417
rect 20088 17368 20130 17408
rect 20170 17368 20212 17408
rect 20252 17368 20294 17408
rect 20334 17368 20376 17408
rect 20048 17359 20416 17368
rect 19468 17023 19508 17032
rect 19948 16316 19988 16325
rect 19948 15476 19988 16276
rect 20048 15896 20416 15905
rect 20088 15856 20130 15896
rect 20170 15856 20212 15896
rect 20252 15856 20294 15896
rect 20334 15856 20376 15896
rect 20048 15847 20416 15856
rect 19948 15427 19988 15436
rect 20048 14384 20416 14393
rect 20088 14344 20130 14384
rect 20170 14344 20212 14384
rect 20252 14344 20294 14384
rect 20334 14344 20376 14384
rect 20048 14335 20416 14344
rect 20048 12872 20416 12881
rect 20088 12832 20130 12872
rect 20170 12832 20212 12872
rect 20252 12832 20294 12872
rect 20334 12832 20376 12872
rect 20048 12823 20416 12832
rect 19372 12487 19412 12496
rect 19948 12536 19988 12545
rect 18808 12116 19176 12125
rect 18848 12076 18890 12116
rect 18930 12076 18972 12116
rect 19012 12076 19054 12116
rect 19094 12076 19136 12116
rect 18808 12067 19176 12076
rect 18808 10604 19176 10613
rect 18848 10564 18890 10604
rect 18930 10564 18972 10604
rect 19012 10564 19054 10604
rect 19094 10564 19136 10604
rect 18808 10555 19176 10564
rect 18808 9092 19176 9101
rect 18848 9052 18890 9092
rect 18930 9052 18972 9092
rect 19012 9052 19054 9092
rect 19094 9052 19136 9092
rect 18808 9043 19176 9052
rect 19948 8420 19988 12496
rect 20048 11360 20416 11369
rect 20088 11320 20130 11360
rect 20170 11320 20212 11360
rect 20252 11320 20294 11360
rect 20334 11320 20376 11360
rect 20048 11311 20416 11320
rect 20048 9848 20416 9857
rect 20088 9808 20130 9848
rect 20170 9808 20212 9848
rect 20252 9808 20294 9848
rect 20334 9808 20376 9848
rect 20048 9799 20416 9808
rect 19948 8371 19988 8380
rect 20048 8336 20416 8345
rect 20088 8296 20130 8336
rect 20170 8296 20212 8336
rect 20252 8296 20294 8336
rect 20334 8296 20376 8336
rect 20048 8287 20416 8296
rect 19276 7832 19316 7841
rect 18808 7580 19176 7589
rect 18848 7540 18890 7580
rect 18930 7540 18972 7580
rect 19012 7540 19054 7580
rect 19094 7540 19136 7580
rect 18808 7531 19176 7540
rect 18808 6068 19176 6077
rect 18848 6028 18890 6068
rect 18930 6028 18972 6068
rect 19012 6028 19054 6068
rect 19094 6028 19136 6068
rect 18808 6019 19176 6028
rect 19276 5648 19316 7792
rect 20048 6824 20416 6833
rect 20088 6784 20130 6824
rect 20170 6784 20212 6824
rect 20252 6784 20294 6824
rect 20334 6784 20376 6824
rect 20048 6775 20416 6784
rect 19276 5599 19316 5608
rect 20048 5312 20416 5321
rect 20088 5272 20130 5312
rect 20170 5272 20212 5312
rect 20252 5272 20294 5312
rect 20334 5272 20376 5312
rect 20048 5263 20416 5272
rect 18808 4556 19176 4565
rect 18848 4516 18890 4556
rect 18930 4516 18972 4556
rect 19012 4516 19054 4556
rect 19094 4516 19136 4556
rect 18808 4507 19176 4516
rect 20048 3800 20416 3809
rect 20088 3760 20130 3800
rect 20170 3760 20212 3800
rect 20252 3760 20294 3800
rect 20334 3760 20376 3800
rect 20048 3751 20416 3760
rect 18808 3044 19176 3053
rect 18848 3004 18890 3044
rect 18930 3004 18972 3044
rect 19012 3004 19054 3044
rect 19094 3004 19136 3044
rect 18808 2995 19176 3004
rect 20048 2288 20416 2297
rect 20088 2248 20130 2288
rect 20170 2248 20212 2288
rect 20252 2248 20294 2288
rect 20334 2248 20376 2288
rect 20048 2239 20416 2248
rect 18808 1532 19176 1541
rect 18848 1492 18890 1532
rect 18930 1492 18972 1532
rect 19012 1492 19054 1532
rect 19094 1492 19136 1532
rect 18808 1483 19176 1492
rect 18700 1231 18740 1240
rect 18316 979 18356 988
rect 20524 860 20564 49288
rect 20620 41432 20660 62812
rect 20716 61424 20756 61433
rect 20716 57392 20756 61384
rect 20716 57343 20756 57352
rect 20716 49664 20756 49673
rect 20716 47312 20756 49624
rect 20716 47263 20756 47272
rect 20812 42188 20852 71464
rect 20908 68480 20948 68489
rect 20908 63701 20948 68440
rect 21196 65120 21236 65129
rect 21004 64784 21044 64793
rect 20907 63692 20949 63701
rect 20907 63652 20908 63692
rect 20948 63652 20949 63692
rect 20907 63643 20949 63652
rect 20908 51932 20948 51941
rect 20908 48656 20948 51892
rect 21004 51512 21044 64744
rect 21004 51463 21044 51472
rect 20908 48607 20948 48616
rect 20812 42139 20852 42148
rect 20908 43280 20948 43289
rect 20908 41600 20948 43240
rect 21196 42860 21236 65080
rect 21196 42811 21236 42820
rect 21388 42776 21428 71800
rect 21388 42727 21428 42736
rect 20620 41383 20660 41392
rect 20812 41560 20948 41600
rect 21004 42608 21044 42617
rect 20620 40592 20660 40601
rect 20620 37652 20660 40552
rect 20620 37603 20660 37612
rect 20716 39248 20756 39257
rect 20620 34712 20660 34721
rect 20620 31520 20660 34672
rect 20716 34628 20756 39208
rect 20812 38324 20852 41560
rect 20812 38275 20852 38284
rect 20716 34579 20756 34588
rect 20715 32108 20757 32117
rect 20715 32068 20716 32108
rect 20756 32068 20757 32108
rect 20715 32059 20757 32068
rect 20620 31471 20660 31480
rect 20619 26648 20661 26657
rect 20619 26608 20620 26648
rect 20660 26608 20661 26648
rect 20619 26599 20661 26608
rect 20620 26480 20660 26599
rect 20620 26431 20660 26440
rect 20716 26312 20756 32059
rect 20716 26263 20756 26272
rect 20619 24632 20661 24641
rect 20619 24592 20620 24632
rect 20660 24592 20661 24632
rect 20619 24583 20661 24592
rect 20620 19760 20660 24583
rect 20811 24548 20853 24557
rect 20811 24508 20812 24548
rect 20852 24508 20853 24548
rect 20811 24499 20853 24508
rect 20620 19711 20660 19720
rect 20812 19424 20852 24499
rect 21004 20180 21044 42568
rect 21388 34376 21428 34385
rect 21388 24128 21428 34336
rect 21388 24079 21428 24088
rect 21004 20131 21044 20140
rect 20812 19375 20852 19384
rect 20620 17408 20660 17417
rect 20620 10520 20660 17368
rect 20620 10471 20660 10480
rect 21388 17072 21428 17081
rect 21388 8756 21428 17032
rect 21388 8707 21428 8716
rect 20524 811 20564 820
rect 20048 776 20416 785
rect 20088 736 20130 776
rect 20170 736 20212 776
rect 20252 736 20294 776
rect 20334 736 20376 776
rect 20048 727 20416 736
rect 18891 692 18933 701
rect 18891 652 18892 692
rect 18932 652 18933 692
rect 18891 643 18933 652
rect 18892 558 18932 643
rect 17356 223 17396 232
rect 16108 139 16148 148
rect 19467 188 19509 197
rect 19467 148 19468 188
rect 19508 148 19509 188
rect 19467 139 19509 148
rect 19468 54 19508 139
<< via4 >>
rect 556 75832 596 75872
rect 556 73144 596 73184
rect 844 73060 884 73100
rect 364 23752 404 23792
rect 652 27700 692 27740
rect 556 23836 596 23876
rect 460 2836 500 2876
rect 1324 84316 1364 84356
rect 844 26608 884 26648
rect 1132 52732 1172 52772
rect 1420 74992 1460 75032
rect 1324 62140 1364 62180
rect 1228 37612 1268 37652
rect 1708 27448 1748 27488
rect 1228 14512 1268 14552
rect 1036 10900 1076 10940
rect 3052 80620 3092 80660
rect 2476 59452 2516 59492
rect 2284 53236 2324 53276
rect 2380 39040 2420 39080
rect 2380 26020 2420 26060
rect 2092 3592 2132 3632
rect 2764 61048 2804 61088
rect 2860 37276 2900 37316
rect 3688 84652 3728 84692
rect 3770 84652 3810 84692
rect 3852 84652 3892 84692
rect 3934 84652 3974 84692
rect 4016 84652 4056 84692
rect 4684 84316 4724 84356
rect 3688 83140 3728 83180
rect 3770 83140 3810 83180
rect 3852 83140 3892 83180
rect 3934 83140 3974 83180
rect 4016 83140 4056 83180
rect 3820 81964 3860 82004
rect 3688 81628 3728 81668
rect 3770 81628 3810 81668
rect 3852 81628 3892 81668
rect 3934 81628 3974 81668
rect 4016 81628 4056 81668
rect 3916 80620 3956 80660
rect 3688 80116 3728 80156
rect 3770 80116 3810 80156
rect 3852 80116 3892 80156
rect 3934 80116 3974 80156
rect 4016 80116 4056 80156
rect 3688 78604 3728 78644
rect 3770 78604 3810 78644
rect 3852 78604 3892 78644
rect 3934 78604 3974 78644
rect 4016 78604 4056 78644
rect 3688 77092 3728 77132
rect 3770 77092 3810 77132
rect 3852 77092 3892 77132
rect 3934 77092 3974 77132
rect 4016 77092 4056 77132
rect 3688 75580 3728 75620
rect 3770 75580 3810 75620
rect 3852 75580 3892 75620
rect 3934 75580 3974 75620
rect 4016 75580 4056 75620
rect 3688 74068 3728 74108
rect 3770 74068 3810 74108
rect 3852 74068 3892 74108
rect 3934 74068 3974 74108
rect 4016 74068 4056 74108
rect 3688 72556 3728 72596
rect 3770 72556 3810 72596
rect 3852 72556 3892 72596
rect 3934 72556 3974 72596
rect 4016 72556 4056 72596
rect 3688 71044 3728 71084
rect 3770 71044 3810 71084
rect 3852 71044 3892 71084
rect 3934 71044 3974 71084
rect 4016 71044 4056 71084
rect 3244 41896 3284 41936
rect 3148 41392 3188 41432
rect 2764 23752 2804 23792
rect 3052 26860 3092 26900
rect 3688 69532 3728 69572
rect 3770 69532 3810 69572
rect 3852 69532 3892 69572
rect 3934 69532 3974 69572
rect 4016 69532 4056 69572
rect 3688 68020 3728 68060
rect 3770 68020 3810 68060
rect 3852 68020 3892 68060
rect 3934 68020 3974 68060
rect 4016 68020 4056 68060
rect 3688 66508 3728 66548
rect 3770 66508 3810 66548
rect 3852 66508 3892 66548
rect 3934 66508 3974 66548
rect 4016 66508 4056 66548
rect 3688 64996 3728 65036
rect 3770 64996 3810 65036
rect 3852 64996 3892 65036
rect 3934 64996 3974 65036
rect 4016 64996 4056 65036
rect 3688 63484 3728 63524
rect 3770 63484 3810 63524
rect 3852 63484 3892 63524
rect 3934 63484 3974 63524
rect 4016 63484 4056 63524
rect 3688 61972 3728 62012
rect 3770 61972 3810 62012
rect 3852 61972 3892 62012
rect 3934 61972 3974 62012
rect 4016 61972 4056 62012
rect 3688 60460 3728 60500
rect 3770 60460 3810 60500
rect 3852 60460 3892 60500
rect 3934 60460 3974 60500
rect 4016 60460 4056 60500
rect 4928 83896 4968 83936
rect 5010 83896 5050 83936
rect 5092 83896 5132 83936
rect 5174 83896 5214 83936
rect 5256 83896 5296 83936
rect 4928 82384 4968 82424
rect 5010 82384 5050 82424
rect 5092 82384 5132 82424
rect 5174 82384 5214 82424
rect 5256 82384 5296 82424
rect 5452 82804 5492 82844
rect 3688 58948 3728 58988
rect 3770 58948 3810 58988
rect 3852 58948 3892 58988
rect 3934 58948 3974 58988
rect 4016 58948 4056 58988
rect 4204 59200 4244 59240
rect 3688 57436 3728 57476
rect 3770 57436 3810 57476
rect 3852 57436 3892 57476
rect 3934 57436 3974 57476
rect 4016 57436 4056 57476
rect 3688 55924 3728 55964
rect 3770 55924 3810 55964
rect 3852 55924 3892 55964
rect 3934 55924 3974 55964
rect 4016 55924 4056 55964
rect 3688 54412 3728 54452
rect 3770 54412 3810 54452
rect 3852 54412 3892 54452
rect 3934 54412 3974 54452
rect 4016 54412 4056 54452
rect 3688 52900 3728 52940
rect 3770 52900 3810 52940
rect 3852 52900 3892 52940
rect 3934 52900 3974 52940
rect 4016 52900 4056 52940
rect 3688 51388 3728 51428
rect 3770 51388 3810 51428
rect 3852 51388 3892 51428
rect 3934 51388 3974 51428
rect 4016 51388 4056 51428
rect 3688 49876 3728 49916
rect 3770 49876 3810 49916
rect 3852 49876 3892 49916
rect 3934 49876 3974 49916
rect 4016 49876 4056 49916
rect 3688 48364 3728 48404
rect 3770 48364 3810 48404
rect 3852 48364 3892 48404
rect 3934 48364 3974 48404
rect 4016 48364 4056 48404
rect 3688 46852 3728 46892
rect 3770 46852 3810 46892
rect 3852 46852 3892 46892
rect 3934 46852 3974 46892
rect 4016 46852 4056 46892
rect 3688 45340 3728 45380
rect 3770 45340 3810 45380
rect 3852 45340 3892 45380
rect 3934 45340 3974 45380
rect 4016 45340 4056 45380
rect 3688 43828 3728 43868
rect 3770 43828 3810 43868
rect 3852 43828 3892 43868
rect 3934 43828 3974 43868
rect 4016 43828 4056 43868
rect 3688 42316 3728 42356
rect 3770 42316 3810 42356
rect 3852 42316 3892 42356
rect 3934 42316 3974 42356
rect 4016 42316 4056 42356
rect 4928 80872 4968 80912
rect 5010 80872 5050 80912
rect 5092 80872 5132 80912
rect 5174 80872 5214 80912
rect 5256 80872 5296 80912
rect 4588 62140 4628 62180
rect 4928 79360 4968 79400
rect 5010 79360 5050 79400
rect 5092 79360 5132 79400
rect 5174 79360 5214 79400
rect 5256 79360 5296 79400
rect 4928 77848 4968 77888
rect 5010 77848 5050 77888
rect 5092 77848 5132 77888
rect 5174 77848 5214 77888
rect 5256 77848 5296 77888
rect 4928 76336 4968 76376
rect 5010 76336 5050 76376
rect 5092 76336 5132 76376
rect 5174 76336 5214 76376
rect 5256 76336 5296 76376
rect 4928 74824 4968 74864
rect 5010 74824 5050 74864
rect 5092 74824 5132 74864
rect 5174 74824 5214 74864
rect 5256 74824 5296 74864
rect 4928 73312 4968 73352
rect 5010 73312 5050 73352
rect 5092 73312 5132 73352
rect 5174 73312 5214 73352
rect 5256 73312 5296 73352
rect 4928 71800 4968 71840
rect 5010 71800 5050 71840
rect 5092 71800 5132 71840
rect 5174 71800 5214 71840
rect 5256 71800 5296 71840
rect 3688 40804 3728 40844
rect 3770 40804 3810 40844
rect 3852 40804 3892 40844
rect 3934 40804 3974 40844
rect 4016 40804 4056 40844
rect 3688 39292 3728 39332
rect 3770 39292 3810 39332
rect 3852 39292 3892 39332
rect 3934 39292 3974 39332
rect 4016 39292 4056 39332
rect 4928 70288 4968 70328
rect 5010 70288 5050 70328
rect 5092 70288 5132 70328
rect 5174 70288 5214 70328
rect 5256 70288 5296 70328
rect 4928 68776 4968 68816
rect 5010 68776 5050 68816
rect 5092 68776 5132 68816
rect 5174 68776 5214 68816
rect 5256 68776 5296 68816
rect 5164 67768 5204 67808
rect 5356 67768 5396 67808
rect 4928 67264 4968 67304
rect 5010 67264 5050 67304
rect 5092 67264 5132 67304
rect 5174 67264 5214 67304
rect 5256 67264 5296 67304
rect 4928 65752 4968 65792
rect 5010 65752 5050 65792
rect 5092 65752 5132 65792
rect 5174 65752 5214 65792
rect 5256 65752 5296 65792
rect 4928 64240 4968 64280
rect 5010 64240 5050 64280
rect 5092 64240 5132 64280
rect 5174 64240 5214 64280
rect 5256 64240 5296 64280
rect 4928 62728 4968 62768
rect 5010 62728 5050 62768
rect 5092 62728 5132 62768
rect 5174 62728 5214 62768
rect 5256 62728 5296 62768
rect 4928 61216 4968 61256
rect 5010 61216 5050 61256
rect 5092 61216 5132 61256
rect 5174 61216 5214 61256
rect 5256 61216 5296 61256
rect 4928 59704 4968 59744
rect 5010 59704 5050 59744
rect 5092 59704 5132 59744
rect 5174 59704 5214 59744
rect 5256 59704 5296 59744
rect 4928 58192 4968 58232
rect 5010 58192 5050 58232
rect 5092 58192 5132 58232
rect 5174 58192 5214 58232
rect 5256 58192 5296 58232
rect 4928 56680 4968 56720
rect 5010 56680 5050 56720
rect 5092 56680 5132 56720
rect 5174 56680 5214 56720
rect 5256 56680 5296 56720
rect 4928 55168 4968 55208
rect 5010 55168 5050 55208
rect 5092 55168 5132 55208
rect 5174 55168 5214 55208
rect 5256 55168 5296 55208
rect 4928 53656 4968 53696
rect 5010 53656 5050 53696
rect 5092 53656 5132 53696
rect 5174 53656 5214 53696
rect 5256 53656 5296 53696
rect 5068 52732 5108 52772
rect 4928 52144 4968 52184
rect 5010 52144 5050 52184
rect 5092 52144 5132 52184
rect 5174 52144 5214 52184
rect 5256 52144 5296 52184
rect 4928 50632 4968 50672
rect 5010 50632 5050 50672
rect 5092 50632 5132 50672
rect 5174 50632 5214 50672
rect 5256 50632 5296 50672
rect 4928 49120 4968 49160
rect 5010 49120 5050 49160
rect 5092 49120 5132 49160
rect 5174 49120 5214 49160
rect 5256 49120 5296 49160
rect 4928 47608 4968 47648
rect 5010 47608 5050 47648
rect 5092 47608 5132 47648
rect 5174 47608 5214 47648
rect 5256 47608 5296 47648
rect 4928 46096 4968 46136
rect 5010 46096 5050 46136
rect 5092 46096 5132 46136
rect 5174 46096 5214 46136
rect 5256 46096 5296 46136
rect 4928 44584 4968 44624
rect 5010 44584 5050 44624
rect 5092 44584 5132 44624
rect 5174 44584 5214 44624
rect 5256 44584 5296 44624
rect 4928 43072 4968 43112
rect 5010 43072 5050 43112
rect 5092 43072 5132 43112
rect 5174 43072 5214 43112
rect 5256 43072 5296 43112
rect 4780 41896 4820 41936
rect 4928 41560 4968 41600
rect 5010 41560 5050 41600
rect 5092 41560 5132 41600
rect 5174 41560 5214 41600
rect 5256 41560 5296 41600
rect 4300 39040 4340 39080
rect 3688 37780 3728 37820
rect 3770 37780 3810 37820
rect 3852 37780 3892 37820
rect 3934 37780 3974 37820
rect 4016 37780 4056 37820
rect 3820 37444 3860 37484
rect 4108 37276 4148 37316
rect 4108 36688 4148 36728
rect 3688 36268 3728 36308
rect 3770 36268 3810 36308
rect 3852 36268 3892 36308
rect 3934 36268 3974 36308
rect 4016 36268 4056 36308
rect 3688 34756 3728 34796
rect 3770 34756 3810 34796
rect 3852 34756 3892 34796
rect 3934 34756 3974 34796
rect 4016 34756 4056 34796
rect 4012 33832 4052 33872
rect 3688 33244 3728 33284
rect 3770 33244 3810 33284
rect 3852 33244 3892 33284
rect 3934 33244 3974 33284
rect 4016 33244 4056 33284
rect 3688 31732 3728 31772
rect 3770 31732 3810 31772
rect 3852 31732 3892 31772
rect 3934 31732 3974 31772
rect 4016 31732 4056 31772
rect 3688 30220 3728 30260
rect 3770 30220 3810 30260
rect 3852 30220 3892 30260
rect 3934 30220 3974 30260
rect 4016 30220 4056 30260
rect 4108 29632 4148 29672
rect 3688 28708 3728 28748
rect 3770 28708 3810 28748
rect 3852 28708 3892 28748
rect 3934 28708 3974 28748
rect 4016 28708 4056 28748
rect 4928 40048 4968 40088
rect 5010 40048 5050 40088
rect 5092 40048 5132 40088
rect 5174 40048 5214 40088
rect 5256 40048 5296 40088
rect 4684 35680 4724 35720
rect 3688 27196 3728 27236
rect 3770 27196 3810 27236
rect 3852 27196 3892 27236
rect 3934 27196 3974 27236
rect 4016 27196 4056 27236
rect 3688 25684 3728 25724
rect 3770 25684 3810 25724
rect 3852 25684 3892 25724
rect 3934 25684 3974 25724
rect 4016 25684 4056 25724
rect 4588 27700 4628 27740
rect 4492 25936 4532 25976
rect 3688 24172 3728 24212
rect 3770 24172 3810 24212
rect 3852 24172 3892 24212
rect 3934 24172 3974 24212
rect 4016 24172 4056 24212
rect 3688 22660 3728 22700
rect 3770 22660 3810 22700
rect 3852 22660 3892 22700
rect 3934 22660 3974 22700
rect 4016 22660 4056 22700
rect 3688 21148 3728 21188
rect 3770 21148 3810 21188
rect 3852 21148 3892 21188
rect 3934 21148 3974 21188
rect 4016 21148 4056 21188
rect 3688 19636 3728 19676
rect 3770 19636 3810 19676
rect 3852 19636 3892 19676
rect 3934 19636 3974 19676
rect 4016 19636 4056 19676
rect 3688 18124 3728 18164
rect 3770 18124 3810 18164
rect 3852 18124 3892 18164
rect 3934 18124 3974 18164
rect 4016 18124 4056 18164
rect 3688 16612 3728 16652
rect 3770 16612 3810 16652
rect 3852 16612 3892 16652
rect 3934 16612 3974 16652
rect 4016 16612 4056 16652
rect 3688 15100 3728 15140
rect 3770 15100 3810 15140
rect 3852 15100 3892 15140
rect 3934 15100 3974 15140
rect 4016 15100 4056 15140
rect 3688 13588 3728 13628
rect 3770 13588 3810 13628
rect 3852 13588 3892 13628
rect 3934 13588 3974 13628
rect 4016 13588 4056 13628
rect 3688 12076 3728 12116
rect 3770 12076 3810 12116
rect 3852 12076 3892 12116
rect 3934 12076 3974 12116
rect 4016 12076 4056 12116
rect 3436 10900 3476 10940
rect 2956 568 2996 608
rect 3688 10564 3728 10604
rect 3770 10564 3810 10604
rect 3852 10564 3892 10604
rect 3934 10564 3974 10604
rect 4016 10564 4056 10604
rect 3688 9052 3728 9092
rect 3770 9052 3810 9092
rect 3852 9052 3892 9092
rect 3934 9052 3974 9092
rect 4016 9052 4056 9092
rect 3688 7540 3728 7580
rect 3770 7540 3810 7580
rect 3852 7540 3892 7580
rect 3934 7540 3974 7580
rect 4016 7540 4056 7580
rect 3688 6028 3728 6068
rect 3770 6028 3810 6068
rect 3852 6028 3892 6068
rect 3934 6028 3974 6068
rect 4016 6028 4056 6068
rect 3688 4516 3728 4556
rect 3770 4516 3810 4556
rect 3852 4516 3892 4556
rect 3934 4516 3974 4556
rect 4016 4516 4056 4556
rect 4204 4516 4244 4556
rect 3688 3004 3728 3044
rect 3770 3004 3810 3044
rect 3852 3004 3892 3044
rect 3934 3004 3974 3044
rect 4016 3004 4056 3044
rect 3628 2752 3668 2792
rect 3688 1492 3728 1532
rect 3770 1492 3810 1532
rect 3852 1492 3892 1532
rect 3934 1492 3974 1532
rect 4016 1492 4056 1532
rect 4928 38536 4968 38576
rect 5010 38536 5050 38576
rect 5092 38536 5132 38576
rect 5174 38536 5214 38576
rect 5256 38536 5296 38576
rect 4928 37024 4968 37064
rect 5010 37024 5050 37064
rect 5092 37024 5132 37064
rect 5174 37024 5214 37064
rect 5256 37024 5296 37064
rect 4928 35512 4968 35552
rect 5010 35512 5050 35552
rect 5092 35512 5132 35552
rect 5174 35512 5214 35552
rect 5256 35512 5296 35552
rect 4928 34000 4968 34040
rect 5010 34000 5050 34040
rect 5092 34000 5132 34040
rect 5174 34000 5214 34040
rect 5256 34000 5296 34040
rect 4928 32488 4968 32528
rect 5010 32488 5050 32528
rect 5092 32488 5132 32528
rect 5174 32488 5214 32528
rect 5256 32488 5296 32528
rect 4928 30976 4968 31016
rect 5010 30976 5050 31016
rect 5092 30976 5132 31016
rect 5174 30976 5214 31016
rect 5256 30976 5296 31016
rect 4928 29464 4968 29504
rect 5010 29464 5050 29504
rect 5092 29464 5132 29504
rect 5174 29464 5214 29504
rect 5256 29464 5296 29504
rect 4928 27952 4968 27992
rect 5010 27952 5050 27992
rect 5092 27952 5132 27992
rect 5174 27952 5214 27992
rect 5256 27952 5296 27992
rect 4928 26440 4968 26480
rect 5010 26440 5050 26480
rect 5092 26440 5132 26480
rect 5174 26440 5214 26480
rect 5256 26440 5296 26480
rect 4928 24928 4968 24968
rect 5010 24928 5050 24968
rect 5092 24928 5132 24968
rect 5174 24928 5214 24968
rect 5256 24928 5296 24968
rect 4928 23416 4968 23456
rect 5010 23416 5050 23456
rect 5092 23416 5132 23456
rect 5174 23416 5214 23456
rect 5256 23416 5296 23456
rect 4928 21904 4968 21944
rect 5010 21904 5050 21944
rect 5092 21904 5132 21944
rect 5174 21904 5214 21944
rect 5256 21904 5296 21944
rect 4928 20392 4968 20432
rect 5010 20392 5050 20432
rect 5092 20392 5132 20432
rect 5174 20392 5214 20432
rect 5256 20392 5296 20432
rect 4928 18880 4968 18920
rect 5010 18880 5050 18920
rect 5092 18880 5132 18920
rect 5174 18880 5214 18920
rect 5256 18880 5296 18920
rect 4928 17368 4968 17408
rect 5010 17368 5050 17408
rect 5092 17368 5132 17408
rect 5174 17368 5214 17408
rect 5256 17368 5296 17408
rect 4928 15856 4968 15896
rect 5010 15856 5050 15896
rect 5092 15856 5132 15896
rect 5174 15856 5214 15896
rect 5256 15856 5296 15896
rect 4928 14344 4968 14384
rect 5010 14344 5050 14384
rect 5092 14344 5132 14384
rect 5174 14344 5214 14384
rect 5256 14344 5296 14384
rect 4928 12832 4968 12872
rect 5010 12832 5050 12872
rect 5092 12832 5132 12872
rect 5174 12832 5214 12872
rect 5256 12832 5296 12872
rect 4928 11320 4968 11360
rect 5010 11320 5050 11360
rect 5092 11320 5132 11360
rect 5174 11320 5214 11360
rect 5256 11320 5296 11360
rect 4876 10900 4916 10940
rect 4928 9808 4968 9848
rect 5010 9808 5050 9848
rect 5092 9808 5132 9848
rect 5174 9808 5214 9848
rect 5256 9808 5296 9848
rect 4928 8296 4968 8336
rect 5010 8296 5050 8336
rect 5092 8296 5132 8336
rect 5174 8296 5214 8336
rect 5256 8296 5296 8336
rect 4928 6784 4968 6824
rect 5010 6784 5050 6824
rect 5092 6784 5132 6824
rect 5174 6784 5214 6824
rect 5256 6784 5296 6824
rect 4928 5272 4968 5312
rect 5010 5272 5050 5312
rect 5092 5272 5132 5312
rect 5174 5272 5214 5312
rect 5256 5272 5296 5312
rect 5548 74992 5588 75032
rect 5644 36520 5684 36560
rect 5836 35680 5876 35720
rect 5836 29128 5876 29168
rect 4972 4516 5012 4556
rect 4928 3760 4968 3800
rect 5010 3760 5050 3800
rect 5092 3760 5132 3800
rect 5174 3760 5214 3800
rect 5256 3760 5296 3800
rect 4928 2248 4968 2288
rect 5010 2248 5050 2288
rect 5092 2248 5132 2288
rect 5174 2248 5214 2288
rect 5256 2248 5296 2288
rect 6028 30808 6068 30848
rect 6412 76840 6452 76880
rect 6220 67432 6260 67472
rect 6316 37612 6356 37652
rect 6316 37444 6356 37484
rect 6508 41644 6548 41684
rect 6508 37612 6548 37652
rect 6412 33832 6452 33872
rect 6220 30808 6260 30848
rect 6412 26860 6452 26900
rect 6412 25936 6452 25976
rect 6988 80620 7028 80660
rect 6700 75832 6740 75872
rect 6892 59200 6932 59240
rect 6892 41644 6932 41684
rect 6988 41560 7028 41600
rect 6988 36688 7028 36728
rect 6796 29632 6836 29672
rect 6988 12580 7028 12620
rect 7468 80788 7508 80828
rect 7276 41392 7316 41432
rect 7180 39040 7220 39080
rect 7180 36520 7220 36560
rect 8140 82804 8180 82844
rect 7756 79444 7796 79484
rect 7660 73060 7700 73100
rect 7564 61804 7604 61844
rect 7852 61804 7892 61844
rect 7564 41560 7604 41600
rect 7852 37696 7892 37736
rect 7180 27364 7220 27404
rect 7564 27448 7604 27488
rect 6796 4768 6836 4808
rect 7276 2752 7316 2792
rect 5740 1828 5780 1868
rect 6796 1072 6836 1112
rect 4928 736 4968 776
rect 5010 736 5050 776
rect 5092 736 5132 776
rect 5174 736 5214 776
rect 5256 736 5296 776
rect 7756 26020 7796 26060
rect 7756 23920 7796 23960
rect 7660 4516 7700 4556
rect 7564 2836 7604 2876
rect 8524 65836 8564 65876
rect 8428 64828 8468 64868
rect 8140 22408 8180 22448
rect 8524 49708 8564 49748
rect 8524 37696 8564 37736
rect 8716 48028 8756 48068
rect 8812 23920 8852 23960
rect 8812 14512 8852 14552
rect 8812 12580 8852 12620
rect 9004 23668 9044 23708
rect 7084 568 7124 608
rect 9964 83140 10004 83180
rect 9772 68608 9812 68648
rect 9676 67768 9716 67808
rect 9676 49456 9716 49496
rect 9868 64408 9908 64448
rect 10540 83476 10580 83516
rect 10060 82048 10100 82088
rect 9964 29128 10004 29168
rect 9772 27616 9812 27656
rect 10252 63148 10292 63188
rect 9580 7372 9620 7412
rect 10540 39880 10580 39920
rect 10636 30892 10676 30932
rect 11116 78100 11156 78140
rect 11020 63148 11060 63188
rect 10924 61384 10964 61424
rect 10828 53992 10868 54032
rect 12460 84064 12500 84104
rect 11212 59368 11252 59408
rect 11020 42484 11060 42524
rect 11116 42316 11156 42356
rect 11116 39880 11156 39920
rect 11020 33664 11060 33704
rect 10828 24844 10868 24884
rect 10732 5608 10772 5648
rect 11116 24508 11156 24548
rect 11788 59452 11828 59492
rect 11500 33664 11540 33704
rect 10540 2836 10580 2876
rect 11020 1828 11060 1868
rect 6988 316 7028 356
rect 8716 316 8756 356
rect 11308 1072 11348 1112
rect 11980 22660 12020 22700
rect 12076 15016 12116 15056
rect 12364 63652 12404 63692
rect 12268 44920 12308 44960
rect 12460 54580 12500 54620
rect 12652 54580 12692 54620
rect 12364 25180 12404 25220
rect 12460 24592 12500 24632
rect 18808 84652 18848 84692
rect 18890 84652 18930 84692
rect 18972 84652 19012 84692
rect 19054 84652 19094 84692
rect 19136 84652 19176 84692
rect 12940 20224 12980 20264
rect 13036 1828 13076 1868
rect 12748 1240 12788 1280
rect 13612 83308 13652 83348
rect 13228 53992 13268 54032
rect 13228 28876 13268 28916
rect 13228 20056 13268 20096
rect 13516 29632 13556 29672
rect 13708 55084 13748 55124
rect 13996 55084 14036 55124
rect 14284 64744 14324 64784
rect 14284 63148 14324 63188
rect 14476 69028 14516 69068
rect 14860 69028 14900 69068
rect 16012 83140 16052 83180
rect 16396 81040 16436 81080
rect 15052 77260 15092 77300
rect 14764 68944 14804 68984
rect 14956 68944 14996 68984
rect 14572 64744 14612 64784
rect 14284 53236 14324 53276
rect 14188 29632 14228 29672
rect 14860 56512 14900 56552
rect 14668 49456 14708 49496
rect 15052 56680 15092 56720
rect 15052 56512 15092 56552
rect 14764 47944 14804 47984
rect 14956 47944 14996 47984
rect 14476 27616 14516 27656
rect 14860 28876 14900 28916
rect 14764 23668 14804 23708
rect 15052 21736 15092 21776
rect 16684 66928 16724 66968
rect 16492 23416 16532 23456
rect 16396 22660 16436 22700
rect 16108 15016 16148 15056
rect 15628 736 15668 776
rect 12652 148 12692 188
rect 16876 30892 16916 30932
rect 18028 78100 18068 78140
rect 17548 42316 17588 42356
rect 17164 27364 17204 27404
rect 17260 23416 17300 23456
rect 17836 24844 17876 24884
rect 18808 83140 18848 83180
rect 18890 83140 18930 83180
rect 18972 83140 19012 83180
rect 19054 83140 19094 83180
rect 19136 83140 19176 83180
rect 18808 81628 18848 81668
rect 18890 81628 18930 81668
rect 18972 81628 19012 81668
rect 19054 81628 19094 81668
rect 19136 81628 19176 81668
rect 18808 80116 18848 80156
rect 18890 80116 18930 80156
rect 18972 80116 19012 80156
rect 19054 80116 19094 80156
rect 19136 80116 19176 80156
rect 18808 78604 18848 78644
rect 18890 78604 18930 78644
rect 18972 78604 19012 78644
rect 19054 78604 19094 78644
rect 19136 78604 19176 78644
rect 18808 77092 18848 77132
rect 18890 77092 18930 77132
rect 18972 77092 19012 77132
rect 19054 77092 19094 77132
rect 19136 77092 19176 77132
rect 20048 83896 20088 83936
rect 20130 83896 20170 83936
rect 20212 83896 20252 83936
rect 20294 83896 20334 83936
rect 20376 83896 20416 83936
rect 20048 82384 20088 82424
rect 20130 82384 20170 82424
rect 20212 82384 20252 82424
rect 20294 82384 20334 82424
rect 20376 82384 20416 82424
rect 20048 80872 20088 80912
rect 20130 80872 20170 80912
rect 20212 80872 20252 80912
rect 20294 80872 20334 80912
rect 20376 80872 20416 80912
rect 20048 79360 20088 79400
rect 20130 79360 20170 79400
rect 20212 79360 20252 79400
rect 20294 79360 20334 79400
rect 20376 79360 20416 79400
rect 20048 77848 20088 77888
rect 20130 77848 20170 77888
rect 20212 77848 20252 77888
rect 20294 77848 20334 77888
rect 20376 77848 20416 77888
rect 20048 76336 20088 76376
rect 20130 76336 20170 76376
rect 20212 76336 20252 76376
rect 20294 76336 20334 76376
rect 20376 76336 20416 76376
rect 18808 75580 18848 75620
rect 18890 75580 18930 75620
rect 18972 75580 19012 75620
rect 19054 75580 19094 75620
rect 19136 75580 19176 75620
rect 20048 74824 20088 74864
rect 20130 74824 20170 74864
rect 20212 74824 20252 74864
rect 20294 74824 20334 74864
rect 20376 74824 20416 74864
rect 18808 74068 18848 74108
rect 18890 74068 18930 74108
rect 18972 74068 19012 74108
rect 19054 74068 19094 74108
rect 19136 74068 19176 74108
rect 20048 73312 20088 73352
rect 20130 73312 20170 73352
rect 20212 73312 20252 73352
rect 20294 73312 20334 73352
rect 20376 73312 20416 73352
rect 18808 72556 18848 72596
rect 18890 72556 18930 72596
rect 18972 72556 19012 72596
rect 19054 72556 19094 72596
rect 19136 72556 19176 72596
rect 18808 71044 18848 71084
rect 18890 71044 18930 71084
rect 18972 71044 19012 71084
rect 19054 71044 19094 71084
rect 19136 71044 19176 71084
rect 18808 69532 18848 69572
rect 18890 69532 18930 69572
rect 18972 69532 19012 69572
rect 19054 69532 19094 69572
rect 19136 69532 19176 69572
rect 20048 71800 20088 71840
rect 20130 71800 20170 71840
rect 20212 71800 20252 71840
rect 20294 71800 20334 71840
rect 20376 71800 20416 71840
rect 18808 68020 18848 68060
rect 18890 68020 18930 68060
rect 18972 68020 19012 68060
rect 19054 68020 19094 68060
rect 19136 68020 19176 68060
rect 18808 66508 18848 66548
rect 18890 66508 18930 66548
rect 18972 66508 19012 66548
rect 19054 66508 19094 66548
rect 19136 66508 19176 66548
rect 18808 64996 18848 65036
rect 18890 64996 18930 65036
rect 18972 64996 19012 65036
rect 19054 64996 19094 65036
rect 19136 64996 19176 65036
rect 19276 64828 19316 64868
rect 19276 64408 19316 64448
rect 18808 63484 18848 63524
rect 18890 63484 18930 63524
rect 18972 63484 19012 63524
rect 19054 63484 19094 63524
rect 19136 63484 19176 63524
rect 18808 61972 18848 62012
rect 18890 61972 18930 62012
rect 18972 61972 19012 62012
rect 19054 61972 19094 62012
rect 19136 61972 19176 62012
rect 18808 60460 18848 60500
rect 18890 60460 18930 60500
rect 18972 60460 19012 60500
rect 19054 60460 19094 60500
rect 19136 60460 19176 60500
rect 18808 58948 18848 58988
rect 18890 58948 18930 58988
rect 18972 58948 19012 58988
rect 19054 58948 19094 58988
rect 19136 58948 19176 58988
rect 18808 57436 18848 57476
rect 18890 57436 18930 57476
rect 18972 57436 19012 57476
rect 19054 57436 19094 57476
rect 19136 57436 19176 57476
rect 18808 55924 18848 55964
rect 18890 55924 18930 55964
rect 18972 55924 19012 55964
rect 19054 55924 19094 55964
rect 19136 55924 19176 55964
rect 18808 54412 18848 54452
rect 18890 54412 18930 54452
rect 18972 54412 19012 54452
rect 19054 54412 19094 54452
rect 19136 54412 19176 54452
rect 18808 52900 18848 52940
rect 18890 52900 18930 52940
rect 18972 52900 19012 52940
rect 19054 52900 19094 52940
rect 19136 52900 19176 52940
rect 18808 51388 18848 51428
rect 18890 51388 18930 51428
rect 18972 51388 19012 51428
rect 19054 51388 19094 51428
rect 19136 51388 19176 51428
rect 18808 49876 18848 49916
rect 18890 49876 18930 49916
rect 18972 49876 19012 49916
rect 19054 49876 19094 49916
rect 19136 49876 19176 49916
rect 18808 48364 18848 48404
rect 18890 48364 18930 48404
rect 18972 48364 19012 48404
rect 19054 48364 19094 48404
rect 19136 48364 19176 48404
rect 18808 46852 18848 46892
rect 18890 46852 18930 46892
rect 18972 46852 19012 46892
rect 19054 46852 19094 46892
rect 19136 46852 19176 46892
rect 18808 45340 18848 45380
rect 18890 45340 18930 45380
rect 18972 45340 19012 45380
rect 19054 45340 19094 45380
rect 19136 45340 19176 45380
rect 18808 43828 18848 43868
rect 18890 43828 18930 43868
rect 18972 43828 19012 43868
rect 19054 43828 19094 43868
rect 19136 43828 19176 43868
rect 18808 42316 18848 42356
rect 18890 42316 18930 42356
rect 18972 42316 19012 42356
rect 19054 42316 19094 42356
rect 19136 42316 19176 42356
rect 19564 59452 19604 59492
rect 18808 40804 18848 40844
rect 18890 40804 18930 40844
rect 18972 40804 19012 40844
rect 19054 40804 19094 40844
rect 19136 40804 19176 40844
rect 18808 39292 18848 39332
rect 18890 39292 18930 39332
rect 18972 39292 19012 39332
rect 19054 39292 19094 39332
rect 19136 39292 19176 39332
rect 18808 37780 18848 37820
rect 18890 37780 18930 37820
rect 18972 37780 19012 37820
rect 19054 37780 19094 37820
rect 19136 37780 19176 37820
rect 18808 36268 18848 36308
rect 18890 36268 18930 36308
rect 18972 36268 19012 36308
rect 19054 36268 19094 36308
rect 19136 36268 19176 36308
rect 18808 34756 18848 34796
rect 18890 34756 18930 34796
rect 18972 34756 19012 34796
rect 19054 34756 19094 34796
rect 19136 34756 19176 34796
rect 18808 33244 18848 33284
rect 18890 33244 18930 33284
rect 18972 33244 19012 33284
rect 19054 33244 19094 33284
rect 19136 33244 19176 33284
rect 18808 31732 18848 31772
rect 18890 31732 18930 31772
rect 18972 31732 19012 31772
rect 19054 31732 19094 31772
rect 19136 31732 19176 31772
rect 18808 30220 18848 30260
rect 18890 30220 18930 30260
rect 18972 30220 19012 30260
rect 19054 30220 19094 30260
rect 19136 30220 19176 30260
rect 18808 28708 18848 28748
rect 18890 28708 18930 28748
rect 18972 28708 19012 28748
rect 19054 28708 19094 28748
rect 19136 28708 19176 28748
rect 18808 27196 18848 27236
rect 18890 27196 18930 27236
rect 18972 27196 19012 27236
rect 19054 27196 19094 27236
rect 19136 27196 19176 27236
rect 18808 25684 18848 25724
rect 18890 25684 18930 25724
rect 18972 25684 19012 25724
rect 19054 25684 19094 25724
rect 19136 25684 19176 25724
rect 18808 24172 18848 24212
rect 18890 24172 18930 24212
rect 18972 24172 19012 24212
rect 19054 24172 19094 24212
rect 19136 24172 19176 24212
rect 18808 22660 18848 22700
rect 18890 22660 18930 22700
rect 18972 22660 19012 22700
rect 19054 22660 19094 22700
rect 19136 22660 19176 22700
rect 18808 21148 18848 21188
rect 18890 21148 18930 21188
rect 18972 21148 19012 21188
rect 19054 21148 19094 21188
rect 19136 21148 19176 21188
rect 18808 19636 18848 19676
rect 18890 19636 18930 19676
rect 18972 19636 19012 19676
rect 19054 19636 19094 19676
rect 19136 19636 19176 19676
rect 20048 70288 20088 70328
rect 20130 70288 20170 70328
rect 20212 70288 20252 70328
rect 20294 70288 20334 70328
rect 20376 70288 20416 70328
rect 20048 68776 20088 68816
rect 20130 68776 20170 68816
rect 20212 68776 20252 68816
rect 20294 68776 20334 68816
rect 20376 68776 20416 68816
rect 19948 68608 19988 68648
rect 20620 67432 20660 67472
rect 20048 67264 20088 67304
rect 20130 67264 20170 67304
rect 20212 67264 20252 67304
rect 20294 67264 20334 67304
rect 20376 67264 20416 67304
rect 20048 65752 20088 65792
rect 20130 65752 20170 65792
rect 20212 65752 20252 65792
rect 20294 65752 20334 65792
rect 20376 65752 20416 65792
rect 20048 64240 20088 64280
rect 20130 64240 20170 64280
rect 20212 64240 20252 64280
rect 20294 64240 20334 64280
rect 20376 64240 20416 64280
rect 20048 62728 20088 62768
rect 20130 62728 20170 62768
rect 20212 62728 20252 62768
rect 20294 62728 20334 62768
rect 20376 62728 20416 62768
rect 20236 61384 20276 61424
rect 20048 61216 20088 61256
rect 20130 61216 20170 61256
rect 20212 61216 20252 61256
rect 20294 61216 20334 61256
rect 20376 61216 20416 61256
rect 20048 59704 20088 59744
rect 20130 59704 20170 59744
rect 20212 59704 20252 59744
rect 20294 59704 20334 59744
rect 20376 59704 20416 59744
rect 20048 58192 20088 58232
rect 20130 58192 20170 58232
rect 20212 58192 20252 58232
rect 20294 58192 20334 58232
rect 20376 58192 20416 58232
rect 20048 56680 20088 56720
rect 20130 56680 20170 56720
rect 20212 56680 20252 56720
rect 20294 56680 20334 56720
rect 20376 56680 20416 56720
rect 20048 55168 20088 55208
rect 20130 55168 20170 55208
rect 20212 55168 20252 55208
rect 20294 55168 20334 55208
rect 20376 55168 20416 55208
rect 20048 53656 20088 53696
rect 20130 53656 20170 53696
rect 20212 53656 20252 53696
rect 20294 53656 20334 53696
rect 20376 53656 20416 53696
rect 20048 52144 20088 52184
rect 20130 52144 20170 52184
rect 20212 52144 20252 52184
rect 20294 52144 20334 52184
rect 20376 52144 20416 52184
rect 20048 50632 20088 50672
rect 20130 50632 20170 50672
rect 20212 50632 20252 50672
rect 20294 50632 20334 50672
rect 20376 50632 20416 50672
rect 20140 49876 20180 49916
rect 20048 49120 20088 49160
rect 20130 49120 20170 49160
rect 20212 49120 20252 49160
rect 20294 49120 20334 49160
rect 20376 49120 20416 49160
rect 20048 47608 20088 47648
rect 20130 47608 20170 47648
rect 20212 47608 20252 47648
rect 20294 47608 20334 47648
rect 20376 47608 20416 47648
rect 20048 46096 20088 46136
rect 20130 46096 20170 46136
rect 20212 46096 20252 46136
rect 20294 46096 20334 46136
rect 20376 46096 20416 46136
rect 20140 44920 20180 44960
rect 20048 44584 20088 44624
rect 20130 44584 20170 44624
rect 20212 44584 20252 44624
rect 20294 44584 20334 44624
rect 20376 44584 20416 44624
rect 20048 43072 20088 43112
rect 20130 43072 20170 43112
rect 20212 43072 20252 43112
rect 20294 43072 20334 43112
rect 20376 43072 20416 43112
rect 19948 42484 19988 42524
rect 20048 41560 20088 41600
rect 20130 41560 20170 41600
rect 20212 41560 20252 41600
rect 20294 41560 20334 41600
rect 20376 41560 20416 41600
rect 20048 40048 20088 40088
rect 20130 40048 20170 40088
rect 20212 40048 20252 40088
rect 20294 40048 20334 40088
rect 20376 40048 20416 40088
rect 20048 38536 20088 38576
rect 20130 38536 20170 38576
rect 20212 38536 20252 38576
rect 20294 38536 20334 38576
rect 20376 38536 20416 38576
rect 20048 37024 20088 37064
rect 20130 37024 20170 37064
rect 20212 37024 20252 37064
rect 20294 37024 20334 37064
rect 20376 37024 20416 37064
rect 20048 35512 20088 35552
rect 20130 35512 20170 35552
rect 20212 35512 20252 35552
rect 20294 35512 20334 35552
rect 20376 35512 20416 35552
rect 20048 34000 20088 34040
rect 20130 34000 20170 34040
rect 20212 34000 20252 34040
rect 20294 34000 20334 34040
rect 20376 34000 20416 34040
rect 20048 32488 20088 32528
rect 20130 32488 20170 32528
rect 20212 32488 20252 32528
rect 20294 32488 20334 32528
rect 20376 32488 20416 32528
rect 20048 30976 20088 31016
rect 20130 30976 20170 31016
rect 20212 30976 20252 31016
rect 20294 30976 20334 31016
rect 20376 30976 20416 31016
rect 20048 29464 20088 29504
rect 20130 29464 20170 29504
rect 20212 29464 20252 29504
rect 20294 29464 20334 29504
rect 20376 29464 20416 29504
rect 20048 27952 20088 27992
rect 20130 27952 20170 27992
rect 20212 27952 20252 27992
rect 20294 27952 20334 27992
rect 20376 27952 20416 27992
rect 20048 26440 20088 26480
rect 20130 26440 20170 26480
rect 20212 26440 20252 26480
rect 20294 26440 20334 26480
rect 20376 26440 20416 26480
rect 20048 24928 20088 24968
rect 20130 24928 20170 24968
rect 20212 24928 20252 24968
rect 20294 24928 20334 24968
rect 20376 24928 20416 24968
rect 20140 23752 20180 23792
rect 20048 23416 20088 23456
rect 20130 23416 20170 23456
rect 20212 23416 20252 23456
rect 20294 23416 20334 23456
rect 20376 23416 20416 23456
rect 18808 18124 18848 18164
rect 18890 18124 18930 18164
rect 18972 18124 19012 18164
rect 19054 18124 19094 18164
rect 19136 18124 19176 18164
rect 18808 16612 18848 16652
rect 18890 16612 18930 16652
rect 18972 16612 19012 16652
rect 19054 16612 19094 16652
rect 19136 16612 19176 16652
rect 18808 15100 18848 15140
rect 18890 15100 18930 15140
rect 18972 15100 19012 15140
rect 19054 15100 19094 15140
rect 19136 15100 19176 15140
rect 18808 13588 18848 13628
rect 18890 13588 18930 13628
rect 18972 13588 19012 13628
rect 19054 13588 19094 13628
rect 19136 13588 19176 13628
rect 20140 22408 20180 22448
rect 20048 21904 20088 21944
rect 20130 21904 20170 21944
rect 20212 21904 20252 21944
rect 20294 21904 20334 21944
rect 20376 21904 20416 21944
rect 20140 21736 20180 21776
rect 20048 20392 20088 20432
rect 20130 20392 20170 20432
rect 20212 20392 20252 20432
rect 20294 20392 20334 20432
rect 20376 20392 20416 20432
rect 20048 18880 20088 18920
rect 20130 18880 20170 18920
rect 20212 18880 20252 18920
rect 20294 18880 20334 18920
rect 20376 18880 20416 18920
rect 20048 17368 20088 17408
rect 20130 17368 20170 17408
rect 20212 17368 20252 17408
rect 20294 17368 20334 17408
rect 20376 17368 20416 17408
rect 20048 15856 20088 15896
rect 20130 15856 20170 15896
rect 20212 15856 20252 15896
rect 20294 15856 20334 15896
rect 20376 15856 20416 15896
rect 20048 14344 20088 14384
rect 20130 14344 20170 14384
rect 20212 14344 20252 14384
rect 20294 14344 20334 14384
rect 20376 14344 20416 14384
rect 20048 12832 20088 12872
rect 20130 12832 20170 12872
rect 20212 12832 20252 12872
rect 20294 12832 20334 12872
rect 20376 12832 20416 12872
rect 18808 12076 18848 12116
rect 18890 12076 18930 12116
rect 18972 12076 19012 12116
rect 19054 12076 19094 12116
rect 19136 12076 19176 12116
rect 18808 10564 18848 10604
rect 18890 10564 18930 10604
rect 18972 10564 19012 10604
rect 19054 10564 19094 10604
rect 19136 10564 19176 10604
rect 18808 9052 18848 9092
rect 18890 9052 18930 9092
rect 18972 9052 19012 9092
rect 19054 9052 19094 9092
rect 19136 9052 19176 9092
rect 20048 11320 20088 11360
rect 20130 11320 20170 11360
rect 20212 11320 20252 11360
rect 20294 11320 20334 11360
rect 20376 11320 20416 11360
rect 20048 9808 20088 9848
rect 20130 9808 20170 9848
rect 20212 9808 20252 9848
rect 20294 9808 20334 9848
rect 20376 9808 20416 9848
rect 20048 8296 20088 8336
rect 20130 8296 20170 8336
rect 20212 8296 20252 8336
rect 20294 8296 20334 8336
rect 20376 8296 20416 8336
rect 18808 7540 18848 7580
rect 18890 7540 18930 7580
rect 18972 7540 19012 7580
rect 19054 7540 19094 7580
rect 19136 7540 19176 7580
rect 18808 6028 18848 6068
rect 18890 6028 18930 6068
rect 18972 6028 19012 6068
rect 19054 6028 19094 6068
rect 19136 6028 19176 6068
rect 20048 6784 20088 6824
rect 20130 6784 20170 6824
rect 20212 6784 20252 6824
rect 20294 6784 20334 6824
rect 20376 6784 20416 6824
rect 20048 5272 20088 5312
rect 20130 5272 20170 5312
rect 20212 5272 20252 5312
rect 20294 5272 20334 5312
rect 20376 5272 20416 5312
rect 18808 4516 18848 4556
rect 18890 4516 18930 4556
rect 18972 4516 19012 4556
rect 19054 4516 19094 4556
rect 19136 4516 19176 4556
rect 20048 3760 20088 3800
rect 20130 3760 20170 3800
rect 20212 3760 20252 3800
rect 20294 3760 20334 3800
rect 20376 3760 20416 3800
rect 18808 3004 18848 3044
rect 18890 3004 18930 3044
rect 18972 3004 19012 3044
rect 19054 3004 19094 3044
rect 19136 3004 19176 3044
rect 20048 2248 20088 2288
rect 20130 2248 20170 2288
rect 20212 2248 20252 2288
rect 20294 2248 20334 2288
rect 20376 2248 20416 2288
rect 18808 1492 18848 1532
rect 18890 1492 18930 1532
rect 18972 1492 19012 1532
rect 19054 1492 19094 1532
rect 19136 1492 19176 1532
rect 20908 63652 20948 63692
rect 20716 32068 20756 32108
rect 20620 26608 20660 26648
rect 20620 24592 20660 24632
rect 20812 24508 20852 24548
rect 20048 736 20088 776
rect 20130 736 20170 776
rect 20212 736 20252 776
rect 20294 736 20334 776
rect 20376 736 20416 776
rect 18892 652 18932 692
rect 19468 148 19508 188
<< metal5 >>
rect 3679 84715 4065 84734
rect 3679 84692 3745 84715
rect 3831 84692 3913 84715
rect 3999 84692 4065 84715
rect 3679 84652 3688 84692
rect 3728 84652 3745 84692
rect 3831 84652 3852 84692
rect 3892 84652 3913 84692
rect 3999 84652 4016 84692
rect 4056 84652 4065 84692
rect 3679 84629 3745 84652
rect 3831 84629 3913 84652
rect 3999 84629 4065 84652
rect 3679 84610 4065 84629
rect 18799 84715 19185 84734
rect 18799 84692 18865 84715
rect 18951 84692 19033 84715
rect 19119 84692 19185 84715
rect 18799 84652 18808 84692
rect 18848 84652 18865 84692
rect 18951 84652 18972 84692
rect 19012 84652 19033 84692
rect 19119 84652 19136 84692
rect 19176 84652 19185 84692
rect 18799 84629 18865 84652
rect 18951 84629 19033 84652
rect 19119 84629 19185 84652
rect 18799 84610 19185 84629
rect 1315 84316 1324 84356
rect 1364 84316 4684 84356
rect 4724 84316 4733 84356
rect 12122 84127 12246 84146
rect 12122 84041 12141 84127
rect 12227 84104 12246 84127
rect 12227 84064 12460 84104
rect 12500 84064 12509 84104
rect 12227 84041 12246 84064
rect 12122 84022 12246 84041
rect 4919 83959 5305 83978
rect 4919 83936 4985 83959
rect 5071 83936 5153 83959
rect 5239 83936 5305 83959
rect 4919 83896 4928 83936
rect 4968 83896 4985 83936
rect 5071 83896 5092 83936
rect 5132 83896 5153 83936
rect 5239 83896 5256 83936
rect 5296 83896 5305 83936
rect 4919 83873 4985 83896
rect 5071 83873 5153 83896
rect 5239 83873 5305 83896
rect 4919 83854 5305 83873
rect 20039 83959 20425 83978
rect 20039 83936 20105 83959
rect 20191 83936 20273 83959
rect 20359 83936 20425 83959
rect 20039 83896 20048 83936
rect 20088 83896 20105 83936
rect 20191 83896 20212 83936
rect 20252 83896 20273 83936
rect 20359 83896 20376 83936
rect 20416 83896 20425 83936
rect 20039 83873 20105 83896
rect 20191 83873 20273 83896
rect 20359 83873 20425 83896
rect 20039 83854 20425 83873
rect 10754 83539 10878 83558
rect 10754 83516 10773 83539
rect 10531 83476 10540 83516
rect 10580 83476 10773 83516
rect 10754 83453 10773 83476
rect 10859 83453 10878 83539
rect 10754 83434 10878 83453
rect 13034 83371 13158 83390
rect 13034 83285 13053 83371
rect 13139 83348 13158 83371
rect 13139 83308 13612 83348
rect 13652 83308 13661 83348
rect 13139 83285 13158 83308
rect 13034 83266 13158 83285
rect 3679 83203 4065 83222
rect 3679 83180 3745 83203
rect 3831 83180 3913 83203
rect 3999 83180 4065 83203
rect 18799 83203 19185 83222
rect 18799 83180 18865 83203
rect 18951 83180 19033 83203
rect 19119 83180 19185 83203
rect 3679 83140 3688 83180
rect 3728 83140 3745 83180
rect 3831 83140 3852 83180
rect 3892 83140 3913 83180
rect 3999 83140 4016 83180
rect 4056 83140 4065 83180
rect 9955 83140 9964 83180
rect 10004 83140 16012 83180
rect 16052 83140 16061 83180
rect 18799 83140 18808 83180
rect 18848 83140 18865 83180
rect 18951 83140 18972 83180
rect 19012 83140 19033 83180
rect 19119 83140 19136 83180
rect 19176 83140 19185 83180
rect 3679 83117 3745 83140
rect 3831 83117 3913 83140
rect 3999 83117 4065 83140
rect 3679 83098 4065 83117
rect 18799 83117 18865 83140
rect 18951 83117 19033 83140
rect 19119 83117 19185 83140
rect 18799 83098 19185 83117
rect 5443 82804 5452 82844
rect 5492 82804 8140 82844
rect 8180 82804 8189 82844
rect 4919 82447 5305 82466
rect 4919 82424 4985 82447
rect 5071 82424 5153 82447
rect 5239 82424 5305 82447
rect 4919 82384 4928 82424
rect 4968 82384 4985 82424
rect 5071 82384 5092 82424
rect 5132 82384 5153 82424
rect 5239 82384 5256 82424
rect 5296 82384 5305 82424
rect 4919 82361 4985 82384
rect 5071 82361 5153 82384
rect 5239 82361 5305 82384
rect 4919 82342 5305 82361
rect 20039 82447 20425 82466
rect 20039 82424 20105 82447
rect 20191 82424 20273 82447
rect 20359 82424 20425 82447
rect 20039 82384 20048 82424
rect 20088 82384 20105 82424
rect 20191 82384 20212 82424
rect 20252 82384 20273 82424
rect 20359 82384 20376 82424
rect 20416 82384 20425 82424
rect 20039 82361 20105 82384
rect 20191 82361 20273 82384
rect 20359 82361 20425 82384
rect 20039 82342 20425 82361
rect 8060 82048 10060 82088
rect 10100 82048 10109 82088
rect 8060 82004 8100 82048
rect 3811 81964 3820 82004
rect 3860 81964 8100 82004
rect 3679 81691 4065 81710
rect 3679 81668 3745 81691
rect 3831 81668 3913 81691
rect 3999 81668 4065 81691
rect 3679 81628 3688 81668
rect 3728 81628 3745 81668
rect 3831 81628 3852 81668
rect 3892 81628 3913 81668
rect 3999 81628 4016 81668
rect 4056 81628 4065 81668
rect 3679 81605 3745 81628
rect 3831 81605 3913 81628
rect 3999 81605 4065 81628
rect 3679 81586 4065 81605
rect 18799 81691 19185 81710
rect 18799 81668 18865 81691
rect 18951 81668 19033 81691
rect 19119 81668 19185 81691
rect 18799 81628 18808 81668
rect 18848 81628 18865 81668
rect 18951 81628 18972 81668
rect 19012 81628 19033 81668
rect 19119 81628 19136 81668
rect 19176 81628 19185 81668
rect 18799 81605 18865 81628
rect 18951 81605 19033 81628
rect 19119 81605 19185 81628
rect 18799 81586 19185 81605
rect 16682 81103 16806 81122
rect 16682 81080 16701 81103
rect 16387 81040 16396 81080
rect 16436 81040 16701 81080
rect 16682 81017 16701 81040
rect 16787 81017 16806 81103
rect 16682 80998 16806 81017
rect 4919 80935 5305 80954
rect 4919 80912 4985 80935
rect 5071 80912 5153 80935
rect 5239 80912 5305 80935
rect 4919 80872 4928 80912
rect 4968 80872 4985 80912
rect 5071 80872 5092 80912
rect 5132 80872 5153 80912
rect 5239 80872 5256 80912
rect 5296 80872 5305 80912
rect 4919 80849 4985 80872
rect 5071 80849 5153 80872
rect 5239 80849 5305 80872
rect 20039 80935 20425 80954
rect 20039 80912 20105 80935
rect 20191 80912 20273 80935
rect 20359 80912 20425 80935
rect 20039 80872 20048 80912
rect 20088 80872 20105 80912
rect 20191 80872 20212 80912
rect 20252 80872 20273 80912
rect 20359 80872 20376 80912
rect 20416 80872 20425 80912
rect 4919 80830 5305 80849
rect 8474 80851 8598 80870
rect 8474 80828 8493 80851
rect 7459 80788 7468 80828
rect 7508 80788 8493 80828
rect 8474 80765 8493 80788
rect 8579 80765 8598 80851
rect 20039 80849 20105 80872
rect 20191 80849 20273 80872
rect 20359 80849 20425 80872
rect 20039 80830 20425 80849
rect 8474 80746 8598 80765
rect 3043 80620 3052 80660
rect 3092 80620 3916 80660
rect 3956 80620 6988 80660
rect 7028 80620 7037 80660
rect 3679 80179 4065 80198
rect 3679 80156 3745 80179
rect 3831 80156 3913 80179
rect 3999 80156 4065 80179
rect 3679 80116 3688 80156
rect 3728 80116 3745 80156
rect 3831 80116 3852 80156
rect 3892 80116 3913 80156
rect 3999 80116 4016 80156
rect 4056 80116 4065 80156
rect 3679 80093 3745 80116
rect 3831 80093 3913 80116
rect 3999 80093 4065 80116
rect 3679 80074 4065 80093
rect 18799 80179 19185 80198
rect 18799 80156 18865 80179
rect 18951 80156 19033 80179
rect 19119 80156 19185 80179
rect 18799 80116 18808 80156
rect 18848 80116 18865 80156
rect 18951 80116 18972 80156
rect 19012 80116 19033 80156
rect 19119 80116 19136 80156
rect 19176 80116 19185 80156
rect 18799 80093 18865 80116
rect 18951 80093 19033 80116
rect 19119 80093 19185 80116
rect 18799 80074 19185 80093
rect 9842 79507 9966 79526
rect 9842 79484 9861 79507
rect 7747 79444 7756 79484
rect 7796 79444 9861 79484
rect 4919 79423 5305 79442
rect 4919 79400 4985 79423
rect 5071 79400 5153 79423
rect 5239 79400 5305 79423
rect 9842 79421 9861 79444
rect 9947 79421 9966 79507
rect 9842 79402 9966 79421
rect 20039 79423 20425 79442
rect 4919 79360 4928 79400
rect 4968 79360 4985 79400
rect 5071 79360 5092 79400
rect 5132 79360 5153 79400
rect 5239 79360 5256 79400
rect 5296 79360 5305 79400
rect 4919 79337 4985 79360
rect 5071 79337 5153 79360
rect 5239 79337 5305 79360
rect 4919 79318 5305 79337
rect 20039 79400 20105 79423
rect 20191 79400 20273 79423
rect 20359 79400 20425 79423
rect 20039 79360 20048 79400
rect 20088 79360 20105 79400
rect 20191 79360 20212 79400
rect 20252 79360 20273 79400
rect 20359 79360 20376 79400
rect 20416 79360 20425 79400
rect 20039 79337 20105 79360
rect 20191 79337 20273 79360
rect 20359 79337 20425 79360
rect 20039 79318 20425 79337
rect 3679 78667 4065 78686
rect 3679 78644 3745 78667
rect 3831 78644 3913 78667
rect 3999 78644 4065 78667
rect 3679 78604 3688 78644
rect 3728 78604 3745 78644
rect 3831 78604 3852 78644
rect 3892 78604 3913 78644
rect 3999 78604 4016 78644
rect 4056 78604 4065 78644
rect 3679 78581 3745 78604
rect 3831 78581 3913 78604
rect 3999 78581 4065 78604
rect 3679 78562 4065 78581
rect 18799 78667 19185 78686
rect 18799 78644 18865 78667
rect 18951 78644 19033 78667
rect 19119 78644 19185 78667
rect 18799 78604 18808 78644
rect 18848 78604 18865 78644
rect 18951 78604 18972 78644
rect 19012 78604 19033 78644
rect 19119 78604 19136 78644
rect 19176 78604 19185 78644
rect 18799 78581 18865 78604
rect 18951 78581 19033 78604
rect 19119 78581 19185 78604
rect 18799 78562 19185 78581
rect 11107 78100 11116 78140
rect 11156 78100 18028 78140
rect 18068 78100 18077 78140
rect 4919 77911 5305 77930
rect 4919 77888 4985 77911
rect 5071 77888 5153 77911
rect 5239 77888 5305 77911
rect 4919 77848 4928 77888
rect 4968 77848 4985 77888
rect 5071 77848 5092 77888
rect 5132 77848 5153 77888
rect 5239 77848 5256 77888
rect 5296 77848 5305 77888
rect 4919 77825 4985 77848
rect 5071 77825 5153 77848
rect 5239 77825 5305 77848
rect 4919 77806 5305 77825
rect 20039 77911 20425 77930
rect 20039 77888 20105 77911
rect 20191 77888 20273 77911
rect 20359 77888 20425 77911
rect 20039 77848 20048 77888
rect 20088 77848 20105 77888
rect 20191 77848 20212 77888
rect 20252 77848 20273 77888
rect 20359 77848 20376 77888
rect 20416 77848 20425 77888
rect 20039 77825 20105 77848
rect 20191 77825 20273 77848
rect 20359 77825 20425 77848
rect 20039 77806 20425 77825
rect 13946 77323 14070 77342
rect 13946 77237 13965 77323
rect 14051 77300 14070 77323
rect 14051 77260 15052 77300
rect 15092 77260 15101 77300
rect 14051 77237 14070 77260
rect 13946 77218 14070 77237
rect 3679 77155 4065 77174
rect 3679 77132 3745 77155
rect 3831 77132 3913 77155
rect 3999 77132 4065 77155
rect 3679 77092 3688 77132
rect 3728 77092 3745 77132
rect 3831 77092 3852 77132
rect 3892 77092 3913 77132
rect 3999 77092 4016 77132
rect 4056 77092 4065 77132
rect 3679 77069 3745 77092
rect 3831 77069 3913 77092
rect 3999 77069 4065 77092
rect 3679 77050 4065 77069
rect 18799 77155 19185 77174
rect 18799 77132 18865 77155
rect 18951 77132 19033 77155
rect 19119 77132 19185 77155
rect 18799 77092 18808 77132
rect 18848 77092 18865 77132
rect 18951 77092 18972 77132
rect 19012 77092 19033 77132
rect 19119 77092 19136 77132
rect 19176 77092 19185 77132
rect 18799 77069 18865 77092
rect 18951 77069 19033 77092
rect 19119 77069 19185 77092
rect 18799 77050 19185 77069
rect 2090 76903 2214 76922
rect 2090 76817 2109 76903
rect 2195 76880 2214 76903
rect 2195 76840 6412 76880
rect 6452 76840 6461 76880
rect 2195 76817 2214 76840
rect 2090 76798 2214 76817
rect 4919 76399 5305 76418
rect 4919 76376 4985 76399
rect 5071 76376 5153 76399
rect 5239 76376 5305 76399
rect 4919 76336 4928 76376
rect 4968 76336 4985 76376
rect 5071 76336 5092 76376
rect 5132 76336 5153 76376
rect 5239 76336 5256 76376
rect 5296 76336 5305 76376
rect 4919 76313 4985 76336
rect 5071 76313 5153 76336
rect 5239 76313 5305 76336
rect 4919 76294 5305 76313
rect 20039 76399 20425 76418
rect 20039 76376 20105 76399
rect 20191 76376 20273 76399
rect 20359 76376 20425 76399
rect 20039 76336 20048 76376
rect 20088 76336 20105 76376
rect 20191 76336 20212 76376
rect 20252 76336 20273 76376
rect 20359 76336 20376 76376
rect 20416 76336 20425 76376
rect 20039 76313 20105 76336
rect 20191 76313 20273 76336
rect 20359 76313 20425 76336
rect 20039 76294 20425 76313
rect 547 75832 556 75872
rect 596 75832 6700 75872
rect 6740 75832 6749 75872
rect 3679 75643 4065 75662
rect 3679 75620 3745 75643
rect 3831 75620 3913 75643
rect 3999 75620 4065 75643
rect 3679 75580 3688 75620
rect 3728 75580 3745 75620
rect 3831 75580 3852 75620
rect 3892 75580 3913 75620
rect 3999 75580 4016 75620
rect 4056 75580 4065 75620
rect 3679 75557 3745 75580
rect 3831 75557 3913 75580
rect 3999 75557 4065 75580
rect 3679 75538 4065 75557
rect 18799 75643 19185 75662
rect 18799 75620 18865 75643
rect 18951 75620 19033 75643
rect 19119 75620 19185 75643
rect 18799 75580 18808 75620
rect 18848 75580 18865 75620
rect 18951 75580 18972 75620
rect 19012 75580 19033 75620
rect 19119 75580 19136 75620
rect 19176 75580 19185 75620
rect 18799 75557 18865 75580
rect 18951 75557 19033 75580
rect 19119 75557 19185 75580
rect 18799 75538 19185 75557
rect 1411 74992 1420 75032
rect 1460 74992 5548 75032
rect 5588 74992 5597 75032
rect 4919 74887 5305 74906
rect 4919 74864 4985 74887
rect 5071 74864 5153 74887
rect 5239 74864 5305 74887
rect 4919 74824 4928 74864
rect 4968 74824 4985 74864
rect 5071 74824 5092 74864
rect 5132 74824 5153 74864
rect 5239 74824 5256 74864
rect 5296 74824 5305 74864
rect 4919 74801 4985 74824
rect 5071 74801 5153 74824
rect 5239 74801 5305 74824
rect 4919 74782 5305 74801
rect 20039 74887 20425 74906
rect 20039 74864 20105 74887
rect 20191 74864 20273 74887
rect 20359 74864 20425 74887
rect 20039 74824 20048 74864
rect 20088 74824 20105 74864
rect 20191 74824 20212 74864
rect 20252 74824 20273 74864
rect 20359 74824 20376 74864
rect 20416 74824 20425 74864
rect 20039 74801 20105 74824
rect 20191 74801 20273 74824
rect 20359 74801 20425 74824
rect 20039 74782 20425 74801
rect 3679 74131 4065 74150
rect 3679 74108 3745 74131
rect 3831 74108 3913 74131
rect 3999 74108 4065 74131
rect 3679 74068 3688 74108
rect 3728 74068 3745 74108
rect 3831 74068 3852 74108
rect 3892 74068 3913 74108
rect 3999 74068 4016 74108
rect 4056 74068 4065 74108
rect 3679 74045 3745 74068
rect 3831 74045 3913 74068
rect 3999 74045 4065 74068
rect 3679 74026 4065 74045
rect 18799 74131 19185 74150
rect 18799 74108 18865 74131
rect 18951 74108 19033 74131
rect 19119 74108 19185 74131
rect 18799 74068 18808 74108
rect 18848 74068 18865 74108
rect 18951 74068 18972 74108
rect 19012 74068 19033 74108
rect 19119 74068 19136 74108
rect 19176 74068 19185 74108
rect 18799 74045 18865 74068
rect 18951 74045 19033 74068
rect 19119 74045 19185 74068
rect 18799 74026 19185 74045
rect 4919 73375 5305 73394
rect 4919 73352 4985 73375
rect 5071 73352 5153 73375
rect 5239 73352 5305 73375
rect 4919 73312 4928 73352
rect 4968 73312 4985 73352
rect 5071 73312 5092 73352
rect 5132 73312 5153 73352
rect 5239 73312 5256 73352
rect 5296 73312 5305 73352
rect 4919 73289 4985 73312
rect 5071 73289 5153 73312
rect 5239 73289 5305 73312
rect 4919 73270 5305 73289
rect 20039 73375 20425 73394
rect 20039 73352 20105 73375
rect 20191 73352 20273 73375
rect 20359 73352 20425 73375
rect 20039 73312 20048 73352
rect 20088 73312 20105 73352
rect 20191 73312 20212 73352
rect 20252 73312 20273 73352
rect 20359 73312 20376 73352
rect 20416 73312 20425 73352
rect 20039 73289 20105 73312
rect 20191 73289 20273 73312
rect 20359 73289 20425 73312
rect 20039 73270 20425 73289
rect 547 73144 556 73184
rect 596 73144 804 73184
rect 764 73100 804 73144
rect 764 73060 844 73100
rect 884 73060 893 73100
rect 7604 73060 7660 73100
rect 7700 73060 7709 73100
rect 1178 73039 1302 73058
rect 1178 72953 1197 73039
rect 1283 73016 1302 73039
rect 7604 73016 7644 73060
rect 1283 72976 7644 73016
rect 1283 72953 1302 72976
rect 1178 72934 1302 72953
rect 3679 72619 4065 72638
rect 3679 72596 3745 72619
rect 3831 72596 3913 72619
rect 3999 72596 4065 72619
rect 3679 72556 3688 72596
rect 3728 72556 3745 72596
rect 3831 72556 3852 72596
rect 3892 72556 3913 72596
rect 3999 72556 4016 72596
rect 4056 72556 4065 72596
rect 3679 72533 3745 72556
rect 3831 72533 3913 72556
rect 3999 72533 4065 72556
rect 3679 72514 4065 72533
rect 18799 72619 19185 72638
rect 18799 72596 18865 72619
rect 18951 72596 19033 72619
rect 19119 72596 19185 72619
rect 18799 72556 18808 72596
rect 18848 72556 18865 72596
rect 18951 72556 18972 72596
rect 19012 72556 19033 72596
rect 19119 72556 19136 72596
rect 19176 72556 19185 72596
rect 18799 72533 18865 72556
rect 18951 72533 19033 72556
rect 19119 72533 19185 72556
rect 18799 72514 19185 72533
rect 4919 71863 5305 71882
rect 4919 71840 4985 71863
rect 5071 71840 5153 71863
rect 5239 71840 5305 71863
rect 4919 71800 4928 71840
rect 4968 71800 4985 71840
rect 5071 71800 5092 71840
rect 5132 71800 5153 71840
rect 5239 71800 5256 71840
rect 5296 71800 5305 71840
rect 4919 71777 4985 71800
rect 5071 71777 5153 71800
rect 5239 71777 5305 71800
rect 4919 71758 5305 71777
rect 20039 71863 20425 71882
rect 20039 71840 20105 71863
rect 20191 71840 20273 71863
rect 20359 71840 20425 71863
rect 20039 71800 20048 71840
rect 20088 71800 20105 71840
rect 20191 71800 20212 71840
rect 20252 71800 20273 71840
rect 20359 71800 20376 71840
rect 20416 71800 20425 71840
rect 20039 71777 20105 71800
rect 20191 71777 20273 71800
rect 20359 71777 20425 71800
rect 20039 71758 20425 71777
rect 3679 71107 4065 71126
rect 3679 71084 3745 71107
rect 3831 71084 3913 71107
rect 3999 71084 4065 71107
rect 3679 71044 3688 71084
rect 3728 71044 3745 71084
rect 3831 71044 3852 71084
rect 3892 71044 3913 71084
rect 3999 71044 4016 71084
rect 4056 71044 4065 71084
rect 3679 71021 3745 71044
rect 3831 71021 3913 71044
rect 3999 71021 4065 71044
rect 3679 71002 4065 71021
rect 18799 71107 19185 71126
rect 18799 71084 18865 71107
rect 18951 71084 19033 71107
rect 19119 71084 19185 71107
rect 18799 71044 18808 71084
rect 18848 71044 18865 71084
rect 18951 71044 18972 71084
rect 19012 71044 19033 71084
rect 19119 71044 19136 71084
rect 19176 71044 19185 71084
rect 18799 71021 18865 71044
rect 18951 71021 19033 71044
rect 19119 71021 19185 71044
rect 18799 71002 19185 71021
rect 4919 70351 5305 70370
rect 4919 70328 4985 70351
rect 5071 70328 5153 70351
rect 5239 70328 5305 70351
rect 4919 70288 4928 70328
rect 4968 70288 4985 70328
rect 5071 70288 5092 70328
rect 5132 70288 5153 70328
rect 5239 70288 5256 70328
rect 5296 70288 5305 70328
rect 4919 70265 4985 70288
rect 5071 70265 5153 70288
rect 5239 70265 5305 70288
rect 4919 70246 5305 70265
rect 20039 70351 20425 70370
rect 20039 70328 20105 70351
rect 20191 70328 20273 70351
rect 20359 70328 20425 70351
rect 20039 70288 20048 70328
rect 20088 70288 20105 70328
rect 20191 70288 20212 70328
rect 20252 70288 20273 70328
rect 20359 70288 20376 70328
rect 20416 70288 20425 70328
rect 20039 70265 20105 70288
rect 20191 70265 20273 70288
rect 20359 70265 20425 70288
rect 20039 70246 20425 70265
rect 3679 69595 4065 69614
rect 3679 69572 3745 69595
rect 3831 69572 3913 69595
rect 3999 69572 4065 69595
rect 3679 69532 3688 69572
rect 3728 69532 3745 69572
rect 3831 69532 3852 69572
rect 3892 69532 3913 69572
rect 3999 69532 4016 69572
rect 4056 69532 4065 69572
rect 3679 69509 3745 69532
rect 3831 69509 3913 69532
rect 3999 69509 4065 69532
rect 3679 69490 4065 69509
rect 18799 69595 19185 69614
rect 18799 69572 18865 69595
rect 18951 69572 19033 69595
rect 19119 69572 19185 69595
rect 18799 69532 18808 69572
rect 18848 69532 18865 69572
rect 18951 69532 18972 69572
rect 19012 69532 19033 69572
rect 19119 69532 19136 69572
rect 19176 69532 19185 69572
rect 18799 69509 18865 69532
rect 18951 69509 19033 69532
rect 19119 69509 19185 69532
rect 18799 69490 19185 69509
rect 14467 69028 14476 69068
rect 14516 69028 14860 69068
rect 14900 69028 14909 69068
rect 14755 68944 14764 68984
rect 14804 68944 14956 68984
rect 14996 68944 15005 68984
rect 4919 68839 5305 68858
rect 4919 68816 4985 68839
rect 5071 68816 5153 68839
rect 5239 68816 5305 68839
rect 4919 68776 4928 68816
rect 4968 68776 4985 68816
rect 5071 68776 5092 68816
rect 5132 68776 5153 68816
rect 5239 68776 5256 68816
rect 5296 68776 5305 68816
rect 4919 68753 4985 68776
rect 5071 68753 5153 68776
rect 5239 68753 5305 68776
rect 4919 68734 5305 68753
rect 20039 68839 20425 68858
rect 20039 68816 20105 68839
rect 20191 68816 20273 68839
rect 20359 68816 20425 68839
rect 20039 68776 20048 68816
rect 20088 68776 20105 68816
rect 20191 68776 20212 68816
rect 20252 68776 20273 68816
rect 20359 68776 20376 68816
rect 20416 68776 20425 68816
rect 20039 68753 20105 68776
rect 20191 68753 20273 68776
rect 20359 68753 20425 68776
rect 20039 68734 20425 68753
rect 9763 68608 9772 68648
rect 9812 68608 19948 68648
rect 19988 68608 19997 68648
rect 3679 68083 4065 68102
rect 3679 68060 3745 68083
rect 3831 68060 3913 68083
rect 3999 68060 4065 68083
rect 3679 68020 3688 68060
rect 3728 68020 3745 68060
rect 3831 68020 3852 68060
rect 3892 68020 3913 68060
rect 3999 68020 4016 68060
rect 4056 68020 4065 68060
rect 3679 67997 3745 68020
rect 3831 67997 3913 68020
rect 3999 67997 4065 68020
rect 3679 67978 4065 67997
rect 18799 68083 19185 68102
rect 18799 68060 18865 68083
rect 18951 68060 19033 68083
rect 19119 68060 19185 68083
rect 18799 68020 18808 68060
rect 18848 68020 18865 68060
rect 18951 68020 18972 68060
rect 19012 68020 19033 68060
rect 19119 68020 19136 68060
rect 19176 68020 19185 68060
rect 18799 67997 18865 68020
rect 18951 67997 19033 68020
rect 19119 67997 19185 68020
rect 18799 67978 19185 67997
rect 5155 67768 5164 67808
rect 5204 67768 5356 67808
rect 5396 67768 9676 67808
rect 9716 67768 9725 67808
rect 6211 67432 6220 67472
rect 6260 67432 20620 67472
rect 20660 67432 20669 67472
rect 4919 67327 5305 67346
rect 4919 67304 4985 67327
rect 5071 67304 5153 67327
rect 5239 67304 5305 67327
rect 4919 67264 4928 67304
rect 4968 67264 4985 67304
rect 5071 67264 5092 67304
rect 5132 67264 5153 67304
rect 5239 67264 5256 67304
rect 5296 67264 5305 67304
rect 4919 67241 4985 67264
rect 5071 67241 5153 67264
rect 5239 67241 5305 67264
rect 4919 67222 5305 67241
rect 20039 67327 20425 67346
rect 20039 67304 20105 67327
rect 20191 67304 20273 67327
rect 20359 67304 20425 67327
rect 20039 67264 20048 67304
rect 20088 67264 20105 67304
rect 20191 67264 20212 67304
rect 20252 67264 20273 67304
rect 20359 67264 20376 67304
rect 20416 67264 20425 67304
rect 20039 67241 20105 67264
rect 20191 67241 20273 67264
rect 20359 67241 20425 67264
rect 20039 67222 20425 67241
rect 15770 66991 15894 67010
rect 15770 66905 15789 66991
rect 15875 66968 15894 66991
rect 15875 66928 16684 66968
rect 16724 66928 16733 66968
rect 15875 66905 15894 66928
rect 15770 66886 15894 66905
rect 3679 66571 4065 66590
rect 3679 66548 3745 66571
rect 3831 66548 3913 66571
rect 3999 66548 4065 66571
rect 3679 66508 3688 66548
rect 3728 66508 3745 66548
rect 3831 66508 3852 66548
rect 3892 66508 3913 66548
rect 3999 66508 4016 66548
rect 4056 66508 4065 66548
rect 3679 66485 3745 66508
rect 3831 66485 3913 66508
rect 3999 66485 4065 66508
rect 3679 66466 4065 66485
rect 18799 66571 19185 66590
rect 18799 66548 18865 66571
rect 18951 66548 19033 66571
rect 19119 66548 19185 66571
rect 18799 66508 18808 66548
rect 18848 66508 18865 66548
rect 18951 66508 18972 66548
rect 19012 66508 19033 66548
rect 19119 66508 19136 66548
rect 19176 66508 19185 66548
rect 18799 66485 18865 66508
rect 18951 66485 19033 66508
rect 19119 66485 19185 66508
rect 18799 66466 19185 66485
rect 6650 65899 6774 65918
rect 4919 65815 5305 65834
rect 4919 65792 4985 65815
rect 5071 65792 5153 65815
rect 5239 65792 5305 65815
rect 6650 65813 6669 65899
rect 6755 65876 6774 65899
rect 6755 65836 8524 65876
rect 8564 65836 8573 65876
rect 6755 65813 6774 65836
rect 6650 65794 6774 65813
rect 20039 65815 20425 65834
rect 4919 65752 4928 65792
rect 4968 65752 4985 65792
rect 5071 65752 5092 65792
rect 5132 65752 5153 65792
rect 5239 65752 5256 65792
rect 5296 65752 5305 65792
rect 4919 65729 4985 65752
rect 5071 65729 5153 65752
rect 5239 65729 5305 65752
rect 4919 65710 5305 65729
rect 20039 65792 20105 65815
rect 20191 65792 20273 65815
rect 20359 65792 20425 65815
rect 20039 65752 20048 65792
rect 20088 65752 20105 65792
rect 20191 65752 20212 65792
rect 20252 65752 20273 65792
rect 20359 65752 20376 65792
rect 20416 65752 20425 65792
rect 20039 65729 20105 65752
rect 20191 65729 20273 65752
rect 20359 65729 20425 65752
rect 20039 65710 20425 65729
rect 3679 65059 4065 65078
rect 3679 65036 3745 65059
rect 3831 65036 3913 65059
rect 3999 65036 4065 65059
rect 3679 64996 3688 65036
rect 3728 64996 3745 65036
rect 3831 64996 3852 65036
rect 3892 64996 3913 65036
rect 3999 64996 4016 65036
rect 4056 64996 4065 65036
rect 3679 64973 3745 64996
rect 3831 64973 3913 64996
rect 3999 64973 4065 64996
rect 3679 64954 4065 64973
rect 18799 65059 19185 65078
rect 18799 65036 18865 65059
rect 18951 65036 19033 65059
rect 19119 65036 19185 65059
rect 18799 64996 18808 65036
rect 18848 64996 18865 65036
rect 18951 64996 18972 65036
rect 19012 64996 19033 65036
rect 19119 64996 19136 65036
rect 19176 64996 19185 65036
rect 18799 64973 18865 64996
rect 18951 64973 19033 64996
rect 19119 64973 19185 64996
rect 18799 64954 19185 64973
rect 8419 64828 8428 64868
rect 8468 64828 19276 64868
rect 19316 64828 19325 64868
rect 14275 64744 14284 64784
rect 14324 64744 14572 64784
rect 14612 64744 14621 64784
rect 9859 64408 9868 64448
rect 9908 64408 19276 64448
rect 19316 64408 19325 64448
rect 4919 64303 5305 64322
rect 4919 64280 4985 64303
rect 5071 64280 5153 64303
rect 5239 64280 5305 64303
rect 4919 64240 4928 64280
rect 4968 64240 4985 64280
rect 5071 64240 5092 64280
rect 5132 64240 5153 64280
rect 5239 64240 5256 64280
rect 5296 64240 5305 64280
rect 4919 64217 4985 64240
rect 5071 64217 5153 64240
rect 5239 64217 5305 64240
rect 4919 64198 5305 64217
rect 20039 64303 20425 64322
rect 20039 64280 20105 64303
rect 20191 64280 20273 64303
rect 20359 64280 20425 64303
rect 20039 64240 20048 64280
rect 20088 64240 20105 64280
rect 20191 64240 20212 64280
rect 20252 64240 20273 64280
rect 20359 64240 20376 64280
rect 20416 64240 20425 64280
rect 20039 64217 20105 64240
rect 20191 64217 20273 64240
rect 20359 64217 20425 64240
rect 20039 64198 20425 64217
rect 12355 63652 12364 63692
rect 12404 63652 20908 63692
rect 20948 63652 20957 63692
rect 3679 63547 4065 63566
rect 3679 63524 3745 63547
rect 3831 63524 3913 63547
rect 3999 63524 4065 63547
rect 3679 63484 3688 63524
rect 3728 63484 3745 63524
rect 3831 63484 3852 63524
rect 3892 63484 3913 63524
rect 3999 63484 4016 63524
rect 4056 63484 4065 63524
rect 3679 63461 3745 63484
rect 3831 63461 3913 63484
rect 3999 63461 4065 63484
rect 3679 63442 4065 63461
rect 18799 63547 19185 63566
rect 18799 63524 18865 63547
rect 18951 63524 19033 63547
rect 19119 63524 19185 63547
rect 18799 63484 18808 63524
rect 18848 63484 18865 63524
rect 18951 63484 18972 63524
rect 19012 63484 19033 63524
rect 19119 63484 19136 63524
rect 19176 63484 19185 63524
rect 18799 63461 18865 63484
rect 18951 63461 19033 63484
rect 19119 63461 19185 63484
rect 18799 63442 19185 63461
rect 10243 63148 10252 63188
rect 10292 63148 11020 63188
rect 11060 63148 14284 63188
rect 14324 63148 14333 63188
rect 4919 62791 5305 62810
rect 4919 62768 4985 62791
rect 5071 62768 5153 62791
rect 5239 62768 5305 62791
rect 4919 62728 4928 62768
rect 4968 62728 4985 62768
rect 5071 62728 5092 62768
rect 5132 62728 5153 62768
rect 5239 62728 5256 62768
rect 5296 62728 5305 62768
rect 4919 62705 4985 62728
rect 5071 62705 5153 62728
rect 5239 62705 5305 62728
rect 4919 62686 5305 62705
rect 20039 62791 20425 62810
rect 20039 62768 20105 62791
rect 20191 62768 20273 62791
rect 20359 62768 20425 62791
rect 20039 62728 20048 62768
rect 20088 62728 20105 62768
rect 20191 62728 20212 62768
rect 20252 62728 20273 62768
rect 20359 62728 20376 62768
rect 20416 62728 20425 62768
rect 20039 62705 20105 62728
rect 20191 62705 20273 62728
rect 20359 62705 20425 62728
rect 20039 62686 20425 62705
rect 1315 62140 1324 62180
rect 1364 62140 4588 62180
rect 4628 62140 4637 62180
rect 3679 62035 4065 62054
rect 3679 62012 3745 62035
rect 3831 62012 3913 62035
rect 3999 62012 4065 62035
rect 3679 61972 3688 62012
rect 3728 61972 3745 62012
rect 3831 61972 3852 62012
rect 3892 61972 3913 62012
rect 3999 61972 4016 62012
rect 4056 61972 4065 62012
rect 3679 61949 3745 61972
rect 3831 61949 3913 61972
rect 3999 61949 4065 61972
rect 3679 61930 4065 61949
rect 18799 62035 19185 62054
rect 18799 62012 18865 62035
rect 18951 62012 19033 62035
rect 19119 62012 19185 62035
rect 18799 61972 18808 62012
rect 18848 61972 18865 62012
rect 18951 61972 18972 62012
rect 19012 61972 19033 62012
rect 19119 61972 19136 62012
rect 19176 61972 19185 62012
rect 18799 61949 18865 61972
rect 18951 61949 19033 61972
rect 19119 61949 19185 61972
rect 18799 61930 19185 61949
rect 7555 61804 7564 61844
rect 7604 61804 7852 61844
rect 7892 61804 7901 61844
rect 10915 61384 10924 61424
rect 10964 61384 20236 61424
rect 20276 61384 20285 61424
rect 4919 61279 5305 61298
rect 4919 61256 4985 61279
rect 5071 61256 5153 61279
rect 5239 61256 5305 61279
rect 4919 61216 4928 61256
rect 4968 61216 4985 61256
rect 5071 61216 5092 61256
rect 5132 61216 5153 61256
rect 5239 61216 5256 61256
rect 5296 61216 5305 61256
rect 4919 61193 4985 61216
rect 5071 61193 5153 61216
rect 5239 61193 5305 61216
rect 4919 61174 5305 61193
rect 20039 61279 20425 61298
rect 20039 61256 20105 61279
rect 20191 61256 20273 61279
rect 20359 61256 20425 61279
rect 20039 61216 20048 61256
rect 20088 61216 20105 61256
rect 20191 61216 20212 61256
rect 20252 61216 20273 61256
rect 20359 61216 20376 61256
rect 20416 61216 20425 61256
rect 20039 61193 20105 61216
rect 20191 61193 20273 61216
rect 20359 61193 20425 61216
rect 20039 61174 20425 61193
rect 13946 61111 14070 61130
rect 13946 61088 13965 61111
rect 2755 61048 2764 61088
rect 2804 61048 13965 61088
rect 13946 61025 13965 61048
rect 14051 61025 14070 61111
rect 13946 61006 14070 61025
rect 3679 60523 4065 60542
rect 3679 60500 3745 60523
rect 3831 60500 3913 60523
rect 3999 60500 4065 60523
rect 3679 60460 3688 60500
rect 3728 60460 3745 60500
rect 3831 60460 3852 60500
rect 3892 60460 3913 60500
rect 3999 60460 4016 60500
rect 4056 60460 4065 60500
rect 3679 60437 3745 60460
rect 3831 60437 3913 60460
rect 3999 60437 4065 60460
rect 3679 60418 4065 60437
rect 18799 60523 19185 60542
rect 18799 60500 18865 60523
rect 18951 60500 19033 60523
rect 19119 60500 19185 60523
rect 18799 60460 18808 60500
rect 18848 60460 18865 60500
rect 18951 60460 18972 60500
rect 19012 60460 19033 60500
rect 19119 60460 19136 60500
rect 19176 60460 19185 60500
rect 18799 60437 18865 60460
rect 18951 60437 19033 60460
rect 19119 60437 19185 60460
rect 18799 60418 19185 60437
rect 4919 59767 5305 59786
rect 4919 59744 4985 59767
rect 5071 59744 5153 59767
rect 5239 59744 5305 59767
rect 4919 59704 4928 59744
rect 4968 59704 4985 59744
rect 5071 59704 5092 59744
rect 5132 59704 5153 59744
rect 5239 59704 5256 59744
rect 5296 59704 5305 59744
rect 4919 59681 4985 59704
rect 5071 59681 5153 59704
rect 5239 59681 5305 59704
rect 4919 59662 5305 59681
rect 20039 59767 20425 59786
rect 20039 59744 20105 59767
rect 20191 59744 20273 59767
rect 20359 59744 20425 59767
rect 20039 59704 20048 59744
rect 20088 59704 20105 59744
rect 20191 59704 20212 59744
rect 20252 59704 20273 59744
rect 20359 59704 20376 59744
rect 20416 59704 20425 59744
rect 20039 59681 20105 59704
rect 20191 59681 20273 59704
rect 20359 59681 20425 59704
rect 20039 59662 20425 59681
rect 2467 59452 2476 59492
rect 2516 59452 11788 59492
rect 11828 59452 11837 59492
rect 15356 59452 19564 59492
rect 19604 59452 19613 59492
rect 15356 59408 15396 59452
rect 11203 59368 11212 59408
rect 11252 59368 15396 59408
rect 4195 59200 4204 59240
rect 4244 59200 6892 59240
rect 6932 59200 6941 59240
rect 3679 59011 4065 59030
rect 3679 58988 3745 59011
rect 3831 58988 3913 59011
rect 3999 58988 4065 59011
rect 3679 58948 3688 58988
rect 3728 58948 3745 58988
rect 3831 58948 3852 58988
rect 3892 58948 3913 58988
rect 3999 58948 4016 58988
rect 4056 58948 4065 58988
rect 3679 58925 3745 58948
rect 3831 58925 3913 58948
rect 3999 58925 4065 58948
rect 3679 58906 4065 58925
rect 18799 59011 19185 59030
rect 18799 58988 18865 59011
rect 18951 58988 19033 59011
rect 19119 58988 19185 59011
rect 18799 58948 18808 58988
rect 18848 58948 18865 58988
rect 18951 58948 18972 58988
rect 19012 58948 19033 58988
rect 19119 58948 19136 58988
rect 19176 58948 19185 58988
rect 18799 58925 18865 58948
rect 18951 58925 19033 58948
rect 19119 58925 19185 58948
rect 18799 58906 19185 58925
rect 4919 58255 5305 58274
rect 4919 58232 4985 58255
rect 5071 58232 5153 58255
rect 5239 58232 5305 58255
rect 4919 58192 4928 58232
rect 4968 58192 4985 58232
rect 5071 58192 5092 58232
rect 5132 58192 5153 58232
rect 5239 58192 5256 58232
rect 5296 58192 5305 58232
rect 4919 58169 4985 58192
rect 5071 58169 5153 58192
rect 5239 58169 5305 58192
rect 4919 58150 5305 58169
rect 20039 58255 20425 58274
rect 20039 58232 20105 58255
rect 20191 58232 20273 58255
rect 20359 58232 20425 58255
rect 20039 58192 20048 58232
rect 20088 58192 20105 58232
rect 20191 58192 20212 58232
rect 20252 58192 20273 58232
rect 20359 58192 20376 58232
rect 20416 58192 20425 58232
rect 20039 58169 20105 58192
rect 20191 58169 20273 58192
rect 20359 58169 20425 58192
rect 20039 58150 20425 58169
rect 3679 57499 4065 57518
rect 3679 57476 3745 57499
rect 3831 57476 3913 57499
rect 3999 57476 4065 57499
rect 3679 57436 3688 57476
rect 3728 57436 3745 57476
rect 3831 57436 3852 57476
rect 3892 57436 3913 57476
rect 3999 57436 4016 57476
rect 4056 57436 4065 57476
rect 3679 57413 3745 57436
rect 3831 57413 3913 57436
rect 3999 57413 4065 57436
rect 3679 57394 4065 57413
rect 18799 57499 19185 57518
rect 18799 57476 18865 57499
rect 18951 57476 19033 57499
rect 19119 57476 19185 57499
rect 18799 57436 18808 57476
rect 18848 57436 18865 57476
rect 18951 57436 18972 57476
rect 19012 57436 19033 57476
rect 19119 57436 19136 57476
rect 19176 57436 19185 57476
rect 18799 57413 18865 57436
rect 18951 57413 19033 57436
rect 19119 57413 19185 57436
rect 18799 57394 19185 57413
rect 4919 56743 5305 56762
rect 4919 56720 4985 56743
rect 5071 56720 5153 56743
rect 5239 56720 5305 56743
rect 4919 56680 4928 56720
rect 4968 56680 4985 56720
rect 5071 56680 5092 56720
rect 5132 56680 5153 56720
rect 5239 56680 5256 56720
rect 5296 56680 5305 56720
rect 4919 56657 4985 56680
rect 5071 56657 5153 56680
rect 5239 56657 5305 56680
rect 4919 56638 5305 56657
rect 13946 56743 14070 56762
rect 13946 56657 13965 56743
rect 14051 56720 14070 56743
rect 20039 56743 20425 56762
rect 20039 56720 20105 56743
rect 20191 56720 20273 56743
rect 20359 56720 20425 56743
rect 14051 56680 15052 56720
rect 15092 56680 15101 56720
rect 20039 56680 20048 56720
rect 20088 56680 20105 56720
rect 20191 56680 20212 56720
rect 20252 56680 20273 56720
rect 20359 56680 20376 56720
rect 20416 56680 20425 56720
rect 14051 56657 14070 56680
rect 13946 56638 14070 56657
rect 20039 56657 20105 56680
rect 20191 56657 20273 56680
rect 20359 56657 20425 56680
rect 20039 56638 20425 56657
rect 14851 56512 14860 56552
rect 14900 56512 15052 56552
rect 15092 56512 15101 56552
rect 3679 55987 4065 56006
rect 3679 55964 3745 55987
rect 3831 55964 3913 55987
rect 3999 55964 4065 55987
rect 3679 55924 3688 55964
rect 3728 55924 3745 55964
rect 3831 55924 3852 55964
rect 3892 55924 3913 55964
rect 3999 55924 4016 55964
rect 4056 55924 4065 55964
rect 3679 55901 3745 55924
rect 3831 55901 3913 55924
rect 3999 55901 4065 55924
rect 3679 55882 4065 55901
rect 18799 55987 19185 56006
rect 18799 55964 18865 55987
rect 18951 55964 19033 55987
rect 19119 55964 19185 55987
rect 18799 55924 18808 55964
rect 18848 55924 18865 55964
rect 18951 55924 18972 55964
rect 19012 55924 19033 55964
rect 19119 55924 19136 55964
rect 19176 55924 19185 55964
rect 18799 55901 18865 55924
rect 18951 55901 19033 55924
rect 19119 55901 19185 55924
rect 18799 55882 19185 55901
rect 4919 55231 5305 55250
rect 4919 55208 4985 55231
rect 5071 55208 5153 55231
rect 5239 55208 5305 55231
rect 4919 55168 4928 55208
rect 4968 55168 4985 55208
rect 5071 55168 5092 55208
rect 5132 55168 5153 55208
rect 5239 55168 5256 55208
rect 5296 55168 5305 55208
rect 4919 55145 4985 55168
rect 5071 55145 5153 55168
rect 5239 55145 5305 55168
rect 4919 55126 5305 55145
rect 20039 55231 20425 55250
rect 20039 55208 20105 55231
rect 20191 55208 20273 55231
rect 20359 55208 20425 55231
rect 20039 55168 20048 55208
rect 20088 55168 20105 55208
rect 20191 55168 20212 55208
rect 20252 55168 20273 55208
rect 20359 55168 20376 55208
rect 20416 55168 20425 55208
rect 20039 55145 20105 55168
rect 20191 55145 20273 55168
rect 20359 55145 20425 55168
rect 20039 55126 20425 55145
rect 13699 55084 13708 55124
rect 13748 55084 13996 55124
rect 14036 55084 14045 55124
rect 12451 54580 12460 54620
rect 12500 54580 12652 54620
rect 12692 54580 12701 54620
rect 3679 54475 4065 54494
rect 3679 54452 3745 54475
rect 3831 54452 3913 54475
rect 3999 54452 4065 54475
rect 3679 54412 3688 54452
rect 3728 54412 3745 54452
rect 3831 54412 3852 54452
rect 3892 54412 3913 54452
rect 3999 54412 4016 54452
rect 4056 54412 4065 54452
rect 3679 54389 3745 54412
rect 3831 54389 3913 54412
rect 3999 54389 4065 54412
rect 3679 54370 4065 54389
rect 18799 54475 19185 54494
rect 18799 54452 18865 54475
rect 18951 54452 19033 54475
rect 19119 54452 19185 54475
rect 18799 54412 18808 54452
rect 18848 54412 18865 54452
rect 18951 54412 18972 54452
rect 19012 54412 19033 54452
rect 19119 54412 19136 54452
rect 19176 54412 19185 54452
rect 18799 54389 18865 54412
rect 18951 54389 19033 54412
rect 19119 54389 19185 54412
rect 18799 54370 19185 54389
rect 10819 53992 10828 54032
rect 10868 53992 13228 54032
rect 13268 53992 13277 54032
rect 4919 53719 5305 53738
rect 4919 53696 4985 53719
rect 5071 53696 5153 53719
rect 5239 53696 5305 53719
rect 4919 53656 4928 53696
rect 4968 53656 4985 53696
rect 5071 53656 5092 53696
rect 5132 53656 5153 53696
rect 5239 53656 5256 53696
rect 5296 53656 5305 53696
rect 4919 53633 4985 53656
rect 5071 53633 5153 53656
rect 5239 53633 5305 53656
rect 4919 53614 5305 53633
rect 20039 53719 20425 53738
rect 20039 53696 20105 53719
rect 20191 53696 20273 53719
rect 20359 53696 20425 53719
rect 20039 53656 20048 53696
rect 20088 53656 20105 53696
rect 20191 53656 20212 53696
rect 20252 53656 20273 53696
rect 20359 53656 20376 53696
rect 20416 53656 20425 53696
rect 20039 53633 20105 53656
rect 20191 53633 20273 53656
rect 20359 53633 20425 53656
rect 20039 53614 20425 53633
rect 2275 53236 2284 53276
rect 2324 53236 14284 53276
rect 14324 53236 14333 53276
rect 3679 52963 4065 52982
rect 3679 52940 3745 52963
rect 3831 52940 3913 52963
rect 3999 52940 4065 52963
rect 3679 52900 3688 52940
rect 3728 52900 3745 52940
rect 3831 52900 3852 52940
rect 3892 52900 3913 52940
rect 3999 52900 4016 52940
rect 4056 52900 4065 52940
rect 3679 52877 3745 52900
rect 3831 52877 3913 52900
rect 3999 52877 4065 52900
rect 3679 52858 4065 52877
rect 18799 52963 19185 52982
rect 18799 52940 18865 52963
rect 18951 52940 19033 52963
rect 19119 52940 19185 52963
rect 18799 52900 18808 52940
rect 18848 52900 18865 52940
rect 18951 52900 18972 52940
rect 19012 52900 19033 52940
rect 19119 52900 19136 52940
rect 19176 52900 19185 52940
rect 18799 52877 18865 52900
rect 18951 52877 19033 52900
rect 19119 52877 19185 52900
rect 18799 52858 19185 52877
rect 1123 52732 1132 52772
rect 1172 52732 5068 52772
rect 5108 52732 5117 52772
rect 4919 52207 5305 52226
rect 4919 52184 4985 52207
rect 5071 52184 5153 52207
rect 5239 52184 5305 52207
rect 4919 52144 4928 52184
rect 4968 52144 4985 52184
rect 5071 52144 5092 52184
rect 5132 52144 5153 52184
rect 5239 52144 5256 52184
rect 5296 52144 5305 52184
rect 4919 52121 4985 52144
rect 5071 52121 5153 52144
rect 5239 52121 5305 52144
rect 4919 52102 5305 52121
rect 20039 52207 20425 52226
rect 20039 52184 20105 52207
rect 20191 52184 20273 52207
rect 20359 52184 20425 52207
rect 20039 52144 20048 52184
rect 20088 52144 20105 52184
rect 20191 52144 20212 52184
rect 20252 52144 20273 52184
rect 20359 52144 20376 52184
rect 20416 52144 20425 52184
rect 20039 52121 20105 52144
rect 20191 52121 20273 52144
rect 20359 52121 20425 52144
rect 20039 52102 20425 52121
rect 3679 51451 4065 51470
rect 3679 51428 3745 51451
rect 3831 51428 3913 51451
rect 3999 51428 4065 51451
rect 3679 51388 3688 51428
rect 3728 51388 3745 51428
rect 3831 51388 3852 51428
rect 3892 51388 3913 51428
rect 3999 51388 4016 51428
rect 4056 51388 4065 51428
rect 3679 51365 3745 51388
rect 3831 51365 3913 51388
rect 3999 51365 4065 51388
rect 3679 51346 4065 51365
rect 18799 51451 19185 51470
rect 18799 51428 18865 51451
rect 18951 51428 19033 51451
rect 19119 51428 19185 51451
rect 18799 51388 18808 51428
rect 18848 51388 18865 51428
rect 18951 51388 18972 51428
rect 19012 51388 19033 51428
rect 19119 51388 19136 51428
rect 19176 51388 19185 51428
rect 18799 51365 18865 51388
rect 18951 51365 19033 51388
rect 19119 51365 19185 51388
rect 18799 51346 19185 51365
rect 4919 50695 5305 50714
rect 4919 50672 4985 50695
rect 5071 50672 5153 50695
rect 5239 50672 5305 50695
rect 4919 50632 4928 50672
rect 4968 50632 4985 50672
rect 5071 50632 5092 50672
rect 5132 50632 5153 50672
rect 5239 50632 5256 50672
rect 5296 50632 5305 50672
rect 4919 50609 4985 50632
rect 5071 50609 5153 50632
rect 5239 50609 5305 50632
rect 4919 50590 5305 50609
rect 20039 50695 20425 50714
rect 20039 50672 20105 50695
rect 20191 50672 20273 50695
rect 20359 50672 20425 50695
rect 20039 50632 20048 50672
rect 20088 50632 20105 50672
rect 20191 50632 20212 50672
rect 20252 50632 20273 50672
rect 20359 50632 20376 50672
rect 20416 50632 20425 50672
rect 20039 50609 20105 50632
rect 20191 50609 20273 50632
rect 20359 50609 20425 50632
rect 20039 50590 20425 50609
rect 3679 49939 4065 49958
rect 3679 49916 3745 49939
rect 3831 49916 3913 49939
rect 3999 49916 4065 49939
rect 3679 49876 3688 49916
rect 3728 49876 3745 49916
rect 3831 49876 3852 49916
rect 3892 49876 3913 49916
rect 3999 49876 4016 49916
rect 4056 49876 4065 49916
rect 3679 49853 3745 49876
rect 3831 49853 3913 49876
rect 3999 49853 4065 49876
rect 3679 49834 4065 49853
rect 18799 49939 19185 49958
rect 18799 49916 18865 49939
rect 18951 49916 19033 49939
rect 19119 49916 19185 49939
rect 18799 49876 18808 49916
rect 18848 49876 18865 49916
rect 18951 49876 18972 49916
rect 19012 49876 19033 49916
rect 19119 49876 19136 49916
rect 19176 49876 19185 49916
rect 18799 49853 18865 49876
rect 18951 49853 19033 49876
rect 19119 49853 19185 49876
rect 18799 49834 19185 49853
rect 19460 49876 20140 49916
rect 20180 49876 20189 49916
rect 19460 49748 19500 49876
rect 8515 49708 8524 49748
rect 8564 49708 19500 49748
rect 9667 49456 9676 49496
rect 9716 49456 14668 49496
rect 14708 49456 14717 49496
rect 4919 49183 5305 49202
rect 4919 49160 4985 49183
rect 5071 49160 5153 49183
rect 5239 49160 5305 49183
rect 4919 49120 4928 49160
rect 4968 49120 4985 49160
rect 5071 49120 5092 49160
rect 5132 49120 5153 49160
rect 5239 49120 5256 49160
rect 5296 49120 5305 49160
rect 4919 49097 4985 49120
rect 5071 49097 5153 49120
rect 5239 49097 5305 49120
rect 4919 49078 5305 49097
rect 20039 49183 20425 49202
rect 20039 49160 20105 49183
rect 20191 49160 20273 49183
rect 20359 49160 20425 49183
rect 20039 49120 20048 49160
rect 20088 49120 20105 49160
rect 20191 49120 20212 49160
rect 20252 49120 20273 49160
rect 20359 49120 20376 49160
rect 20416 49120 20425 49160
rect 20039 49097 20105 49120
rect 20191 49097 20273 49120
rect 20359 49097 20425 49120
rect 20039 49078 20425 49097
rect 3679 48427 4065 48446
rect 3679 48404 3745 48427
rect 3831 48404 3913 48427
rect 3999 48404 4065 48427
rect 3679 48364 3688 48404
rect 3728 48364 3745 48404
rect 3831 48364 3852 48404
rect 3892 48364 3913 48404
rect 3999 48364 4016 48404
rect 4056 48364 4065 48404
rect 3679 48341 3745 48364
rect 3831 48341 3913 48364
rect 3999 48341 4065 48364
rect 3679 48322 4065 48341
rect 18799 48427 19185 48446
rect 18799 48404 18865 48427
rect 18951 48404 19033 48427
rect 19119 48404 19185 48427
rect 18799 48364 18808 48404
rect 18848 48364 18865 48404
rect 18951 48364 18972 48404
rect 19012 48364 19033 48404
rect 19119 48364 19136 48404
rect 19176 48364 19185 48404
rect 18799 48341 18865 48364
rect 18951 48341 19033 48364
rect 19119 48341 19185 48364
rect 18799 48322 19185 48341
rect 8474 48091 8598 48110
rect 8474 48005 8493 48091
rect 8579 48068 8598 48091
rect 8579 48028 8716 48068
rect 8756 48028 8765 48068
rect 8579 48005 8598 48028
rect 8474 47986 8598 48005
rect 14755 47944 14764 47984
rect 14804 47944 14956 47984
rect 14996 47944 15005 47984
rect 4919 47671 5305 47690
rect 4919 47648 4985 47671
rect 5071 47648 5153 47671
rect 5239 47648 5305 47671
rect 4919 47608 4928 47648
rect 4968 47608 4985 47648
rect 5071 47608 5092 47648
rect 5132 47608 5153 47648
rect 5239 47608 5256 47648
rect 5296 47608 5305 47648
rect 4919 47585 4985 47608
rect 5071 47585 5153 47608
rect 5239 47585 5305 47608
rect 4919 47566 5305 47585
rect 20039 47671 20425 47690
rect 20039 47648 20105 47671
rect 20191 47648 20273 47671
rect 20359 47648 20425 47671
rect 20039 47608 20048 47648
rect 20088 47608 20105 47648
rect 20191 47608 20212 47648
rect 20252 47608 20273 47648
rect 20359 47608 20376 47648
rect 20416 47608 20425 47648
rect 20039 47585 20105 47608
rect 20191 47585 20273 47608
rect 20359 47585 20425 47608
rect 20039 47566 20425 47585
rect 3679 46915 4065 46934
rect 3679 46892 3745 46915
rect 3831 46892 3913 46915
rect 3999 46892 4065 46915
rect 3679 46852 3688 46892
rect 3728 46852 3745 46892
rect 3831 46852 3852 46892
rect 3892 46852 3913 46892
rect 3999 46852 4016 46892
rect 4056 46852 4065 46892
rect 3679 46829 3745 46852
rect 3831 46829 3913 46852
rect 3999 46829 4065 46852
rect 3679 46810 4065 46829
rect 18799 46915 19185 46934
rect 18799 46892 18865 46915
rect 18951 46892 19033 46915
rect 19119 46892 19185 46915
rect 18799 46852 18808 46892
rect 18848 46852 18865 46892
rect 18951 46852 18972 46892
rect 19012 46852 19033 46892
rect 19119 46852 19136 46892
rect 19176 46852 19185 46892
rect 18799 46829 18865 46852
rect 18951 46829 19033 46852
rect 19119 46829 19185 46852
rect 18799 46810 19185 46829
rect 4919 46159 5305 46178
rect 4919 46136 4985 46159
rect 5071 46136 5153 46159
rect 5239 46136 5305 46159
rect 4919 46096 4928 46136
rect 4968 46096 4985 46136
rect 5071 46096 5092 46136
rect 5132 46096 5153 46136
rect 5239 46096 5256 46136
rect 5296 46096 5305 46136
rect 4919 46073 4985 46096
rect 5071 46073 5153 46096
rect 5239 46073 5305 46096
rect 4919 46054 5305 46073
rect 20039 46159 20425 46178
rect 20039 46136 20105 46159
rect 20191 46136 20273 46159
rect 20359 46136 20425 46159
rect 20039 46096 20048 46136
rect 20088 46096 20105 46136
rect 20191 46096 20212 46136
rect 20252 46096 20273 46136
rect 20359 46096 20376 46136
rect 20416 46096 20425 46136
rect 20039 46073 20105 46096
rect 20191 46073 20273 46096
rect 20359 46073 20425 46096
rect 20039 46054 20425 46073
rect 3679 45403 4065 45422
rect 3679 45380 3745 45403
rect 3831 45380 3913 45403
rect 3999 45380 4065 45403
rect 3679 45340 3688 45380
rect 3728 45340 3745 45380
rect 3831 45340 3852 45380
rect 3892 45340 3913 45380
rect 3999 45340 4016 45380
rect 4056 45340 4065 45380
rect 3679 45317 3745 45340
rect 3831 45317 3913 45340
rect 3999 45317 4065 45340
rect 3679 45298 4065 45317
rect 18799 45403 19185 45422
rect 18799 45380 18865 45403
rect 18951 45380 19033 45403
rect 19119 45380 19185 45403
rect 18799 45340 18808 45380
rect 18848 45340 18865 45380
rect 18951 45340 18972 45380
rect 19012 45340 19033 45380
rect 19119 45340 19136 45380
rect 19176 45340 19185 45380
rect 18799 45317 18865 45340
rect 18951 45317 19033 45340
rect 19119 45317 19185 45340
rect 18799 45298 19185 45317
rect 12259 44920 12268 44960
rect 12308 44920 20140 44960
rect 20180 44920 20189 44960
rect 4919 44647 5305 44666
rect 4919 44624 4985 44647
rect 5071 44624 5153 44647
rect 5239 44624 5305 44647
rect 4919 44584 4928 44624
rect 4968 44584 4985 44624
rect 5071 44584 5092 44624
rect 5132 44584 5153 44624
rect 5239 44584 5256 44624
rect 5296 44584 5305 44624
rect 4919 44561 4985 44584
rect 5071 44561 5153 44584
rect 5239 44561 5305 44584
rect 4919 44542 5305 44561
rect 20039 44647 20425 44666
rect 20039 44624 20105 44647
rect 20191 44624 20273 44647
rect 20359 44624 20425 44647
rect 20039 44584 20048 44624
rect 20088 44584 20105 44624
rect 20191 44584 20212 44624
rect 20252 44584 20273 44624
rect 20359 44584 20376 44624
rect 20416 44584 20425 44624
rect 20039 44561 20105 44584
rect 20191 44561 20273 44584
rect 20359 44561 20425 44584
rect 20039 44542 20425 44561
rect 3679 43891 4065 43910
rect 3679 43868 3745 43891
rect 3831 43868 3913 43891
rect 3999 43868 4065 43891
rect 3679 43828 3688 43868
rect 3728 43828 3745 43868
rect 3831 43828 3852 43868
rect 3892 43828 3913 43868
rect 3999 43828 4016 43868
rect 4056 43828 4065 43868
rect 3679 43805 3745 43828
rect 3831 43805 3913 43828
rect 3999 43805 4065 43828
rect 3679 43786 4065 43805
rect 18799 43891 19185 43910
rect 18799 43868 18865 43891
rect 18951 43868 19033 43891
rect 19119 43868 19185 43891
rect 18799 43828 18808 43868
rect 18848 43828 18865 43868
rect 18951 43828 18972 43868
rect 19012 43828 19033 43868
rect 19119 43828 19136 43868
rect 19176 43828 19185 43868
rect 18799 43805 18865 43828
rect 18951 43805 19033 43828
rect 19119 43805 19185 43828
rect 18799 43786 19185 43805
rect 4919 43135 5305 43154
rect 4919 43112 4985 43135
rect 5071 43112 5153 43135
rect 5239 43112 5305 43135
rect 4919 43072 4928 43112
rect 4968 43072 4985 43112
rect 5071 43072 5092 43112
rect 5132 43072 5153 43112
rect 5239 43072 5256 43112
rect 5296 43072 5305 43112
rect 4919 43049 4985 43072
rect 5071 43049 5153 43072
rect 5239 43049 5305 43072
rect 4919 43030 5305 43049
rect 20039 43135 20425 43154
rect 20039 43112 20105 43135
rect 20191 43112 20273 43135
rect 20359 43112 20425 43135
rect 20039 43072 20048 43112
rect 20088 43072 20105 43112
rect 20191 43072 20212 43112
rect 20252 43072 20273 43112
rect 20359 43072 20376 43112
rect 20416 43072 20425 43112
rect 20039 43049 20105 43072
rect 20191 43049 20273 43072
rect 20359 43049 20425 43072
rect 20039 43030 20425 43049
rect 11011 42484 11020 42524
rect 11060 42484 19948 42524
rect 19988 42484 19997 42524
rect 3679 42379 4065 42398
rect 3679 42356 3745 42379
rect 3831 42356 3913 42379
rect 3999 42356 4065 42379
rect 18799 42379 19185 42398
rect 18799 42356 18865 42379
rect 18951 42356 19033 42379
rect 19119 42356 19185 42379
rect 3679 42316 3688 42356
rect 3728 42316 3745 42356
rect 3831 42316 3852 42356
rect 3892 42316 3913 42356
rect 3999 42316 4016 42356
rect 4056 42316 4065 42356
rect 11107 42316 11116 42356
rect 11156 42316 17548 42356
rect 17588 42316 17597 42356
rect 18799 42316 18808 42356
rect 18848 42316 18865 42356
rect 18951 42316 18972 42356
rect 19012 42316 19033 42356
rect 19119 42316 19136 42356
rect 19176 42316 19185 42356
rect 3679 42293 3745 42316
rect 3831 42293 3913 42316
rect 3999 42293 4065 42316
rect 3679 42274 4065 42293
rect 18799 42293 18865 42316
rect 18951 42293 19033 42316
rect 19119 42293 19185 42316
rect 18799 42274 19185 42293
rect 3235 41896 3244 41936
rect 3284 41896 4780 41936
rect 4820 41896 4829 41936
rect 6499 41644 6508 41684
rect 6548 41644 6892 41684
rect 6932 41644 6941 41684
rect 4919 41623 5305 41642
rect 4919 41600 4985 41623
rect 5071 41600 5153 41623
rect 5239 41600 5305 41623
rect 20039 41623 20425 41642
rect 20039 41600 20105 41623
rect 20191 41600 20273 41623
rect 20359 41600 20425 41623
rect 4919 41560 4928 41600
rect 4968 41560 4985 41600
rect 5071 41560 5092 41600
rect 5132 41560 5153 41600
rect 5239 41560 5256 41600
rect 5296 41560 5305 41600
rect 6979 41560 6988 41600
rect 7028 41560 7564 41600
rect 7604 41560 7613 41600
rect 20039 41560 20048 41600
rect 20088 41560 20105 41600
rect 20191 41560 20212 41600
rect 20252 41560 20273 41600
rect 20359 41560 20376 41600
rect 20416 41560 20425 41600
rect 4919 41537 4985 41560
rect 5071 41537 5153 41560
rect 5239 41537 5305 41560
rect 4919 41518 5305 41537
rect 20039 41537 20105 41560
rect 20191 41537 20273 41560
rect 20359 41537 20425 41560
rect 20039 41518 20425 41537
rect 3139 41392 3148 41432
rect 3188 41392 7276 41432
rect 7316 41392 7325 41432
rect 3679 40867 4065 40886
rect 3679 40844 3745 40867
rect 3831 40844 3913 40867
rect 3999 40844 4065 40867
rect 3679 40804 3688 40844
rect 3728 40804 3745 40844
rect 3831 40804 3852 40844
rect 3892 40804 3913 40844
rect 3999 40804 4016 40844
rect 4056 40804 4065 40844
rect 3679 40781 3745 40804
rect 3831 40781 3913 40804
rect 3999 40781 4065 40804
rect 3679 40762 4065 40781
rect 18799 40867 19185 40886
rect 18799 40844 18865 40867
rect 18951 40844 19033 40867
rect 19119 40844 19185 40867
rect 18799 40804 18808 40844
rect 18848 40804 18865 40844
rect 18951 40804 18972 40844
rect 19012 40804 19033 40844
rect 19119 40804 19136 40844
rect 19176 40804 19185 40844
rect 18799 40781 18865 40804
rect 18951 40781 19033 40804
rect 19119 40781 19185 40804
rect 18799 40762 19185 40781
rect 4919 40111 5305 40130
rect 4919 40088 4985 40111
rect 5071 40088 5153 40111
rect 5239 40088 5305 40111
rect 4919 40048 4928 40088
rect 4968 40048 4985 40088
rect 5071 40048 5092 40088
rect 5132 40048 5153 40088
rect 5239 40048 5256 40088
rect 5296 40048 5305 40088
rect 4919 40025 4985 40048
rect 5071 40025 5153 40048
rect 5239 40025 5305 40048
rect 4919 40006 5305 40025
rect 20039 40111 20425 40130
rect 20039 40088 20105 40111
rect 20191 40088 20273 40111
rect 20359 40088 20425 40111
rect 20039 40048 20048 40088
rect 20088 40048 20105 40088
rect 20191 40048 20212 40088
rect 20252 40048 20273 40088
rect 20359 40048 20376 40088
rect 20416 40048 20425 40088
rect 20039 40025 20105 40048
rect 20191 40025 20273 40048
rect 20359 40025 20425 40048
rect 20039 40006 20425 40025
rect 10531 39880 10540 39920
rect 10580 39880 11116 39920
rect 11156 39880 11165 39920
rect 3679 39355 4065 39374
rect 3679 39332 3745 39355
rect 3831 39332 3913 39355
rect 3999 39332 4065 39355
rect 3679 39292 3688 39332
rect 3728 39292 3745 39332
rect 3831 39292 3852 39332
rect 3892 39292 3913 39332
rect 3999 39292 4016 39332
rect 4056 39292 4065 39332
rect 3679 39269 3745 39292
rect 3831 39269 3913 39292
rect 3999 39269 4065 39292
rect 3679 39250 4065 39269
rect 18799 39355 19185 39374
rect 18799 39332 18865 39355
rect 18951 39332 19033 39355
rect 19119 39332 19185 39355
rect 18799 39292 18808 39332
rect 18848 39292 18865 39332
rect 18951 39292 18972 39332
rect 19012 39292 19033 39332
rect 19119 39292 19136 39332
rect 19176 39292 19185 39332
rect 18799 39269 18865 39292
rect 18951 39269 19033 39292
rect 19119 39269 19185 39292
rect 18799 39250 19185 39269
rect 2371 39040 2380 39080
rect 2420 39040 4300 39080
rect 4340 39040 7180 39080
rect 7220 39040 7229 39080
rect 4919 38599 5305 38618
rect 4919 38576 4985 38599
rect 5071 38576 5153 38599
rect 5239 38576 5305 38599
rect 4919 38536 4928 38576
rect 4968 38536 4985 38576
rect 5071 38536 5092 38576
rect 5132 38536 5153 38576
rect 5239 38536 5256 38576
rect 5296 38536 5305 38576
rect 4919 38513 4985 38536
rect 5071 38513 5153 38536
rect 5239 38513 5305 38536
rect 4919 38494 5305 38513
rect 20039 38599 20425 38618
rect 20039 38576 20105 38599
rect 20191 38576 20273 38599
rect 20359 38576 20425 38599
rect 20039 38536 20048 38576
rect 20088 38536 20105 38576
rect 20191 38536 20212 38576
rect 20252 38536 20273 38576
rect 20359 38536 20376 38576
rect 20416 38536 20425 38576
rect 20039 38513 20105 38536
rect 20191 38513 20273 38536
rect 20359 38513 20425 38536
rect 20039 38494 20425 38513
rect 3679 37843 4065 37862
rect 3679 37820 3745 37843
rect 3831 37820 3913 37843
rect 3999 37820 4065 37843
rect 3679 37780 3688 37820
rect 3728 37780 3745 37820
rect 3831 37780 3852 37820
rect 3892 37780 3913 37820
rect 3999 37780 4016 37820
rect 4056 37780 4065 37820
rect 3679 37757 3745 37780
rect 3831 37757 3913 37780
rect 3999 37757 4065 37780
rect 3679 37738 4065 37757
rect 18799 37843 19185 37862
rect 18799 37820 18865 37843
rect 18951 37820 19033 37843
rect 19119 37820 19185 37843
rect 18799 37780 18808 37820
rect 18848 37780 18865 37820
rect 18951 37780 18972 37820
rect 19012 37780 19033 37820
rect 19119 37780 19136 37820
rect 19176 37780 19185 37820
rect 18799 37757 18865 37780
rect 18951 37757 19033 37780
rect 19119 37757 19185 37780
rect 18799 37738 19185 37757
rect 5780 37696 7852 37736
rect 7892 37696 8524 37736
rect 8564 37696 8573 37736
rect 5780 37652 5820 37696
rect 1219 37612 1228 37652
rect 1268 37612 5820 37652
rect 6307 37612 6316 37652
rect 6356 37612 6508 37652
rect 6548 37612 6557 37652
rect 3811 37444 3820 37484
rect 3860 37444 6316 37484
rect 6356 37444 6365 37484
rect 2851 37276 2860 37316
rect 2900 37276 4108 37316
rect 4148 37276 4157 37316
rect 4919 37087 5305 37106
rect 4919 37064 4985 37087
rect 5071 37064 5153 37087
rect 5239 37064 5305 37087
rect 4919 37024 4928 37064
rect 4968 37024 4985 37064
rect 5071 37024 5092 37064
rect 5132 37024 5153 37064
rect 5239 37024 5256 37064
rect 5296 37024 5305 37064
rect 4919 37001 4985 37024
rect 5071 37001 5153 37024
rect 5239 37001 5305 37024
rect 4919 36982 5305 37001
rect 20039 37087 20425 37106
rect 20039 37064 20105 37087
rect 20191 37064 20273 37087
rect 20359 37064 20425 37087
rect 20039 37024 20048 37064
rect 20088 37024 20105 37064
rect 20191 37024 20212 37064
rect 20252 37024 20273 37064
rect 20359 37024 20376 37064
rect 20416 37024 20425 37064
rect 20039 37001 20105 37024
rect 20191 37001 20273 37024
rect 20359 37001 20425 37024
rect 20039 36982 20425 37001
rect 4099 36688 4108 36728
rect 4148 36688 6988 36728
rect 7028 36688 7037 36728
rect 5635 36520 5644 36560
rect 5684 36520 7180 36560
rect 7220 36520 7229 36560
rect 3679 36331 4065 36350
rect 3679 36308 3745 36331
rect 3831 36308 3913 36331
rect 3999 36308 4065 36331
rect 3679 36268 3688 36308
rect 3728 36268 3745 36308
rect 3831 36268 3852 36308
rect 3892 36268 3913 36308
rect 3999 36268 4016 36308
rect 4056 36268 4065 36308
rect 3679 36245 3745 36268
rect 3831 36245 3913 36268
rect 3999 36245 4065 36268
rect 3679 36226 4065 36245
rect 18799 36331 19185 36350
rect 18799 36308 18865 36331
rect 18951 36308 19033 36331
rect 19119 36308 19185 36331
rect 18799 36268 18808 36308
rect 18848 36268 18865 36308
rect 18951 36268 18972 36308
rect 19012 36268 19033 36308
rect 19119 36268 19136 36308
rect 19176 36268 19185 36308
rect 18799 36245 18865 36268
rect 18951 36245 19033 36268
rect 19119 36245 19185 36268
rect 18799 36226 19185 36245
rect 4675 35680 4684 35720
rect 4724 35680 5836 35720
rect 5876 35680 5885 35720
rect 4919 35575 5305 35594
rect 4919 35552 4985 35575
rect 5071 35552 5153 35575
rect 5239 35552 5305 35575
rect 4919 35512 4928 35552
rect 4968 35512 4985 35552
rect 5071 35512 5092 35552
rect 5132 35512 5153 35552
rect 5239 35512 5256 35552
rect 5296 35512 5305 35552
rect 4919 35489 4985 35512
rect 5071 35489 5153 35512
rect 5239 35489 5305 35512
rect 4919 35470 5305 35489
rect 20039 35575 20425 35594
rect 20039 35552 20105 35575
rect 20191 35552 20273 35575
rect 20359 35552 20425 35575
rect 20039 35512 20048 35552
rect 20088 35512 20105 35552
rect 20191 35512 20212 35552
rect 20252 35512 20273 35552
rect 20359 35512 20376 35552
rect 20416 35512 20425 35552
rect 20039 35489 20105 35512
rect 20191 35489 20273 35512
rect 20359 35489 20425 35512
rect 20039 35470 20425 35489
rect 3679 34819 4065 34838
rect 3679 34796 3745 34819
rect 3831 34796 3913 34819
rect 3999 34796 4065 34819
rect 3679 34756 3688 34796
rect 3728 34756 3745 34796
rect 3831 34756 3852 34796
rect 3892 34756 3913 34796
rect 3999 34756 4016 34796
rect 4056 34756 4065 34796
rect 3679 34733 3745 34756
rect 3831 34733 3913 34756
rect 3999 34733 4065 34756
rect 3679 34714 4065 34733
rect 18799 34819 19185 34838
rect 18799 34796 18865 34819
rect 18951 34796 19033 34819
rect 19119 34796 19185 34819
rect 18799 34756 18808 34796
rect 18848 34756 18865 34796
rect 18951 34756 18972 34796
rect 19012 34756 19033 34796
rect 19119 34756 19136 34796
rect 19176 34756 19185 34796
rect 18799 34733 18865 34756
rect 18951 34733 19033 34756
rect 19119 34733 19185 34756
rect 18799 34714 19185 34733
rect 4919 34063 5305 34082
rect 4919 34040 4985 34063
rect 5071 34040 5153 34063
rect 5239 34040 5305 34063
rect 4919 34000 4928 34040
rect 4968 34000 4985 34040
rect 5071 34000 5092 34040
rect 5132 34000 5153 34040
rect 5239 34000 5256 34040
rect 5296 34000 5305 34040
rect 4919 33977 4985 34000
rect 5071 33977 5153 34000
rect 5239 33977 5305 34000
rect 4919 33958 5305 33977
rect 20039 34063 20425 34082
rect 20039 34040 20105 34063
rect 20191 34040 20273 34063
rect 20359 34040 20425 34063
rect 20039 34000 20048 34040
rect 20088 34000 20105 34040
rect 20191 34000 20212 34040
rect 20252 34000 20273 34040
rect 20359 34000 20376 34040
rect 20416 34000 20425 34040
rect 20039 33977 20105 34000
rect 20191 33977 20273 34000
rect 20359 33977 20425 34000
rect 20039 33958 20425 33977
rect 4003 33832 4012 33872
rect 4052 33832 6412 33872
rect 6452 33832 6461 33872
rect 11011 33664 11020 33704
rect 11060 33664 11500 33704
rect 11540 33664 11549 33704
rect 3679 33307 4065 33326
rect 3679 33284 3745 33307
rect 3831 33284 3913 33307
rect 3999 33284 4065 33307
rect 3679 33244 3688 33284
rect 3728 33244 3745 33284
rect 3831 33244 3852 33284
rect 3892 33244 3913 33284
rect 3999 33244 4016 33284
rect 4056 33244 4065 33284
rect 3679 33221 3745 33244
rect 3831 33221 3913 33244
rect 3999 33221 4065 33244
rect 3679 33202 4065 33221
rect 18799 33307 19185 33326
rect 18799 33284 18865 33307
rect 18951 33284 19033 33307
rect 19119 33284 19185 33307
rect 18799 33244 18808 33284
rect 18848 33244 18865 33284
rect 18951 33244 18972 33284
rect 19012 33244 19033 33284
rect 19119 33244 19136 33284
rect 19176 33244 19185 33284
rect 18799 33221 18865 33244
rect 18951 33221 19033 33244
rect 19119 33221 19185 33244
rect 18799 33202 19185 33221
rect 4919 32551 5305 32570
rect 4919 32528 4985 32551
rect 5071 32528 5153 32551
rect 5239 32528 5305 32551
rect 4919 32488 4928 32528
rect 4968 32488 4985 32528
rect 5071 32488 5092 32528
rect 5132 32488 5153 32528
rect 5239 32488 5256 32528
rect 5296 32488 5305 32528
rect 4919 32465 4985 32488
rect 5071 32465 5153 32488
rect 5239 32465 5305 32488
rect 4919 32446 5305 32465
rect 20039 32551 20425 32570
rect 20039 32528 20105 32551
rect 20191 32528 20273 32551
rect 20359 32528 20425 32551
rect 20039 32488 20048 32528
rect 20088 32488 20105 32528
rect 20191 32488 20212 32528
rect 20252 32488 20273 32528
rect 20359 32488 20376 32528
rect 20416 32488 20425 32528
rect 20039 32465 20105 32488
rect 20191 32465 20273 32488
rect 20359 32465 20425 32488
rect 20039 32446 20425 32465
rect 1178 32131 1302 32150
rect 1178 32045 1197 32131
rect 1283 32108 1302 32131
rect 1283 32068 20716 32108
rect 20756 32068 20765 32108
rect 1283 32045 1302 32068
rect 1178 32026 1302 32045
rect 3679 31795 4065 31814
rect 3679 31772 3745 31795
rect 3831 31772 3913 31795
rect 3999 31772 4065 31795
rect 3679 31732 3688 31772
rect 3728 31732 3745 31772
rect 3831 31732 3852 31772
rect 3892 31732 3913 31772
rect 3999 31732 4016 31772
rect 4056 31732 4065 31772
rect 3679 31709 3745 31732
rect 3831 31709 3913 31732
rect 3999 31709 4065 31732
rect 3679 31690 4065 31709
rect 18799 31795 19185 31814
rect 18799 31772 18865 31795
rect 18951 31772 19033 31795
rect 19119 31772 19185 31795
rect 18799 31732 18808 31772
rect 18848 31732 18865 31772
rect 18951 31732 18972 31772
rect 19012 31732 19033 31772
rect 19119 31732 19136 31772
rect 19176 31732 19185 31772
rect 18799 31709 18865 31732
rect 18951 31709 19033 31732
rect 19119 31709 19185 31732
rect 18799 31690 19185 31709
rect 4919 31039 5305 31058
rect 4919 31016 4985 31039
rect 5071 31016 5153 31039
rect 5239 31016 5305 31039
rect 4919 30976 4928 31016
rect 4968 30976 4985 31016
rect 5071 30976 5092 31016
rect 5132 30976 5153 31016
rect 5239 30976 5256 31016
rect 5296 30976 5305 31016
rect 4919 30953 4985 30976
rect 5071 30953 5153 30976
rect 5239 30953 5305 30976
rect 4919 30934 5305 30953
rect 20039 31039 20425 31058
rect 20039 31016 20105 31039
rect 20191 31016 20273 31039
rect 20359 31016 20425 31039
rect 20039 30976 20048 31016
rect 20088 30976 20105 31016
rect 20191 30976 20212 31016
rect 20252 30976 20273 31016
rect 20359 30976 20376 31016
rect 20416 30976 20425 31016
rect 20039 30953 20105 30976
rect 20191 30953 20273 30976
rect 20359 30953 20425 30976
rect 20039 30934 20425 30953
rect 10627 30892 10636 30932
rect 10676 30892 16876 30932
rect 16916 30892 16925 30932
rect 6019 30808 6028 30848
rect 6068 30808 6220 30848
rect 6260 30808 6269 30848
rect 3679 30283 4065 30302
rect 3679 30260 3745 30283
rect 3831 30260 3913 30283
rect 3999 30260 4065 30283
rect 3679 30220 3688 30260
rect 3728 30220 3745 30260
rect 3831 30220 3852 30260
rect 3892 30220 3913 30260
rect 3999 30220 4016 30260
rect 4056 30220 4065 30260
rect 3679 30197 3745 30220
rect 3831 30197 3913 30220
rect 3999 30197 4065 30220
rect 3679 30178 4065 30197
rect 18799 30283 19185 30302
rect 18799 30260 18865 30283
rect 18951 30260 19033 30283
rect 19119 30260 19185 30283
rect 18799 30220 18808 30260
rect 18848 30220 18865 30260
rect 18951 30220 18972 30260
rect 19012 30220 19033 30260
rect 19119 30220 19136 30260
rect 19176 30220 19185 30260
rect 18799 30197 18865 30220
rect 18951 30197 19033 30220
rect 19119 30197 19185 30220
rect 18799 30178 19185 30197
rect 4099 29632 4108 29672
rect 4148 29632 6796 29672
rect 6836 29632 6845 29672
rect 13507 29632 13516 29672
rect 13556 29632 14188 29672
rect 14228 29632 14237 29672
rect 4919 29527 5305 29546
rect 4919 29504 4985 29527
rect 5071 29504 5153 29527
rect 5239 29504 5305 29527
rect 4919 29464 4928 29504
rect 4968 29464 4985 29504
rect 5071 29464 5092 29504
rect 5132 29464 5153 29504
rect 5239 29464 5256 29504
rect 5296 29464 5305 29504
rect 4919 29441 4985 29464
rect 5071 29441 5153 29464
rect 5239 29441 5305 29464
rect 4919 29422 5305 29441
rect 20039 29527 20425 29546
rect 20039 29504 20105 29527
rect 20191 29504 20273 29527
rect 20359 29504 20425 29527
rect 20039 29464 20048 29504
rect 20088 29464 20105 29504
rect 20191 29464 20212 29504
rect 20252 29464 20273 29504
rect 20359 29464 20376 29504
rect 20416 29464 20425 29504
rect 20039 29441 20105 29464
rect 20191 29441 20273 29464
rect 20359 29441 20425 29464
rect 20039 29422 20425 29441
rect 5827 29128 5836 29168
rect 5876 29128 9964 29168
rect 10004 29128 10013 29168
rect 13219 28876 13228 28916
rect 13268 28876 14860 28916
rect 14900 28876 14909 28916
rect 3679 28771 4065 28790
rect 3679 28748 3745 28771
rect 3831 28748 3913 28771
rect 3999 28748 4065 28771
rect 3679 28708 3688 28748
rect 3728 28708 3745 28748
rect 3831 28708 3852 28748
rect 3892 28708 3913 28748
rect 3999 28708 4016 28748
rect 4056 28708 4065 28748
rect 3679 28685 3745 28708
rect 3831 28685 3913 28708
rect 3999 28685 4065 28708
rect 3679 28666 4065 28685
rect 18799 28771 19185 28790
rect 18799 28748 18865 28771
rect 18951 28748 19033 28771
rect 19119 28748 19185 28771
rect 18799 28708 18808 28748
rect 18848 28708 18865 28748
rect 18951 28708 18972 28748
rect 19012 28708 19033 28748
rect 19119 28708 19136 28748
rect 19176 28708 19185 28748
rect 18799 28685 18865 28708
rect 18951 28685 19033 28708
rect 19119 28685 19185 28708
rect 18799 28666 19185 28685
rect 4919 28015 5305 28034
rect 4919 27992 4985 28015
rect 5071 27992 5153 28015
rect 5239 27992 5305 28015
rect 4919 27952 4928 27992
rect 4968 27952 4985 27992
rect 5071 27952 5092 27992
rect 5132 27952 5153 27992
rect 5239 27952 5256 27992
rect 5296 27952 5305 27992
rect 4919 27929 4985 27952
rect 5071 27929 5153 27952
rect 5239 27929 5305 27952
rect 4919 27910 5305 27929
rect 20039 28015 20425 28034
rect 20039 27992 20105 28015
rect 20191 27992 20273 28015
rect 20359 27992 20425 28015
rect 20039 27952 20048 27992
rect 20088 27952 20105 27992
rect 20191 27952 20212 27992
rect 20252 27952 20273 27992
rect 20359 27952 20376 27992
rect 20416 27952 20425 27992
rect 20039 27929 20105 27952
rect 20191 27929 20273 27952
rect 20359 27929 20425 27952
rect 20039 27910 20425 27929
rect 643 27700 652 27740
rect 692 27700 4588 27740
rect 4628 27700 4637 27740
rect 9763 27616 9772 27656
rect 9812 27616 14476 27656
rect 14516 27616 14525 27656
rect 1699 27448 1708 27488
rect 1748 27448 7564 27488
rect 7604 27448 7613 27488
rect 7171 27364 7180 27404
rect 7220 27364 17164 27404
rect 17204 27364 17213 27404
rect 3679 27259 4065 27278
rect 3679 27236 3745 27259
rect 3831 27236 3913 27259
rect 3999 27236 4065 27259
rect 3679 27196 3688 27236
rect 3728 27196 3745 27236
rect 3831 27196 3852 27236
rect 3892 27196 3913 27236
rect 3999 27196 4016 27236
rect 4056 27196 4065 27236
rect 3679 27173 3745 27196
rect 3831 27173 3913 27196
rect 3999 27173 4065 27196
rect 3679 27154 4065 27173
rect 18799 27259 19185 27278
rect 18799 27236 18865 27259
rect 18951 27236 19033 27259
rect 19119 27236 19185 27259
rect 18799 27196 18808 27236
rect 18848 27196 18865 27236
rect 18951 27196 18972 27236
rect 19012 27196 19033 27236
rect 19119 27196 19136 27236
rect 19176 27196 19185 27236
rect 18799 27173 18865 27196
rect 18951 27173 19033 27196
rect 19119 27173 19185 27196
rect 18799 27154 19185 27173
rect 3043 26860 3052 26900
rect 3092 26860 6412 26900
rect 6452 26860 6461 26900
rect 835 26608 844 26648
rect 884 26608 20620 26648
rect 20660 26608 20669 26648
rect 4919 26503 5305 26522
rect 4919 26480 4985 26503
rect 5071 26480 5153 26503
rect 5239 26480 5305 26503
rect 4919 26440 4928 26480
rect 4968 26440 4985 26480
rect 5071 26440 5092 26480
rect 5132 26440 5153 26480
rect 5239 26440 5256 26480
rect 5296 26440 5305 26480
rect 4919 26417 4985 26440
rect 5071 26417 5153 26440
rect 5239 26417 5305 26440
rect 4919 26398 5305 26417
rect 20039 26503 20425 26522
rect 20039 26480 20105 26503
rect 20191 26480 20273 26503
rect 20359 26480 20425 26503
rect 20039 26440 20048 26480
rect 20088 26440 20105 26480
rect 20191 26440 20212 26480
rect 20252 26440 20273 26480
rect 20359 26440 20376 26480
rect 20416 26440 20425 26480
rect 20039 26417 20105 26440
rect 20191 26417 20273 26440
rect 20359 26417 20425 26440
rect 20039 26398 20425 26417
rect 2371 26020 2380 26060
rect 2420 26020 7756 26060
rect 7796 26020 7805 26060
rect 4483 25936 4492 25976
rect 4532 25936 6412 25976
rect 6452 25936 6461 25976
rect 3679 25747 4065 25766
rect 3679 25724 3745 25747
rect 3831 25724 3913 25747
rect 3999 25724 4065 25747
rect 3679 25684 3688 25724
rect 3728 25684 3745 25724
rect 3831 25684 3852 25724
rect 3892 25684 3913 25724
rect 3999 25684 4016 25724
rect 4056 25684 4065 25724
rect 3679 25661 3745 25684
rect 3831 25661 3913 25684
rect 3999 25661 4065 25684
rect 3679 25642 4065 25661
rect 18799 25747 19185 25766
rect 18799 25724 18865 25747
rect 18951 25724 19033 25747
rect 19119 25724 19185 25747
rect 18799 25684 18808 25724
rect 18848 25684 18865 25724
rect 18951 25684 18972 25724
rect 19012 25684 19033 25724
rect 19119 25684 19136 25724
rect 19176 25684 19185 25724
rect 18799 25661 18865 25684
rect 18951 25661 19033 25684
rect 19119 25661 19185 25684
rect 18799 25642 19185 25661
rect 13946 25243 14070 25262
rect 13946 25220 13965 25243
rect 12355 25180 12364 25220
rect 12404 25180 13965 25220
rect 13946 25157 13965 25180
rect 14051 25157 14070 25243
rect 13946 25138 14070 25157
rect 4919 24991 5305 25010
rect 4919 24968 4985 24991
rect 5071 24968 5153 24991
rect 5239 24968 5305 24991
rect 4919 24928 4928 24968
rect 4968 24928 4985 24968
rect 5071 24928 5092 24968
rect 5132 24928 5153 24968
rect 5239 24928 5256 24968
rect 5296 24928 5305 24968
rect 4919 24905 4985 24928
rect 5071 24905 5153 24928
rect 5239 24905 5305 24928
rect 4919 24886 5305 24905
rect 20039 24991 20425 25010
rect 20039 24968 20105 24991
rect 20191 24968 20273 24991
rect 20359 24968 20425 24991
rect 20039 24928 20048 24968
rect 20088 24928 20105 24968
rect 20191 24928 20212 24968
rect 20252 24928 20273 24968
rect 20359 24928 20376 24968
rect 20416 24928 20425 24968
rect 20039 24905 20105 24928
rect 20191 24905 20273 24928
rect 20359 24905 20425 24928
rect 20039 24886 20425 24905
rect 10819 24844 10828 24884
rect 10868 24844 17836 24884
rect 17876 24844 17885 24884
rect 12451 24592 12460 24632
rect 12500 24592 20620 24632
rect 20660 24592 20669 24632
rect 11107 24508 11116 24548
rect 11156 24508 20812 24548
rect 20852 24508 20861 24548
rect 3679 24235 4065 24254
rect 3679 24212 3745 24235
rect 3831 24212 3913 24235
rect 3999 24212 4065 24235
rect 3679 24172 3688 24212
rect 3728 24172 3745 24212
rect 3831 24172 3852 24212
rect 3892 24172 3913 24212
rect 3999 24172 4016 24212
rect 4056 24172 4065 24212
rect 3679 24149 3745 24172
rect 3831 24149 3913 24172
rect 3999 24149 4065 24172
rect 3679 24130 4065 24149
rect 18799 24235 19185 24254
rect 18799 24212 18865 24235
rect 18951 24212 19033 24235
rect 19119 24212 19185 24235
rect 18799 24172 18808 24212
rect 18848 24172 18865 24212
rect 18951 24172 18972 24212
rect 19012 24172 19033 24212
rect 19119 24172 19136 24212
rect 19176 24172 19185 24212
rect 18799 24149 18865 24172
rect 18951 24149 19033 24172
rect 19119 24149 19185 24172
rect 18799 24130 19185 24149
rect 7747 23920 7756 23960
rect 7796 23920 8812 23960
rect 8852 23920 8861 23960
rect 547 23836 556 23876
rect 596 23836 11360 23876
rect 11320 23792 11360 23836
rect 355 23752 364 23792
rect 404 23752 2764 23792
rect 2804 23752 2813 23792
rect 11320 23752 20140 23792
rect 20180 23752 20189 23792
rect 8995 23668 9004 23708
rect 9044 23668 14764 23708
rect 14804 23668 14813 23708
rect 4919 23479 5305 23498
rect 4919 23456 4985 23479
rect 5071 23456 5153 23479
rect 5239 23456 5305 23479
rect 20039 23479 20425 23498
rect 20039 23456 20105 23479
rect 20191 23456 20273 23479
rect 20359 23456 20425 23479
rect 4919 23416 4928 23456
rect 4968 23416 4985 23456
rect 5071 23416 5092 23456
rect 5132 23416 5153 23456
rect 5239 23416 5256 23456
rect 5296 23416 5305 23456
rect 16483 23416 16492 23456
rect 16532 23416 17260 23456
rect 17300 23416 17309 23456
rect 20039 23416 20048 23456
rect 20088 23416 20105 23456
rect 20191 23416 20212 23456
rect 20252 23416 20273 23456
rect 20359 23416 20376 23456
rect 20416 23416 20425 23456
rect 4919 23393 4985 23416
rect 5071 23393 5153 23416
rect 5239 23393 5305 23416
rect 4919 23374 5305 23393
rect 20039 23393 20105 23416
rect 20191 23393 20273 23416
rect 20359 23393 20425 23416
rect 20039 23374 20425 23393
rect 3679 22723 4065 22742
rect 3679 22700 3745 22723
rect 3831 22700 3913 22723
rect 3999 22700 4065 22723
rect 18799 22723 19185 22742
rect 18799 22700 18865 22723
rect 18951 22700 19033 22723
rect 19119 22700 19185 22723
rect 3679 22660 3688 22700
rect 3728 22660 3745 22700
rect 3831 22660 3852 22700
rect 3892 22660 3913 22700
rect 3999 22660 4016 22700
rect 4056 22660 4065 22700
rect 11971 22660 11980 22700
rect 12020 22660 16396 22700
rect 16436 22660 16445 22700
rect 18799 22660 18808 22700
rect 18848 22660 18865 22700
rect 18951 22660 18972 22700
rect 19012 22660 19033 22700
rect 19119 22660 19136 22700
rect 19176 22660 19185 22700
rect 3679 22637 3745 22660
rect 3831 22637 3913 22660
rect 3999 22637 4065 22660
rect 3679 22618 4065 22637
rect 18799 22637 18865 22660
rect 18951 22637 19033 22660
rect 19119 22637 19185 22660
rect 18799 22618 19185 22637
rect 8131 22408 8140 22448
rect 8180 22408 20140 22448
rect 20180 22408 20189 22448
rect 4919 21967 5305 21986
rect 4919 21944 4985 21967
rect 5071 21944 5153 21967
rect 5239 21944 5305 21967
rect 4919 21904 4928 21944
rect 4968 21904 4985 21944
rect 5071 21904 5092 21944
rect 5132 21904 5153 21944
rect 5239 21904 5256 21944
rect 5296 21904 5305 21944
rect 4919 21881 4985 21904
rect 5071 21881 5153 21904
rect 5239 21881 5305 21904
rect 4919 21862 5305 21881
rect 20039 21967 20425 21986
rect 20039 21944 20105 21967
rect 20191 21944 20273 21967
rect 20359 21944 20425 21967
rect 20039 21904 20048 21944
rect 20088 21904 20105 21944
rect 20191 21904 20212 21944
rect 20252 21904 20273 21944
rect 20359 21904 20376 21944
rect 20416 21904 20425 21944
rect 20039 21881 20105 21904
rect 20191 21881 20273 21904
rect 20359 21881 20425 21904
rect 20039 21862 20425 21881
rect 15043 21736 15052 21776
rect 15092 21736 20140 21776
rect 20180 21736 20189 21776
rect 3679 21211 4065 21230
rect 3679 21188 3745 21211
rect 3831 21188 3913 21211
rect 3999 21188 4065 21211
rect 3679 21148 3688 21188
rect 3728 21148 3745 21188
rect 3831 21148 3852 21188
rect 3892 21148 3913 21188
rect 3999 21148 4016 21188
rect 4056 21148 4065 21188
rect 3679 21125 3745 21148
rect 3831 21125 3913 21148
rect 3999 21125 4065 21148
rect 3679 21106 4065 21125
rect 18799 21211 19185 21230
rect 18799 21188 18865 21211
rect 18951 21188 19033 21211
rect 19119 21188 19185 21211
rect 18799 21148 18808 21188
rect 18848 21148 18865 21188
rect 18951 21148 18972 21188
rect 19012 21148 19033 21188
rect 19119 21148 19136 21188
rect 19176 21148 19185 21188
rect 18799 21125 18865 21148
rect 18951 21125 19033 21148
rect 19119 21125 19185 21148
rect 18799 21106 19185 21125
rect 4919 20455 5305 20474
rect 4919 20432 4985 20455
rect 5071 20432 5153 20455
rect 5239 20432 5305 20455
rect 4919 20392 4928 20432
rect 4968 20392 4985 20432
rect 5071 20392 5092 20432
rect 5132 20392 5153 20432
rect 5239 20392 5256 20432
rect 5296 20392 5305 20432
rect 4919 20369 4985 20392
rect 5071 20369 5153 20392
rect 5239 20369 5305 20392
rect 4919 20350 5305 20369
rect 20039 20455 20425 20474
rect 20039 20432 20105 20455
rect 20191 20432 20273 20455
rect 20359 20432 20425 20455
rect 20039 20392 20048 20432
rect 20088 20392 20105 20432
rect 20191 20392 20212 20432
rect 20252 20392 20273 20432
rect 20359 20392 20376 20432
rect 20416 20392 20425 20432
rect 20039 20369 20105 20392
rect 20191 20369 20273 20392
rect 20359 20369 20425 20392
rect 20039 20350 20425 20369
rect 12931 20224 12940 20264
rect 12980 20224 13116 20264
rect 13076 20096 13116 20224
rect 13076 20056 13228 20096
rect 13268 20056 13277 20096
rect 3679 19699 4065 19718
rect 3679 19676 3745 19699
rect 3831 19676 3913 19699
rect 3999 19676 4065 19699
rect 3679 19636 3688 19676
rect 3728 19636 3745 19676
rect 3831 19636 3852 19676
rect 3892 19636 3913 19676
rect 3999 19636 4016 19676
rect 4056 19636 4065 19676
rect 3679 19613 3745 19636
rect 3831 19613 3913 19636
rect 3999 19613 4065 19636
rect 3679 19594 4065 19613
rect 18799 19699 19185 19718
rect 18799 19676 18865 19699
rect 18951 19676 19033 19699
rect 19119 19676 19185 19699
rect 18799 19636 18808 19676
rect 18848 19636 18865 19676
rect 18951 19636 18972 19676
rect 19012 19636 19033 19676
rect 19119 19636 19136 19676
rect 19176 19636 19185 19676
rect 18799 19613 18865 19636
rect 18951 19613 19033 19636
rect 19119 19613 19185 19636
rect 18799 19594 19185 19613
rect 4919 18943 5305 18962
rect 4919 18920 4985 18943
rect 5071 18920 5153 18943
rect 5239 18920 5305 18943
rect 4919 18880 4928 18920
rect 4968 18880 4985 18920
rect 5071 18880 5092 18920
rect 5132 18880 5153 18920
rect 5239 18880 5256 18920
rect 5296 18880 5305 18920
rect 4919 18857 4985 18880
rect 5071 18857 5153 18880
rect 5239 18857 5305 18880
rect 4919 18838 5305 18857
rect 20039 18943 20425 18962
rect 20039 18920 20105 18943
rect 20191 18920 20273 18943
rect 20359 18920 20425 18943
rect 20039 18880 20048 18920
rect 20088 18880 20105 18920
rect 20191 18880 20212 18920
rect 20252 18880 20273 18920
rect 20359 18880 20376 18920
rect 20416 18880 20425 18920
rect 20039 18857 20105 18880
rect 20191 18857 20273 18880
rect 20359 18857 20425 18880
rect 20039 18838 20425 18857
rect 3679 18187 4065 18206
rect 3679 18164 3745 18187
rect 3831 18164 3913 18187
rect 3999 18164 4065 18187
rect 3679 18124 3688 18164
rect 3728 18124 3745 18164
rect 3831 18124 3852 18164
rect 3892 18124 3913 18164
rect 3999 18124 4016 18164
rect 4056 18124 4065 18164
rect 3679 18101 3745 18124
rect 3831 18101 3913 18124
rect 3999 18101 4065 18124
rect 3679 18082 4065 18101
rect 18799 18187 19185 18206
rect 18799 18164 18865 18187
rect 18951 18164 19033 18187
rect 19119 18164 19185 18187
rect 18799 18124 18808 18164
rect 18848 18124 18865 18164
rect 18951 18124 18972 18164
rect 19012 18124 19033 18164
rect 19119 18124 19136 18164
rect 19176 18124 19185 18164
rect 18799 18101 18865 18124
rect 18951 18101 19033 18124
rect 19119 18101 19185 18124
rect 18799 18082 19185 18101
rect 4919 17431 5305 17450
rect 4919 17408 4985 17431
rect 5071 17408 5153 17431
rect 5239 17408 5305 17431
rect 4919 17368 4928 17408
rect 4968 17368 4985 17408
rect 5071 17368 5092 17408
rect 5132 17368 5153 17408
rect 5239 17368 5256 17408
rect 5296 17368 5305 17408
rect 4919 17345 4985 17368
rect 5071 17345 5153 17368
rect 5239 17345 5305 17368
rect 4919 17326 5305 17345
rect 20039 17431 20425 17450
rect 20039 17408 20105 17431
rect 20191 17408 20273 17431
rect 20359 17408 20425 17431
rect 20039 17368 20048 17408
rect 20088 17368 20105 17408
rect 20191 17368 20212 17408
rect 20252 17368 20273 17408
rect 20359 17368 20376 17408
rect 20416 17368 20425 17408
rect 20039 17345 20105 17368
rect 20191 17345 20273 17368
rect 20359 17345 20425 17368
rect 20039 17326 20425 17345
rect 3679 16675 4065 16694
rect 3679 16652 3745 16675
rect 3831 16652 3913 16675
rect 3999 16652 4065 16675
rect 3679 16612 3688 16652
rect 3728 16612 3745 16652
rect 3831 16612 3852 16652
rect 3892 16612 3913 16652
rect 3999 16612 4016 16652
rect 4056 16612 4065 16652
rect 3679 16589 3745 16612
rect 3831 16589 3913 16612
rect 3999 16589 4065 16612
rect 3679 16570 4065 16589
rect 18799 16675 19185 16694
rect 18799 16652 18865 16675
rect 18951 16652 19033 16675
rect 19119 16652 19185 16675
rect 18799 16612 18808 16652
rect 18848 16612 18865 16652
rect 18951 16612 18972 16652
rect 19012 16612 19033 16652
rect 19119 16612 19136 16652
rect 19176 16612 19185 16652
rect 18799 16589 18865 16612
rect 18951 16589 19033 16612
rect 19119 16589 19185 16612
rect 18799 16570 19185 16589
rect 4919 15919 5305 15938
rect 4919 15896 4985 15919
rect 5071 15896 5153 15919
rect 5239 15896 5305 15919
rect 4919 15856 4928 15896
rect 4968 15856 4985 15896
rect 5071 15856 5092 15896
rect 5132 15856 5153 15896
rect 5239 15856 5256 15896
rect 5296 15856 5305 15896
rect 4919 15833 4985 15856
rect 5071 15833 5153 15856
rect 5239 15833 5305 15856
rect 4919 15814 5305 15833
rect 20039 15919 20425 15938
rect 20039 15896 20105 15919
rect 20191 15896 20273 15919
rect 20359 15896 20425 15919
rect 20039 15856 20048 15896
rect 20088 15856 20105 15896
rect 20191 15856 20212 15896
rect 20252 15856 20273 15896
rect 20359 15856 20376 15896
rect 20416 15856 20425 15896
rect 20039 15833 20105 15856
rect 20191 15833 20273 15856
rect 20359 15833 20425 15856
rect 20039 15814 20425 15833
rect 3679 15163 4065 15182
rect 3679 15140 3745 15163
rect 3831 15140 3913 15163
rect 3999 15140 4065 15163
rect 3679 15100 3688 15140
rect 3728 15100 3745 15140
rect 3831 15100 3852 15140
rect 3892 15100 3913 15140
rect 3999 15100 4016 15140
rect 4056 15100 4065 15140
rect 3679 15077 3745 15100
rect 3831 15077 3913 15100
rect 3999 15077 4065 15100
rect 3679 15058 4065 15077
rect 18799 15163 19185 15182
rect 18799 15140 18865 15163
rect 18951 15140 19033 15163
rect 19119 15140 19185 15163
rect 18799 15100 18808 15140
rect 18848 15100 18865 15140
rect 18951 15100 18972 15140
rect 19012 15100 19033 15140
rect 19119 15100 19136 15140
rect 19176 15100 19185 15140
rect 18799 15077 18865 15100
rect 18951 15077 19033 15100
rect 19119 15077 19185 15100
rect 18799 15058 19185 15077
rect 12067 15016 12076 15056
rect 12116 15016 16108 15056
rect 16148 15016 16157 15056
rect 1219 14512 1228 14552
rect 1268 14512 8812 14552
rect 8852 14512 8861 14552
rect 4919 14407 5305 14426
rect 4919 14384 4985 14407
rect 5071 14384 5153 14407
rect 5239 14384 5305 14407
rect 4919 14344 4928 14384
rect 4968 14344 4985 14384
rect 5071 14344 5092 14384
rect 5132 14344 5153 14384
rect 5239 14344 5256 14384
rect 5296 14344 5305 14384
rect 4919 14321 4985 14344
rect 5071 14321 5153 14344
rect 5239 14321 5305 14344
rect 4919 14302 5305 14321
rect 20039 14407 20425 14426
rect 20039 14384 20105 14407
rect 20191 14384 20273 14407
rect 20359 14384 20425 14407
rect 20039 14344 20048 14384
rect 20088 14344 20105 14384
rect 20191 14344 20212 14384
rect 20252 14344 20273 14384
rect 20359 14344 20376 14384
rect 20416 14344 20425 14384
rect 20039 14321 20105 14344
rect 20191 14321 20273 14344
rect 20359 14321 20425 14344
rect 20039 14302 20425 14321
rect 3679 13651 4065 13670
rect 3679 13628 3745 13651
rect 3831 13628 3913 13651
rect 3999 13628 4065 13651
rect 3679 13588 3688 13628
rect 3728 13588 3745 13628
rect 3831 13588 3852 13628
rect 3892 13588 3913 13628
rect 3999 13588 4016 13628
rect 4056 13588 4065 13628
rect 3679 13565 3745 13588
rect 3831 13565 3913 13588
rect 3999 13565 4065 13588
rect 3679 13546 4065 13565
rect 18799 13651 19185 13670
rect 18799 13628 18865 13651
rect 18951 13628 19033 13651
rect 19119 13628 19185 13651
rect 18799 13588 18808 13628
rect 18848 13588 18865 13628
rect 18951 13588 18972 13628
rect 19012 13588 19033 13628
rect 19119 13588 19136 13628
rect 19176 13588 19185 13628
rect 18799 13565 18865 13588
rect 18951 13565 19033 13588
rect 19119 13565 19185 13588
rect 18799 13546 19185 13565
rect 4919 12895 5305 12914
rect 4919 12872 4985 12895
rect 5071 12872 5153 12895
rect 5239 12872 5305 12895
rect 4919 12832 4928 12872
rect 4968 12832 4985 12872
rect 5071 12832 5092 12872
rect 5132 12832 5153 12872
rect 5239 12832 5256 12872
rect 5296 12832 5305 12872
rect 4919 12809 4985 12832
rect 5071 12809 5153 12832
rect 5239 12809 5305 12832
rect 4919 12790 5305 12809
rect 20039 12895 20425 12914
rect 20039 12872 20105 12895
rect 20191 12872 20273 12895
rect 20359 12872 20425 12895
rect 20039 12832 20048 12872
rect 20088 12832 20105 12872
rect 20191 12832 20212 12872
rect 20252 12832 20273 12872
rect 20359 12832 20376 12872
rect 20416 12832 20425 12872
rect 20039 12809 20105 12832
rect 20191 12809 20273 12832
rect 20359 12809 20425 12832
rect 20039 12790 20425 12809
rect 6979 12580 6988 12620
rect 7028 12580 8812 12620
rect 8852 12580 8861 12620
rect 3679 12139 4065 12158
rect 3679 12116 3745 12139
rect 3831 12116 3913 12139
rect 3999 12116 4065 12139
rect 3679 12076 3688 12116
rect 3728 12076 3745 12116
rect 3831 12076 3852 12116
rect 3892 12076 3913 12116
rect 3999 12076 4016 12116
rect 4056 12076 4065 12116
rect 3679 12053 3745 12076
rect 3831 12053 3913 12076
rect 3999 12053 4065 12076
rect 3679 12034 4065 12053
rect 18799 12139 19185 12158
rect 18799 12116 18865 12139
rect 18951 12116 19033 12139
rect 19119 12116 19185 12139
rect 18799 12076 18808 12116
rect 18848 12076 18865 12116
rect 18951 12076 18972 12116
rect 19012 12076 19033 12116
rect 19119 12076 19136 12116
rect 19176 12076 19185 12116
rect 18799 12053 18865 12076
rect 18951 12053 19033 12076
rect 19119 12053 19185 12076
rect 18799 12034 19185 12053
rect 4919 11383 5305 11402
rect 4919 11360 4985 11383
rect 5071 11360 5153 11383
rect 5239 11360 5305 11383
rect 4919 11320 4928 11360
rect 4968 11320 4985 11360
rect 5071 11320 5092 11360
rect 5132 11320 5153 11360
rect 5239 11320 5256 11360
rect 5296 11320 5305 11360
rect 4919 11297 4985 11320
rect 5071 11297 5153 11320
rect 5239 11297 5305 11320
rect 4919 11278 5305 11297
rect 20039 11383 20425 11402
rect 20039 11360 20105 11383
rect 20191 11360 20273 11383
rect 20359 11360 20425 11383
rect 20039 11320 20048 11360
rect 20088 11320 20105 11360
rect 20191 11320 20212 11360
rect 20252 11320 20273 11360
rect 20359 11320 20376 11360
rect 20416 11320 20425 11360
rect 20039 11297 20105 11320
rect 20191 11297 20273 11320
rect 20359 11297 20425 11320
rect 20039 11278 20425 11297
rect 1027 10900 1036 10940
rect 1076 10900 3436 10940
rect 3476 10900 4876 10940
rect 4916 10900 4925 10940
rect 3679 10627 4065 10646
rect 3679 10604 3745 10627
rect 3831 10604 3913 10627
rect 3999 10604 4065 10627
rect 3679 10564 3688 10604
rect 3728 10564 3745 10604
rect 3831 10564 3852 10604
rect 3892 10564 3913 10604
rect 3999 10564 4016 10604
rect 4056 10564 4065 10604
rect 3679 10541 3745 10564
rect 3831 10541 3913 10564
rect 3999 10541 4065 10564
rect 3679 10522 4065 10541
rect 18799 10627 19185 10646
rect 18799 10604 18865 10627
rect 18951 10604 19033 10627
rect 19119 10604 19185 10627
rect 18799 10564 18808 10604
rect 18848 10564 18865 10604
rect 18951 10564 18972 10604
rect 19012 10564 19033 10604
rect 19119 10564 19136 10604
rect 19176 10564 19185 10604
rect 18799 10541 18865 10564
rect 18951 10541 19033 10564
rect 19119 10541 19185 10564
rect 18799 10522 19185 10541
rect 4919 9871 5305 9890
rect 4919 9848 4985 9871
rect 5071 9848 5153 9871
rect 5239 9848 5305 9871
rect 4919 9808 4928 9848
rect 4968 9808 4985 9848
rect 5071 9808 5092 9848
rect 5132 9808 5153 9848
rect 5239 9808 5256 9848
rect 5296 9808 5305 9848
rect 4919 9785 4985 9808
rect 5071 9785 5153 9808
rect 5239 9785 5305 9808
rect 4919 9766 5305 9785
rect 20039 9871 20425 9890
rect 20039 9848 20105 9871
rect 20191 9848 20273 9871
rect 20359 9848 20425 9871
rect 20039 9808 20048 9848
rect 20088 9808 20105 9848
rect 20191 9808 20212 9848
rect 20252 9808 20273 9848
rect 20359 9808 20376 9848
rect 20416 9808 20425 9848
rect 20039 9785 20105 9808
rect 20191 9785 20273 9808
rect 20359 9785 20425 9808
rect 20039 9766 20425 9785
rect 3679 9115 4065 9134
rect 3679 9092 3745 9115
rect 3831 9092 3913 9115
rect 3999 9092 4065 9115
rect 3679 9052 3688 9092
rect 3728 9052 3745 9092
rect 3831 9052 3852 9092
rect 3892 9052 3913 9092
rect 3999 9052 4016 9092
rect 4056 9052 4065 9092
rect 3679 9029 3745 9052
rect 3831 9029 3913 9052
rect 3999 9029 4065 9052
rect 3679 9010 4065 9029
rect 18799 9115 19185 9134
rect 18799 9092 18865 9115
rect 18951 9092 19033 9115
rect 19119 9092 19185 9115
rect 18799 9052 18808 9092
rect 18848 9052 18865 9092
rect 18951 9052 18972 9092
rect 19012 9052 19033 9092
rect 19119 9052 19136 9092
rect 19176 9052 19185 9092
rect 18799 9029 18865 9052
rect 18951 9029 19033 9052
rect 19119 9029 19185 9052
rect 18799 9010 19185 9029
rect 4919 8359 5305 8378
rect 4919 8336 4985 8359
rect 5071 8336 5153 8359
rect 5239 8336 5305 8359
rect 4919 8296 4928 8336
rect 4968 8296 4985 8336
rect 5071 8296 5092 8336
rect 5132 8296 5153 8336
rect 5239 8296 5256 8336
rect 5296 8296 5305 8336
rect 4919 8273 4985 8296
rect 5071 8273 5153 8296
rect 5239 8273 5305 8296
rect 4919 8254 5305 8273
rect 20039 8359 20425 8378
rect 20039 8336 20105 8359
rect 20191 8336 20273 8359
rect 20359 8336 20425 8359
rect 20039 8296 20048 8336
rect 20088 8296 20105 8336
rect 20191 8296 20212 8336
rect 20252 8296 20273 8336
rect 20359 8296 20376 8336
rect 20416 8296 20425 8336
rect 20039 8273 20105 8296
rect 20191 8273 20273 8296
rect 20359 8273 20425 8296
rect 20039 8254 20425 8273
rect 3679 7603 4065 7622
rect 3679 7580 3745 7603
rect 3831 7580 3913 7603
rect 3999 7580 4065 7603
rect 3679 7540 3688 7580
rect 3728 7540 3745 7580
rect 3831 7540 3852 7580
rect 3892 7540 3913 7580
rect 3999 7540 4016 7580
rect 4056 7540 4065 7580
rect 3679 7517 3745 7540
rect 3831 7517 3913 7540
rect 3999 7517 4065 7540
rect 3679 7498 4065 7517
rect 18799 7603 19185 7622
rect 18799 7580 18865 7603
rect 18951 7580 19033 7603
rect 19119 7580 19185 7603
rect 18799 7540 18808 7580
rect 18848 7540 18865 7580
rect 18951 7540 18972 7580
rect 19012 7540 19033 7580
rect 19119 7540 19136 7580
rect 19176 7540 19185 7580
rect 18799 7517 18865 7540
rect 18951 7517 19033 7540
rect 19119 7517 19185 7540
rect 18799 7498 19185 7517
rect 9842 7435 9966 7454
rect 9842 7412 9861 7435
rect 9571 7372 9580 7412
rect 9620 7372 9861 7412
rect 9842 7349 9861 7372
rect 9947 7349 9966 7435
rect 9842 7330 9966 7349
rect 4919 6847 5305 6866
rect 4919 6824 4985 6847
rect 5071 6824 5153 6847
rect 5239 6824 5305 6847
rect 4919 6784 4928 6824
rect 4968 6784 4985 6824
rect 5071 6784 5092 6824
rect 5132 6784 5153 6824
rect 5239 6784 5256 6824
rect 5296 6784 5305 6824
rect 4919 6761 4985 6784
rect 5071 6761 5153 6784
rect 5239 6761 5305 6784
rect 4919 6742 5305 6761
rect 20039 6847 20425 6866
rect 20039 6824 20105 6847
rect 20191 6824 20273 6847
rect 20359 6824 20425 6847
rect 20039 6784 20048 6824
rect 20088 6784 20105 6824
rect 20191 6784 20212 6824
rect 20252 6784 20273 6824
rect 20359 6784 20376 6824
rect 20416 6784 20425 6824
rect 20039 6761 20105 6784
rect 20191 6761 20273 6784
rect 20359 6761 20425 6784
rect 20039 6742 20425 6761
rect 3679 6091 4065 6110
rect 3679 6068 3745 6091
rect 3831 6068 3913 6091
rect 3999 6068 4065 6091
rect 3679 6028 3688 6068
rect 3728 6028 3745 6068
rect 3831 6028 3852 6068
rect 3892 6028 3913 6068
rect 3999 6028 4016 6068
rect 4056 6028 4065 6068
rect 3679 6005 3745 6028
rect 3831 6005 3913 6028
rect 3999 6005 4065 6028
rect 3679 5986 4065 6005
rect 18799 6091 19185 6110
rect 18799 6068 18865 6091
rect 18951 6068 19033 6091
rect 19119 6068 19185 6091
rect 18799 6028 18808 6068
rect 18848 6028 18865 6068
rect 18951 6028 18972 6068
rect 19012 6028 19033 6068
rect 19119 6028 19136 6068
rect 19176 6028 19185 6068
rect 18799 6005 18865 6028
rect 18951 6005 19033 6028
rect 19119 6005 19185 6028
rect 18799 5986 19185 6005
rect 10754 5671 10878 5690
rect 10754 5648 10773 5671
rect 10723 5608 10732 5648
rect 10772 5608 10773 5648
rect 10754 5585 10773 5608
rect 10859 5585 10878 5671
rect 10754 5566 10878 5585
rect 4919 5335 5305 5354
rect 4919 5312 4985 5335
rect 5071 5312 5153 5335
rect 5239 5312 5305 5335
rect 4919 5272 4928 5312
rect 4968 5272 4985 5312
rect 5071 5272 5092 5312
rect 5132 5272 5153 5312
rect 5239 5272 5256 5312
rect 5296 5272 5305 5312
rect 4919 5249 4985 5272
rect 5071 5249 5153 5272
rect 5239 5249 5305 5272
rect 4919 5230 5305 5249
rect 20039 5335 20425 5354
rect 20039 5312 20105 5335
rect 20191 5312 20273 5335
rect 20359 5312 20425 5335
rect 20039 5272 20048 5312
rect 20088 5272 20105 5312
rect 20191 5272 20212 5312
rect 20252 5272 20273 5312
rect 20359 5272 20376 5312
rect 20416 5272 20425 5312
rect 20039 5249 20105 5272
rect 20191 5249 20273 5272
rect 20359 5249 20425 5272
rect 20039 5230 20425 5249
rect 6650 4831 6774 4850
rect 6650 4745 6669 4831
rect 6755 4808 6774 4831
rect 6755 4768 6796 4808
rect 6836 4768 6845 4808
rect 6755 4745 6774 4768
rect 6650 4726 6774 4745
rect 3679 4579 4065 4598
rect 3679 4556 3745 4579
rect 3831 4556 3913 4579
rect 3999 4556 4065 4579
rect 18799 4579 19185 4598
rect 18799 4556 18865 4579
rect 18951 4556 19033 4579
rect 19119 4556 19185 4579
rect 3679 4516 3688 4556
rect 3728 4516 3745 4556
rect 3831 4516 3852 4556
rect 3892 4516 3913 4556
rect 3999 4516 4016 4556
rect 4056 4516 4065 4556
rect 4195 4516 4204 4556
rect 4244 4516 4972 4556
rect 5012 4516 7660 4556
rect 7700 4516 7709 4556
rect 18799 4516 18808 4556
rect 18848 4516 18865 4556
rect 18951 4516 18972 4556
rect 19012 4516 19033 4556
rect 19119 4516 19136 4556
rect 19176 4516 19185 4556
rect 3679 4493 3745 4516
rect 3831 4493 3913 4516
rect 3999 4493 4065 4516
rect 3679 4474 4065 4493
rect 18799 4493 18865 4516
rect 18951 4493 19033 4516
rect 19119 4493 19185 4516
rect 18799 4474 19185 4493
rect 4919 3823 5305 3842
rect 4919 3800 4985 3823
rect 5071 3800 5153 3823
rect 5239 3800 5305 3823
rect 4919 3760 4928 3800
rect 4968 3760 4985 3800
rect 5071 3760 5092 3800
rect 5132 3760 5153 3800
rect 5239 3760 5256 3800
rect 5296 3760 5305 3800
rect 4919 3737 4985 3760
rect 5071 3737 5153 3760
rect 5239 3737 5305 3760
rect 4919 3718 5305 3737
rect 20039 3823 20425 3842
rect 20039 3800 20105 3823
rect 20191 3800 20273 3823
rect 20359 3800 20425 3823
rect 20039 3760 20048 3800
rect 20088 3760 20105 3800
rect 20191 3760 20212 3800
rect 20252 3760 20273 3800
rect 20359 3760 20376 3800
rect 20416 3760 20425 3800
rect 20039 3737 20105 3760
rect 20191 3737 20273 3760
rect 20359 3737 20425 3760
rect 20039 3718 20425 3737
rect 2090 3655 2214 3674
rect 2090 3632 2109 3655
rect 2083 3592 2092 3632
rect 2090 3569 2109 3592
rect 2195 3569 2214 3655
rect 2090 3550 2214 3569
rect 3679 3067 4065 3086
rect 3679 3044 3745 3067
rect 3831 3044 3913 3067
rect 3999 3044 4065 3067
rect 3679 3004 3688 3044
rect 3728 3004 3745 3044
rect 3831 3004 3852 3044
rect 3892 3004 3913 3044
rect 3999 3004 4016 3044
rect 4056 3004 4065 3044
rect 3679 2981 3745 3004
rect 3831 2981 3913 3004
rect 3999 2981 4065 3004
rect 3679 2962 4065 2981
rect 18799 3067 19185 3086
rect 18799 3044 18865 3067
rect 18951 3044 19033 3067
rect 19119 3044 19185 3067
rect 18799 3004 18808 3044
rect 18848 3004 18865 3044
rect 18951 3004 18972 3044
rect 19012 3004 19033 3044
rect 19119 3004 19136 3044
rect 19176 3004 19185 3044
rect 18799 2981 18865 3004
rect 18951 2981 19033 3004
rect 19119 2981 19185 3004
rect 18799 2962 19185 2981
rect 451 2836 460 2876
rect 500 2836 7564 2876
rect 7604 2836 10540 2876
rect 10580 2836 10589 2876
rect 3619 2752 3628 2792
rect 3668 2752 7276 2792
rect 7316 2752 7325 2792
rect 4919 2311 5305 2330
rect 4919 2288 4985 2311
rect 5071 2288 5153 2311
rect 5239 2288 5305 2311
rect 4919 2248 4928 2288
rect 4968 2248 4985 2288
rect 5071 2248 5092 2288
rect 5132 2248 5153 2288
rect 5239 2248 5256 2288
rect 5296 2248 5305 2288
rect 4919 2225 4985 2248
rect 5071 2225 5153 2248
rect 5239 2225 5305 2248
rect 4919 2206 5305 2225
rect 20039 2311 20425 2330
rect 20039 2288 20105 2311
rect 20191 2288 20273 2311
rect 20359 2288 20425 2311
rect 20039 2248 20048 2288
rect 20088 2248 20105 2288
rect 20191 2248 20212 2288
rect 20252 2248 20273 2288
rect 20359 2248 20376 2288
rect 20416 2248 20425 2288
rect 20039 2225 20105 2248
rect 20191 2225 20273 2248
rect 20359 2225 20425 2248
rect 20039 2206 20425 2225
rect 12122 1891 12246 1910
rect 5731 1828 5740 1868
rect 5780 1828 11020 1868
rect 11060 1828 11069 1868
rect 12122 1805 12141 1891
rect 12227 1868 12246 1891
rect 12227 1828 13036 1868
rect 13076 1828 13085 1868
rect 12227 1805 12246 1828
rect 12122 1786 12246 1805
rect 3679 1555 4065 1574
rect 3679 1532 3745 1555
rect 3831 1532 3913 1555
rect 3999 1532 4065 1555
rect 3679 1492 3688 1532
rect 3728 1492 3745 1532
rect 3831 1492 3852 1532
rect 3892 1492 3913 1532
rect 3999 1492 4016 1532
rect 4056 1492 4065 1532
rect 3679 1469 3745 1492
rect 3831 1469 3913 1492
rect 3999 1469 4065 1492
rect 3679 1450 4065 1469
rect 18799 1555 19185 1574
rect 18799 1532 18865 1555
rect 18951 1532 19033 1555
rect 19119 1532 19185 1555
rect 18799 1492 18808 1532
rect 18848 1492 18865 1532
rect 18951 1492 18972 1532
rect 19012 1492 19033 1532
rect 19119 1492 19136 1532
rect 19176 1492 19185 1532
rect 18799 1469 18865 1492
rect 18951 1469 19033 1492
rect 19119 1469 19185 1492
rect 18799 1450 19185 1469
rect 13034 1303 13158 1322
rect 13034 1280 13053 1303
rect 12739 1240 12748 1280
rect 12788 1240 13053 1280
rect 13034 1217 13053 1240
rect 13139 1217 13158 1303
rect 13034 1198 13158 1217
rect 6787 1072 6796 1112
rect 6836 1072 11308 1112
rect 11348 1072 11357 1112
rect 4919 799 5305 818
rect 4919 776 4985 799
rect 5071 776 5153 799
rect 5239 776 5305 799
rect 15770 799 15894 818
rect 15770 776 15789 799
rect 4919 736 4928 776
rect 4968 736 4985 776
rect 5071 736 5092 776
rect 5132 736 5153 776
rect 5239 736 5256 776
rect 5296 736 5305 776
rect 15619 736 15628 776
rect 15668 736 15789 776
rect 4919 713 4985 736
rect 5071 713 5153 736
rect 5239 713 5305 736
rect 4919 694 5305 713
rect 15770 713 15789 736
rect 15875 713 15894 799
rect 20039 799 20425 818
rect 20039 776 20105 799
rect 20191 776 20273 799
rect 20359 776 20425 799
rect 20039 736 20048 776
rect 20088 736 20105 776
rect 20191 736 20212 776
rect 20252 736 20273 776
rect 20359 736 20376 776
rect 20416 736 20425 776
rect 15770 694 15894 713
rect 16682 715 16806 734
rect 16682 629 16701 715
rect 16787 692 16806 715
rect 20039 713 20105 736
rect 20191 713 20273 736
rect 20359 713 20425 736
rect 20039 694 20425 713
rect 16787 652 18892 692
rect 18932 652 18941 692
rect 16787 629 16806 652
rect 16682 610 16806 629
rect 2947 568 2956 608
rect 2996 568 7084 608
rect 7124 568 7133 608
rect 6979 316 6988 356
rect 7028 316 8716 356
rect 8756 316 8765 356
rect 12643 148 12652 188
rect 12692 148 19468 188
rect 19508 148 19517 188
<< via5 >>
rect 3745 84692 3831 84715
rect 3913 84692 3999 84715
rect 3745 84652 3770 84692
rect 3770 84652 3810 84692
rect 3810 84652 3831 84692
rect 3913 84652 3934 84692
rect 3934 84652 3974 84692
rect 3974 84652 3999 84692
rect 3745 84629 3831 84652
rect 3913 84629 3999 84652
rect 18865 84692 18951 84715
rect 19033 84692 19119 84715
rect 18865 84652 18890 84692
rect 18890 84652 18930 84692
rect 18930 84652 18951 84692
rect 19033 84652 19054 84692
rect 19054 84652 19094 84692
rect 19094 84652 19119 84692
rect 18865 84629 18951 84652
rect 19033 84629 19119 84652
rect 12141 84041 12227 84127
rect 4985 83936 5071 83959
rect 5153 83936 5239 83959
rect 4985 83896 5010 83936
rect 5010 83896 5050 83936
rect 5050 83896 5071 83936
rect 5153 83896 5174 83936
rect 5174 83896 5214 83936
rect 5214 83896 5239 83936
rect 4985 83873 5071 83896
rect 5153 83873 5239 83896
rect 20105 83936 20191 83959
rect 20273 83936 20359 83959
rect 20105 83896 20130 83936
rect 20130 83896 20170 83936
rect 20170 83896 20191 83936
rect 20273 83896 20294 83936
rect 20294 83896 20334 83936
rect 20334 83896 20359 83936
rect 20105 83873 20191 83896
rect 20273 83873 20359 83896
rect 10773 83453 10859 83539
rect 13053 83285 13139 83371
rect 3745 83180 3831 83203
rect 3913 83180 3999 83203
rect 18865 83180 18951 83203
rect 19033 83180 19119 83203
rect 3745 83140 3770 83180
rect 3770 83140 3810 83180
rect 3810 83140 3831 83180
rect 3913 83140 3934 83180
rect 3934 83140 3974 83180
rect 3974 83140 3999 83180
rect 18865 83140 18890 83180
rect 18890 83140 18930 83180
rect 18930 83140 18951 83180
rect 19033 83140 19054 83180
rect 19054 83140 19094 83180
rect 19094 83140 19119 83180
rect 3745 83117 3831 83140
rect 3913 83117 3999 83140
rect 18865 83117 18951 83140
rect 19033 83117 19119 83140
rect 4985 82424 5071 82447
rect 5153 82424 5239 82447
rect 4985 82384 5010 82424
rect 5010 82384 5050 82424
rect 5050 82384 5071 82424
rect 5153 82384 5174 82424
rect 5174 82384 5214 82424
rect 5214 82384 5239 82424
rect 4985 82361 5071 82384
rect 5153 82361 5239 82384
rect 20105 82424 20191 82447
rect 20273 82424 20359 82447
rect 20105 82384 20130 82424
rect 20130 82384 20170 82424
rect 20170 82384 20191 82424
rect 20273 82384 20294 82424
rect 20294 82384 20334 82424
rect 20334 82384 20359 82424
rect 20105 82361 20191 82384
rect 20273 82361 20359 82384
rect 3745 81668 3831 81691
rect 3913 81668 3999 81691
rect 3745 81628 3770 81668
rect 3770 81628 3810 81668
rect 3810 81628 3831 81668
rect 3913 81628 3934 81668
rect 3934 81628 3974 81668
rect 3974 81628 3999 81668
rect 3745 81605 3831 81628
rect 3913 81605 3999 81628
rect 18865 81668 18951 81691
rect 19033 81668 19119 81691
rect 18865 81628 18890 81668
rect 18890 81628 18930 81668
rect 18930 81628 18951 81668
rect 19033 81628 19054 81668
rect 19054 81628 19094 81668
rect 19094 81628 19119 81668
rect 18865 81605 18951 81628
rect 19033 81605 19119 81628
rect 16701 81017 16787 81103
rect 4985 80912 5071 80935
rect 5153 80912 5239 80935
rect 4985 80872 5010 80912
rect 5010 80872 5050 80912
rect 5050 80872 5071 80912
rect 5153 80872 5174 80912
rect 5174 80872 5214 80912
rect 5214 80872 5239 80912
rect 4985 80849 5071 80872
rect 5153 80849 5239 80872
rect 20105 80912 20191 80935
rect 20273 80912 20359 80935
rect 20105 80872 20130 80912
rect 20130 80872 20170 80912
rect 20170 80872 20191 80912
rect 20273 80872 20294 80912
rect 20294 80872 20334 80912
rect 20334 80872 20359 80912
rect 8493 80765 8579 80851
rect 20105 80849 20191 80872
rect 20273 80849 20359 80872
rect 3745 80156 3831 80179
rect 3913 80156 3999 80179
rect 3745 80116 3770 80156
rect 3770 80116 3810 80156
rect 3810 80116 3831 80156
rect 3913 80116 3934 80156
rect 3934 80116 3974 80156
rect 3974 80116 3999 80156
rect 3745 80093 3831 80116
rect 3913 80093 3999 80116
rect 18865 80156 18951 80179
rect 19033 80156 19119 80179
rect 18865 80116 18890 80156
rect 18890 80116 18930 80156
rect 18930 80116 18951 80156
rect 19033 80116 19054 80156
rect 19054 80116 19094 80156
rect 19094 80116 19119 80156
rect 18865 80093 18951 80116
rect 19033 80093 19119 80116
rect 4985 79400 5071 79423
rect 5153 79400 5239 79423
rect 9861 79421 9947 79507
rect 4985 79360 5010 79400
rect 5010 79360 5050 79400
rect 5050 79360 5071 79400
rect 5153 79360 5174 79400
rect 5174 79360 5214 79400
rect 5214 79360 5239 79400
rect 4985 79337 5071 79360
rect 5153 79337 5239 79360
rect 20105 79400 20191 79423
rect 20273 79400 20359 79423
rect 20105 79360 20130 79400
rect 20130 79360 20170 79400
rect 20170 79360 20191 79400
rect 20273 79360 20294 79400
rect 20294 79360 20334 79400
rect 20334 79360 20359 79400
rect 20105 79337 20191 79360
rect 20273 79337 20359 79360
rect 3745 78644 3831 78667
rect 3913 78644 3999 78667
rect 3745 78604 3770 78644
rect 3770 78604 3810 78644
rect 3810 78604 3831 78644
rect 3913 78604 3934 78644
rect 3934 78604 3974 78644
rect 3974 78604 3999 78644
rect 3745 78581 3831 78604
rect 3913 78581 3999 78604
rect 18865 78644 18951 78667
rect 19033 78644 19119 78667
rect 18865 78604 18890 78644
rect 18890 78604 18930 78644
rect 18930 78604 18951 78644
rect 19033 78604 19054 78644
rect 19054 78604 19094 78644
rect 19094 78604 19119 78644
rect 18865 78581 18951 78604
rect 19033 78581 19119 78604
rect 4985 77888 5071 77911
rect 5153 77888 5239 77911
rect 4985 77848 5010 77888
rect 5010 77848 5050 77888
rect 5050 77848 5071 77888
rect 5153 77848 5174 77888
rect 5174 77848 5214 77888
rect 5214 77848 5239 77888
rect 4985 77825 5071 77848
rect 5153 77825 5239 77848
rect 20105 77888 20191 77911
rect 20273 77888 20359 77911
rect 20105 77848 20130 77888
rect 20130 77848 20170 77888
rect 20170 77848 20191 77888
rect 20273 77848 20294 77888
rect 20294 77848 20334 77888
rect 20334 77848 20359 77888
rect 20105 77825 20191 77848
rect 20273 77825 20359 77848
rect 13965 77237 14051 77323
rect 3745 77132 3831 77155
rect 3913 77132 3999 77155
rect 3745 77092 3770 77132
rect 3770 77092 3810 77132
rect 3810 77092 3831 77132
rect 3913 77092 3934 77132
rect 3934 77092 3974 77132
rect 3974 77092 3999 77132
rect 3745 77069 3831 77092
rect 3913 77069 3999 77092
rect 18865 77132 18951 77155
rect 19033 77132 19119 77155
rect 18865 77092 18890 77132
rect 18890 77092 18930 77132
rect 18930 77092 18951 77132
rect 19033 77092 19054 77132
rect 19054 77092 19094 77132
rect 19094 77092 19119 77132
rect 18865 77069 18951 77092
rect 19033 77069 19119 77092
rect 2109 76817 2195 76903
rect 4985 76376 5071 76399
rect 5153 76376 5239 76399
rect 4985 76336 5010 76376
rect 5010 76336 5050 76376
rect 5050 76336 5071 76376
rect 5153 76336 5174 76376
rect 5174 76336 5214 76376
rect 5214 76336 5239 76376
rect 4985 76313 5071 76336
rect 5153 76313 5239 76336
rect 20105 76376 20191 76399
rect 20273 76376 20359 76399
rect 20105 76336 20130 76376
rect 20130 76336 20170 76376
rect 20170 76336 20191 76376
rect 20273 76336 20294 76376
rect 20294 76336 20334 76376
rect 20334 76336 20359 76376
rect 20105 76313 20191 76336
rect 20273 76313 20359 76336
rect 3745 75620 3831 75643
rect 3913 75620 3999 75643
rect 3745 75580 3770 75620
rect 3770 75580 3810 75620
rect 3810 75580 3831 75620
rect 3913 75580 3934 75620
rect 3934 75580 3974 75620
rect 3974 75580 3999 75620
rect 3745 75557 3831 75580
rect 3913 75557 3999 75580
rect 18865 75620 18951 75643
rect 19033 75620 19119 75643
rect 18865 75580 18890 75620
rect 18890 75580 18930 75620
rect 18930 75580 18951 75620
rect 19033 75580 19054 75620
rect 19054 75580 19094 75620
rect 19094 75580 19119 75620
rect 18865 75557 18951 75580
rect 19033 75557 19119 75580
rect 4985 74864 5071 74887
rect 5153 74864 5239 74887
rect 4985 74824 5010 74864
rect 5010 74824 5050 74864
rect 5050 74824 5071 74864
rect 5153 74824 5174 74864
rect 5174 74824 5214 74864
rect 5214 74824 5239 74864
rect 4985 74801 5071 74824
rect 5153 74801 5239 74824
rect 20105 74864 20191 74887
rect 20273 74864 20359 74887
rect 20105 74824 20130 74864
rect 20130 74824 20170 74864
rect 20170 74824 20191 74864
rect 20273 74824 20294 74864
rect 20294 74824 20334 74864
rect 20334 74824 20359 74864
rect 20105 74801 20191 74824
rect 20273 74801 20359 74824
rect 3745 74108 3831 74131
rect 3913 74108 3999 74131
rect 3745 74068 3770 74108
rect 3770 74068 3810 74108
rect 3810 74068 3831 74108
rect 3913 74068 3934 74108
rect 3934 74068 3974 74108
rect 3974 74068 3999 74108
rect 3745 74045 3831 74068
rect 3913 74045 3999 74068
rect 18865 74108 18951 74131
rect 19033 74108 19119 74131
rect 18865 74068 18890 74108
rect 18890 74068 18930 74108
rect 18930 74068 18951 74108
rect 19033 74068 19054 74108
rect 19054 74068 19094 74108
rect 19094 74068 19119 74108
rect 18865 74045 18951 74068
rect 19033 74045 19119 74068
rect 4985 73352 5071 73375
rect 5153 73352 5239 73375
rect 4985 73312 5010 73352
rect 5010 73312 5050 73352
rect 5050 73312 5071 73352
rect 5153 73312 5174 73352
rect 5174 73312 5214 73352
rect 5214 73312 5239 73352
rect 4985 73289 5071 73312
rect 5153 73289 5239 73312
rect 20105 73352 20191 73375
rect 20273 73352 20359 73375
rect 20105 73312 20130 73352
rect 20130 73312 20170 73352
rect 20170 73312 20191 73352
rect 20273 73312 20294 73352
rect 20294 73312 20334 73352
rect 20334 73312 20359 73352
rect 20105 73289 20191 73312
rect 20273 73289 20359 73312
rect 1197 72953 1283 73039
rect 3745 72596 3831 72619
rect 3913 72596 3999 72619
rect 3745 72556 3770 72596
rect 3770 72556 3810 72596
rect 3810 72556 3831 72596
rect 3913 72556 3934 72596
rect 3934 72556 3974 72596
rect 3974 72556 3999 72596
rect 3745 72533 3831 72556
rect 3913 72533 3999 72556
rect 18865 72596 18951 72619
rect 19033 72596 19119 72619
rect 18865 72556 18890 72596
rect 18890 72556 18930 72596
rect 18930 72556 18951 72596
rect 19033 72556 19054 72596
rect 19054 72556 19094 72596
rect 19094 72556 19119 72596
rect 18865 72533 18951 72556
rect 19033 72533 19119 72556
rect 4985 71840 5071 71863
rect 5153 71840 5239 71863
rect 4985 71800 5010 71840
rect 5010 71800 5050 71840
rect 5050 71800 5071 71840
rect 5153 71800 5174 71840
rect 5174 71800 5214 71840
rect 5214 71800 5239 71840
rect 4985 71777 5071 71800
rect 5153 71777 5239 71800
rect 20105 71840 20191 71863
rect 20273 71840 20359 71863
rect 20105 71800 20130 71840
rect 20130 71800 20170 71840
rect 20170 71800 20191 71840
rect 20273 71800 20294 71840
rect 20294 71800 20334 71840
rect 20334 71800 20359 71840
rect 20105 71777 20191 71800
rect 20273 71777 20359 71800
rect 3745 71084 3831 71107
rect 3913 71084 3999 71107
rect 3745 71044 3770 71084
rect 3770 71044 3810 71084
rect 3810 71044 3831 71084
rect 3913 71044 3934 71084
rect 3934 71044 3974 71084
rect 3974 71044 3999 71084
rect 3745 71021 3831 71044
rect 3913 71021 3999 71044
rect 18865 71084 18951 71107
rect 19033 71084 19119 71107
rect 18865 71044 18890 71084
rect 18890 71044 18930 71084
rect 18930 71044 18951 71084
rect 19033 71044 19054 71084
rect 19054 71044 19094 71084
rect 19094 71044 19119 71084
rect 18865 71021 18951 71044
rect 19033 71021 19119 71044
rect 4985 70328 5071 70351
rect 5153 70328 5239 70351
rect 4985 70288 5010 70328
rect 5010 70288 5050 70328
rect 5050 70288 5071 70328
rect 5153 70288 5174 70328
rect 5174 70288 5214 70328
rect 5214 70288 5239 70328
rect 4985 70265 5071 70288
rect 5153 70265 5239 70288
rect 20105 70328 20191 70351
rect 20273 70328 20359 70351
rect 20105 70288 20130 70328
rect 20130 70288 20170 70328
rect 20170 70288 20191 70328
rect 20273 70288 20294 70328
rect 20294 70288 20334 70328
rect 20334 70288 20359 70328
rect 20105 70265 20191 70288
rect 20273 70265 20359 70288
rect 3745 69572 3831 69595
rect 3913 69572 3999 69595
rect 3745 69532 3770 69572
rect 3770 69532 3810 69572
rect 3810 69532 3831 69572
rect 3913 69532 3934 69572
rect 3934 69532 3974 69572
rect 3974 69532 3999 69572
rect 3745 69509 3831 69532
rect 3913 69509 3999 69532
rect 18865 69572 18951 69595
rect 19033 69572 19119 69595
rect 18865 69532 18890 69572
rect 18890 69532 18930 69572
rect 18930 69532 18951 69572
rect 19033 69532 19054 69572
rect 19054 69532 19094 69572
rect 19094 69532 19119 69572
rect 18865 69509 18951 69532
rect 19033 69509 19119 69532
rect 4985 68816 5071 68839
rect 5153 68816 5239 68839
rect 4985 68776 5010 68816
rect 5010 68776 5050 68816
rect 5050 68776 5071 68816
rect 5153 68776 5174 68816
rect 5174 68776 5214 68816
rect 5214 68776 5239 68816
rect 4985 68753 5071 68776
rect 5153 68753 5239 68776
rect 20105 68816 20191 68839
rect 20273 68816 20359 68839
rect 20105 68776 20130 68816
rect 20130 68776 20170 68816
rect 20170 68776 20191 68816
rect 20273 68776 20294 68816
rect 20294 68776 20334 68816
rect 20334 68776 20359 68816
rect 20105 68753 20191 68776
rect 20273 68753 20359 68776
rect 3745 68060 3831 68083
rect 3913 68060 3999 68083
rect 3745 68020 3770 68060
rect 3770 68020 3810 68060
rect 3810 68020 3831 68060
rect 3913 68020 3934 68060
rect 3934 68020 3974 68060
rect 3974 68020 3999 68060
rect 3745 67997 3831 68020
rect 3913 67997 3999 68020
rect 18865 68060 18951 68083
rect 19033 68060 19119 68083
rect 18865 68020 18890 68060
rect 18890 68020 18930 68060
rect 18930 68020 18951 68060
rect 19033 68020 19054 68060
rect 19054 68020 19094 68060
rect 19094 68020 19119 68060
rect 18865 67997 18951 68020
rect 19033 67997 19119 68020
rect 4985 67304 5071 67327
rect 5153 67304 5239 67327
rect 4985 67264 5010 67304
rect 5010 67264 5050 67304
rect 5050 67264 5071 67304
rect 5153 67264 5174 67304
rect 5174 67264 5214 67304
rect 5214 67264 5239 67304
rect 4985 67241 5071 67264
rect 5153 67241 5239 67264
rect 20105 67304 20191 67327
rect 20273 67304 20359 67327
rect 20105 67264 20130 67304
rect 20130 67264 20170 67304
rect 20170 67264 20191 67304
rect 20273 67264 20294 67304
rect 20294 67264 20334 67304
rect 20334 67264 20359 67304
rect 20105 67241 20191 67264
rect 20273 67241 20359 67264
rect 15789 66905 15875 66991
rect 3745 66548 3831 66571
rect 3913 66548 3999 66571
rect 3745 66508 3770 66548
rect 3770 66508 3810 66548
rect 3810 66508 3831 66548
rect 3913 66508 3934 66548
rect 3934 66508 3974 66548
rect 3974 66508 3999 66548
rect 3745 66485 3831 66508
rect 3913 66485 3999 66508
rect 18865 66548 18951 66571
rect 19033 66548 19119 66571
rect 18865 66508 18890 66548
rect 18890 66508 18930 66548
rect 18930 66508 18951 66548
rect 19033 66508 19054 66548
rect 19054 66508 19094 66548
rect 19094 66508 19119 66548
rect 18865 66485 18951 66508
rect 19033 66485 19119 66508
rect 4985 65792 5071 65815
rect 5153 65792 5239 65815
rect 6669 65813 6755 65899
rect 4985 65752 5010 65792
rect 5010 65752 5050 65792
rect 5050 65752 5071 65792
rect 5153 65752 5174 65792
rect 5174 65752 5214 65792
rect 5214 65752 5239 65792
rect 4985 65729 5071 65752
rect 5153 65729 5239 65752
rect 20105 65792 20191 65815
rect 20273 65792 20359 65815
rect 20105 65752 20130 65792
rect 20130 65752 20170 65792
rect 20170 65752 20191 65792
rect 20273 65752 20294 65792
rect 20294 65752 20334 65792
rect 20334 65752 20359 65792
rect 20105 65729 20191 65752
rect 20273 65729 20359 65752
rect 3745 65036 3831 65059
rect 3913 65036 3999 65059
rect 3745 64996 3770 65036
rect 3770 64996 3810 65036
rect 3810 64996 3831 65036
rect 3913 64996 3934 65036
rect 3934 64996 3974 65036
rect 3974 64996 3999 65036
rect 3745 64973 3831 64996
rect 3913 64973 3999 64996
rect 18865 65036 18951 65059
rect 19033 65036 19119 65059
rect 18865 64996 18890 65036
rect 18890 64996 18930 65036
rect 18930 64996 18951 65036
rect 19033 64996 19054 65036
rect 19054 64996 19094 65036
rect 19094 64996 19119 65036
rect 18865 64973 18951 64996
rect 19033 64973 19119 64996
rect 4985 64280 5071 64303
rect 5153 64280 5239 64303
rect 4985 64240 5010 64280
rect 5010 64240 5050 64280
rect 5050 64240 5071 64280
rect 5153 64240 5174 64280
rect 5174 64240 5214 64280
rect 5214 64240 5239 64280
rect 4985 64217 5071 64240
rect 5153 64217 5239 64240
rect 20105 64280 20191 64303
rect 20273 64280 20359 64303
rect 20105 64240 20130 64280
rect 20130 64240 20170 64280
rect 20170 64240 20191 64280
rect 20273 64240 20294 64280
rect 20294 64240 20334 64280
rect 20334 64240 20359 64280
rect 20105 64217 20191 64240
rect 20273 64217 20359 64240
rect 3745 63524 3831 63547
rect 3913 63524 3999 63547
rect 3745 63484 3770 63524
rect 3770 63484 3810 63524
rect 3810 63484 3831 63524
rect 3913 63484 3934 63524
rect 3934 63484 3974 63524
rect 3974 63484 3999 63524
rect 3745 63461 3831 63484
rect 3913 63461 3999 63484
rect 18865 63524 18951 63547
rect 19033 63524 19119 63547
rect 18865 63484 18890 63524
rect 18890 63484 18930 63524
rect 18930 63484 18951 63524
rect 19033 63484 19054 63524
rect 19054 63484 19094 63524
rect 19094 63484 19119 63524
rect 18865 63461 18951 63484
rect 19033 63461 19119 63484
rect 4985 62768 5071 62791
rect 5153 62768 5239 62791
rect 4985 62728 5010 62768
rect 5010 62728 5050 62768
rect 5050 62728 5071 62768
rect 5153 62728 5174 62768
rect 5174 62728 5214 62768
rect 5214 62728 5239 62768
rect 4985 62705 5071 62728
rect 5153 62705 5239 62728
rect 20105 62768 20191 62791
rect 20273 62768 20359 62791
rect 20105 62728 20130 62768
rect 20130 62728 20170 62768
rect 20170 62728 20191 62768
rect 20273 62728 20294 62768
rect 20294 62728 20334 62768
rect 20334 62728 20359 62768
rect 20105 62705 20191 62728
rect 20273 62705 20359 62728
rect 3745 62012 3831 62035
rect 3913 62012 3999 62035
rect 3745 61972 3770 62012
rect 3770 61972 3810 62012
rect 3810 61972 3831 62012
rect 3913 61972 3934 62012
rect 3934 61972 3974 62012
rect 3974 61972 3999 62012
rect 3745 61949 3831 61972
rect 3913 61949 3999 61972
rect 18865 62012 18951 62035
rect 19033 62012 19119 62035
rect 18865 61972 18890 62012
rect 18890 61972 18930 62012
rect 18930 61972 18951 62012
rect 19033 61972 19054 62012
rect 19054 61972 19094 62012
rect 19094 61972 19119 62012
rect 18865 61949 18951 61972
rect 19033 61949 19119 61972
rect 4985 61256 5071 61279
rect 5153 61256 5239 61279
rect 4985 61216 5010 61256
rect 5010 61216 5050 61256
rect 5050 61216 5071 61256
rect 5153 61216 5174 61256
rect 5174 61216 5214 61256
rect 5214 61216 5239 61256
rect 4985 61193 5071 61216
rect 5153 61193 5239 61216
rect 20105 61256 20191 61279
rect 20273 61256 20359 61279
rect 20105 61216 20130 61256
rect 20130 61216 20170 61256
rect 20170 61216 20191 61256
rect 20273 61216 20294 61256
rect 20294 61216 20334 61256
rect 20334 61216 20359 61256
rect 20105 61193 20191 61216
rect 20273 61193 20359 61216
rect 13965 61025 14051 61111
rect 3745 60500 3831 60523
rect 3913 60500 3999 60523
rect 3745 60460 3770 60500
rect 3770 60460 3810 60500
rect 3810 60460 3831 60500
rect 3913 60460 3934 60500
rect 3934 60460 3974 60500
rect 3974 60460 3999 60500
rect 3745 60437 3831 60460
rect 3913 60437 3999 60460
rect 18865 60500 18951 60523
rect 19033 60500 19119 60523
rect 18865 60460 18890 60500
rect 18890 60460 18930 60500
rect 18930 60460 18951 60500
rect 19033 60460 19054 60500
rect 19054 60460 19094 60500
rect 19094 60460 19119 60500
rect 18865 60437 18951 60460
rect 19033 60437 19119 60460
rect 4985 59744 5071 59767
rect 5153 59744 5239 59767
rect 4985 59704 5010 59744
rect 5010 59704 5050 59744
rect 5050 59704 5071 59744
rect 5153 59704 5174 59744
rect 5174 59704 5214 59744
rect 5214 59704 5239 59744
rect 4985 59681 5071 59704
rect 5153 59681 5239 59704
rect 20105 59744 20191 59767
rect 20273 59744 20359 59767
rect 20105 59704 20130 59744
rect 20130 59704 20170 59744
rect 20170 59704 20191 59744
rect 20273 59704 20294 59744
rect 20294 59704 20334 59744
rect 20334 59704 20359 59744
rect 20105 59681 20191 59704
rect 20273 59681 20359 59704
rect 3745 58988 3831 59011
rect 3913 58988 3999 59011
rect 3745 58948 3770 58988
rect 3770 58948 3810 58988
rect 3810 58948 3831 58988
rect 3913 58948 3934 58988
rect 3934 58948 3974 58988
rect 3974 58948 3999 58988
rect 3745 58925 3831 58948
rect 3913 58925 3999 58948
rect 18865 58988 18951 59011
rect 19033 58988 19119 59011
rect 18865 58948 18890 58988
rect 18890 58948 18930 58988
rect 18930 58948 18951 58988
rect 19033 58948 19054 58988
rect 19054 58948 19094 58988
rect 19094 58948 19119 58988
rect 18865 58925 18951 58948
rect 19033 58925 19119 58948
rect 4985 58232 5071 58255
rect 5153 58232 5239 58255
rect 4985 58192 5010 58232
rect 5010 58192 5050 58232
rect 5050 58192 5071 58232
rect 5153 58192 5174 58232
rect 5174 58192 5214 58232
rect 5214 58192 5239 58232
rect 4985 58169 5071 58192
rect 5153 58169 5239 58192
rect 20105 58232 20191 58255
rect 20273 58232 20359 58255
rect 20105 58192 20130 58232
rect 20130 58192 20170 58232
rect 20170 58192 20191 58232
rect 20273 58192 20294 58232
rect 20294 58192 20334 58232
rect 20334 58192 20359 58232
rect 20105 58169 20191 58192
rect 20273 58169 20359 58192
rect 3745 57476 3831 57499
rect 3913 57476 3999 57499
rect 3745 57436 3770 57476
rect 3770 57436 3810 57476
rect 3810 57436 3831 57476
rect 3913 57436 3934 57476
rect 3934 57436 3974 57476
rect 3974 57436 3999 57476
rect 3745 57413 3831 57436
rect 3913 57413 3999 57436
rect 18865 57476 18951 57499
rect 19033 57476 19119 57499
rect 18865 57436 18890 57476
rect 18890 57436 18930 57476
rect 18930 57436 18951 57476
rect 19033 57436 19054 57476
rect 19054 57436 19094 57476
rect 19094 57436 19119 57476
rect 18865 57413 18951 57436
rect 19033 57413 19119 57436
rect 4985 56720 5071 56743
rect 5153 56720 5239 56743
rect 4985 56680 5010 56720
rect 5010 56680 5050 56720
rect 5050 56680 5071 56720
rect 5153 56680 5174 56720
rect 5174 56680 5214 56720
rect 5214 56680 5239 56720
rect 4985 56657 5071 56680
rect 5153 56657 5239 56680
rect 13965 56657 14051 56743
rect 20105 56720 20191 56743
rect 20273 56720 20359 56743
rect 20105 56680 20130 56720
rect 20130 56680 20170 56720
rect 20170 56680 20191 56720
rect 20273 56680 20294 56720
rect 20294 56680 20334 56720
rect 20334 56680 20359 56720
rect 20105 56657 20191 56680
rect 20273 56657 20359 56680
rect 3745 55964 3831 55987
rect 3913 55964 3999 55987
rect 3745 55924 3770 55964
rect 3770 55924 3810 55964
rect 3810 55924 3831 55964
rect 3913 55924 3934 55964
rect 3934 55924 3974 55964
rect 3974 55924 3999 55964
rect 3745 55901 3831 55924
rect 3913 55901 3999 55924
rect 18865 55964 18951 55987
rect 19033 55964 19119 55987
rect 18865 55924 18890 55964
rect 18890 55924 18930 55964
rect 18930 55924 18951 55964
rect 19033 55924 19054 55964
rect 19054 55924 19094 55964
rect 19094 55924 19119 55964
rect 18865 55901 18951 55924
rect 19033 55901 19119 55924
rect 4985 55208 5071 55231
rect 5153 55208 5239 55231
rect 4985 55168 5010 55208
rect 5010 55168 5050 55208
rect 5050 55168 5071 55208
rect 5153 55168 5174 55208
rect 5174 55168 5214 55208
rect 5214 55168 5239 55208
rect 4985 55145 5071 55168
rect 5153 55145 5239 55168
rect 20105 55208 20191 55231
rect 20273 55208 20359 55231
rect 20105 55168 20130 55208
rect 20130 55168 20170 55208
rect 20170 55168 20191 55208
rect 20273 55168 20294 55208
rect 20294 55168 20334 55208
rect 20334 55168 20359 55208
rect 20105 55145 20191 55168
rect 20273 55145 20359 55168
rect 3745 54452 3831 54475
rect 3913 54452 3999 54475
rect 3745 54412 3770 54452
rect 3770 54412 3810 54452
rect 3810 54412 3831 54452
rect 3913 54412 3934 54452
rect 3934 54412 3974 54452
rect 3974 54412 3999 54452
rect 3745 54389 3831 54412
rect 3913 54389 3999 54412
rect 18865 54452 18951 54475
rect 19033 54452 19119 54475
rect 18865 54412 18890 54452
rect 18890 54412 18930 54452
rect 18930 54412 18951 54452
rect 19033 54412 19054 54452
rect 19054 54412 19094 54452
rect 19094 54412 19119 54452
rect 18865 54389 18951 54412
rect 19033 54389 19119 54412
rect 4985 53696 5071 53719
rect 5153 53696 5239 53719
rect 4985 53656 5010 53696
rect 5010 53656 5050 53696
rect 5050 53656 5071 53696
rect 5153 53656 5174 53696
rect 5174 53656 5214 53696
rect 5214 53656 5239 53696
rect 4985 53633 5071 53656
rect 5153 53633 5239 53656
rect 20105 53696 20191 53719
rect 20273 53696 20359 53719
rect 20105 53656 20130 53696
rect 20130 53656 20170 53696
rect 20170 53656 20191 53696
rect 20273 53656 20294 53696
rect 20294 53656 20334 53696
rect 20334 53656 20359 53696
rect 20105 53633 20191 53656
rect 20273 53633 20359 53656
rect 3745 52940 3831 52963
rect 3913 52940 3999 52963
rect 3745 52900 3770 52940
rect 3770 52900 3810 52940
rect 3810 52900 3831 52940
rect 3913 52900 3934 52940
rect 3934 52900 3974 52940
rect 3974 52900 3999 52940
rect 3745 52877 3831 52900
rect 3913 52877 3999 52900
rect 18865 52940 18951 52963
rect 19033 52940 19119 52963
rect 18865 52900 18890 52940
rect 18890 52900 18930 52940
rect 18930 52900 18951 52940
rect 19033 52900 19054 52940
rect 19054 52900 19094 52940
rect 19094 52900 19119 52940
rect 18865 52877 18951 52900
rect 19033 52877 19119 52900
rect 4985 52184 5071 52207
rect 5153 52184 5239 52207
rect 4985 52144 5010 52184
rect 5010 52144 5050 52184
rect 5050 52144 5071 52184
rect 5153 52144 5174 52184
rect 5174 52144 5214 52184
rect 5214 52144 5239 52184
rect 4985 52121 5071 52144
rect 5153 52121 5239 52144
rect 20105 52184 20191 52207
rect 20273 52184 20359 52207
rect 20105 52144 20130 52184
rect 20130 52144 20170 52184
rect 20170 52144 20191 52184
rect 20273 52144 20294 52184
rect 20294 52144 20334 52184
rect 20334 52144 20359 52184
rect 20105 52121 20191 52144
rect 20273 52121 20359 52144
rect 3745 51428 3831 51451
rect 3913 51428 3999 51451
rect 3745 51388 3770 51428
rect 3770 51388 3810 51428
rect 3810 51388 3831 51428
rect 3913 51388 3934 51428
rect 3934 51388 3974 51428
rect 3974 51388 3999 51428
rect 3745 51365 3831 51388
rect 3913 51365 3999 51388
rect 18865 51428 18951 51451
rect 19033 51428 19119 51451
rect 18865 51388 18890 51428
rect 18890 51388 18930 51428
rect 18930 51388 18951 51428
rect 19033 51388 19054 51428
rect 19054 51388 19094 51428
rect 19094 51388 19119 51428
rect 18865 51365 18951 51388
rect 19033 51365 19119 51388
rect 4985 50672 5071 50695
rect 5153 50672 5239 50695
rect 4985 50632 5010 50672
rect 5010 50632 5050 50672
rect 5050 50632 5071 50672
rect 5153 50632 5174 50672
rect 5174 50632 5214 50672
rect 5214 50632 5239 50672
rect 4985 50609 5071 50632
rect 5153 50609 5239 50632
rect 20105 50672 20191 50695
rect 20273 50672 20359 50695
rect 20105 50632 20130 50672
rect 20130 50632 20170 50672
rect 20170 50632 20191 50672
rect 20273 50632 20294 50672
rect 20294 50632 20334 50672
rect 20334 50632 20359 50672
rect 20105 50609 20191 50632
rect 20273 50609 20359 50632
rect 3745 49916 3831 49939
rect 3913 49916 3999 49939
rect 3745 49876 3770 49916
rect 3770 49876 3810 49916
rect 3810 49876 3831 49916
rect 3913 49876 3934 49916
rect 3934 49876 3974 49916
rect 3974 49876 3999 49916
rect 3745 49853 3831 49876
rect 3913 49853 3999 49876
rect 18865 49916 18951 49939
rect 19033 49916 19119 49939
rect 18865 49876 18890 49916
rect 18890 49876 18930 49916
rect 18930 49876 18951 49916
rect 19033 49876 19054 49916
rect 19054 49876 19094 49916
rect 19094 49876 19119 49916
rect 18865 49853 18951 49876
rect 19033 49853 19119 49876
rect 4985 49160 5071 49183
rect 5153 49160 5239 49183
rect 4985 49120 5010 49160
rect 5010 49120 5050 49160
rect 5050 49120 5071 49160
rect 5153 49120 5174 49160
rect 5174 49120 5214 49160
rect 5214 49120 5239 49160
rect 4985 49097 5071 49120
rect 5153 49097 5239 49120
rect 20105 49160 20191 49183
rect 20273 49160 20359 49183
rect 20105 49120 20130 49160
rect 20130 49120 20170 49160
rect 20170 49120 20191 49160
rect 20273 49120 20294 49160
rect 20294 49120 20334 49160
rect 20334 49120 20359 49160
rect 20105 49097 20191 49120
rect 20273 49097 20359 49120
rect 3745 48404 3831 48427
rect 3913 48404 3999 48427
rect 3745 48364 3770 48404
rect 3770 48364 3810 48404
rect 3810 48364 3831 48404
rect 3913 48364 3934 48404
rect 3934 48364 3974 48404
rect 3974 48364 3999 48404
rect 3745 48341 3831 48364
rect 3913 48341 3999 48364
rect 18865 48404 18951 48427
rect 19033 48404 19119 48427
rect 18865 48364 18890 48404
rect 18890 48364 18930 48404
rect 18930 48364 18951 48404
rect 19033 48364 19054 48404
rect 19054 48364 19094 48404
rect 19094 48364 19119 48404
rect 18865 48341 18951 48364
rect 19033 48341 19119 48364
rect 8493 48005 8579 48091
rect 4985 47648 5071 47671
rect 5153 47648 5239 47671
rect 4985 47608 5010 47648
rect 5010 47608 5050 47648
rect 5050 47608 5071 47648
rect 5153 47608 5174 47648
rect 5174 47608 5214 47648
rect 5214 47608 5239 47648
rect 4985 47585 5071 47608
rect 5153 47585 5239 47608
rect 20105 47648 20191 47671
rect 20273 47648 20359 47671
rect 20105 47608 20130 47648
rect 20130 47608 20170 47648
rect 20170 47608 20191 47648
rect 20273 47608 20294 47648
rect 20294 47608 20334 47648
rect 20334 47608 20359 47648
rect 20105 47585 20191 47608
rect 20273 47585 20359 47608
rect 3745 46892 3831 46915
rect 3913 46892 3999 46915
rect 3745 46852 3770 46892
rect 3770 46852 3810 46892
rect 3810 46852 3831 46892
rect 3913 46852 3934 46892
rect 3934 46852 3974 46892
rect 3974 46852 3999 46892
rect 3745 46829 3831 46852
rect 3913 46829 3999 46852
rect 18865 46892 18951 46915
rect 19033 46892 19119 46915
rect 18865 46852 18890 46892
rect 18890 46852 18930 46892
rect 18930 46852 18951 46892
rect 19033 46852 19054 46892
rect 19054 46852 19094 46892
rect 19094 46852 19119 46892
rect 18865 46829 18951 46852
rect 19033 46829 19119 46852
rect 4985 46136 5071 46159
rect 5153 46136 5239 46159
rect 4985 46096 5010 46136
rect 5010 46096 5050 46136
rect 5050 46096 5071 46136
rect 5153 46096 5174 46136
rect 5174 46096 5214 46136
rect 5214 46096 5239 46136
rect 4985 46073 5071 46096
rect 5153 46073 5239 46096
rect 20105 46136 20191 46159
rect 20273 46136 20359 46159
rect 20105 46096 20130 46136
rect 20130 46096 20170 46136
rect 20170 46096 20191 46136
rect 20273 46096 20294 46136
rect 20294 46096 20334 46136
rect 20334 46096 20359 46136
rect 20105 46073 20191 46096
rect 20273 46073 20359 46096
rect 3745 45380 3831 45403
rect 3913 45380 3999 45403
rect 3745 45340 3770 45380
rect 3770 45340 3810 45380
rect 3810 45340 3831 45380
rect 3913 45340 3934 45380
rect 3934 45340 3974 45380
rect 3974 45340 3999 45380
rect 3745 45317 3831 45340
rect 3913 45317 3999 45340
rect 18865 45380 18951 45403
rect 19033 45380 19119 45403
rect 18865 45340 18890 45380
rect 18890 45340 18930 45380
rect 18930 45340 18951 45380
rect 19033 45340 19054 45380
rect 19054 45340 19094 45380
rect 19094 45340 19119 45380
rect 18865 45317 18951 45340
rect 19033 45317 19119 45340
rect 4985 44624 5071 44647
rect 5153 44624 5239 44647
rect 4985 44584 5010 44624
rect 5010 44584 5050 44624
rect 5050 44584 5071 44624
rect 5153 44584 5174 44624
rect 5174 44584 5214 44624
rect 5214 44584 5239 44624
rect 4985 44561 5071 44584
rect 5153 44561 5239 44584
rect 20105 44624 20191 44647
rect 20273 44624 20359 44647
rect 20105 44584 20130 44624
rect 20130 44584 20170 44624
rect 20170 44584 20191 44624
rect 20273 44584 20294 44624
rect 20294 44584 20334 44624
rect 20334 44584 20359 44624
rect 20105 44561 20191 44584
rect 20273 44561 20359 44584
rect 3745 43868 3831 43891
rect 3913 43868 3999 43891
rect 3745 43828 3770 43868
rect 3770 43828 3810 43868
rect 3810 43828 3831 43868
rect 3913 43828 3934 43868
rect 3934 43828 3974 43868
rect 3974 43828 3999 43868
rect 3745 43805 3831 43828
rect 3913 43805 3999 43828
rect 18865 43868 18951 43891
rect 19033 43868 19119 43891
rect 18865 43828 18890 43868
rect 18890 43828 18930 43868
rect 18930 43828 18951 43868
rect 19033 43828 19054 43868
rect 19054 43828 19094 43868
rect 19094 43828 19119 43868
rect 18865 43805 18951 43828
rect 19033 43805 19119 43828
rect 4985 43112 5071 43135
rect 5153 43112 5239 43135
rect 4985 43072 5010 43112
rect 5010 43072 5050 43112
rect 5050 43072 5071 43112
rect 5153 43072 5174 43112
rect 5174 43072 5214 43112
rect 5214 43072 5239 43112
rect 4985 43049 5071 43072
rect 5153 43049 5239 43072
rect 20105 43112 20191 43135
rect 20273 43112 20359 43135
rect 20105 43072 20130 43112
rect 20130 43072 20170 43112
rect 20170 43072 20191 43112
rect 20273 43072 20294 43112
rect 20294 43072 20334 43112
rect 20334 43072 20359 43112
rect 20105 43049 20191 43072
rect 20273 43049 20359 43072
rect 3745 42356 3831 42379
rect 3913 42356 3999 42379
rect 18865 42356 18951 42379
rect 19033 42356 19119 42379
rect 3745 42316 3770 42356
rect 3770 42316 3810 42356
rect 3810 42316 3831 42356
rect 3913 42316 3934 42356
rect 3934 42316 3974 42356
rect 3974 42316 3999 42356
rect 18865 42316 18890 42356
rect 18890 42316 18930 42356
rect 18930 42316 18951 42356
rect 19033 42316 19054 42356
rect 19054 42316 19094 42356
rect 19094 42316 19119 42356
rect 3745 42293 3831 42316
rect 3913 42293 3999 42316
rect 18865 42293 18951 42316
rect 19033 42293 19119 42316
rect 4985 41600 5071 41623
rect 5153 41600 5239 41623
rect 20105 41600 20191 41623
rect 20273 41600 20359 41623
rect 4985 41560 5010 41600
rect 5010 41560 5050 41600
rect 5050 41560 5071 41600
rect 5153 41560 5174 41600
rect 5174 41560 5214 41600
rect 5214 41560 5239 41600
rect 20105 41560 20130 41600
rect 20130 41560 20170 41600
rect 20170 41560 20191 41600
rect 20273 41560 20294 41600
rect 20294 41560 20334 41600
rect 20334 41560 20359 41600
rect 4985 41537 5071 41560
rect 5153 41537 5239 41560
rect 20105 41537 20191 41560
rect 20273 41537 20359 41560
rect 3745 40844 3831 40867
rect 3913 40844 3999 40867
rect 3745 40804 3770 40844
rect 3770 40804 3810 40844
rect 3810 40804 3831 40844
rect 3913 40804 3934 40844
rect 3934 40804 3974 40844
rect 3974 40804 3999 40844
rect 3745 40781 3831 40804
rect 3913 40781 3999 40804
rect 18865 40844 18951 40867
rect 19033 40844 19119 40867
rect 18865 40804 18890 40844
rect 18890 40804 18930 40844
rect 18930 40804 18951 40844
rect 19033 40804 19054 40844
rect 19054 40804 19094 40844
rect 19094 40804 19119 40844
rect 18865 40781 18951 40804
rect 19033 40781 19119 40804
rect 4985 40088 5071 40111
rect 5153 40088 5239 40111
rect 4985 40048 5010 40088
rect 5010 40048 5050 40088
rect 5050 40048 5071 40088
rect 5153 40048 5174 40088
rect 5174 40048 5214 40088
rect 5214 40048 5239 40088
rect 4985 40025 5071 40048
rect 5153 40025 5239 40048
rect 20105 40088 20191 40111
rect 20273 40088 20359 40111
rect 20105 40048 20130 40088
rect 20130 40048 20170 40088
rect 20170 40048 20191 40088
rect 20273 40048 20294 40088
rect 20294 40048 20334 40088
rect 20334 40048 20359 40088
rect 20105 40025 20191 40048
rect 20273 40025 20359 40048
rect 3745 39332 3831 39355
rect 3913 39332 3999 39355
rect 3745 39292 3770 39332
rect 3770 39292 3810 39332
rect 3810 39292 3831 39332
rect 3913 39292 3934 39332
rect 3934 39292 3974 39332
rect 3974 39292 3999 39332
rect 3745 39269 3831 39292
rect 3913 39269 3999 39292
rect 18865 39332 18951 39355
rect 19033 39332 19119 39355
rect 18865 39292 18890 39332
rect 18890 39292 18930 39332
rect 18930 39292 18951 39332
rect 19033 39292 19054 39332
rect 19054 39292 19094 39332
rect 19094 39292 19119 39332
rect 18865 39269 18951 39292
rect 19033 39269 19119 39292
rect 4985 38576 5071 38599
rect 5153 38576 5239 38599
rect 4985 38536 5010 38576
rect 5010 38536 5050 38576
rect 5050 38536 5071 38576
rect 5153 38536 5174 38576
rect 5174 38536 5214 38576
rect 5214 38536 5239 38576
rect 4985 38513 5071 38536
rect 5153 38513 5239 38536
rect 20105 38576 20191 38599
rect 20273 38576 20359 38599
rect 20105 38536 20130 38576
rect 20130 38536 20170 38576
rect 20170 38536 20191 38576
rect 20273 38536 20294 38576
rect 20294 38536 20334 38576
rect 20334 38536 20359 38576
rect 20105 38513 20191 38536
rect 20273 38513 20359 38536
rect 3745 37820 3831 37843
rect 3913 37820 3999 37843
rect 3745 37780 3770 37820
rect 3770 37780 3810 37820
rect 3810 37780 3831 37820
rect 3913 37780 3934 37820
rect 3934 37780 3974 37820
rect 3974 37780 3999 37820
rect 3745 37757 3831 37780
rect 3913 37757 3999 37780
rect 18865 37820 18951 37843
rect 19033 37820 19119 37843
rect 18865 37780 18890 37820
rect 18890 37780 18930 37820
rect 18930 37780 18951 37820
rect 19033 37780 19054 37820
rect 19054 37780 19094 37820
rect 19094 37780 19119 37820
rect 18865 37757 18951 37780
rect 19033 37757 19119 37780
rect 4985 37064 5071 37087
rect 5153 37064 5239 37087
rect 4985 37024 5010 37064
rect 5010 37024 5050 37064
rect 5050 37024 5071 37064
rect 5153 37024 5174 37064
rect 5174 37024 5214 37064
rect 5214 37024 5239 37064
rect 4985 37001 5071 37024
rect 5153 37001 5239 37024
rect 20105 37064 20191 37087
rect 20273 37064 20359 37087
rect 20105 37024 20130 37064
rect 20130 37024 20170 37064
rect 20170 37024 20191 37064
rect 20273 37024 20294 37064
rect 20294 37024 20334 37064
rect 20334 37024 20359 37064
rect 20105 37001 20191 37024
rect 20273 37001 20359 37024
rect 3745 36308 3831 36331
rect 3913 36308 3999 36331
rect 3745 36268 3770 36308
rect 3770 36268 3810 36308
rect 3810 36268 3831 36308
rect 3913 36268 3934 36308
rect 3934 36268 3974 36308
rect 3974 36268 3999 36308
rect 3745 36245 3831 36268
rect 3913 36245 3999 36268
rect 18865 36308 18951 36331
rect 19033 36308 19119 36331
rect 18865 36268 18890 36308
rect 18890 36268 18930 36308
rect 18930 36268 18951 36308
rect 19033 36268 19054 36308
rect 19054 36268 19094 36308
rect 19094 36268 19119 36308
rect 18865 36245 18951 36268
rect 19033 36245 19119 36268
rect 4985 35552 5071 35575
rect 5153 35552 5239 35575
rect 4985 35512 5010 35552
rect 5010 35512 5050 35552
rect 5050 35512 5071 35552
rect 5153 35512 5174 35552
rect 5174 35512 5214 35552
rect 5214 35512 5239 35552
rect 4985 35489 5071 35512
rect 5153 35489 5239 35512
rect 20105 35552 20191 35575
rect 20273 35552 20359 35575
rect 20105 35512 20130 35552
rect 20130 35512 20170 35552
rect 20170 35512 20191 35552
rect 20273 35512 20294 35552
rect 20294 35512 20334 35552
rect 20334 35512 20359 35552
rect 20105 35489 20191 35512
rect 20273 35489 20359 35512
rect 3745 34796 3831 34819
rect 3913 34796 3999 34819
rect 3745 34756 3770 34796
rect 3770 34756 3810 34796
rect 3810 34756 3831 34796
rect 3913 34756 3934 34796
rect 3934 34756 3974 34796
rect 3974 34756 3999 34796
rect 3745 34733 3831 34756
rect 3913 34733 3999 34756
rect 18865 34796 18951 34819
rect 19033 34796 19119 34819
rect 18865 34756 18890 34796
rect 18890 34756 18930 34796
rect 18930 34756 18951 34796
rect 19033 34756 19054 34796
rect 19054 34756 19094 34796
rect 19094 34756 19119 34796
rect 18865 34733 18951 34756
rect 19033 34733 19119 34756
rect 4985 34040 5071 34063
rect 5153 34040 5239 34063
rect 4985 34000 5010 34040
rect 5010 34000 5050 34040
rect 5050 34000 5071 34040
rect 5153 34000 5174 34040
rect 5174 34000 5214 34040
rect 5214 34000 5239 34040
rect 4985 33977 5071 34000
rect 5153 33977 5239 34000
rect 20105 34040 20191 34063
rect 20273 34040 20359 34063
rect 20105 34000 20130 34040
rect 20130 34000 20170 34040
rect 20170 34000 20191 34040
rect 20273 34000 20294 34040
rect 20294 34000 20334 34040
rect 20334 34000 20359 34040
rect 20105 33977 20191 34000
rect 20273 33977 20359 34000
rect 3745 33284 3831 33307
rect 3913 33284 3999 33307
rect 3745 33244 3770 33284
rect 3770 33244 3810 33284
rect 3810 33244 3831 33284
rect 3913 33244 3934 33284
rect 3934 33244 3974 33284
rect 3974 33244 3999 33284
rect 3745 33221 3831 33244
rect 3913 33221 3999 33244
rect 18865 33284 18951 33307
rect 19033 33284 19119 33307
rect 18865 33244 18890 33284
rect 18890 33244 18930 33284
rect 18930 33244 18951 33284
rect 19033 33244 19054 33284
rect 19054 33244 19094 33284
rect 19094 33244 19119 33284
rect 18865 33221 18951 33244
rect 19033 33221 19119 33244
rect 4985 32528 5071 32551
rect 5153 32528 5239 32551
rect 4985 32488 5010 32528
rect 5010 32488 5050 32528
rect 5050 32488 5071 32528
rect 5153 32488 5174 32528
rect 5174 32488 5214 32528
rect 5214 32488 5239 32528
rect 4985 32465 5071 32488
rect 5153 32465 5239 32488
rect 20105 32528 20191 32551
rect 20273 32528 20359 32551
rect 20105 32488 20130 32528
rect 20130 32488 20170 32528
rect 20170 32488 20191 32528
rect 20273 32488 20294 32528
rect 20294 32488 20334 32528
rect 20334 32488 20359 32528
rect 20105 32465 20191 32488
rect 20273 32465 20359 32488
rect 1197 32045 1283 32131
rect 3745 31772 3831 31795
rect 3913 31772 3999 31795
rect 3745 31732 3770 31772
rect 3770 31732 3810 31772
rect 3810 31732 3831 31772
rect 3913 31732 3934 31772
rect 3934 31732 3974 31772
rect 3974 31732 3999 31772
rect 3745 31709 3831 31732
rect 3913 31709 3999 31732
rect 18865 31772 18951 31795
rect 19033 31772 19119 31795
rect 18865 31732 18890 31772
rect 18890 31732 18930 31772
rect 18930 31732 18951 31772
rect 19033 31732 19054 31772
rect 19054 31732 19094 31772
rect 19094 31732 19119 31772
rect 18865 31709 18951 31732
rect 19033 31709 19119 31732
rect 4985 31016 5071 31039
rect 5153 31016 5239 31039
rect 4985 30976 5010 31016
rect 5010 30976 5050 31016
rect 5050 30976 5071 31016
rect 5153 30976 5174 31016
rect 5174 30976 5214 31016
rect 5214 30976 5239 31016
rect 4985 30953 5071 30976
rect 5153 30953 5239 30976
rect 20105 31016 20191 31039
rect 20273 31016 20359 31039
rect 20105 30976 20130 31016
rect 20130 30976 20170 31016
rect 20170 30976 20191 31016
rect 20273 30976 20294 31016
rect 20294 30976 20334 31016
rect 20334 30976 20359 31016
rect 20105 30953 20191 30976
rect 20273 30953 20359 30976
rect 3745 30260 3831 30283
rect 3913 30260 3999 30283
rect 3745 30220 3770 30260
rect 3770 30220 3810 30260
rect 3810 30220 3831 30260
rect 3913 30220 3934 30260
rect 3934 30220 3974 30260
rect 3974 30220 3999 30260
rect 3745 30197 3831 30220
rect 3913 30197 3999 30220
rect 18865 30260 18951 30283
rect 19033 30260 19119 30283
rect 18865 30220 18890 30260
rect 18890 30220 18930 30260
rect 18930 30220 18951 30260
rect 19033 30220 19054 30260
rect 19054 30220 19094 30260
rect 19094 30220 19119 30260
rect 18865 30197 18951 30220
rect 19033 30197 19119 30220
rect 4985 29504 5071 29527
rect 5153 29504 5239 29527
rect 4985 29464 5010 29504
rect 5010 29464 5050 29504
rect 5050 29464 5071 29504
rect 5153 29464 5174 29504
rect 5174 29464 5214 29504
rect 5214 29464 5239 29504
rect 4985 29441 5071 29464
rect 5153 29441 5239 29464
rect 20105 29504 20191 29527
rect 20273 29504 20359 29527
rect 20105 29464 20130 29504
rect 20130 29464 20170 29504
rect 20170 29464 20191 29504
rect 20273 29464 20294 29504
rect 20294 29464 20334 29504
rect 20334 29464 20359 29504
rect 20105 29441 20191 29464
rect 20273 29441 20359 29464
rect 3745 28748 3831 28771
rect 3913 28748 3999 28771
rect 3745 28708 3770 28748
rect 3770 28708 3810 28748
rect 3810 28708 3831 28748
rect 3913 28708 3934 28748
rect 3934 28708 3974 28748
rect 3974 28708 3999 28748
rect 3745 28685 3831 28708
rect 3913 28685 3999 28708
rect 18865 28748 18951 28771
rect 19033 28748 19119 28771
rect 18865 28708 18890 28748
rect 18890 28708 18930 28748
rect 18930 28708 18951 28748
rect 19033 28708 19054 28748
rect 19054 28708 19094 28748
rect 19094 28708 19119 28748
rect 18865 28685 18951 28708
rect 19033 28685 19119 28708
rect 4985 27992 5071 28015
rect 5153 27992 5239 28015
rect 4985 27952 5010 27992
rect 5010 27952 5050 27992
rect 5050 27952 5071 27992
rect 5153 27952 5174 27992
rect 5174 27952 5214 27992
rect 5214 27952 5239 27992
rect 4985 27929 5071 27952
rect 5153 27929 5239 27952
rect 20105 27992 20191 28015
rect 20273 27992 20359 28015
rect 20105 27952 20130 27992
rect 20130 27952 20170 27992
rect 20170 27952 20191 27992
rect 20273 27952 20294 27992
rect 20294 27952 20334 27992
rect 20334 27952 20359 27992
rect 20105 27929 20191 27952
rect 20273 27929 20359 27952
rect 3745 27236 3831 27259
rect 3913 27236 3999 27259
rect 3745 27196 3770 27236
rect 3770 27196 3810 27236
rect 3810 27196 3831 27236
rect 3913 27196 3934 27236
rect 3934 27196 3974 27236
rect 3974 27196 3999 27236
rect 3745 27173 3831 27196
rect 3913 27173 3999 27196
rect 18865 27236 18951 27259
rect 19033 27236 19119 27259
rect 18865 27196 18890 27236
rect 18890 27196 18930 27236
rect 18930 27196 18951 27236
rect 19033 27196 19054 27236
rect 19054 27196 19094 27236
rect 19094 27196 19119 27236
rect 18865 27173 18951 27196
rect 19033 27173 19119 27196
rect 4985 26480 5071 26503
rect 5153 26480 5239 26503
rect 4985 26440 5010 26480
rect 5010 26440 5050 26480
rect 5050 26440 5071 26480
rect 5153 26440 5174 26480
rect 5174 26440 5214 26480
rect 5214 26440 5239 26480
rect 4985 26417 5071 26440
rect 5153 26417 5239 26440
rect 20105 26480 20191 26503
rect 20273 26480 20359 26503
rect 20105 26440 20130 26480
rect 20130 26440 20170 26480
rect 20170 26440 20191 26480
rect 20273 26440 20294 26480
rect 20294 26440 20334 26480
rect 20334 26440 20359 26480
rect 20105 26417 20191 26440
rect 20273 26417 20359 26440
rect 3745 25724 3831 25747
rect 3913 25724 3999 25747
rect 3745 25684 3770 25724
rect 3770 25684 3810 25724
rect 3810 25684 3831 25724
rect 3913 25684 3934 25724
rect 3934 25684 3974 25724
rect 3974 25684 3999 25724
rect 3745 25661 3831 25684
rect 3913 25661 3999 25684
rect 18865 25724 18951 25747
rect 19033 25724 19119 25747
rect 18865 25684 18890 25724
rect 18890 25684 18930 25724
rect 18930 25684 18951 25724
rect 19033 25684 19054 25724
rect 19054 25684 19094 25724
rect 19094 25684 19119 25724
rect 18865 25661 18951 25684
rect 19033 25661 19119 25684
rect 13965 25157 14051 25243
rect 4985 24968 5071 24991
rect 5153 24968 5239 24991
rect 4985 24928 5010 24968
rect 5010 24928 5050 24968
rect 5050 24928 5071 24968
rect 5153 24928 5174 24968
rect 5174 24928 5214 24968
rect 5214 24928 5239 24968
rect 4985 24905 5071 24928
rect 5153 24905 5239 24928
rect 20105 24968 20191 24991
rect 20273 24968 20359 24991
rect 20105 24928 20130 24968
rect 20130 24928 20170 24968
rect 20170 24928 20191 24968
rect 20273 24928 20294 24968
rect 20294 24928 20334 24968
rect 20334 24928 20359 24968
rect 20105 24905 20191 24928
rect 20273 24905 20359 24928
rect 3745 24212 3831 24235
rect 3913 24212 3999 24235
rect 3745 24172 3770 24212
rect 3770 24172 3810 24212
rect 3810 24172 3831 24212
rect 3913 24172 3934 24212
rect 3934 24172 3974 24212
rect 3974 24172 3999 24212
rect 3745 24149 3831 24172
rect 3913 24149 3999 24172
rect 18865 24212 18951 24235
rect 19033 24212 19119 24235
rect 18865 24172 18890 24212
rect 18890 24172 18930 24212
rect 18930 24172 18951 24212
rect 19033 24172 19054 24212
rect 19054 24172 19094 24212
rect 19094 24172 19119 24212
rect 18865 24149 18951 24172
rect 19033 24149 19119 24172
rect 4985 23456 5071 23479
rect 5153 23456 5239 23479
rect 20105 23456 20191 23479
rect 20273 23456 20359 23479
rect 4985 23416 5010 23456
rect 5010 23416 5050 23456
rect 5050 23416 5071 23456
rect 5153 23416 5174 23456
rect 5174 23416 5214 23456
rect 5214 23416 5239 23456
rect 20105 23416 20130 23456
rect 20130 23416 20170 23456
rect 20170 23416 20191 23456
rect 20273 23416 20294 23456
rect 20294 23416 20334 23456
rect 20334 23416 20359 23456
rect 4985 23393 5071 23416
rect 5153 23393 5239 23416
rect 20105 23393 20191 23416
rect 20273 23393 20359 23416
rect 3745 22700 3831 22723
rect 3913 22700 3999 22723
rect 18865 22700 18951 22723
rect 19033 22700 19119 22723
rect 3745 22660 3770 22700
rect 3770 22660 3810 22700
rect 3810 22660 3831 22700
rect 3913 22660 3934 22700
rect 3934 22660 3974 22700
rect 3974 22660 3999 22700
rect 18865 22660 18890 22700
rect 18890 22660 18930 22700
rect 18930 22660 18951 22700
rect 19033 22660 19054 22700
rect 19054 22660 19094 22700
rect 19094 22660 19119 22700
rect 3745 22637 3831 22660
rect 3913 22637 3999 22660
rect 18865 22637 18951 22660
rect 19033 22637 19119 22660
rect 4985 21944 5071 21967
rect 5153 21944 5239 21967
rect 4985 21904 5010 21944
rect 5010 21904 5050 21944
rect 5050 21904 5071 21944
rect 5153 21904 5174 21944
rect 5174 21904 5214 21944
rect 5214 21904 5239 21944
rect 4985 21881 5071 21904
rect 5153 21881 5239 21904
rect 20105 21944 20191 21967
rect 20273 21944 20359 21967
rect 20105 21904 20130 21944
rect 20130 21904 20170 21944
rect 20170 21904 20191 21944
rect 20273 21904 20294 21944
rect 20294 21904 20334 21944
rect 20334 21904 20359 21944
rect 20105 21881 20191 21904
rect 20273 21881 20359 21904
rect 3745 21188 3831 21211
rect 3913 21188 3999 21211
rect 3745 21148 3770 21188
rect 3770 21148 3810 21188
rect 3810 21148 3831 21188
rect 3913 21148 3934 21188
rect 3934 21148 3974 21188
rect 3974 21148 3999 21188
rect 3745 21125 3831 21148
rect 3913 21125 3999 21148
rect 18865 21188 18951 21211
rect 19033 21188 19119 21211
rect 18865 21148 18890 21188
rect 18890 21148 18930 21188
rect 18930 21148 18951 21188
rect 19033 21148 19054 21188
rect 19054 21148 19094 21188
rect 19094 21148 19119 21188
rect 18865 21125 18951 21148
rect 19033 21125 19119 21148
rect 4985 20432 5071 20455
rect 5153 20432 5239 20455
rect 4985 20392 5010 20432
rect 5010 20392 5050 20432
rect 5050 20392 5071 20432
rect 5153 20392 5174 20432
rect 5174 20392 5214 20432
rect 5214 20392 5239 20432
rect 4985 20369 5071 20392
rect 5153 20369 5239 20392
rect 20105 20432 20191 20455
rect 20273 20432 20359 20455
rect 20105 20392 20130 20432
rect 20130 20392 20170 20432
rect 20170 20392 20191 20432
rect 20273 20392 20294 20432
rect 20294 20392 20334 20432
rect 20334 20392 20359 20432
rect 20105 20369 20191 20392
rect 20273 20369 20359 20392
rect 3745 19676 3831 19699
rect 3913 19676 3999 19699
rect 3745 19636 3770 19676
rect 3770 19636 3810 19676
rect 3810 19636 3831 19676
rect 3913 19636 3934 19676
rect 3934 19636 3974 19676
rect 3974 19636 3999 19676
rect 3745 19613 3831 19636
rect 3913 19613 3999 19636
rect 18865 19676 18951 19699
rect 19033 19676 19119 19699
rect 18865 19636 18890 19676
rect 18890 19636 18930 19676
rect 18930 19636 18951 19676
rect 19033 19636 19054 19676
rect 19054 19636 19094 19676
rect 19094 19636 19119 19676
rect 18865 19613 18951 19636
rect 19033 19613 19119 19636
rect 4985 18920 5071 18943
rect 5153 18920 5239 18943
rect 4985 18880 5010 18920
rect 5010 18880 5050 18920
rect 5050 18880 5071 18920
rect 5153 18880 5174 18920
rect 5174 18880 5214 18920
rect 5214 18880 5239 18920
rect 4985 18857 5071 18880
rect 5153 18857 5239 18880
rect 20105 18920 20191 18943
rect 20273 18920 20359 18943
rect 20105 18880 20130 18920
rect 20130 18880 20170 18920
rect 20170 18880 20191 18920
rect 20273 18880 20294 18920
rect 20294 18880 20334 18920
rect 20334 18880 20359 18920
rect 20105 18857 20191 18880
rect 20273 18857 20359 18880
rect 3745 18164 3831 18187
rect 3913 18164 3999 18187
rect 3745 18124 3770 18164
rect 3770 18124 3810 18164
rect 3810 18124 3831 18164
rect 3913 18124 3934 18164
rect 3934 18124 3974 18164
rect 3974 18124 3999 18164
rect 3745 18101 3831 18124
rect 3913 18101 3999 18124
rect 18865 18164 18951 18187
rect 19033 18164 19119 18187
rect 18865 18124 18890 18164
rect 18890 18124 18930 18164
rect 18930 18124 18951 18164
rect 19033 18124 19054 18164
rect 19054 18124 19094 18164
rect 19094 18124 19119 18164
rect 18865 18101 18951 18124
rect 19033 18101 19119 18124
rect 4985 17408 5071 17431
rect 5153 17408 5239 17431
rect 4985 17368 5010 17408
rect 5010 17368 5050 17408
rect 5050 17368 5071 17408
rect 5153 17368 5174 17408
rect 5174 17368 5214 17408
rect 5214 17368 5239 17408
rect 4985 17345 5071 17368
rect 5153 17345 5239 17368
rect 20105 17408 20191 17431
rect 20273 17408 20359 17431
rect 20105 17368 20130 17408
rect 20130 17368 20170 17408
rect 20170 17368 20191 17408
rect 20273 17368 20294 17408
rect 20294 17368 20334 17408
rect 20334 17368 20359 17408
rect 20105 17345 20191 17368
rect 20273 17345 20359 17368
rect 3745 16652 3831 16675
rect 3913 16652 3999 16675
rect 3745 16612 3770 16652
rect 3770 16612 3810 16652
rect 3810 16612 3831 16652
rect 3913 16612 3934 16652
rect 3934 16612 3974 16652
rect 3974 16612 3999 16652
rect 3745 16589 3831 16612
rect 3913 16589 3999 16612
rect 18865 16652 18951 16675
rect 19033 16652 19119 16675
rect 18865 16612 18890 16652
rect 18890 16612 18930 16652
rect 18930 16612 18951 16652
rect 19033 16612 19054 16652
rect 19054 16612 19094 16652
rect 19094 16612 19119 16652
rect 18865 16589 18951 16612
rect 19033 16589 19119 16612
rect 4985 15896 5071 15919
rect 5153 15896 5239 15919
rect 4985 15856 5010 15896
rect 5010 15856 5050 15896
rect 5050 15856 5071 15896
rect 5153 15856 5174 15896
rect 5174 15856 5214 15896
rect 5214 15856 5239 15896
rect 4985 15833 5071 15856
rect 5153 15833 5239 15856
rect 20105 15896 20191 15919
rect 20273 15896 20359 15919
rect 20105 15856 20130 15896
rect 20130 15856 20170 15896
rect 20170 15856 20191 15896
rect 20273 15856 20294 15896
rect 20294 15856 20334 15896
rect 20334 15856 20359 15896
rect 20105 15833 20191 15856
rect 20273 15833 20359 15856
rect 3745 15140 3831 15163
rect 3913 15140 3999 15163
rect 3745 15100 3770 15140
rect 3770 15100 3810 15140
rect 3810 15100 3831 15140
rect 3913 15100 3934 15140
rect 3934 15100 3974 15140
rect 3974 15100 3999 15140
rect 3745 15077 3831 15100
rect 3913 15077 3999 15100
rect 18865 15140 18951 15163
rect 19033 15140 19119 15163
rect 18865 15100 18890 15140
rect 18890 15100 18930 15140
rect 18930 15100 18951 15140
rect 19033 15100 19054 15140
rect 19054 15100 19094 15140
rect 19094 15100 19119 15140
rect 18865 15077 18951 15100
rect 19033 15077 19119 15100
rect 4985 14384 5071 14407
rect 5153 14384 5239 14407
rect 4985 14344 5010 14384
rect 5010 14344 5050 14384
rect 5050 14344 5071 14384
rect 5153 14344 5174 14384
rect 5174 14344 5214 14384
rect 5214 14344 5239 14384
rect 4985 14321 5071 14344
rect 5153 14321 5239 14344
rect 20105 14384 20191 14407
rect 20273 14384 20359 14407
rect 20105 14344 20130 14384
rect 20130 14344 20170 14384
rect 20170 14344 20191 14384
rect 20273 14344 20294 14384
rect 20294 14344 20334 14384
rect 20334 14344 20359 14384
rect 20105 14321 20191 14344
rect 20273 14321 20359 14344
rect 3745 13628 3831 13651
rect 3913 13628 3999 13651
rect 3745 13588 3770 13628
rect 3770 13588 3810 13628
rect 3810 13588 3831 13628
rect 3913 13588 3934 13628
rect 3934 13588 3974 13628
rect 3974 13588 3999 13628
rect 3745 13565 3831 13588
rect 3913 13565 3999 13588
rect 18865 13628 18951 13651
rect 19033 13628 19119 13651
rect 18865 13588 18890 13628
rect 18890 13588 18930 13628
rect 18930 13588 18951 13628
rect 19033 13588 19054 13628
rect 19054 13588 19094 13628
rect 19094 13588 19119 13628
rect 18865 13565 18951 13588
rect 19033 13565 19119 13588
rect 4985 12872 5071 12895
rect 5153 12872 5239 12895
rect 4985 12832 5010 12872
rect 5010 12832 5050 12872
rect 5050 12832 5071 12872
rect 5153 12832 5174 12872
rect 5174 12832 5214 12872
rect 5214 12832 5239 12872
rect 4985 12809 5071 12832
rect 5153 12809 5239 12832
rect 20105 12872 20191 12895
rect 20273 12872 20359 12895
rect 20105 12832 20130 12872
rect 20130 12832 20170 12872
rect 20170 12832 20191 12872
rect 20273 12832 20294 12872
rect 20294 12832 20334 12872
rect 20334 12832 20359 12872
rect 20105 12809 20191 12832
rect 20273 12809 20359 12832
rect 3745 12116 3831 12139
rect 3913 12116 3999 12139
rect 3745 12076 3770 12116
rect 3770 12076 3810 12116
rect 3810 12076 3831 12116
rect 3913 12076 3934 12116
rect 3934 12076 3974 12116
rect 3974 12076 3999 12116
rect 3745 12053 3831 12076
rect 3913 12053 3999 12076
rect 18865 12116 18951 12139
rect 19033 12116 19119 12139
rect 18865 12076 18890 12116
rect 18890 12076 18930 12116
rect 18930 12076 18951 12116
rect 19033 12076 19054 12116
rect 19054 12076 19094 12116
rect 19094 12076 19119 12116
rect 18865 12053 18951 12076
rect 19033 12053 19119 12076
rect 4985 11360 5071 11383
rect 5153 11360 5239 11383
rect 4985 11320 5010 11360
rect 5010 11320 5050 11360
rect 5050 11320 5071 11360
rect 5153 11320 5174 11360
rect 5174 11320 5214 11360
rect 5214 11320 5239 11360
rect 4985 11297 5071 11320
rect 5153 11297 5239 11320
rect 20105 11360 20191 11383
rect 20273 11360 20359 11383
rect 20105 11320 20130 11360
rect 20130 11320 20170 11360
rect 20170 11320 20191 11360
rect 20273 11320 20294 11360
rect 20294 11320 20334 11360
rect 20334 11320 20359 11360
rect 20105 11297 20191 11320
rect 20273 11297 20359 11320
rect 3745 10604 3831 10627
rect 3913 10604 3999 10627
rect 3745 10564 3770 10604
rect 3770 10564 3810 10604
rect 3810 10564 3831 10604
rect 3913 10564 3934 10604
rect 3934 10564 3974 10604
rect 3974 10564 3999 10604
rect 3745 10541 3831 10564
rect 3913 10541 3999 10564
rect 18865 10604 18951 10627
rect 19033 10604 19119 10627
rect 18865 10564 18890 10604
rect 18890 10564 18930 10604
rect 18930 10564 18951 10604
rect 19033 10564 19054 10604
rect 19054 10564 19094 10604
rect 19094 10564 19119 10604
rect 18865 10541 18951 10564
rect 19033 10541 19119 10564
rect 4985 9848 5071 9871
rect 5153 9848 5239 9871
rect 4985 9808 5010 9848
rect 5010 9808 5050 9848
rect 5050 9808 5071 9848
rect 5153 9808 5174 9848
rect 5174 9808 5214 9848
rect 5214 9808 5239 9848
rect 4985 9785 5071 9808
rect 5153 9785 5239 9808
rect 20105 9848 20191 9871
rect 20273 9848 20359 9871
rect 20105 9808 20130 9848
rect 20130 9808 20170 9848
rect 20170 9808 20191 9848
rect 20273 9808 20294 9848
rect 20294 9808 20334 9848
rect 20334 9808 20359 9848
rect 20105 9785 20191 9808
rect 20273 9785 20359 9808
rect 3745 9092 3831 9115
rect 3913 9092 3999 9115
rect 3745 9052 3770 9092
rect 3770 9052 3810 9092
rect 3810 9052 3831 9092
rect 3913 9052 3934 9092
rect 3934 9052 3974 9092
rect 3974 9052 3999 9092
rect 3745 9029 3831 9052
rect 3913 9029 3999 9052
rect 18865 9092 18951 9115
rect 19033 9092 19119 9115
rect 18865 9052 18890 9092
rect 18890 9052 18930 9092
rect 18930 9052 18951 9092
rect 19033 9052 19054 9092
rect 19054 9052 19094 9092
rect 19094 9052 19119 9092
rect 18865 9029 18951 9052
rect 19033 9029 19119 9052
rect 4985 8336 5071 8359
rect 5153 8336 5239 8359
rect 4985 8296 5010 8336
rect 5010 8296 5050 8336
rect 5050 8296 5071 8336
rect 5153 8296 5174 8336
rect 5174 8296 5214 8336
rect 5214 8296 5239 8336
rect 4985 8273 5071 8296
rect 5153 8273 5239 8296
rect 20105 8336 20191 8359
rect 20273 8336 20359 8359
rect 20105 8296 20130 8336
rect 20130 8296 20170 8336
rect 20170 8296 20191 8336
rect 20273 8296 20294 8336
rect 20294 8296 20334 8336
rect 20334 8296 20359 8336
rect 20105 8273 20191 8296
rect 20273 8273 20359 8296
rect 3745 7580 3831 7603
rect 3913 7580 3999 7603
rect 3745 7540 3770 7580
rect 3770 7540 3810 7580
rect 3810 7540 3831 7580
rect 3913 7540 3934 7580
rect 3934 7540 3974 7580
rect 3974 7540 3999 7580
rect 3745 7517 3831 7540
rect 3913 7517 3999 7540
rect 18865 7580 18951 7603
rect 19033 7580 19119 7603
rect 18865 7540 18890 7580
rect 18890 7540 18930 7580
rect 18930 7540 18951 7580
rect 19033 7540 19054 7580
rect 19054 7540 19094 7580
rect 19094 7540 19119 7580
rect 18865 7517 18951 7540
rect 19033 7517 19119 7540
rect 9861 7349 9947 7435
rect 4985 6824 5071 6847
rect 5153 6824 5239 6847
rect 4985 6784 5010 6824
rect 5010 6784 5050 6824
rect 5050 6784 5071 6824
rect 5153 6784 5174 6824
rect 5174 6784 5214 6824
rect 5214 6784 5239 6824
rect 4985 6761 5071 6784
rect 5153 6761 5239 6784
rect 20105 6824 20191 6847
rect 20273 6824 20359 6847
rect 20105 6784 20130 6824
rect 20130 6784 20170 6824
rect 20170 6784 20191 6824
rect 20273 6784 20294 6824
rect 20294 6784 20334 6824
rect 20334 6784 20359 6824
rect 20105 6761 20191 6784
rect 20273 6761 20359 6784
rect 3745 6068 3831 6091
rect 3913 6068 3999 6091
rect 3745 6028 3770 6068
rect 3770 6028 3810 6068
rect 3810 6028 3831 6068
rect 3913 6028 3934 6068
rect 3934 6028 3974 6068
rect 3974 6028 3999 6068
rect 3745 6005 3831 6028
rect 3913 6005 3999 6028
rect 18865 6068 18951 6091
rect 19033 6068 19119 6091
rect 18865 6028 18890 6068
rect 18890 6028 18930 6068
rect 18930 6028 18951 6068
rect 19033 6028 19054 6068
rect 19054 6028 19094 6068
rect 19094 6028 19119 6068
rect 18865 6005 18951 6028
rect 19033 6005 19119 6028
rect 10773 5585 10859 5671
rect 4985 5312 5071 5335
rect 5153 5312 5239 5335
rect 4985 5272 5010 5312
rect 5010 5272 5050 5312
rect 5050 5272 5071 5312
rect 5153 5272 5174 5312
rect 5174 5272 5214 5312
rect 5214 5272 5239 5312
rect 4985 5249 5071 5272
rect 5153 5249 5239 5272
rect 20105 5312 20191 5335
rect 20273 5312 20359 5335
rect 20105 5272 20130 5312
rect 20130 5272 20170 5312
rect 20170 5272 20191 5312
rect 20273 5272 20294 5312
rect 20294 5272 20334 5312
rect 20334 5272 20359 5312
rect 20105 5249 20191 5272
rect 20273 5249 20359 5272
rect 6669 4745 6755 4831
rect 3745 4556 3831 4579
rect 3913 4556 3999 4579
rect 18865 4556 18951 4579
rect 19033 4556 19119 4579
rect 3745 4516 3770 4556
rect 3770 4516 3810 4556
rect 3810 4516 3831 4556
rect 3913 4516 3934 4556
rect 3934 4516 3974 4556
rect 3974 4516 3999 4556
rect 18865 4516 18890 4556
rect 18890 4516 18930 4556
rect 18930 4516 18951 4556
rect 19033 4516 19054 4556
rect 19054 4516 19094 4556
rect 19094 4516 19119 4556
rect 3745 4493 3831 4516
rect 3913 4493 3999 4516
rect 18865 4493 18951 4516
rect 19033 4493 19119 4516
rect 4985 3800 5071 3823
rect 5153 3800 5239 3823
rect 4985 3760 5010 3800
rect 5010 3760 5050 3800
rect 5050 3760 5071 3800
rect 5153 3760 5174 3800
rect 5174 3760 5214 3800
rect 5214 3760 5239 3800
rect 4985 3737 5071 3760
rect 5153 3737 5239 3760
rect 20105 3800 20191 3823
rect 20273 3800 20359 3823
rect 20105 3760 20130 3800
rect 20130 3760 20170 3800
rect 20170 3760 20191 3800
rect 20273 3760 20294 3800
rect 20294 3760 20334 3800
rect 20334 3760 20359 3800
rect 20105 3737 20191 3760
rect 20273 3737 20359 3760
rect 2109 3632 2195 3655
rect 2109 3592 2132 3632
rect 2132 3592 2195 3632
rect 2109 3569 2195 3592
rect 3745 3044 3831 3067
rect 3913 3044 3999 3067
rect 3745 3004 3770 3044
rect 3770 3004 3810 3044
rect 3810 3004 3831 3044
rect 3913 3004 3934 3044
rect 3934 3004 3974 3044
rect 3974 3004 3999 3044
rect 3745 2981 3831 3004
rect 3913 2981 3999 3004
rect 18865 3044 18951 3067
rect 19033 3044 19119 3067
rect 18865 3004 18890 3044
rect 18890 3004 18930 3044
rect 18930 3004 18951 3044
rect 19033 3004 19054 3044
rect 19054 3004 19094 3044
rect 19094 3004 19119 3044
rect 18865 2981 18951 3004
rect 19033 2981 19119 3004
rect 4985 2288 5071 2311
rect 5153 2288 5239 2311
rect 4985 2248 5010 2288
rect 5010 2248 5050 2288
rect 5050 2248 5071 2288
rect 5153 2248 5174 2288
rect 5174 2248 5214 2288
rect 5214 2248 5239 2288
rect 4985 2225 5071 2248
rect 5153 2225 5239 2248
rect 20105 2288 20191 2311
rect 20273 2288 20359 2311
rect 20105 2248 20130 2288
rect 20130 2248 20170 2288
rect 20170 2248 20191 2288
rect 20273 2248 20294 2288
rect 20294 2248 20334 2288
rect 20334 2248 20359 2288
rect 20105 2225 20191 2248
rect 20273 2225 20359 2248
rect 12141 1805 12227 1891
rect 3745 1532 3831 1555
rect 3913 1532 3999 1555
rect 3745 1492 3770 1532
rect 3770 1492 3810 1532
rect 3810 1492 3831 1532
rect 3913 1492 3934 1532
rect 3934 1492 3974 1532
rect 3974 1492 3999 1532
rect 3745 1469 3831 1492
rect 3913 1469 3999 1492
rect 18865 1532 18951 1555
rect 19033 1532 19119 1555
rect 18865 1492 18890 1532
rect 18890 1492 18930 1532
rect 18930 1492 18951 1532
rect 19033 1492 19054 1532
rect 19054 1492 19094 1532
rect 19094 1492 19119 1532
rect 18865 1469 18951 1492
rect 19033 1469 19119 1492
rect 13053 1217 13139 1303
rect 4985 776 5071 799
rect 5153 776 5239 799
rect 4985 736 5010 776
rect 5010 736 5050 776
rect 5050 736 5071 776
rect 5153 736 5174 776
rect 5174 736 5214 776
rect 5214 736 5239 776
rect 4985 713 5071 736
rect 5153 713 5239 736
rect 15789 713 15875 799
rect 20105 776 20191 799
rect 20273 776 20359 799
rect 20105 736 20130 776
rect 20130 736 20170 776
rect 20170 736 20191 776
rect 20273 736 20294 776
rect 20294 736 20334 776
rect 20334 736 20359 776
rect 16701 629 16787 715
rect 20105 713 20191 736
rect 20273 713 20359 736
<< metal6 >>
rect 3652 84715 4092 86016
rect 3652 84629 3745 84715
rect 3831 84629 3913 84715
rect 3999 84629 4092 84715
rect 3652 83203 4092 84629
rect 3652 83117 3745 83203
rect 3831 83117 3913 83203
rect 3999 83117 4092 83203
rect 3652 81691 4092 83117
rect 3652 81605 3745 81691
rect 3831 81605 3913 81691
rect 3999 81605 4092 81691
rect 3652 80179 4092 81605
rect 3652 80093 3745 80179
rect 3831 80093 3913 80179
rect 3999 80093 4092 80179
rect 3652 78667 4092 80093
rect 3652 78581 3745 78667
rect 3831 78581 3913 78667
rect 3999 78581 4092 78667
rect 3652 77155 4092 78581
rect 3652 77069 3745 77155
rect 3831 77069 3913 77155
rect 3999 77069 4092 77155
rect 1988 76903 2316 77024
rect 1988 76817 2109 76903
rect 2195 76817 2316 76903
rect 1076 73039 1404 73160
rect 1076 72953 1197 73039
rect 1283 72953 1404 73039
rect 1076 32131 1404 72953
rect 1076 32045 1197 32131
rect 1283 32045 1404 32131
rect 1076 31924 1404 32045
rect 1988 3655 2316 76817
rect 1988 3569 2109 3655
rect 2195 3569 2316 3655
rect 1988 3448 2316 3569
rect 3652 75643 4092 77069
rect 3652 75557 3745 75643
rect 3831 75557 3913 75643
rect 3999 75557 4092 75643
rect 3652 74131 4092 75557
rect 3652 74045 3745 74131
rect 3831 74045 3913 74131
rect 3999 74045 4092 74131
rect 3652 72619 4092 74045
rect 3652 72533 3745 72619
rect 3831 72533 3913 72619
rect 3999 72533 4092 72619
rect 3652 71107 4092 72533
rect 3652 71021 3745 71107
rect 3831 71021 3913 71107
rect 3999 71021 4092 71107
rect 3652 69595 4092 71021
rect 3652 69509 3745 69595
rect 3831 69509 3913 69595
rect 3999 69509 4092 69595
rect 3652 68083 4092 69509
rect 3652 67997 3745 68083
rect 3831 67997 3913 68083
rect 3999 67997 4092 68083
rect 3652 66571 4092 67997
rect 3652 66485 3745 66571
rect 3831 66485 3913 66571
rect 3999 66485 4092 66571
rect 3652 65059 4092 66485
rect 3652 64973 3745 65059
rect 3831 64973 3913 65059
rect 3999 64973 4092 65059
rect 3652 63547 4092 64973
rect 3652 63461 3745 63547
rect 3831 63461 3913 63547
rect 3999 63461 4092 63547
rect 3652 62035 4092 63461
rect 3652 61949 3745 62035
rect 3831 61949 3913 62035
rect 3999 61949 4092 62035
rect 3652 60523 4092 61949
rect 3652 60437 3745 60523
rect 3831 60437 3913 60523
rect 3999 60437 4092 60523
rect 3652 59011 4092 60437
rect 3652 58925 3745 59011
rect 3831 58925 3913 59011
rect 3999 58925 4092 59011
rect 3652 57499 4092 58925
rect 3652 57413 3745 57499
rect 3831 57413 3913 57499
rect 3999 57413 4092 57499
rect 3652 55987 4092 57413
rect 3652 55901 3745 55987
rect 3831 55901 3913 55987
rect 3999 55901 4092 55987
rect 3652 54475 4092 55901
rect 3652 54389 3745 54475
rect 3831 54389 3913 54475
rect 3999 54389 4092 54475
rect 3652 52963 4092 54389
rect 3652 52877 3745 52963
rect 3831 52877 3913 52963
rect 3999 52877 4092 52963
rect 3652 51451 4092 52877
rect 3652 51365 3745 51451
rect 3831 51365 3913 51451
rect 3999 51365 4092 51451
rect 3652 49939 4092 51365
rect 3652 49853 3745 49939
rect 3831 49853 3913 49939
rect 3999 49853 4092 49939
rect 3652 48427 4092 49853
rect 3652 48341 3745 48427
rect 3831 48341 3913 48427
rect 3999 48341 4092 48427
rect 3652 46915 4092 48341
rect 3652 46829 3745 46915
rect 3831 46829 3913 46915
rect 3999 46829 4092 46915
rect 3652 45403 4092 46829
rect 3652 45317 3745 45403
rect 3831 45317 3913 45403
rect 3999 45317 4092 45403
rect 3652 43891 4092 45317
rect 3652 43805 3745 43891
rect 3831 43805 3913 43891
rect 3999 43805 4092 43891
rect 3652 42379 4092 43805
rect 3652 42293 3745 42379
rect 3831 42293 3913 42379
rect 3999 42293 4092 42379
rect 3652 40867 4092 42293
rect 3652 40781 3745 40867
rect 3831 40781 3913 40867
rect 3999 40781 4092 40867
rect 3652 39355 4092 40781
rect 3652 39269 3745 39355
rect 3831 39269 3913 39355
rect 3999 39269 4092 39355
rect 3652 37843 4092 39269
rect 3652 37757 3745 37843
rect 3831 37757 3913 37843
rect 3999 37757 4092 37843
rect 3652 36331 4092 37757
rect 3652 36245 3745 36331
rect 3831 36245 3913 36331
rect 3999 36245 4092 36331
rect 3652 34819 4092 36245
rect 3652 34733 3745 34819
rect 3831 34733 3913 34819
rect 3999 34733 4092 34819
rect 3652 33307 4092 34733
rect 3652 33221 3745 33307
rect 3831 33221 3913 33307
rect 3999 33221 4092 33307
rect 3652 31795 4092 33221
rect 3652 31709 3745 31795
rect 3831 31709 3913 31795
rect 3999 31709 4092 31795
rect 3652 30283 4092 31709
rect 3652 30197 3745 30283
rect 3831 30197 3913 30283
rect 3999 30197 4092 30283
rect 3652 28771 4092 30197
rect 3652 28685 3745 28771
rect 3831 28685 3913 28771
rect 3999 28685 4092 28771
rect 3652 27259 4092 28685
rect 3652 27173 3745 27259
rect 3831 27173 3913 27259
rect 3999 27173 4092 27259
rect 3652 25747 4092 27173
rect 3652 25661 3745 25747
rect 3831 25661 3913 25747
rect 3999 25661 4092 25747
rect 3652 24235 4092 25661
rect 3652 24149 3745 24235
rect 3831 24149 3913 24235
rect 3999 24149 4092 24235
rect 3652 22723 4092 24149
rect 3652 22637 3745 22723
rect 3831 22637 3913 22723
rect 3999 22637 4092 22723
rect 3652 21211 4092 22637
rect 3652 21125 3745 21211
rect 3831 21125 3913 21211
rect 3999 21125 4092 21211
rect 3652 19699 4092 21125
rect 3652 19613 3745 19699
rect 3831 19613 3913 19699
rect 3999 19613 4092 19699
rect 3652 18187 4092 19613
rect 3652 18101 3745 18187
rect 3831 18101 3913 18187
rect 3999 18101 4092 18187
rect 3652 16675 4092 18101
rect 3652 16589 3745 16675
rect 3831 16589 3913 16675
rect 3999 16589 4092 16675
rect 3652 15163 4092 16589
rect 3652 15077 3745 15163
rect 3831 15077 3913 15163
rect 3999 15077 4092 15163
rect 3652 13651 4092 15077
rect 3652 13565 3745 13651
rect 3831 13565 3913 13651
rect 3999 13565 4092 13651
rect 3652 12139 4092 13565
rect 3652 12053 3745 12139
rect 3831 12053 3913 12139
rect 3999 12053 4092 12139
rect 3652 10627 4092 12053
rect 3652 10541 3745 10627
rect 3831 10541 3913 10627
rect 3999 10541 4092 10627
rect 3652 9115 4092 10541
rect 3652 9029 3745 9115
rect 3831 9029 3913 9115
rect 3999 9029 4092 9115
rect 3652 7603 4092 9029
rect 3652 7517 3745 7603
rect 3831 7517 3913 7603
rect 3999 7517 4092 7603
rect 3652 6091 4092 7517
rect 3652 6005 3745 6091
rect 3831 6005 3913 6091
rect 3999 6005 4092 6091
rect 3652 4579 4092 6005
rect 3652 4493 3745 4579
rect 3831 4493 3913 4579
rect 3999 4493 4092 4579
rect 3652 3067 4092 4493
rect 3652 2981 3745 3067
rect 3831 2981 3913 3067
rect 3999 2981 4092 3067
rect 3652 1555 4092 2981
rect 3652 1469 3745 1555
rect 3831 1469 3913 1555
rect 3999 1469 4092 1555
rect 3652 0 4092 1469
rect 4892 83959 5332 86016
rect 18772 84715 19212 86016
rect 18772 84629 18865 84715
rect 18951 84629 19033 84715
rect 19119 84629 19212 84715
rect 4892 83873 4985 83959
rect 5071 83873 5153 83959
rect 5239 83873 5332 83959
rect 4892 82447 5332 83873
rect 12020 84127 12348 84248
rect 12020 84041 12141 84127
rect 12227 84041 12348 84127
rect 4892 82361 4985 82447
rect 5071 82361 5153 82447
rect 5239 82361 5332 82447
rect 4892 80935 5332 82361
rect 10652 83539 10980 83660
rect 10652 83453 10773 83539
rect 10859 83453 10980 83539
rect 4892 80849 4985 80935
rect 5071 80849 5153 80935
rect 5239 80849 5332 80935
rect 4892 79423 5332 80849
rect 4892 79337 4985 79423
rect 5071 79337 5153 79423
rect 5239 79337 5332 79423
rect 4892 77911 5332 79337
rect 4892 77825 4985 77911
rect 5071 77825 5153 77911
rect 5239 77825 5332 77911
rect 4892 76399 5332 77825
rect 4892 76313 4985 76399
rect 5071 76313 5153 76399
rect 5239 76313 5332 76399
rect 4892 74887 5332 76313
rect 4892 74801 4985 74887
rect 5071 74801 5153 74887
rect 5239 74801 5332 74887
rect 4892 73375 5332 74801
rect 4892 73289 4985 73375
rect 5071 73289 5153 73375
rect 5239 73289 5332 73375
rect 4892 71863 5332 73289
rect 4892 71777 4985 71863
rect 5071 71777 5153 71863
rect 5239 71777 5332 71863
rect 4892 70351 5332 71777
rect 4892 70265 4985 70351
rect 5071 70265 5153 70351
rect 5239 70265 5332 70351
rect 4892 68839 5332 70265
rect 4892 68753 4985 68839
rect 5071 68753 5153 68839
rect 5239 68753 5332 68839
rect 4892 67327 5332 68753
rect 4892 67241 4985 67327
rect 5071 67241 5153 67327
rect 5239 67241 5332 67327
rect 4892 65815 5332 67241
rect 8372 80851 8700 80972
rect 8372 80765 8493 80851
rect 8579 80765 8700 80851
rect 4892 65729 4985 65815
rect 5071 65729 5153 65815
rect 5239 65729 5332 65815
rect 4892 64303 5332 65729
rect 4892 64217 4985 64303
rect 5071 64217 5153 64303
rect 5239 64217 5332 64303
rect 4892 62791 5332 64217
rect 4892 62705 4985 62791
rect 5071 62705 5153 62791
rect 5239 62705 5332 62791
rect 4892 61279 5332 62705
rect 4892 61193 4985 61279
rect 5071 61193 5153 61279
rect 5239 61193 5332 61279
rect 4892 59767 5332 61193
rect 4892 59681 4985 59767
rect 5071 59681 5153 59767
rect 5239 59681 5332 59767
rect 4892 58255 5332 59681
rect 4892 58169 4985 58255
rect 5071 58169 5153 58255
rect 5239 58169 5332 58255
rect 4892 56743 5332 58169
rect 4892 56657 4985 56743
rect 5071 56657 5153 56743
rect 5239 56657 5332 56743
rect 4892 55231 5332 56657
rect 4892 55145 4985 55231
rect 5071 55145 5153 55231
rect 5239 55145 5332 55231
rect 4892 53719 5332 55145
rect 4892 53633 4985 53719
rect 5071 53633 5153 53719
rect 5239 53633 5332 53719
rect 4892 52207 5332 53633
rect 4892 52121 4985 52207
rect 5071 52121 5153 52207
rect 5239 52121 5332 52207
rect 4892 50695 5332 52121
rect 4892 50609 4985 50695
rect 5071 50609 5153 50695
rect 5239 50609 5332 50695
rect 4892 49183 5332 50609
rect 4892 49097 4985 49183
rect 5071 49097 5153 49183
rect 5239 49097 5332 49183
rect 4892 47671 5332 49097
rect 4892 47585 4985 47671
rect 5071 47585 5153 47671
rect 5239 47585 5332 47671
rect 4892 46159 5332 47585
rect 4892 46073 4985 46159
rect 5071 46073 5153 46159
rect 5239 46073 5332 46159
rect 4892 44647 5332 46073
rect 4892 44561 4985 44647
rect 5071 44561 5153 44647
rect 5239 44561 5332 44647
rect 4892 43135 5332 44561
rect 4892 43049 4985 43135
rect 5071 43049 5153 43135
rect 5239 43049 5332 43135
rect 4892 41623 5332 43049
rect 4892 41537 4985 41623
rect 5071 41537 5153 41623
rect 5239 41537 5332 41623
rect 4892 40111 5332 41537
rect 4892 40025 4985 40111
rect 5071 40025 5153 40111
rect 5239 40025 5332 40111
rect 4892 38599 5332 40025
rect 4892 38513 4985 38599
rect 5071 38513 5153 38599
rect 5239 38513 5332 38599
rect 4892 37087 5332 38513
rect 4892 37001 4985 37087
rect 5071 37001 5153 37087
rect 5239 37001 5332 37087
rect 4892 35575 5332 37001
rect 4892 35489 4985 35575
rect 5071 35489 5153 35575
rect 5239 35489 5332 35575
rect 4892 34063 5332 35489
rect 4892 33977 4985 34063
rect 5071 33977 5153 34063
rect 5239 33977 5332 34063
rect 4892 32551 5332 33977
rect 4892 32465 4985 32551
rect 5071 32465 5153 32551
rect 5239 32465 5332 32551
rect 4892 31039 5332 32465
rect 4892 30953 4985 31039
rect 5071 30953 5153 31039
rect 5239 30953 5332 31039
rect 4892 29527 5332 30953
rect 4892 29441 4985 29527
rect 5071 29441 5153 29527
rect 5239 29441 5332 29527
rect 4892 28015 5332 29441
rect 4892 27929 4985 28015
rect 5071 27929 5153 28015
rect 5239 27929 5332 28015
rect 4892 26503 5332 27929
rect 4892 26417 4985 26503
rect 5071 26417 5153 26503
rect 5239 26417 5332 26503
rect 4892 24991 5332 26417
rect 4892 24905 4985 24991
rect 5071 24905 5153 24991
rect 5239 24905 5332 24991
rect 4892 23479 5332 24905
rect 4892 23393 4985 23479
rect 5071 23393 5153 23479
rect 5239 23393 5332 23479
rect 4892 21967 5332 23393
rect 4892 21881 4985 21967
rect 5071 21881 5153 21967
rect 5239 21881 5332 21967
rect 4892 20455 5332 21881
rect 4892 20369 4985 20455
rect 5071 20369 5153 20455
rect 5239 20369 5332 20455
rect 4892 18943 5332 20369
rect 4892 18857 4985 18943
rect 5071 18857 5153 18943
rect 5239 18857 5332 18943
rect 4892 17431 5332 18857
rect 4892 17345 4985 17431
rect 5071 17345 5153 17431
rect 5239 17345 5332 17431
rect 4892 15919 5332 17345
rect 4892 15833 4985 15919
rect 5071 15833 5153 15919
rect 5239 15833 5332 15919
rect 4892 14407 5332 15833
rect 4892 14321 4985 14407
rect 5071 14321 5153 14407
rect 5239 14321 5332 14407
rect 4892 12895 5332 14321
rect 4892 12809 4985 12895
rect 5071 12809 5153 12895
rect 5239 12809 5332 12895
rect 4892 11383 5332 12809
rect 4892 11297 4985 11383
rect 5071 11297 5153 11383
rect 5239 11297 5332 11383
rect 4892 9871 5332 11297
rect 4892 9785 4985 9871
rect 5071 9785 5153 9871
rect 5239 9785 5332 9871
rect 4892 8359 5332 9785
rect 4892 8273 4985 8359
rect 5071 8273 5153 8359
rect 5239 8273 5332 8359
rect 4892 6847 5332 8273
rect 4892 6761 4985 6847
rect 5071 6761 5153 6847
rect 5239 6761 5332 6847
rect 4892 5335 5332 6761
rect 4892 5249 4985 5335
rect 5071 5249 5153 5335
rect 5239 5249 5332 5335
rect 4892 3823 5332 5249
rect 6548 65899 6876 66020
rect 6548 65813 6669 65899
rect 6755 65813 6876 65899
rect 6548 4831 6876 65813
rect 8372 48091 8700 80765
rect 8372 48005 8493 48091
rect 8579 48005 8700 48091
rect 8372 47884 8700 48005
rect 9740 79507 10068 79628
rect 9740 79421 9861 79507
rect 9947 79421 10068 79507
rect 9740 7435 10068 79421
rect 9740 7349 9861 7435
rect 9947 7349 10068 7435
rect 9740 7228 10068 7349
rect 10652 5671 10980 83453
rect 10652 5585 10773 5671
rect 10859 5585 10980 5671
rect 10652 5464 10980 5585
rect 6548 4745 6669 4831
rect 6755 4745 6876 4831
rect 6548 4624 6876 4745
rect 4892 3737 4985 3823
rect 5071 3737 5153 3823
rect 5239 3737 5332 3823
rect 4892 2311 5332 3737
rect 4892 2225 4985 2311
rect 5071 2225 5153 2311
rect 5239 2225 5332 2311
rect 4892 799 5332 2225
rect 12020 1891 12348 84041
rect 12020 1805 12141 1891
rect 12227 1805 12348 1891
rect 12020 1684 12348 1805
rect 12932 83371 13260 83492
rect 12932 83285 13053 83371
rect 13139 83285 13260 83371
rect 12932 1303 13260 83285
rect 18772 83203 19212 84629
rect 18772 83117 18865 83203
rect 18951 83117 19033 83203
rect 19119 83117 19212 83203
rect 18772 81691 19212 83117
rect 18772 81605 18865 81691
rect 18951 81605 19033 81691
rect 19119 81605 19212 81691
rect 16580 81103 16908 81224
rect 16580 81017 16701 81103
rect 16787 81017 16908 81103
rect 13844 77323 14172 77444
rect 13844 77237 13965 77323
rect 14051 77237 14172 77323
rect 13844 61111 14172 77237
rect 13844 61025 13965 61111
rect 14051 61025 14172 61111
rect 13844 60904 14172 61025
rect 15668 66991 15996 67112
rect 15668 66905 15789 66991
rect 15875 66905 15996 66991
rect 13844 56743 14172 56864
rect 13844 56657 13965 56743
rect 14051 56657 14172 56743
rect 13844 25243 14172 56657
rect 13844 25157 13965 25243
rect 14051 25157 14172 25243
rect 13844 25036 14172 25157
rect 12932 1217 13053 1303
rect 13139 1217 13260 1303
rect 12932 1096 13260 1217
rect 4892 713 4985 799
rect 5071 713 5153 799
rect 5239 713 5332 799
rect 4892 0 5332 713
rect 15668 799 15996 66905
rect 15668 713 15789 799
rect 15875 713 15996 799
rect 15668 592 15996 713
rect 16580 715 16908 81017
rect 16580 629 16701 715
rect 16787 629 16908 715
rect 16580 508 16908 629
rect 18772 80179 19212 81605
rect 18772 80093 18865 80179
rect 18951 80093 19033 80179
rect 19119 80093 19212 80179
rect 18772 78667 19212 80093
rect 18772 78581 18865 78667
rect 18951 78581 19033 78667
rect 19119 78581 19212 78667
rect 18772 77155 19212 78581
rect 18772 77069 18865 77155
rect 18951 77069 19033 77155
rect 19119 77069 19212 77155
rect 18772 75643 19212 77069
rect 18772 75557 18865 75643
rect 18951 75557 19033 75643
rect 19119 75557 19212 75643
rect 18772 74131 19212 75557
rect 18772 74045 18865 74131
rect 18951 74045 19033 74131
rect 19119 74045 19212 74131
rect 18772 72619 19212 74045
rect 18772 72533 18865 72619
rect 18951 72533 19033 72619
rect 19119 72533 19212 72619
rect 18772 71107 19212 72533
rect 18772 71021 18865 71107
rect 18951 71021 19033 71107
rect 19119 71021 19212 71107
rect 18772 69595 19212 71021
rect 18772 69509 18865 69595
rect 18951 69509 19033 69595
rect 19119 69509 19212 69595
rect 18772 68083 19212 69509
rect 18772 67997 18865 68083
rect 18951 67997 19033 68083
rect 19119 67997 19212 68083
rect 18772 66571 19212 67997
rect 18772 66485 18865 66571
rect 18951 66485 19033 66571
rect 19119 66485 19212 66571
rect 18772 65059 19212 66485
rect 18772 64973 18865 65059
rect 18951 64973 19033 65059
rect 19119 64973 19212 65059
rect 18772 63547 19212 64973
rect 18772 63461 18865 63547
rect 18951 63461 19033 63547
rect 19119 63461 19212 63547
rect 18772 62035 19212 63461
rect 18772 61949 18865 62035
rect 18951 61949 19033 62035
rect 19119 61949 19212 62035
rect 18772 60523 19212 61949
rect 18772 60437 18865 60523
rect 18951 60437 19033 60523
rect 19119 60437 19212 60523
rect 18772 59011 19212 60437
rect 18772 58925 18865 59011
rect 18951 58925 19033 59011
rect 19119 58925 19212 59011
rect 18772 57499 19212 58925
rect 18772 57413 18865 57499
rect 18951 57413 19033 57499
rect 19119 57413 19212 57499
rect 18772 55987 19212 57413
rect 18772 55901 18865 55987
rect 18951 55901 19033 55987
rect 19119 55901 19212 55987
rect 18772 54475 19212 55901
rect 18772 54389 18865 54475
rect 18951 54389 19033 54475
rect 19119 54389 19212 54475
rect 18772 52963 19212 54389
rect 18772 52877 18865 52963
rect 18951 52877 19033 52963
rect 19119 52877 19212 52963
rect 18772 51451 19212 52877
rect 18772 51365 18865 51451
rect 18951 51365 19033 51451
rect 19119 51365 19212 51451
rect 18772 49939 19212 51365
rect 18772 49853 18865 49939
rect 18951 49853 19033 49939
rect 19119 49853 19212 49939
rect 18772 48427 19212 49853
rect 18772 48341 18865 48427
rect 18951 48341 19033 48427
rect 19119 48341 19212 48427
rect 18772 46915 19212 48341
rect 18772 46829 18865 46915
rect 18951 46829 19033 46915
rect 19119 46829 19212 46915
rect 18772 45403 19212 46829
rect 18772 45317 18865 45403
rect 18951 45317 19033 45403
rect 19119 45317 19212 45403
rect 18772 43891 19212 45317
rect 18772 43805 18865 43891
rect 18951 43805 19033 43891
rect 19119 43805 19212 43891
rect 18772 42379 19212 43805
rect 18772 42293 18865 42379
rect 18951 42293 19033 42379
rect 19119 42293 19212 42379
rect 18772 40867 19212 42293
rect 18772 40781 18865 40867
rect 18951 40781 19033 40867
rect 19119 40781 19212 40867
rect 18772 39355 19212 40781
rect 18772 39269 18865 39355
rect 18951 39269 19033 39355
rect 19119 39269 19212 39355
rect 18772 37843 19212 39269
rect 18772 37757 18865 37843
rect 18951 37757 19033 37843
rect 19119 37757 19212 37843
rect 18772 36331 19212 37757
rect 18772 36245 18865 36331
rect 18951 36245 19033 36331
rect 19119 36245 19212 36331
rect 18772 34819 19212 36245
rect 18772 34733 18865 34819
rect 18951 34733 19033 34819
rect 19119 34733 19212 34819
rect 18772 33307 19212 34733
rect 18772 33221 18865 33307
rect 18951 33221 19033 33307
rect 19119 33221 19212 33307
rect 18772 31795 19212 33221
rect 18772 31709 18865 31795
rect 18951 31709 19033 31795
rect 19119 31709 19212 31795
rect 18772 30283 19212 31709
rect 18772 30197 18865 30283
rect 18951 30197 19033 30283
rect 19119 30197 19212 30283
rect 18772 28771 19212 30197
rect 18772 28685 18865 28771
rect 18951 28685 19033 28771
rect 19119 28685 19212 28771
rect 18772 27259 19212 28685
rect 18772 27173 18865 27259
rect 18951 27173 19033 27259
rect 19119 27173 19212 27259
rect 18772 25747 19212 27173
rect 18772 25661 18865 25747
rect 18951 25661 19033 25747
rect 19119 25661 19212 25747
rect 18772 24235 19212 25661
rect 18772 24149 18865 24235
rect 18951 24149 19033 24235
rect 19119 24149 19212 24235
rect 18772 22723 19212 24149
rect 18772 22637 18865 22723
rect 18951 22637 19033 22723
rect 19119 22637 19212 22723
rect 18772 21211 19212 22637
rect 18772 21125 18865 21211
rect 18951 21125 19033 21211
rect 19119 21125 19212 21211
rect 18772 19699 19212 21125
rect 18772 19613 18865 19699
rect 18951 19613 19033 19699
rect 19119 19613 19212 19699
rect 18772 18187 19212 19613
rect 18772 18101 18865 18187
rect 18951 18101 19033 18187
rect 19119 18101 19212 18187
rect 18772 16675 19212 18101
rect 18772 16589 18865 16675
rect 18951 16589 19033 16675
rect 19119 16589 19212 16675
rect 18772 15163 19212 16589
rect 18772 15077 18865 15163
rect 18951 15077 19033 15163
rect 19119 15077 19212 15163
rect 18772 13651 19212 15077
rect 18772 13565 18865 13651
rect 18951 13565 19033 13651
rect 19119 13565 19212 13651
rect 18772 12139 19212 13565
rect 18772 12053 18865 12139
rect 18951 12053 19033 12139
rect 19119 12053 19212 12139
rect 18772 10627 19212 12053
rect 18772 10541 18865 10627
rect 18951 10541 19033 10627
rect 19119 10541 19212 10627
rect 18772 9115 19212 10541
rect 18772 9029 18865 9115
rect 18951 9029 19033 9115
rect 19119 9029 19212 9115
rect 18772 7603 19212 9029
rect 18772 7517 18865 7603
rect 18951 7517 19033 7603
rect 19119 7517 19212 7603
rect 18772 6091 19212 7517
rect 18772 6005 18865 6091
rect 18951 6005 19033 6091
rect 19119 6005 19212 6091
rect 18772 4579 19212 6005
rect 18772 4493 18865 4579
rect 18951 4493 19033 4579
rect 19119 4493 19212 4579
rect 18772 3067 19212 4493
rect 18772 2981 18865 3067
rect 18951 2981 19033 3067
rect 19119 2981 19212 3067
rect 18772 1555 19212 2981
rect 18772 1469 18865 1555
rect 18951 1469 19033 1555
rect 19119 1469 19212 1555
rect 18772 0 19212 1469
rect 20012 83959 20452 86016
rect 20012 83873 20105 83959
rect 20191 83873 20273 83959
rect 20359 83873 20452 83959
rect 20012 82447 20452 83873
rect 20012 82361 20105 82447
rect 20191 82361 20273 82447
rect 20359 82361 20452 82447
rect 20012 80935 20452 82361
rect 20012 80849 20105 80935
rect 20191 80849 20273 80935
rect 20359 80849 20452 80935
rect 20012 79423 20452 80849
rect 20012 79337 20105 79423
rect 20191 79337 20273 79423
rect 20359 79337 20452 79423
rect 20012 77911 20452 79337
rect 20012 77825 20105 77911
rect 20191 77825 20273 77911
rect 20359 77825 20452 77911
rect 20012 76399 20452 77825
rect 20012 76313 20105 76399
rect 20191 76313 20273 76399
rect 20359 76313 20452 76399
rect 20012 74887 20452 76313
rect 20012 74801 20105 74887
rect 20191 74801 20273 74887
rect 20359 74801 20452 74887
rect 20012 73375 20452 74801
rect 20012 73289 20105 73375
rect 20191 73289 20273 73375
rect 20359 73289 20452 73375
rect 20012 71863 20452 73289
rect 20012 71777 20105 71863
rect 20191 71777 20273 71863
rect 20359 71777 20452 71863
rect 20012 70351 20452 71777
rect 20012 70265 20105 70351
rect 20191 70265 20273 70351
rect 20359 70265 20452 70351
rect 20012 68839 20452 70265
rect 20012 68753 20105 68839
rect 20191 68753 20273 68839
rect 20359 68753 20452 68839
rect 20012 67327 20452 68753
rect 20012 67241 20105 67327
rect 20191 67241 20273 67327
rect 20359 67241 20452 67327
rect 20012 65815 20452 67241
rect 20012 65729 20105 65815
rect 20191 65729 20273 65815
rect 20359 65729 20452 65815
rect 20012 64303 20452 65729
rect 20012 64217 20105 64303
rect 20191 64217 20273 64303
rect 20359 64217 20452 64303
rect 20012 62791 20452 64217
rect 20012 62705 20105 62791
rect 20191 62705 20273 62791
rect 20359 62705 20452 62791
rect 20012 61279 20452 62705
rect 20012 61193 20105 61279
rect 20191 61193 20273 61279
rect 20359 61193 20452 61279
rect 20012 59767 20452 61193
rect 20012 59681 20105 59767
rect 20191 59681 20273 59767
rect 20359 59681 20452 59767
rect 20012 58255 20452 59681
rect 20012 58169 20105 58255
rect 20191 58169 20273 58255
rect 20359 58169 20452 58255
rect 20012 56743 20452 58169
rect 20012 56657 20105 56743
rect 20191 56657 20273 56743
rect 20359 56657 20452 56743
rect 20012 55231 20452 56657
rect 20012 55145 20105 55231
rect 20191 55145 20273 55231
rect 20359 55145 20452 55231
rect 20012 53719 20452 55145
rect 20012 53633 20105 53719
rect 20191 53633 20273 53719
rect 20359 53633 20452 53719
rect 20012 52207 20452 53633
rect 20012 52121 20105 52207
rect 20191 52121 20273 52207
rect 20359 52121 20452 52207
rect 20012 50695 20452 52121
rect 20012 50609 20105 50695
rect 20191 50609 20273 50695
rect 20359 50609 20452 50695
rect 20012 49183 20452 50609
rect 20012 49097 20105 49183
rect 20191 49097 20273 49183
rect 20359 49097 20452 49183
rect 20012 47671 20452 49097
rect 20012 47585 20105 47671
rect 20191 47585 20273 47671
rect 20359 47585 20452 47671
rect 20012 46159 20452 47585
rect 20012 46073 20105 46159
rect 20191 46073 20273 46159
rect 20359 46073 20452 46159
rect 20012 44647 20452 46073
rect 20012 44561 20105 44647
rect 20191 44561 20273 44647
rect 20359 44561 20452 44647
rect 20012 43135 20452 44561
rect 20012 43049 20105 43135
rect 20191 43049 20273 43135
rect 20359 43049 20452 43135
rect 20012 41623 20452 43049
rect 20012 41537 20105 41623
rect 20191 41537 20273 41623
rect 20359 41537 20452 41623
rect 20012 40111 20452 41537
rect 20012 40025 20105 40111
rect 20191 40025 20273 40111
rect 20359 40025 20452 40111
rect 20012 38599 20452 40025
rect 20012 38513 20105 38599
rect 20191 38513 20273 38599
rect 20359 38513 20452 38599
rect 20012 37087 20452 38513
rect 20012 37001 20105 37087
rect 20191 37001 20273 37087
rect 20359 37001 20452 37087
rect 20012 35575 20452 37001
rect 20012 35489 20105 35575
rect 20191 35489 20273 35575
rect 20359 35489 20452 35575
rect 20012 34063 20452 35489
rect 20012 33977 20105 34063
rect 20191 33977 20273 34063
rect 20359 33977 20452 34063
rect 20012 32551 20452 33977
rect 20012 32465 20105 32551
rect 20191 32465 20273 32551
rect 20359 32465 20452 32551
rect 20012 31039 20452 32465
rect 20012 30953 20105 31039
rect 20191 30953 20273 31039
rect 20359 30953 20452 31039
rect 20012 29527 20452 30953
rect 20012 29441 20105 29527
rect 20191 29441 20273 29527
rect 20359 29441 20452 29527
rect 20012 28015 20452 29441
rect 20012 27929 20105 28015
rect 20191 27929 20273 28015
rect 20359 27929 20452 28015
rect 20012 26503 20452 27929
rect 20012 26417 20105 26503
rect 20191 26417 20273 26503
rect 20359 26417 20452 26503
rect 20012 24991 20452 26417
rect 20012 24905 20105 24991
rect 20191 24905 20273 24991
rect 20359 24905 20452 24991
rect 20012 23479 20452 24905
rect 20012 23393 20105 23479
rect 20191 23393 20273 23479
rect 20359 23393 20452 23479
rect 20012 21967 20452 23393
rect 20012 21881 20105 21967
rect 20191 21881 20273 21967
rect 20359 21881 20452 21967
rect 20012 20455 20452 21881
rect 20012 20369 20105 20455
rect 20191 20369 20273 20455
rect 20359 20369 20452 20455
rect 20012 18943 20452 20369
rect 20012 18857 20105 18943
rect 20191 18857 20273 18943
rect 20359 18857 20452 18943
rect 20012 17431 20452 18857
rect 20012 17345 20105 17431
rect 20191 17345 20273 17431
rect 20359 17345 20452 17431
rect 20012 15919 20452 17345
rect 20012 15833 20105 15919
rect 20191 15833 20273 15919
rect 20359 15833 20452 15919
rect 20012 14407 20452 15833
rect 20012 14321 20105 14407
rect 20191 14321 20273 14407
rect 20359 14321 20452 14407
rect 20012 12895 20452 14321
rect 20012 12809 20105 12895
rect 20191 12809 20273 12895
rect 20359 12809 20452 12895
rect 20012 11383 20452 12809
rect 20012 11297 20105 11383
rect 20191 11297 20273 11383
rect 20359 11297 20452 11383
rect 20012 9871 20452 11297
rect 20012 9785 20105 9871
rect 20191 9785 20273 9871
rect 20359 9785 20452 9871
rect 20012 8359 20452 9785
rect 20012 8273 20105 8359
rect 20191 8273 20273 8359
rect 20359 8273 20452 8359
rect 20012 6847 20452 8273
rect 20012 6761 20105 6847
rect 20191 6761 20273 6847
rect 20359 6761 20452 6847
rect 20012 5335 20452 6761
rect 20012 5249 20105 5335
rect 20191 5249 20273 5335
rect 20359 5249 20452 5335
rect 20012 3823 20452 5249
rect 20012 3737 20105 3823
rect 20191 3737 20273 3823
rect 20359 3737 20452 3823
rect 20012 2311 20452 3737
rect 20012 2225 20105 2311
rect 20191 2225 20273 2311
rect 20359 2225 20452 2311
rect 20012 799 20452 2225
rect 20012 713 20105 799
rect 20191 713 20273 799
rect 20359 713 20452 799
rect 20012 0 20452 713
use sg13g2_inv_1  _0297_
timestamp 1676382929
transform 1 0 6816 0 -1 40068
box -48 -56 336 834
use sg13g2_inv_1  _0298_
timestamp 1676382929
transform 1 0 2400 0 -1 40068
box -48 -56 336 834
use sg13g2_inv_1  _0299_
timestamp 1676382929
transform -1 0 9504 0 1 43092
box -48 -56 336 834
use sg13g2_inv_1  _0300_
timestamp 1676382929
transform 1 0 14592 0 -1 59724
box -48 -56 336 834
use sg13g2_inv_1  _0301_
timestamp 1676382929
transform -1 0 11328 0 1 70308
box -48 -56 336 834
use sg13g2_inv_1  _0302_
timestamp 1676382929
transform 1 0 15936 0 1 73332
box -48 -56 336 834
use sg13g2_inv_1  _0303_
timestamp 1676382929
transform -1 0 10656 0 -1 73332
box -48 -56 336 834
use sg13g2_inv_1  _0304_
timestamp 1676382929
transform -1 0 15936 0 -1 26460
box -48 -56 336 834
use sg13g2_inv_1  _0305_
timestamp 1676382929
transform 1 0 9984 0 -1 32508
box -48 -56 336 834
use sg13g2_inv_1  _0306_
timestamp 1676382929
transform 1 0 11424 0 -1 27972
box -48 -56 336 834
use sg13g2_inv_1  _0307_
timestamp 1676382929
transform 1 0 14304 0 1 21924
box -48 -56 336 834
use sg13g2_inv_1  _0308_
timestamp 1676382929
transform 1 0 8448 0 -1 77868
box -48 -56 336 834
use sg13g2_inv_1  _0309_
timestamp 1676382929
transform -1 0 9600 0 -1 50652
box -48 -56 336 834
use sg13g2_inv_1  _0310_
timestamp 1676382929
transform 1 0 9120 0 1 65772
box -48 -56 336 834
use sg13g2_inv_1  _0311_
timestamp 1676382929
transform 1 0 11712 0 -1 80892
box -48 -56 336 834
use sg13g2_inv_1  _0312_
timestamp 1676382929
transform -1 0 11808 0 1 71820
box -48 -56 336 834
use sg13g2_inv_1  _0313_
timestamp 1676382929
transform 1 0 15552 0 1 56700
box -48 -56 336 834
use sg13g2_inv_1  _0314_
timestamp 1676382929
transform 1 0 15552 0 -1 53676
box -48 -56 336 834
use sg13g2_inv_1  _0315_
timestamp 1676382929
transform -1 0 17760 0 -1 79380
box -48 -56 336 834
use sg13g2_inv_1  _0316_
timestamp 1676382929
transform 1 0 14688 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0317_
timestamp 1676382929
transform 1 0 17856 0 -1 23436
box -48 -56 336 834
use sg13g2_inv_1  _0318_
timestamp 1676382929
transform 1 0 7104 0 -1 35532
box -48 -56 336 834
use sg13g2_inv_1  _0319_
timestamp 1676382929
transform 1 0 5856 0 -1 34020
box -48 -56 336 834
use sg13g2_inv_1  _0320_
timestamp 1676382929
transform 1 0 5376 0 1 37044
box -48 -56 336 834
use sg13g2_inv_1  _0321_
timestamp 1676382929
transform 1 0 7104 0 1 35532
box -48 -56 336 834
use sg13g2_inv_1  _0322_
timestamp 1676382929
transform -1 0 12768 0 1 38556
box -48 -56 336 834
use sg13g2_inv_1  _0323_
timestamp 1676382929
transform 1 0 12864 0 -1 40068
box -48 -56 336 834
use sg13g2_inv_1  _0324_
timestamp 1676382929
transform -1 0 17856 0 1 17388
box -48 -56 336 834
use sg13g2_inv_1  _0325_
timestamp 1676382929
transform -1 0 19872 0 1 14364
box -48 -56 336 834
use sg13g2_inv_1  _0326_
timestamp 1676382929
transform -1 0 12576 0 1 27972
box -48 -56 336 834
use sg13g2_inv_1  _0327_
timestamp 1676382929
transform -1 0 14496 0 1 30996
box -48 -56 336 834
use sg13g2_inv_1  _0328_
timestamp 1676382929
transform 1 0 6624 0 1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0329_
timestamp 1676382929
transform 1 0 7200 0 -1 29484
box -48 -56 336 834
use sg13g2_inv_1  _0330_
timestamp 1676382929
transform -1 0 16224 0 1 20412
box -48 -56 336 834
use sg13g2_inv_1  _0331_
timestamp 1676382929
transform 1 0 17568 0 -1 18900
box -48 -56 336 834
use sg13g2_inv_1  _0332_
timestamp 1676382929
transform 1 0 6624 0 -1 41580
box -48 -56 336 834
use sg13g2_inv_1  _0333_
timestamp 1676382929
transform 1 0 7680 0 1 43092
box -48 -56 336 834
use sg13g2_inv_1  _0334_
timestamp 1676382929
transform 1 0 2784 0 -1 41580
box -48 -56 336 834
use sg13g2_inv_1  _0335_
timestamp 1676382929
transform -1 0 8256 0 1 73332
box -48 -56 336 834
use sg13g2_inv_1  _0336_
timestamp 1676382929
transform 1 0 6816 0 -1 67284
box -48 -56 336 834
use sg13g2_inv_1  _0337_
timestamp 1676382929
transform 1 0 10176 0 1 64260
box -48 -56 336 834
use sg13g2_inv_1  _0338_
timestamp 1676382929
transform 1 0 6144 0 1 74844
box -48 -56 336 834
use sg13g2_inv_1  _0339_
timestamp 1676382929
transform -1 0 5568 0 1 77868
box -48 -56 336 834
use sg13g2_mux4_1  _0340_
timestamp 1677257233
transform 1 0 1440 0 1 73332
box -48 -56 2064 834
use sg13g2_mux4_1  _0341_
timestamp 1677257233
transform 1 0 3168 0 -1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0342_
timestamp 1677257233
transform 1 0 2016 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0343_
timestamp 1677257233
transform -1 0 5664 0 -1 80892
box -48 -56 2064 834
use sg13g2_o21ai_1  _0344_
timestamp 1685175443
transform -1 0 10560 0 1 40068
box -48 -56 538 834
use sg13g2_nor2_1  _0345_
timestamp 1676627187
transform 1 0 8832 0 1 40068
box -48 -56 432 834
use sg13g2_a22oi_1  _0346_
timestamp 1685173987
transform -1 0 10080 0 1 40068
box -48 -56 624 834
use sg13g2_nand3_1  _0347_
timestamp 1683988354
transform -1 0 9696 0 -1 41580
box -48 -56 528 834
use sg13g2_nand2_1  _0348_
timestamp 1676557249
transform 1 0 9024 0 -1 43092
box -48 -56 432 834
use sg13g2_o21ai_1  _0349_
timestamp 1685175443
transform 1 0 9120 0 1 41580
box -48 -56 538 834
use sg13g2_nand3b_1  _0350_
timestamp 1676573470
transform 1 0 9696 0 -1 41580
box -48 -56 720 834
use sg13g2_o21ai_1  _0351_
timestamp 1685175443
transform 1 0 10368 0 -1 41580
box -48 -56 538 834
use sg13g2_o21ai_1  _0352_
timestamp 1685175443
transform 1 0 10848 0 -1 41580
box -48 -56 538 834
use sg13g2_mux4_1  _0353_
timestamp 1677257233
transform 1 0 7104 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0354_
timestamp 1677257233
transform 1 0 7104 0 1 38556
box -48 -56 2064 834
use sg13g2_mux2_1  _0355_
timestamp 1677247768
transform 1 0 9216 0 -1 40068
box -48 -56 1008 834
use sg13g2_o21ai_1  _0356_
timestamp 1685175443
transform 1 0 19776 0 1 40068
box -48 -56 538 834
use sg13g2_a21oi_1  _0357_
timestamp 1683973020
transform -1 0 19968 0 -1 41580
box -48 -56 528 834
use sg13g2_nand2b_1  _0358_
timestamp 1676567195
transform 1 0 15168 0 -1 61236
box -48 -56 528 834
use sg13g2_nor3_1  _0359_
timestamp 1676639442
transform -1 0 12960 0 -1 59724
box -48 -56 528 834
use sg13g2_a221oi_1  _0360_
timestamp 1685197497
transform 1 0 14400 0 -1 61236
box -48 -56 816 834
use sg13g2_mux4_1  _0361_
timestamp 1677257233
transform 1 0 14208 0 1 59724
box -48 -56 2064 834
use sg13g2_nand2b_1  _0362_
timestamp 1676567195
transform 1 0 12480 0 -1 27972
box -48 -56 528 834
use sg13g2_nor3_1  _0363_
timestamp 1676639442
transform -1 0 12672 0 1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  _0364_
timestamp 1685197497
transform -1 0 12480 0 -1 27972
box -48 -56 816 834
use sg13g2_mux4_1  _0365_
timestamp 1677257233
transform 1 0 10752 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0366_
timestamp 1677257233
transform 1 0 12480 0 1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0367_
timestamp 1677257233
transform 1 0 14208 0 -1 62748
box -48 -56 2064 834
use sg13g2_nand2b_1  _0368_
timestamp 1676567195
transform -1 0 11424 0 1 71820
box -48 -56 528 834
use sg13g2_nor3_1  _0369_
timestamp 1676639442
transform -1 0 11904 0 -1 71820
box -48 -56 528 834
use sg13g2_a221oi_1  _0370_
timestamp 1685197497
transform -1 0 11040 0 1 70308
box -48 -56 816 834
use sg13g2_mux4_1  _0371_
timestamp 1677257233
transform 1 0 8160 0 1 70308
box -48 -56 2064 834
use sg13g2_nor3_1  _0372_
timestamp 1676639442
transform 1 0 8160 0 -1 34020
box -48 -56 528 834
use sg13g2_nand2b_1  _0373_
timestamp 1676567195
transform 1 0 8640 0 -1 34020
box -48 -56 528 834
use sg13g2_a221oi_1  _0374_
timestamp 1685197497
transform 1 0 9216 0 -1 32508
box -48 -56 816 834
use sg13g2_mux4_1  _0375_
timestamp 1677257233
transform 1 0 8160 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0376_
timestamp 1677257233
transform 1 0 10944 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0377_
timestamp 1677257233
transform 1 0 7776 0 -1 71820
box -48 -56 2064 834
use sg13g2_nand2b_1  _0378_
timestamp 1676567195
transform 1 0 15168 0 1 74844
box -48 -56 528 834
use sg13g2_nor3_1  _0379_
timestamp 1676639442
transform -1 0 16032 0 -1 76356
box -48 -56 528 834
use sg13g2_a221oi_1  _0380_
timestamp 1685197497
transform 1 0 15648 0 1 74844
box -48 -56 816 834
use sg13g2_mux4_1  _0381_
timestamp 1677257233
transform 1 0 16512 0 1 74844
box -48 -56 2064 834
use sg13g2_nor3_1  _0382_
timestamp 1676639442
transform -1 0 15360 0 1 26460
box -48 -56 528 834
use sg13g2_nand2b_1  _0383_
timestamp 1676567195
transform 1 0 15168 0 -1 26460
box -48 -56 528 834
use sg13g2_a221oi_1  _0384_
timestamp 1685197497
transform -1 0 15072 0 -1 27972
box -48 -56 816 834
use sg13g2_mux4_1  _0385_
timestamp 1677257233
transform 1 0 12864 0 1 41580
box -48 -56 2064 834
use sg13g2_mux4_1  _0386_
timestamp 1677257233
transform 1 0 15168 0 1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0387_
timestamp 1677257233
transform 1 0 15648 0 1 79380
box -48 -56 2064 834
use sg13g2_mux4_1  _0388_
timestamp 1677257233
transform 1 0 1152 0 -1 80892
box -48 -56 2064 834
use sg13g2_mux4_1  _0389_
timestamp 1677257233
transform 1 0 2688 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0390_
timestamp 1677257233
transform 1 0 3936 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0391_
timestamp 1677257233
transform 1 0 2112 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0392_
timestamp 1677257233
transform 1 0 4512 0 1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0393_
timestamp 1677257233
transform 1 0 2304 0 -1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0394_
timestamp 1677257233
transform 1 0 1536 0 -1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0395_
timestamp 1677257233
transform -1 0 4800 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0396_
timestamp 1677257233
transform 1 0 1824 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0397_
timestamp 1677257233
transform 1 0 4128 0 -1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0398_
timestamp 1677257233
transform 1 0 1344 0 -1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0399_
timestamp 1677257233
transform 1 0 2784 0 1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0400_
timestamp 1677257233
transform 1 0 2880 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0401_
timestamp 1677257233
transform 1 0 2688 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0402_
timestamp 1677257233
transform 1 0 3264 0 1 80892
box -48 -56 2064 834
use sg13g2_mux4_1  _0403_
timestamp 1677257233
transform 1 0 2496 0 1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0404_
timestamp 1677257233
transform 1 0 5856 0 -1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0405_
timestamp 1677257233
transform 1 0 6816 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0406_
timestamp 1677257233
transform 1 0 5088 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0407_
timestamp 1677257233
transform 1 0 7296 0 -1 80892
box -48 -56 2064 834
use sg13g2_mux4_1  _0408_
timestamp 1677257233
transform 1 0 2496 0 1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0409_
timestamp 1677257233
transform 1 0 8064 0 -1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0410_
timestamp 1677257233
transform -1 0 6720 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0411_
timestamp 1677257233
transform 1 0 2208 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0412_
timestamp 1677257233
transform 1 0 4512 0 -1 82404
box -48 -56 2064 834
use sg13g2_mux4_1  _0413_
timestamp 1677257233
transform 1 0 1920 0 1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0414_
timestamp 1677257233
transform 1 0 5568 0 1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0415_
timestamp 1677257233
transform 1 0 5376 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0416_
timestamp 1677257233
transform 1 0 3168 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0417_
timestamp 1677257233
transform 1 0 6528 0 1 82404
box -48 -56 2064 834
use sg13g2_mux4_1  _0418_
timestamp 1677257233
transform 1 0 3264 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0419_
timestamp 1677257233
transform 1 0 6048 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0420_
timestamp 1677257233
transform 1 0 9504 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0421_
timestamp 1677257233
transform 1 0 8160 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _0422_
timestamp 1677257233
transform 1 0 9888 0 -1 83916
box -48 -56 2064 834
use sg13g2_mux4_1  _0423_
timestamp 1677257233
transform -1 0 5568 0 -1 73332
box -48 -56 2064 834
use sg13g2_nand2b_1  _0424_
timestamp 1676567195
transform 1 0 9600 0 -1 74844
box -48 -56 528 834
use sg13g2_nor3_1  _0425_
timestamp 1676639442
transform 1 0 9888 0 -1 73332
box -48 -56 528 834
use sg13g2_a221oi_1  _0426_
timestamp 1685197497
transform 1 0 9984 0 1 73332
box -48 -56 816 834
use sg13g2_mux4_1  _0427_
timestamp 1677257233
transform 1 0 13248 0 -1 74844
box -48 -56 2064 834
use sg13g2_nor3_1  _0428_
timestamp 1676639442
transform 1 0 14592 0 1 21924
box -48 -56 528 834
use sg13g2_nand2b_1  _0429_
timestamp 1676567195
transform 1 0 15264 0 1 20412
box -48 -56 528 834
use sg13g2_a221oi_1  _0430_
timestamp 1685197497
transform 1 0 15456 0 -1 21924
box -48 -56 816 834
use sg13g2_mux4_1  _0431_
timestamp 1677257233
transform 1 0 12480 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _0432_
timestamp 1677257233
transform 1 0 10368 0 -1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0433_
timestamp 1677257233
transform 1 0 11808 0 -1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0434_
timestamp 1677257233
transform 1 0 9984 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0435_
timestamp 1677257233
transform 1 0 14208 0 -1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0436_
timestamp 1677257233
transform 1 0 5856 0 -1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0437_
timestamp 1677257233
transform 1 0 7680 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0438_
timestamp 1677257233
transform 1 0 2592 0 1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0439_
timestamp 1677257233
transform 1 0 3360 0 -1 58212
box -48 -56 2064 834
use sg13g2_mux4_1  _0440_
timestamp 1677257233
transform 1 0 9888 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0441_
timestamp 1677257233
transform 1 0 5760 0 -1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0442_
timestamp 1677257233
transform 1 0 3648 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0443_
timestamp 1677257233
transform -1 0 4320 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0444_
timestamp 1677257233
transform 1 0 6048 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0445_
timestamp 1677257233
transform 1 0 7968 0 1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0446_
timestamp 1677257233
transform 1 0 2592 0 1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0447_
timestamp 1677257233
transform 1 0 3072 0 1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0448_
timestamp 1677257233
transform 1 0 10368 0 1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0449_
timestamp 1677257233
transform 1 0 6048 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0450_
timestamp 1677257233
transform 1 0 3552 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0451_
timestamp 1677257233
transform -1 0 4416 0 -1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0452_
timestamp 1677257233
transform 1 0 13824 0 -1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0453_
timestamp 1677257233
transform 1 0 9792 0 -1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0454_
timestamp 1677257233
transform 1 0 10176 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0455_
timestamp 1677257233
transform 1 0 10080 0 -1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0456_
timestamp 1677257233
transform 1 0 5856 0 1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0457_
timestamp 1677257233
transform 1 0 14304 0 -1 82404
box -48 -56 2064 834
use sg13g2_mux4_1  _0458_
timestamp 1677257233
transform -1 0 12096 0 -1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0459_
timestamp 1677257233
transform 1 0 10944 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0460_
timestamp 1677257233
transform 1 0 6336 0 -1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0461_
timestamp 1677257233
transform 1 0 12384 0 -1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0462_
timestamp 1677257233
transform 1 0 3840 0 1 50652
box -48 -56 2064 834
use sg13g2_mux4_1  _0463_
timestamp 1677257233
transform 1 0 10464 0 -1 79380
box -48 -56 2064 834
use sg13g2_mux4_1  _0464_
timestamp 1677257233
transform 1 0 6144 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0465_
timestamp 1677257233
transform 1 0 13728 0 1 82404
box -48 -56 2064 834
use sg13g2_mux4_1  _0466_
timestamp 1677257233
transform 1 0 13344 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0467_
timestamp 1677257233
transform 1 0 11328 0 1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0468_
timestamp 1677257233
transform 1 0 8160 0 1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0469_
timestamp 1677257233
transform 1 0 12576 0 1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0470_
timestamp 1677257233
transform 1 0 3072 0 1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0471_
timestamp 1677257233
transform 1 0 10368 0 1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0472_
timestamp 1677257233
transform -1 0 4896 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0473_
timestamp 1677257233
transform 1 0 13632 0 -1 80892
box -48 -56 2064 834
use sg13g2_mux4_1  _0474_
timestamp 1677257233
transform 1 0 9600 0 1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0475_
timestamp 1677257233
transform 1 0 11328 0 -1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0476_
timestamp 1677257233
transform 1 0 7872 0 1 53676
box -48 -56 2064 834
use sg13g2_mux4_1  _0477_
timestamp 1677257233
transform 1 0 12768 0 1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0478_
timestamp 1677257233
transform 1 0 3648 0 -1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0479_
timestamp 1677257233
transform 1 0 10560 0 -1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0480_
timestamp 1677257233
transform -1 0 4896 0 1 61236
box -48 -56 2064 834
use sg13g2_mux4_1  _0481_
timestamp 1677257233
transform 1 0 11328 0 1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0482_
timestamp 1677257233
transform 1 0 11424 0 -1 53676
box -48 -56 2064 834
use sg13g2_mux4_1  _0483_
timestamp 1677257233
transform 1 0 11328 0 1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0484_
timestamp 1677257233
transform 1 0 13152 0 1 77868
box -48 -56 2064 834
use sg13g2_mux4_1  _0485_
timestamp 1677257233
transform 1 0 11328 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0486_
timestamp 1677257233
transform 1 0 8064 0 1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0487_
timestamp 1677257233
transform 1 0 3840 0 -1 53676
box -48 -56 2064 834
use sg13g2_mux4_1  _0488_
timestamp 1677257233
transform 1 0 6432 0 1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0489_
timestamp 1677257233
transform 1 0 11616 0 1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0490_
timestamp 1677257233
transform 1 0 7776 0 -1 58212
box -48 -56 2064 834
use sg13g2_mux4_1  _0491_
timestamp 1677257233
transform 1 0 3456 0 -1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0492_
timestamp 1677257233
transform 1 0 3168 0 -1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0493_
timestamp 1677257233
transform 1 0 14784 0 1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0494_
timestamp 1677257233
transform 1 0 18144 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0495_
timestamp 1677257233
transform 1 0 17760 0 -1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0496_
timestamp 1677257233
transform 1 0 18336 0 1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0497_
timestamp 1677257233
transform 1 0 17376 0 1 64260
box -48 -56 2064 834
use sg13g2_mux4_1  _0498_
timestamp 1677257233
transform 1 0 15264 0 1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0499_
timestamp 1677257233
transform 1 0 17664 0 -1 55188
box -48 -56 2064 834
use sg13g2_mux4_1  _0500_
timestamp 1677257233
transform 1 0 18144 0 1 68796
box -48 -56 2064 834
use sg13g2_mux4_1  _0501_
timestamp 1677257233
transform 1 0 15552 0 1 71820
box -48 -56 2064 834
use sg13g2_mux4_1  _0502_
timestamp 1677257233
transform 1 0 17856 0 -1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0503_
timestamp 1677257233
transform 1 0 17664 0 -1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0504_
timestamp 1677257233
transform 1 0 18240 0 -1 79380
box -48 -56 2064 834
use sg13g2_mux4_1  _0505_
timestamp 1677257233
transform 1 0 14208 0 -1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0506_
timestamp 1677257233
transform 1 0 15264 0 -1 47628
box -48 -56 2064 834
use sg13g2_mux4_1  _0507_
timestamp 1677257233
transform 1 0 17280 0 1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0508_
timestamp 1677257233
transform 1 0 17760 0 -1 67284
box -48 -56 2064 834
use sg13g2_mux4_1  _0509_
timestamp 1677257233
transform 1 0 14784 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0510_
timestamp 1677257233
transform 1 0 18240 0 1 46116
box -48 -56 2064 834
use sg13g2_mux4_1  _0511_
timestamp 1677257233
transform 1 0 17760 0 1 62748
box -48 -56 2064 834
use sg13g2_mux4_1  _0512_
timestamp 1677257233
transform 1 0 18336 0 -1 74844
box -48 -56 2064 834
use sg13g2_mux4_1  _0513_
timestamp 1677257233
transform 1 0 17280 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0514_
timestamp 1677257233
transform 1 0 15264 0 -1 44604
box -48 -56 2064 834
use sg13g2_mux4_1  _0515_
timestamp 1677257233
transform 1 0 17664 0 1 56700
box -48 -56 2064 834
use sg13g2_mux4_1  _0516_
timestamp 1677257233
transform 1 0 18048 0 -1 70308
box -48 -56 2064 834
use sg13g2_mux4_1  _0517_
timestamp 1677257233
transform 1 0 15552 0 -1 73332
box -48 -56 2064 834
use sg13g2_mux4_1  _0518_
timestamp 1677257233
transform 1 0 17856 0 1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0519_
timestamp 1677257233
transform 1 0 17664 0 1 59724
box -48 -56 2064 834
use sg13g2_mux4_1  _0520_
timestamp 1677257233
transform 1 0 18240 0 1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0521_
timestamp 1677257233
transform 1 0 14112 0 -1 65772
box -48 -56 2064 834
use sg13g2_mux4_1  _0522_
timestamp 1677257233
transform 1 0 15360 0 -1 49140
box -48 -56 2064 834
use sg13g2_mux4_1  _0523_
timestamp 1677257233
transform 1 0 17184 0 -1 52164
box -48 -56 2064 834
use sg13g2_mux4_1  _0524_
timestamp 1677257233
transform 1 0 17760 0 1 67284
box -48 -56 2064 834
use sg13g2_nor3_1  _0525_
timestamp 1676639442
transform 1 0 6720 0 1 73332
box -48 -56 528 834
use sg13g2_nand2b_1  _0526_
timestamp 1676567195
transform 1 0 7584 0 -1 73332
box -48 -56 528 834
use sg13g2_a221oi_1  _0527_
timestamp 1685197497
transform 1 0 7200 0 1 73332
box -48 -56 816 834
use sg13g2_nor3_1  _0528_
timestamp 1676639442
transform 1 0 5568 0 -1 65772
box -48 -56 528 834
use sg13g2_nand2b_1  _0529_
timestamp 1676567195
transform 1 0 7392 0 1 65772
box -48 -56 528 834
use sg13g2_a221oi_1  _0530_
timestamp 1685197497
transform 1 0 6624 0 1 65772
box -48 -56 816 834
use sg13g2_nor3_1  _0531_
timestamp 1676639442
transform 1 0 8640 0 1 65772
box -48 -56 528 834
use sg13g2_nand2b_1  _0532_
timestamp 1676567195
transform -1 0 8640 0 -1 64260
box -48 -56 528 834
use sg13g2_a221oi_1  _0533_
timestamp 1685197497
transform 1 0 9408 0 1 64260
box -48 -56 816 834
use sg13g2_nor3_1  _0534_
timestamp 1676639442
transform -1 0 8256 0 -1 76356
box -48 -56 528 834
use sg13g2_nand2b_1  _0535_
timestamp 1676567195
transform -1 0 7776 0 -1 76356
box -48 -56 528 834
use sg13g2_a221oi_1  _0536_
timestamp 1685197497
transform -1 0 7296 0 -1 76356
box -48 -56 816 834
use sg13g2_nor3_1  _0537_
timestamp 1676639442
transform -1 0 2496 0 1 76356
box -48 -56 528 834
use sg13g2_nand2b_1  _0538_
timestamp 1676567195
transform 1 0 4800 0 1 77868
box -48 -56 528 834
use sg13g2_a221oi_1  _0539_
timestamp 1685197497
transform -1 0 2016 0 1 79380
box -48 -56 816 834
use sg13g2_mux2_1  _0540_
timestamp 1677247768
transform 1 0 7200 0 1 77868
box -48 -56 1008 834
use sg13g2_nor2b_1  _0541_
timestamp 1685181386
transform 1 0 6528 0 -1 80892
box -54 -56 528 834
use sg13g2_o21ai_1  _0542_
timestamp 1685175443
transform 1 0 6816 0 -1 79380
box -48 -56 538 834
use sg13g2_o21ai_1  _0543_
timestamp 1685175443
transform 1 0 7968 0 -1 77868
box -48 -56 538 834
use sg13g2_a21oi_1  _0544_
timestamp 1683973020
transform 1 0 7680 0 -1 79380
box -48 -56 528 834
use sg13g2_mux4_1  _0545_
timestamp 1677257233
transform 1 0 5952 0 -1 77868
box -48 -56 2064 834
use sg13g2_nor2_1  _0546_
timestamp 1676627187
transform -1 0 8544 0 -1 79380
box -48 -56 432 834
use sg13g2_nor2_1  _0547_
timestamp 1676627187
transform -1 0 6336 0 -1 80892
box -48 -56 432 834
use sg13g2_mux2_1  _0548_
timestamp 1677247768
transform -1 0 10560 0 -1 50652
box -48 -56 1008 834
use sg13g2_nor2b_1  _0549_
timestamp 1685181386
transform -1 0 9696 0 -1 52164
box -54 -56 528 834
use sg13g2_o21ai_1  _0550_
timestamp 1685175443
transform 1 0 9984 0 -1 49140
box -48 -56 538 834
use sg13g2_o21ai_1  _0551_
timestamp 1685175443
transform 1 0 10272 0 1 49140
box -48 -56 538 834
use sg13g2_a21oi_1  _0552_
timestamp 1683973020
transform -1 0 8352 0 -1 49140
box -48 -56 528 834
use sg13g2_mux4_1  _0553_
timestamp 1677257233
transform 1 0 8256 0 1 49140
box -48 -56 2064 834
use sg13g2_nor2_1  _0554_
timestamp 1676627187
transform -1 0 11136 0 1 49140
box -48 -56 432 834
use sg13g2_nor2_1  _0555_
timestamp 1676627187
transform 1 0 8544 0 1 47628
box -48 -56 432 834
use sg13g2_mux2_1  _0556_
timestamp 1677247768
transform 1 0 8736 0 -1 67284
box -48 -56 1008 834
use sg13g2_nor2b_1  _0557_
timestamp 1685181386
transform -1 0 7776 0 1 67284
box -54 -56 528 834
use sg13g2_o21ai_1  _0558_
timestamp 1685175443
transform 1 0 8736 0 1 68796
box -48 -56 538 834
use sg13g2_o21ai_1  _0559_
timestamp 1685175443
transform 1 0 9792 0 1 67284
box -48 -56 538 834
use sg13g2_a21oi_1  _0560_
timestamp 1683973020
transform 1 0 10272 0 1 67284
box -48 -56 528 834
use sg13g2_mux4_1  _0561_
timestamp 1677257233
transform 1 0 7776 0 1 67284
box -48 -56 2064 834
use sg13g2_nor2_1  _0562_
timestamp 1676627187
transform -1 0 10080 0 -1 68796
box -48 -56 432 834
use sg13g2_nor2_1  _0563_
timestamp 1676627187
transform 1 0 8352 0 1 68796
box -48 -56 432 834
use sg13g2_mux2_1  _0564_
timestamp 1677247768
transform 1 0 11232 0 -1 82404
box -48 -56 1008 834
use sg13g2_nor2b_1  _0565_
timestamp 1685181386
transform 1 0 10752 0 -1 82404
box -54 -56 528 834
use sg13g2_o21ai_1  _0566_
timestamp 1685175443
transform 1 0 11136 0 1 80892
box -48 -56 538 834
use sg13g2_o21ai_1  _0567_
timestamp 1685175443
transform 1 0 12384 0 1 82404
box -48 -56 538 834
use sg13g2_a21oi_1  _0568_
timestamp 1683973020
transform 1 0 11616 0 1 80892
box -48 -56 528 834
use sg13g2_mux4_1  _0569_
timestamp 1677257233
transform 1 0 9600 0 -1 80892
box -48 -56 2064 834
use sg13g2_nor2_1  _0570_
timestamp 1676627187
transform -1 0 12576 0 -1 82404
box -48 -56 432 834
use sg13g2_nor2_1  _0571_
timestamp 1676627187
transform 1 0 11616 0 1 83916
box -48 -56 432 834
use sg13g2_mux2_1  _0572_
timestamp 1677247768
transform -1 0 13344 0 1 70308
box -48 -56 1008 834
use sg13g2_nor2b_1  _0573_
timestamp 1685181386
transform -1 0 13920 0 1 71820
box -54 -56 528 834
use sg13g2_o21ai_1  _0574_
timestamp 1685175443
transform -1 0 13728 0 -1 73332
box -48 -56 538 834
use sg13g2_o21ai_1  _0575_
timestamp 1685175443
transform -1 0 13248 0 -1 74844
box -48 -56 538 834
use sg13g2_a21oi_1  _0576_
timestamp 1683973020
transform -1 0 12384 0 1 70308
box -48 -56 528 834
use sg13g2_mux4_1  _0577_
timestamp 1677257233
transform 1 0 12096 0 -1 71820
box -48 -56 2064 834
use sg13g2_nor2_1  _0578_
timestamp 1676627187
transform 1 0 14112 0 -1 71820
box -48 -56 432 834
use sg13g2_nor2_1  _0579_
timestamp 1676627187
transform -1 0 15360 0 1 70308
box -48 -56 432 834
use sg13g2_mux2_1  _0580_
timestamp 1677247768
transform 1 0 16224 0 -1 55188
box -48 -56 1008 834
use sg13g2_nor2b_1  _0581_
timestamp 1685181386
transform -1 0 16320 0 1 56700
box -54 -56 528 834
use sg13g2_o21ai_1  _0582_
timestamp 1685175443
transform 1 0 17088 0 -1 56700
box -48 -56 538 834
use sg13g2_o21ai_1  _0583_
timestamp 1685175443
transform 1 0 16800 0 1 56700
box -48 -56 538 834
use sg13g2_a21oi_1  _0584_
timestamp 1683973020
transform -1 0 16800 0 1 56700
box -48 -56 528 834
use sg13g2_mux4_1  _0585_
timestamp 1677257233
transform 1 0 15072 0 -1 56700
box -48 -56 2064 834
use sg13g2_nor2_1  _0586_
timestamp 1676627187
transform 1 0 17280 0 1 56700
box -48 -56 432 834
use sg13g2_nor2_1  _0587_
timestamp 1676627187
transform -1 0 17952 0 -1 56700
box -48 -56 432 834
use sg13g2_mux2_1  _0588_
timestamp 1677247768
transform 1 0 14688 0 1 52164
box -48 -56 1008 834
use sg13g2_nor2b_1  _0589_
timestamp 1685181386
transform -1 0 14496 0 -1 52164
box -54 -56 528 834
use sg13g2_o21ai_1  _0590_
timestamp 1685175443
transform 1 0 14400 0 1 50652
box -48 -56 538 834
use sg13g2_o21ai_1  _0591_
timestamp 1685175443
transform 1 0 14880 0 1 50652
box -48 -56 538 834
use sg13g2_a21oi_1  _0592_
timestamp 1683973020
transform 1 0 15360 0 1 50652
box -48 -56 528 834
use sg13g2_mux4_1  _0593_
timestamp 1677257233
transform 1 0 13536 0 -1 53676
box -48 -56 2064 834
use sg13g2_nor2_1  _0594_
timestamp 1676627187
transform -1 0 16896 0 -1 52164
box -48 -56 432 834
use sg13g2_nor2_1  _0595_
timestamp 1676627187
transform 1 0 16128 0 -1 52164
box -48 -56 432 834
use sg13g2_mux2_1  _0596_
timestamp 1677247768
transform -1 0 19968 0 1 82404
box -48 -56 1008 834
use sg13g2_nor2b_1  _0597_
timestamp 1685181386
transform -1 0 16608 0 -1 80892
box -54 -56 528 834
use sg13g2_o21ai_1  _0598_
timestamp 1685175443
transform 1 0 19680 0 1 79380
box -48 -56 538 834
use sg13g2_o21ai_1  _0599_
timestamp 1685175443
transform 1 0 17760 0 -1 79380
box -48 -56 538 834
use sg13g2_a21oi_1  _0600_
timestamp 1683973020
transform 1 0 19008 0 -1 83916
box -48 -56 528 834
use sg13g2_mux4_1  _0601_
timestamp 1677257233
transform -1 0 19680 0 1 79380
box -48 -56 2064 834
use sg13g2_nor2_1  _0602_
timestamp 1676627187
transform 1 0 15264 0 1 79380
box -48 -56 432 834
use sg13g2_nor2_1  _0603_
timestamp 1676627187
transform -1 0 16128 0 -1 80892
box -48 -56 432 834
use sg13g2_mux4_1  _0604_
timestamp 1677257233
transform 1 0 16608 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0605_
timestamp 1677257233
transform 1 0 12576 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0606_
timestamp 1677257233
transform 1 0 8640 0 1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0607_
timestamp 1677257233
transform 1 0 15552 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0608_
timestamp 1677257233
transform 1 0 8256 0 1 76356
box -48 -56 2064 834
use sg13g2_mux4_1  _0609_
timestamp 1677257233
transform 1 0 12096 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0610_
timestamp 1677257233
transform 1 0 9024 0 -1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0611_
timestamp 1677257233
transform 1 0 7392 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0612_
timestamp 1677257233
transform 1 0 12384 0 1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0613_
timestamp 1677257233
transform 1 0 2112 0 1 23436
box -48 -56 2064 834
use sg13g2_mux4_1  _0614_
timestamp 1677257233
transform 1 0 2208 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0615_
timestamp 1677257233
transform 1 0 1824 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0616_
timestamp 1677257233
transform 1 0 7680 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0617_
timestamp 1677257233
transform 1 0 7584 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0618_
timestamp 1677257233
transform 1 0 5568 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0619_
timestamp 1677257233
transform 1 0 4608 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0620_
timestamp 1677257233
transform 1 0 10368 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0621_
timestamp 1677257233
transform -1 0 20256 0 -1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0622_
timestamp 1677257233
transform 1 0 11040 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0623_
timestamp 1677257233
transform 1 0 8448 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0624_
timestamp 1677257233
transform 1 0 18048 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0625_
timestamp 1677257233
transform -1 0 10560 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0626_
timestamp 1677257233
transform 1 0 2496 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0627_
timestamp 1677257233
transform 1 0 2496 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0628_
timestamp 1677257233
transform 1 0 11616 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0629_
timestamp 1677257233
transform -1 0 8736 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0630_
timestamp 1677257233
transform -1 0 4128 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0631_
timestamp 1677257233
transform 1 0 3072 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0632_
timestamp 1677257233
transform 1 0 14304 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0633_
timestamp 1677257233
transform 1 0 8448 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0634_
timestamp 1677257233
transform -1 0 4416 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0635_
timestamp 1677257233
transform 1 0 2400 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0636_
timestamp 1677257233
transform 1 0 11616 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0637_
timestamp 1677257233
transform 1 0 6624 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0638_
timestamp 1677257233
transform 1 0 2112 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0639_
timestamp 1677257233
transform 1 0 2880 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0640_
timestamp 1677257233
transform 1 0 14400 0 1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0641_
timestamp 1677257233
transform 1 0 11904 0 -1 6804
box -48 -56 2064 834
use sg13g2_mux4_1  _0642_
timestamp 1677257233
transform 1 0 5472 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0643_
timestamp 1677257233
transform 1 0 7200 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0644_
timestamp 1677257233
transform 1 0 13824 0 1 5292
box -48 -56 2064 834
use sg13g2_mux4_1  _0645_
timestamp 1677257233
transform 1 0 18144 0 -1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0646_
timestamp 1677257233
transform -1 0 11808 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0647_
timestamp 1677257233
transform 1 0 8064 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0648_
timestamp 1677257233
transform 1 0 5088 0 -1 17388
box -48 -56 2064 834
use sg13g2_mux4_1  _0649_
timestamp 1677257233
transform 1 0 12576 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0650_
timestamp 1677257233
transform 1 0 4992 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0651_
timestamp 1677257233
transform 1 0 17760 0 -1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0652_
timestamp 1677257233
transform -1 0 16800 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0653_
timestamp 1677257233
transform 1 0 18048 0 1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0654_
timestamp 1677257233
transform 1 0 9792 0 -1 9828
box -48 -56 2064 834
use sg13g2_mux4_1  _0655_
timestamp 1677257233
transform 1 0 8544 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0656_
timestamp 1677257233
transform 1 0 2784 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0657_
timestamp 1677257233
transform 1 0 12384 0 1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0658_
timestamp 1677257233
transform 1 0 5280 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0659_
timestamp 1677257233
transform 1 0 17760 0 -1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0660_
timestamp 1677257233
transform 1 0 14976 0 1 2268
box -48 -56 2064 834
use sg13g2_mux4_1  _0661_
timestamp 1677257233
transform 1 0 18240 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0662_
timestamp 1677257233
transform 1 0 12384 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0663_
timestamp 1677257233
transform 1 0 8352 0 1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0664_
timestamp 1677257233
transform 1 0 2784 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0665_
timestamp 1677257233
transform 1 0 12576 0 -1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0666_
timestamp 1677257233
transform 1 0 5664 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0667_
timestamp 1677257233
transform 1 0 17664 0 1 3780
box -48 -56 2064 834
use sg13g2_mux4_1  _0668_
timestamp 1677257233
transform 1 0 14400 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0669_
timestamp 1677257233
transform 1 0 12192 0 1 8316
box -48 -56 2064 834
use sg13g2_mux4_1  _0670_
timestamp 1677257233
transform 1 0 10080 0 1 15876
box -48 -56 2064 834
use sg13g2_mux4_1  _0671_
timestamp 1677257233
transform 1 0 8352 0 1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0672_
timestamp 1677257233
transform 1 0 15840 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0673_
timestamp 1677257233
transform 1 0 10080 0 -1 11340
box -48 -56 2064 834
use sg13g2_mux4_1  _0674_
timestamp 1677257233
transform 1 0 5472 0 -1 18900
box -48 -56 2064 834
use sg13g2_mux4_1  _0675_
timestamp 1677257233
transform 1 0 5280 0 1 12852
box -48 -56 2064 834
use sg13g2_mux4_1  _0676_
timestamp 1677257233
transform 1 0 14976 0 1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0677_
timestamp 1677257233
transform 1 0 13056 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0678_
timestamp 1677257233
transform -1 0 4416 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0679_
timestamp 1677257233
transform 1 0 6048 0 -1 14364
box -48 -56 2064 834
use sg13g2_mux4_1  _0680_
timestamp 1677257233
transform 1 0 15360 0 1 15876
box -48 -56 2064 834
use sg13g2_nand3b_1  _0681_
timestamp 1676573470
transform -1 0 12672 0 -1 24948
box -48 -56 720 834
use sg13g2_nor2b_1  _0682_
timestamp 1685181386
transform 1 0 9888 0 -1 24948
box -54 -56 528 834
use sg13g2_a21oi_1  _0683_
timestamp 1683973020
transform 1 0 10368 0 1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _0684_
timestamp 1685175443
transform 1 0 11712 0 -1 23436
box -48 -56 538 834
use sg13g2_nand3b_1  _0685_
timestamp 1676573470
transform 1 0 5760 0 1 23436
box -48 -56 720 834
use sg13g2_nor2b_1  _0686_
timestamp 1685181386
transform 1 0 1536 0 -1 24948
box -54 -56 528 834
use sg13g2_a21oi_1  _0687_
timestamp 1683973020
transform 1 0 5280 0 -1 23436
box -48 -56 528 834
use sg13g2_o21ai_1  _0688_
timestamp 1685175443
transform 1 0 5760 0 -1 23436
box -48 -56 538 834
use sg13g2_nand3b_1  _0689_
timestamp 1676573470
transform 1 0 6240 0 -1 26460
box -48 -56 720 834
use sg13g2_nor2b_1  _0690_
timestamp 1685181386
transform -1 0 7872 0 1 26460
box -54 -56 528 834
use sg13g2_a21oi_1  _0691_
timestamp 1683973020
transform -1 0 7392 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _0692_
timestamp 1685175443
transform 1 0 6528 0 1 24948
box -48 -56 538 834
use sg13g2_nand3b_1  _0693_
timestamp 1676573470
transform -1 0 12192 0 1 38556
box -48 -56 720 834
use sg13g2_nor2_1  _0694_
timestamp 1676627187
transform 1 0 9504 0 1 38556
box -48 -56 432 834
use sg13g2_a21oi_1  _0695_
timestamp 1683973020
transform 1 0 10272 0 -1 40068
box -48 -56 528 834
use sg13g2_o21ai_1  _0696_
timestamp 1685175443
transform 1 0 11040 0 -1 38556
box -48 -56 538 834
use sg13g2_nand3b_1  _0697_
timestamp 1676573470
transform 1 0 9408 0 -1 26460
box -48 -56 720 834
use sg13g2_nor2b_1  _0698_
timestamp 1685181386
transform 1 0 7296 0 -1 26460
box -54 -56 528 834
use sg13g2_a21oi_1  _0699_
timestamp 1683973020
transform 1 0 8448 0 1 26460
box -48 -56 528 834
use sg13g2_o21ai_1  _0700_
timestamp 1685175443
transform 1 0 10080 0 -1 26460
box -48 -56 538 834
use sg13g2_mux4_1  _0701_
timestamp 1677257233
transform 1 0 17088 0 1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0702_
timestamp 1677257233
transform 1 0 14688 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0703_
timestamp 1677257233
transform 1 0 9120 0 -1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0704_
timestamp 1677257233
transform 1 0 18336 0 1 27972
box -48 -56 2064 834
use sg13g2_mux4_1  _0705_
timestamp 1677257233
transform 1 0 18336 0 -1 24948
box -48 -56 2064 834
use sg13g2_mux4_1  _0706_
timestamp 1677257233
transform 1 0 18240 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0707_
timestamp 1677257233
transform 1 0 12288 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0708_
timestamp 1677257233
transform 1 0 15360 0 -1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0709_
timestamp 1677257233
transform 1 0 17568 0 1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0710_
timestamp 1677257233
transform 1 0 14592 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0711_
timestamp 1677257233
transform 1 0 9408 0 1 30996
box -48 -56 2064 834
use sg13g2_mux4_1  _0712_
timestamp 1677257233
transform 1 0 18144 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0713_
timestamp 1677257233
transform 1 0 18240 0 -1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0714_
timestamp 1677257233
transform 1 0 17568 0 -1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0715_
timestamp 1677257233
transform 1 0 12096 0 -1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0716_
timestamp 1677257233
transform 1 0 15456 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0717_
timestamp 1677257233
transform 1 0 18048 0 -1 26460
box -48 -56 2064 834
use sg13g2_mux4_1  _0718_
timestamp 1677257233
transform 1 0 14592 0 1 32508
box -48 -56 2064 834
use sg13g2_mux4_1  _0719_
timestamp 1677257233
transform 1 0 9120 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0720_
timestamp 1677257233
transform 1 0 18240 0 1 38556
box -48 -56 2064 834
use sg13g2_mux4_1  _0721_
timestamp 1677257233
transform 1 0 18336 0 1 21924
box -48 -56 2064 834
use sg13g2_mux4_1  _0722_
timestamp 1677257233
transform 1 0 18336 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0723_
timestamp 1677257233
transform 1 0 12576 0 -1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0724_
timestamp 1677257233
transform 1 0 15552 0 1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0725_
timestamp 1677257233
transform 1 0 17760 0 -1 29484
box -48 -56 2064 834
use sg13g2_mux4_1  _0726_
timestamp 1677257233
transform 1 0 14496 0 -1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0727_
timestamp 1677257233
transform 1 0 9312 0 1 35532
box -48 -56 2064 834
use sg13g2_mux4_1  _0728_
timestamp 1677257233
transform 1 0 17952 0 -1 40068
box -48 -56 2064 834
use sg13g2_mux4_1  _0729_
timestamp 1677257233
transform 1 0 18336 0 -1 20412
box -48 -56 2064 834
use sg13g2_mux4_1  _0730_
timestamp 1677257233
transform 1 0 17664 0 1 34020
box -48 -56 2064 834
use sg13g2_mux4_1  _0731_
timestamp 1677257233
transform 1 0 12096 0 1 37044
box -48 -56 2064 834
use sg13g2_mux4_1  _0732_
timestamp 1677257233
transform 1 0 15552 0 1 41580
box -48 -56 2064 834
use sg13g2_o21ai_1  _0733_
timestamp 1685175443
transform 1 0 14496 0 1 23436
box -48 -56 538 834
use sg13g2_inv_1  _0734_
timestamp 1676382929
transform 1 0 17568 0 -1 23436
box -48 -56 336 834
use sg13g2_o21ai_1  _0735_
timestamp 1685175443
transform 1 0 15936 0 1 24948
box -48 -56 538 834
use sg13g2_mux2_1  _0736_
timestamp 1677247768
transform 1 0 14976 0 1 23436
box -48 -56 1008 834
use sg13g2_a21oi_1  _0737_
timestamp 1683973020
transform 1 0 16608 0 -1 23436
box -48 -56 528 834
use sg13g2_nor2_1  _0738_
timestamp 1676627187
transform 1 0 15072 0 1 24948
box -48 -56 432 834
use sg13g2_o21ai_1  _0739_
timestamp 1685175443
transform 1 0 17088 0 -1 23436
box -48 -56 538 834
use sg13g2_mux2_1  _0740_
timestamp 1677247768
transform -1 0 16896 0 1 23436
box -48 -56 1008 834
use sg13g2_o21ai_1  _0741_
timestamp 1685175443
transform 1 0 15456 0 1 24948
box -48 -56 538 834
use sg13g2_a21oi_1  _0742_
timestamp 1683973020
transform 1 0 15936 0 -1 26460
box -48 -56 528 834
use sg13g2_a21oi_1  _0743_
timestamp 1683973020
transform 1 0 16224 0 -1 24948
box -48 -56 528 834
use sg13g2_o21ai_1  _0744_
timestamp 1685175443
transform 1 0 5184 0 -1 35532
box -48 -56 538 834
use sg13g2_inv_1  _0745_
timestamp 1676382929
transform 1 0 5664 0 1 34020
box -48 -56 336 834
use sg13g2_o21ai_1  _0746_
timestamp 1685175443
transform -1 0 7392 0 1 34020
box -48 -56 538 834
use sg13g2_mux2_1  _0747_
timestamp 1677247768
transform 1 0 6144 0 1 32508
box -48 -56 1008 834
use sg13g2_a21oi_1  _0748_
timestamp 1683973020
transform 1 0 7584 0 -1 34020
box -48 -56 528 834
use sg13g2_nor2_1  _0749_
timestamp 1676627187
transform -1 0 6144 0 1 32508
box -48 -56 432 834
use sg13g2_o21ai_1  _0750_
timestamp 1685175443
transform -1 0 6432 0 1 34020
box -48 -56 538 834
use sg13g2_mux2_1  _0751_
timestamp 1677247768
transform 1 0 6144 0 -1 34020
box -48 -56 1008 834
use sg13g2_o21ai_1  _0752_
timestamp 1685175443
transform 1 0 7104 0 1 32508
box -48 -56 538 834
use sg13g2_a21oi_1  _0753_
timestamp 1683973020
transform -1 0 7584 0 -1 34020
box -48 -56 528 834
use sg13g2_a21oi_1  _0754_
timestamp 1683973020
transform -1 0 6912 0 1 34020
box -48 -56 528 834
use sg13g2_o21ai_1  _0755_
timestamp 1685175443
transform 1 0 5664 0 -1 35532
box -48 -56 538 834
use sg13g2_inv_1  _0756_
timestamp 1676382929
transform 1 0 7392 0 1 35532
box -48 -56 336 834
use sg13g2_o21ai_1  _0757_
timestamp 1685175443
transform 1 0 5664 0 1 35532
box -48 -56 538 834
use sg13g2_mux2_1  _0758_
timestamp 1677247768
transform 1 0 6144 0 1 35532
box -48 -56 1008 834
use sg13g2_a21oi_1  _0759_
timestamp 1683973020
transform 1 0 6048 0 -1 37044
box -48 -56 528 834
use sg13g2_nor2_1  _0760_
timestamp 1676627187
transform -1 0 7872 0 -1 37044
box -48 -56 432 834
use sg13g2_o21ai_1  _0761_
timestamp 1685175443
transform 1 0 5664 0 1 37044
box -48 -56 538 834
use sg13g2_mux2_1  _0762_
timestamp 1677247768
transform 1 0 6144 0 -1 35532
box -48 -56 1008 834
use sg13g2_o21ai_1  _0763_
timestamp 1685175443
transform -1 0 6624 0 1 37044
box -48 -56 538 834
use sg13g2_a21oi_1  _0764_
timestamp 1683973020
transform 1 0 7008 0 -1 37044
box -48 -56 528 834
use sg13g2_a21oi_1  _0765_
timestamp 1683973020
transform -1 0 7008 0 -1 37044
box -48 -56 528 834
use sg13g2_o21ai_1  _0766_
timestamp 1685175443
transform -1 0 13248 0 1 38556
box -48 -56 538 834
use sg13g2_inv_1  _0767_
timestamp 1676382929
transform -1 0 12480 0 1 38556
box -48 -56 336 834
use sg13g2_o21ai_1  _0768_
timestamp 1685175443
transform 1 0 15072 0 -1 40068
box -48 -56 538 834
use sg13g2_mux2_1  _0769_
timestamp 1677247768
transform 1 0 13248 0 1 38556
box -48 -56 1008 834
use sg13g2_a21oi_1  _0770_
timestamp 1683973020
transform 1 0 13536 0 -1 41580
box -48 -56 528 834
use sg13g2_nor2_1  _0771_
timestamp 1676627187
transform 1 0 13152 0 -1 41580
box -48 -56 432 834
use sg13g2_o21ai_1  _0772_
timestamp 1685175443
transform 1 0 14112 0 -1 40068
box -48 -56 538 834
use sg13g2_mux2_1  _0773_
timestamp 1677247768
transform 1 0 13152 0 -1 40068
box -48 -56 1008 834
use sg13g2_o21ai_1  _0774_
timestamp 1685175443
transform 1 0 14592 0 -1 40068
box -48 -56 538 834
use sg13g2_a21oi_1  _0775_
timestamp 1683973020
transform -1 0 14688 0 1 38556
box -48 -56 528 834
use sg13g2_a21oi_1  _0776_
timestamp 1683973020
transform 1 0 13248 0 1 40068
box -48 -56 528 834
use sg13g2_o21ai_1  _0777_
timestamp 1685175443
transform 1 0 19872 0 -1 17388
box -48 -56 538 834
use sg13g2_inv_1  _0778_
timestamp 1676382929
transform -1 0 20256 0 1 17388
box -48 -56 336 834
use sg13g2_o21ai_1  _0779_
timestamp 1685175443
transform 1 0 19488 0 1 17388
box -48 -56 538 834
use sg13g2_mux2_1  _0780_
timestamp 1677247768
transform 1 0 18912 0 -1 17388
box -48 -56 1008 834
use sg13g2_a21oi_1  _0781_
timestamp 1683973020
transform -1 0 20160 0 -1 15876
box -48 -56 528 834
use sg13g2_nor2_1  _0782_
timestamp 1676627187
transform -1 0 18720 0 -1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _0783_
timestamp 1685175443
transform 1 0 18240 0 1 15876
box -48 -56 538 834
use sg13g2_mux2_1  _0784_
timestamp 1677247768
transform 1 0 18720 0 1 15876
box -48 -56 1008 834
use sg13g2_o21ai_1  _0785_
timestamp 1685175443
transform 1 0 19680 0 1 15876
box -48 -56 538 834
use sg13g2_a21oi_1  _0786_
timestamp 1683973020
transform 1 0 19104 0 1 14364
box -48 -56 528 834
use sg13g2_a21oi_1  _0787_
timestamp 1683973020
transform -1 0 18240 0 1 15876
box -48 -56 528 834
use sg13g2_o21ai_1  _0788_
timestamp 1685175443
transform -1 0 13536 0 -1 30996
box -48 -56 538 834
use sg13g2_inv_1  _0789_
timestamp 1676382929
transform -1 0 11520 0 1 29484
box -48 -56 336 834
use sg13g2_o21ai_1  _0790_
timestamp 1685175443
transform 1 0 14688 0 -1 29484
box -48 -56 538 834
use sg13g2_mux2_1  _0791_
timestamp 1677247768
transform 1 0 13248 0 -1 29484
box -48 -56 1008 834
use sg13g2_a21oi_1  _0792_
timestamp 1683973020
transform 1 0 15168 0 -1 29484
box -48 -56 528 834
use sg13g2_nor2_1  _0793_
timestamp 1676627187
transform -1 0 13248 0 -1 29484
box -48 -56 432 834
use sg13g2_o21ai_1  _0794_
timestamp 1685175443
transform 1 0 14208 0 -1 29484
box -48 -56 538 834
use sg13g2_mux2_1  _0795_
timestamp 1677247768
transform 1 0 13248 0 1 29484
box -48 -56 1008 834
use sg13g2_o21ai_1  _0796_
timestamp 1685175443
transform -1 0 13056 0 1 27972
box -48 -56 538 834
use sg13g2_a21oi_1  _0797_
timestamp 1683973020
transform 1 0 13632 0 -1 27972
box -48 -56 528 834
use sg13g2_a21oi_1  _0798_
timestamp 1683973020
transform -1 0 13632 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _0799_
timestamp 1685175443
transform -1 0 6624 0 1 29484
box -48 -56 538 834
use sg13g2_inv_1  _0800_
timestamp 1676382929
transform -1 0 6240 0 -1 29484
box -48 -56 336 834
use sg13g2_o21ai_1  _0801_
timestamp 1685175443
transform 1 0 7680 0 1 27972
box -48 -56 538 834
use sg13g2_mux2_1  _0802_
timestamp 1677247768
transform -1 0 7200 0 -1 29484
box -48 -56 1008 834
use sg13g2_a21oi_1  _0803_
timestamp 1683973020
transform -1 0 6336 0 1 26460
box -48 -56 528 834
use sg13g2_nor2_1  _0804_
timestamp 1676627187
transform -1 0 6816 0 -1 27972
box -48 -56 432 834
use sg13g2_o21ai_1  _0805_
timestamp 1685175443
transform 1 0 6048 0 1 24948
box -48 -56 538 834
use sg13g2_mux2_1  _0806_
timestamp 1677247768
transform 1 0 6240 0 1 27972
box -48 -56 1008 834
use sg13g2_o21ai_1  _0807_
timestamp 1685175443
transform 1 0 6432 0 1 26460
box -48 -56 538 834
use sg13g2_a21oi_1  _0808_
timestamp 1683973020
transform 1 0 7200 0 1 27972
box -48 -56 528 834
use sg13g2_a21oi_1  _0809_
timestamp 1683973020
transform -1 0 7296 0 -1 27972
box -48 -56 528 834
use sg13g2_o21ai_1  _0810_
timestamp 1685175443
transform 1 0 16224 0 1 20412
box -48 -56 538 834
use sg13g2_inv_1  _0811_
timestamp 1676382929
transform 1 0 17856 0 -1 20412
box -48 -56 336 834
use sg13g2_o21ai_1  _0812_
timestamp 1685175443
transform -1 0 15936 0 1 18900
box -48 -56 538 834
use sg13g2_mux2_1  _0813_
timestamp 1677247768
transform 1 0 16416 0 -1 20412
box -48 -56 1008 834
use sg13g2_a21oi_1  _0814_
timestamp 1683973020
transform 1 0 17376 0 -1 20412
box -48 -56 528 834
use sg13g2_nor2_1  _0815_
timestamp 1676627187
transform -1 0 14976 0 1 18900
box -48 -56 432 834
use sg13g2_o21ai_1  _0816_
timestamp 1685175443
transform 1 0 16608 0 -1 18900
box -48 -56 538 834
use sg13g2_mux2_1  _0817_
timestamp 1677247768
transform 1 0 15936 0 1 18900
box -48 -56 1008 834
use sg13g2_o21ai_1  _0818_
timestamp 1685175443
transform 1 0 17088 0 -1 18900
box -48 -56 538 834
use sg13g2_a21oi_1  _0819_
timestamp 1683973020
transform -1 0 17184 0 1 20412
box -48 -56 528 834
use sg13g2_a21oi_1  _0820_
timestamp 1683973020
transform -1 0 15456 0 1 18900
box -48 -56 528 834
use sg13g2_nor2b_1  _0821_
timestamp 1685181386
transform -1 0 7584 0 1 40068
box -54 -56 528 834
use sg13g2_nand2b_1  _0822_
timestamp 1676567195
transform 1 0 7200 0 1 43092
box -48 -56 528 834
use sg13g2_nand2_1  _0823_
timestamp 1676557249
transform -1 0 4992 0 -1 41580
box -48 -56 432 834
use sg13g2_or2_1  _0824_
timestamp 1684236171
transform 1 0 6624 0 1 40068
box -48 -56 528 834
use sg13g2_a21oi_1  _0825_
timestamp 1683973020
transform -1 0 7200 0 1 43092
box -48 -56 528 834
use sg13g2_nand2_1  _0826_
timestamp 1676557249
transform -1 0 10944 0 1 40068
box -48 -56 432 834
use sg13g2_nand2_1  _0827_
timestamp 1676557249
transform 1 0 6336 0 1 43092
box -48 -56 432 834
use sg13g2_nand4_1  _0828_
timestamp 1685201930
transform 1 0 7680 0 -1 41580
box -48 -56 624 834
use sg13g2_a21oi_1  _0829_
timestamp 1683973020
transform 1 0 8256 0 1 40068
box -48 -56 528 834
use sg13g2_o21ai_1  _0830_
timestamp 1685175443
transform -1 0 9216 0 -1 41580
box -48 -56 538 834
use sg13g2_and2_1  _0831_
timestamp 1676901763
transform 1 0 5664 0 1 40068
box -48 -56 528 834
use sg13g2_a21oi_1  _0832_
timestamp 1683973020
transform 1 0 6144 0 1 40068
box -48 -56 528 834
use sg13g2_a22oi_1  _0833_
timestamp 1685173987
transform -1 0 7488 0 -1 41580
box -48 -56 624 834
use sg13g2_nand3_1  _0834_
timestamp 1683988354
transform 1 0 7776 0 1 40068
box -48 -56 528 834
use sg13g2_nand2b_1  _0835_
timestamp 1676567195
transform 1 0 6816 0 1 41580
box -48 -56 528 834
use sg13g2_or3_1  _0836_
timestamp 1677141922
transform 1 0 7296 0 1 41580
box -48 -56 720 834
use sg13g2_or2_1  _0837_
timestamp 1684236171
transform 1 0 7200 0 -1 43092
box -48 -56 528 834
use sg13g2_nand4_1  _0838_
timestamp 1685201930
transform 1 0 7968 0 1 41580
box -48 -56 624 834
use sg13g2_nand2b_1  _0839_
timestamp 1676567195
transform -1 0 9024 0 1 41580
box -48 -56 528 834
use sg13g2_nor3_1  _0840_
timestamp 1676639442
transform -1 0 8736 0 -1 41580
box -48 -56 528 834
use sg13g2_a221oi_1  _0841_
timestamp 1685197497
transform 1 0 8256 0 -1 43092
box -48 -56 816 834
use sg13g2_a21oi_1  _0842_
timestamp 1683973020
transform 1 0 7968 0 1 43092
box -48 -56 528 834
use sg13g2_a22oi_1  _0843_
timestamp 1685173987
transform 1 0 7680 0 -1 43092
box -48 -56 624 834
use sg13g2_mux4_1  _0844_
timestamp 1677257233
transform 1 0 2400 0 1 40068
box -48 -56 2064 834
use sg13g2_nand2_1  _0845_
timestamp 1676557249
transform -1 0 5184 0 -1 40068
box -48 -56 432 834
use sg13g2_nor2b_1  _0846_
timestamp 1685181386
transform -1 0 5376 0 1 40068
box -54 -56 528 834
use sg13g2_nor3_1  _0847_
timestamp 1676639442
transform 1 0 4320 0 -1 40068
box -48 -56 528 834
use sg13g2_nand2_1  _0848_
timestamp 1676557249
transform -1 0 4992 0 -1 43092
box -48 -56 432 834
use sg13g2_nand2b_1  _0849_
timestamp 1676567195
transform -1 0 2400 0 1 40068
box -48 -56 528 834
use sg13g2_a21oi_1  _0850_
timestamp 1683973020
transform -1 0 4224 0 1 43092
box -48 -56 528 834
use sg13g2_a22oi_1  _0851_
timestamp 1685173987
transform 1 0 3552 0 -1 41580
box -48 -56 624 834
use sg13g2_o21ai_1  _0852_
timestamp 1685175443
transform -1 0 4896 0 1 40068
box -48 -56 538 834
use sg13g2_nor3_1  _0853_
timestamp 1676639442
transform 1 0 3168 0 -1 43092
box -48 -56 528 834
use sg13g2_nor3_1  _0854_
timestamp 1676639442
transform 1 0 3072 0 -1 41580
box -48 -56 528 834
use sg13g2_o21ai_1  _0855_
timestamp 1685175443
transform -1 0 4992 0 1 41580
box -48 -56 538 834
use sg13g2_nor3_1  _0856_
timestamp 1676639442
transform 1 0 3264 0 1 41580
box -48 -56 528 834
use sg13g2_a21oi_1  _0857_
timestamp 1683973020
transform 1 0 2688 0 -1 43092
box -48 -56 528 834
use sg13g2_a21oi_1  _0858_
timestamp 1683973020
transform 1 0 2784 0 1 41580
box -48 -56 528 834
use sg13g2_nor3_1  _0859_
timestamp 1676639442
transform -1 0 4608 0 -1 41580
box -48 -56 528 834
use sg13g2_nor3_1  _0860_
timestamp 1676639442
transform 1 0 3744 0 1 41580
box -48 -56 528 834
use sg13g2_o21ai_1  _0861_
timestamp 1685175443
transform 1 0 3648 0 -1 43092
box -48 -56 538 834
use sg13g2_o21ai_1  _0862_
timestamp 1685175443
transform 1 0 4128 0 -1 43092
box -48 -56 538 834
use sg13g2_dlhq_1  _0863_
timestamp 1678805552
transform 1 0 14496 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0864_
timestamp 1678805552
transform 1 0 13920 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0865_
timestamp 1678805552
transform 1 0 9792 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0866_
timestamp 1678805552
transform 1 0 9312 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0867_
timestamp 1678805552
transform 1 0 12576 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _0868_
timestamp 1678805552
transform -1 0 14592 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _0869_
timestamp 1678805552
transform 1 0 8352 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0870_
timestamp 1678805552
transform 1 0 8256 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0871_
timestamp 1678805552
transform 1 0 8352 0 1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0872_
timestamp 1678805552
transform 1 0 10272 0 1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0873_
timestamp 1678805552
transform 1 0 3264 0 -1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0874_
timestamp 1678805552
transform 1 0 7296 0 -1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0875_
timestamp 1678805552
transform 1 0 3648 0 1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0876_
timestamp 1678805552
transform 1 0 4896 0 -1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0877_
timestamp 1678805552
transform 1 0 5664 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0878_
timestamp 1678805552
transform 1 0 7584 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0879_
timestamp 1678805552
transform 1 0 3360 0 1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0880_
timestamp 1678805552
transform 1 0 1632 0 -1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0881_
timestamp 1678805552
transform 1 0 4224 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0882_
timestamp 1678805552
transform 1 0 3456 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0883_
timestamp 1678805552
transform -1 0 6048 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0884_
timestamp 1678805552
transform 1 0 4704 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0885_
timestamp 1678805552
transform -1 0 10848 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0886_
timestamp 1678805552
transform 1 0 2016 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0887_
timestamp 1678805552
transform -1 0 18240 0 -1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0888_
timestamp 1678805552
transform 1 0 13344 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0889_
timestamp 1678805552
transform 1 0 11136 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0890_
timestamp 1678805552
transform 1 0 9504 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0891_
timestamp 1678805552
transform 1 0 12864 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0892_
timestamp 1678805552
transform 1 0 10848 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _0893_
timestamp 1678805552
transform 1 0 9696 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0894_
timestamp 1678805552
transform 1 0 8064 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0895_
timestamp 1678805552
transform 1 0 15264 0 1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0896_
timestamp 1678805552
transform 1 0 12576 0 -1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0897_
timestamp 1678805552
transform 1 0 11136 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0898_
timestamp 1678805552
transform 1 0 9312 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0899_
timestamp 1678805552
transform 1 0 12672 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0900_
timestamp 1678805552
transform 1 0 10752 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0901_
timestamp 1678805552
transform 1 0 11040 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0902_
timestamp 1678805552
transform 1 0 8736 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0903_
timestamp 1678805552
transform 1 0 13920 0 -1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0904_
timestamp 1678805552
transform 1 0 12096 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0905_
timestamp 1678805552
transform -1 0 13920 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0906_
timestamp 1678805552
transform 1 0 10080 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0907_
timestamp 1678805552
transform 1 0 13056 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _0908_
timestamp 1678805552
transform 1 0 10944 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0909_
timestamp 1678805552
transform 1 0 9408 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0910_
timestamp 1678805552
transform 1 0 7776 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _0911_
timestamp 1678805552
transform 1 0 13728 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0912_
timestamp 1678805552
transform 1 0 12000 0 -1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0913_
timestamp 1678805552
transform -1 0 14976 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0914_
timestamp 1678805552
transform 1 0 9696 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0915_
timestamp 1678805552
transform -1 0 16416 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _0916_
timestamp 1678805552
transform 1 0 11136 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _0917_
timestamp 1678805552
transform 1 0 11040 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0918_
timestamp 1678805552
transform 1 0 8928 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0919_
timestamp 1678805552
transform 1 0 1248 0 1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0920_
timestamp 1678805552
transform 1 0 1152 0 -1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0921_
timestamp 1678805552
transform 1 0 4992 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0922_
timestamp 1678805552
transform 1 0 4896 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0923_
timestamp 1678805552
transform 1 0 7776 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _0924_
timestamp 1678805552
transform 1 0 7680 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0925_
timestamp 1678805552
transform 1 0 5088 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0926_
timestamp 1678805552
transform 1 0 4992 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0927_
timestamp 1678805552
transform 1 0 5952 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0928_
timestamp 1678805552
transform 1 0 5856 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0929_
timestamp 1678805552
transform 1 0 18240 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0930_
timestamp 1678805552
transform 1 0 16128 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0931_
timestamp 1678805552
transform 1 0 17376 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _0932_
timestamp 1678805552
transform 1 0 15840 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0933_
timestamp 1678805552
transform 1 0 16032 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0934_
timestamp 1678805552
transform 1 0 14400 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0935_
timestamp 1678805552
transform 1 0 14400 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0936_
timestamp 1678805552
transform 1 0 12768 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0937_
timestamp 1678805552
transform 1 0 18528 0 -1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0938_
timestamp 1678805552
transform 1 0 16704 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0939_
timestamp 1678805552
transform 1 0 18048 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0940_
timestamp 1678805552
transform 1 0 16224 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0941_
timestamp 1678805552
transform 1 0 18240 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0942_
timestamp 1678805552
transform 1 0 16224 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0943_
timestamp 1678805552
transform 1 0 16128 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0944_
timestamp 1678805552
transform 1 0 13920 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0945_
timestamp 1678805552
transform 1 0 18432 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0946_
timestamp 1678805552
transform 1 0 16800 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0947_
timestamp 1678805552
transform 1 0 17952 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0948_
timestamp 1678805552
transform -1 0 18912 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0949_
timestamp 1678805552
transform 1 0 15648 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _0950_
timestamp 1678805552
transform 1 0 13632 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _0951_
timestamp 1678805552
transform 1 0 18336 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0952_
timestamp 1678805552
transform 1 0 15840 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _0953_
timestamp 1678805552
transform 1 0 18720 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0954_
timestamp 1678805552
transform -1 0 20256 0 -1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _0955_
timestamp 1678805552
transform 1 0 18240 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0956_
timestamp 1678805552
transform 1 0 16224 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _0957_
timestamp 1678805552
transform 1 0 18432 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _0958_
timestamp 1678805552
transform 1 0 17376 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _0959_
timestamp 1678805552
transform 1 0 14496 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0960_
timestamp 1678805552
transform 1 0 13152 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0961_
timestamp 1678805552
transform 1 0 18336 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0962_
timestamp 1678805552
transform 1 0 16128 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0963_
timestamp 1678805552
transform 1 0 17952 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0964_
timestamp 1678805552
transform 1 0 15648 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _0965_
timestamp 1678805552
transform -1 0 17856 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0966_
timestamp 1678805552
transform 1 0 14592 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0967_
timestamp 1678805552
transform 1 0 13152 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0968_
timestamp 1678805552
transform -1 0 15552 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0969_
timestamp 1678805552
transform 1 0 17184 0 1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _0970_
timestamp 1678805552
transform 1 0 16704 0 -1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _0971_
timestamp 1678805552
transform 1 0 18048 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0972_
timestamp 1678805552
transform 1 0 16224 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _0973_
timestamp 1678805552
transform 1 0 18240 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _0974_
timestamp 1678805552
transform -1 0 19296 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _0975_
timestamp 1678805552
transform 1 0 16128 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0976_
timestamp 1678805552
transform 1 0 14208 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _0977_
timestamp 1678805552
transform 1 0 18528 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0978_
timestamp 1678805552
transform 1 0 16704 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _0979_
timestamp 1678805552
transform 1 0 18048 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0980_
timestamp 1678805552
transform 1 0 15744 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _0981_
timestamp 1678805552
transform 1 0 15744 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _0982_
timestamp 1678805552
transform 1 0 13728 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _0983_
timestamp 1678805552
transform 1 0 18432 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0984_
timestamp 1678805552
transform 1 0 15840 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _0985_
timestamp 1678805552
transform 1 0 18624 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _0986_
timestamp 1678805552
transform -1 0 19392 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _0987_
timestamp 1678805552
transform 1 0 16608 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0988_
timestamp 1678805552
transform -1 0 19488 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _0989_
timestamp 1678805552
transform 1 0 18528 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _0990_
timestamp 1678805552
transform -1 0 19488 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _0991_
timestamp 1678805552
transform 1 0 13920 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _0992_
timestamp 1678805552
transform 1 0 13344 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _0993_
timestamp 1678805552
transform 1 0 1344 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _0994_
timestamp 1678805552
transform 1 0 3744 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _0995_
timestamp 1678805552
transform 1 0 1536 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0996_
timestamp 1678805552
transform 1 0 4320 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _0997_
timestamp 1678805552
transform 1 0 6240 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0998_
timestamp 1678805552
transform 1 0 7968 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _0999_
timestamp 1678805552
transform 1 0 10272 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1000_
timestamp 1678805552
transform 1 0 12192 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1001_
timestamp 1678805552
transform 1 0 6816 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1002_
timestamp 1678805552
transform 1 0 5088 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1003_
timestamp 1678805552
transform 1 0 4320 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1004_
timestamp 1678805552
transform 1 0 2016 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1005_
timestamp 1678805552
transform 1 0 6432 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1006_
timestamp 1678805552
transform 1 0 8448 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1007_
timestamp 1678805552
transform 1 0 10080 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1008_
timestamp 1678805552
transform 1 0 11808 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1009_
timestamp 1678805552
transform -1 0 15744 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1010_
timestamp 1678805552
transform 1 0 12480 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1011_
timestamp 1678805552
transform 1 0 11712 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1012_
timestamp 1678805552
transform 1 0 9984 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1013_
timestamp 1678805552
transform 1 0 11520 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1014_
timestamp 1678805552
transform 1 0 9792 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1015_
timestamp 1678805552
transform 1 0 12096 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _1016_
timestamp 1678805552
transform 1 0 10080 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _1017_
timestamp 1678805552
transform -1 0 4224 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1018_
timestamp 1678805552
transform 1 0 1344 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1019_
timestamp 1678805552
transform 1 0 4320 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1020_
timestamp 1678805552
transform 1 0 1920 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1021_
timestamp 1678805552
transform 1 0 8352 0 -1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1022_
timestamp 1678805552
transform 1 0 6240 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1023_
timestamp 1678805552
transform -1 0 12192 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1024_
timestamp 1678805552
transform 1 0 8640 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1025_
timestamp 1678805552
transform 1 0 1824 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1026_
timestamp 1678805552
transform 1 0 1248 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1027_
timestamp 1678805552
transform 1 0 3072 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1028_
timestamp 1678805552
transform 1 0 1440 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1029_
timestamp 1678805552
transform 1 0 8160 0 -1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1030_
timestamp 1678805552
transform 1 0 6528 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1031_
timestamp 1678805552
transform 1 0 13632 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1032_
timestamp 1678805552
transform 1 0 12288 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1033_
timestamp 1678805552
transform 1 0 6432 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1034_
timestamp 1678805552
transform 1 0 3456 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1035_
timestamp 1678805552
transform 1 0 4224 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1036_
timestamp 1678805552
transform 1 0 1440 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1037_
timestamp 1678805552
transform 1 0 6432 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1038_
timestamp 1678805552
transform 1 0 4704 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1039_
timestamp 1678805552
transform 1 0 9696 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1040_
timestamp 1678805552
transform 1 0 8064 0 1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1041_
timestamp 1678805552
transform 1 0 5952 0 -1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1042_
timestamp 1678805552
transform 1 0 4224 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1043_
timestamp 1678805552
transform 1 0 10560 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1044_
timestamp 1678805552
transform 1 0 8928 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1045_
timestamp 1678805552
transform 1 0 10272 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1046_
timestamp 1678805552
transform 1 0 8448 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1047_
timestamp 1678805552
transform 1 0 14400 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1048_
timestamp 1678805552
transform 1 0 12576 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1049_
timestamp 1678805552
transform 1 0 2496 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1050_
timestamp 1678805552
transform 1 0 1152 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1051_
timestamp 1678805552
transform 1 0 4032 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1052_
timestamp 1678805552
transform 1 0 1920 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1053_
timestamp 1678805552
transform 1 0 6336 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1054_
timestamp 1678805552
transform 1 0 4704 0 1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1055_
timestamp 1678805552
transform 1 0 10944 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1056_
timestamp 1678805552
transform 1 0 8832 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1057_
timestamp 1678805552
transform 1 0 1440 0 1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1058_
timestamp 1678805552
transform 1 0 1248 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1059_
timestamp 1678805552
transform 1 0 2592 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1060_
timestamp 1678805552
transform 1 0 1152 0 1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1061_
timestamp 1678805552
transform 1 0 8448 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1062_
timestamp 1678805552
transform 1 0 6336 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1063_
timestamp 1678805552
transform 1 0 6144 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1064_
timestamp 1678805552
transform 1 0 4608 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1065_
timestamp 1678805552
transform 1 0 1344 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1066_
timestamp 1678805552
transform 1 0 1152 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1067_
timestamp 1678805552
transform 1 0 4128 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1068_
timestamp 1678805552
transform 1 0 1824 0 -1 47628
box -50 -56 1692 834
use sg13g2_dlhq_1  _1069_
timestamp 1678805552
transform 1 0 5856 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1070_
timestamp 1678805552
transform 1 0 4608 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1071_
timestamp 1678805552
transform 1 0 9984 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1072_
timestamp 1678805552
transform 1 0 8256 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1073_
timestamp 1678805552
transform 1 0 2976 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1074_
timestamp 1678805552
transform 1 0 1632 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1075_
timestamp 1678805552
transform 1 0 2496 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1076_
timestamp 1678805552
transform 1 0 1152 0 1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1077_
timestamp 1678805552
transform 1 0 8064 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1078_
timestamp 1678805552
transform 1 0 6048 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1079_
timestamp 1678805552
transform 1 0 5952 0 -1 56700
box -50 -56 1692 834
use sg13g2_dlhq_1  _1080_
timestamp 1678805552
transform 1 0 4608 0 1 55188
box -50 -56 1692 834
use sg13g2_dlhq_1  _1081_
timestamp 1678805552
transform 1 0 13152 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1082_
timestamp 1678805552
transform 1 0 14784 0 1 53676
box -50 -56 1692 834
use sg13g2_dlhq_1  _1083_
timestamp 1678805552
transform 1 0 8640 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1084_
timestamp 1678805552
transform 1 0 10272 0 -1 46116
box -50 -56 1692 834
use sg13g2_dlhq_1  _1085_
timestamp 1678805552
transform 1 0 10176 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1086_
timestamp 1678805552
transform 1 0 12096 0 1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1087_
timestamp 1678805552
transform 1 0 8736 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1088_
timestamp 1678805552
transform 1 0 11040 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1089_
timestamp 1678805552
transform 1 0 13632 0 1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _1090_
timestamp 1678805552
transform 1 0 16416 0 -1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _1091_
timestamp 1678805552
transform 1 0 17376 0 1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _1092_
timestamp 1678805552
transform 1 0 14496 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1093_
timestamp 1678805552
transform 1 0 12192 0 -1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1094_
timestamp 1678805552
transform 1 0 12864 0 1 52164
box -50 -56 1692 834
use sg13g2_dlhq_1  _1095_
timestamp 1678805552
transform 1 0 15648 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1096_
timestamp 1678805552
transform 1 0 14016 0 -1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1097_
timestamp 1678805552
transform 1 0 15264 0 1 58212
box -50 -56 1692 834
use sg13g2_dlhq_1  _1098_
timestamp 1678805552
transform 1 0 11808 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1099_
timestamp 1678805552
transform 1 0 11616 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1100_
timestamp 1678805552
transform 1 0 10752 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1101_
timestamp 1678805552
transform 1 0 6144 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1102_
timestamp 1678805552
transform 1 0 4704 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1103_
timestamp 1678805552
transform 1 0 6048 0 -1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1104_
timestamp 1678805552
transform 1 0 3936 0 1 64260
box -50 -56 1692 834
use sg13g2_dlhq_1  _1105_
timestamp 1678805552
transform 1 0 7968 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1106_
timestamp 1678805552
transform 1 0 6432 0 -1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1107_
timestamp 1678805552
transform 1 0 4512 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1108_
timestamp 1678805552
transform 1 0 6432 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1109_
timestamp 1678805552
transform -1 0 5376 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1110_
timestamp 1678805552
transform -1 0 11616 0 1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _1111_
timestamp 1678805552
transform 1 0 1632 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1112_
timestamp 1678805552
transform 1 0 1152 0 -1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1113_
timestamp 1678805552
transform 1 0 3264 0 1 65772
box -50 -56 1692 834
use sg13g2_dlhq_1  _1114_
timestamp 1678805552
transform 1 0 1152 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1115_
timestamp 1678805552
transform -1 0 4800 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _1116_
timestamp 1678805552
transform 1 0 1152 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1117_
timestamp 1678805552
transform 1 0 15840 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1118_
timestamp 1678805552
transform 1 0 15456 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1119_
timestamp 1678805552
transform 1 0 8640 0 -1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1120_
timestamp 1678805552
transform 1 0 6528 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1121_
timestamp 1678805552
transform 1 0 14880 0 -1 59724
box -50 -56 1692 834
use sg13g2_dlhq_1  _1122_
timestamp 1678805552
transform 1 0 12768 0 -1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1123_
timestamp 1678805552
transform 1 0 12384 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1124_
timestamp 1678805552
transform 1 0 13440 0 1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1125_
timestamp 1678805552
transform 1 0 8640 0 1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _1126_
timestamp 1678805552
transform 1 0 7488 0 -1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _1127_
timestamp 1678805552
transform 1 0 9120 0 -1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _1128_
timestamp 1678805552
transform 1 0 8064 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1129_
timestamp 1678805552
transform 1 0 6432 0 -1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1130_
timestamp 1678805552
transform 1 0 7104 0 -1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1131_
timestamp 1678805552
transform 1 0 8352 0 -1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1132_
timestamp 1678805552
transform 1 0 6624 0 1 49140
box -50 -56 1692 834
use sg13g2_dlhq_1  _1133_
timestamp 1678805552
transform 1 0 7680 0 -1 50652
box -50 -56 1692 834
use sg13g2_dlhq_1  _1134_
timestamp 1678805552
transform 1 0 5664 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1135_
timestamp 1678805552
transform 1 0 5568 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1136_
timestamp 1678805552
transform 1 0 4896 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1137_
timestamp 1678805552
transform -1 0 5568 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1138_
timestamp 1678805552
transform -1 0 6720 0 1 73332
box -50 -56 1692 834
use sg13g2_dlhq_1  _1139_
timestamp 1678805552
transform 1 0 3072 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1140_
timestamp 1678805552
transform 1 0 1824 0 -1 74844
box -50 -56 1692 834
use sg13g2_dlhq_1  _1141_
timestamp 1678805552
transform 1 0 1728 0 1 67284
box -50 -56 1692 834
use sg13g2_dlhq_1  _1142_
timestamp 1678805552
transform 1 0 1152 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1143_
timestamp 1678805552
transform 1 0 2880 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1144_
timestamp 1678805552
transform 1 0 1152 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1145_
timestamp 1678805552
transform 1 0 3168 0 -1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1146_
timestamp 1678805552
transform 1 0 1152 0 1 80892
box -50 -56 1692 834
use sg13g2_dlhq_1  _1147_
timestamp 1678805552
transform 1 0 1536 0 -1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _1148_
timestamp 1678805552
transform 1 0 1152 0 -1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1149_
timestamp 1678805552
transform 1 0 2784 0 1 68796
box -50 -56 1692 834
use sg13g2_dlhq_1  _1150_
timestamp 1678805552
transform 1 0 1152 0 1 70308
box -50 -56 1692 834
use sg13g2_dlhq_1  _1151_
timestamp 1678805552
transform 1 0 2016 0 1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _1152_
timestamp 1678805552
transform -1 0 6912 0 1 83916
box -50 -56 1692 834
use sg13g2_dlhq_1  _1153_
timestamp 1678805552
transform 1 0 15744 0 1 82404
box -50 -56 1692 834
use sg13g2_dlhq_1  _1154_
timestamp 1678805552
transform 1 0 13632 0 1 79380
box -50 -56 1692 834
use sg13g2_dlhq_1  _1155_
timestamp 1678805552
transform 1 0 7680 0 1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1156_
timestamp 1678805552
transform 1 0 6144 0 -1 71820
box -50 -56 1692 834
use sg13g2_dlhq_1  _1157_
timestamp 1678805552
transform 1 0 14784 0 1 62748
box -50 -56 1692 834
use sg13g2_dlhq_1  _1158_
timestamp 1678805552
transform 1 0 13152 0 1 61236
box -50 -56 1692 834
use sg13g2_dlhq_1  _1159_
timestamp 1678805552
transform 1 0 6624 0 1 76356
box -50 -56 1692 834
use sg13g2_dlhq_1  _1160_
timestamp 1678805552
transform 1 0 8352 0 1 77868
box -50 -56 1692 834
use sg13g2_dlhq_1  _1161_
timestamp 1678805552
transform 1 0 13248 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1162_
timestamp 1678805552
transform 1 0 13536 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1163_
timestamp 1678805552
transform 1 0 7584 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1164_
timestamp 1678805552
transform 1 0 7680 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1165_
timestamp 1678805552
transform 1 0 10560 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1166_
timestamp 1678805552
transform 1 0 10560 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1167_
timestamp 1678805552
transform 1 0 13824 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1168_
timestamp 1678805552
transform 1 0 13632 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1169_
timestamp 1678805552
transform 1 0 9120 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1170_
timestamp 1678805552
transform 1 0 7488 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1171_
timestamp 1678805552
transform 1 0 5664 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1172_
timestamp 1678805552
transform 1 0 4224 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1173_
timestamp 1678805552
transform 1 0 3552 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1174_
timestamp 1678805552
transform -1 0 7584 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1175_
timestamp 1678805552
transform 1 0 5184 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1176_
timestamp 1678805552
transform 1 0 1344 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1177_
timestamp 1678805552
transform 1 0 1152 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1178_
timestamp 1678805552
transform 1 0 2688 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1179_
timestamp 1678805552
transform 1 0 1152 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1180_
timestamp 1678805552
transform 1 0 1152 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1181_
timestamp 1678805552
transform -1 0 12000 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1182_
timestamp 1678805552
transform -1 0 15264 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1183_
timestamp 1678805552
transform -1 0 16896 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1184_
timestamp 1678805552
transform -1 0 8736 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1185_
timestamp 1678805552
transform 1 0 16320 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1186_
timestamp 1678805552
transform 1 0 14304 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1187_
timestamp 1678805552
transform 1 0 9120 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1188_
timestamp 1678805552
transform 1 0 7008 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1189_
timestamp 1678805552
transform 1 0 13248 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1190_
timestamp 1678805552
transform 1 0 11232 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1191_
timestamp 1678805552
transform 1 0 16416 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1192_
timestamp 1678805552
transform 1 0 15840 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1193_
timestamp 1678805552
transform 1 0 18624 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1194_
timestamp 1678805552
transform 1 0 17184 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1195_
timestamp 1678805552
transform 1 0 8352 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1196_
timestamp 1678805552
transform 1 0 6912 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1197_
timestamp 1678805552
transform 1 0 13344 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1198_
timestamp 1678805552
transform 1 0 10944 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1199_
timestamp 1678805552
transform 1 0 18432 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1200_
timestamp 1678805552
transform 1 0 16512 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1201_
timestamp 1678805552
transform 1 0 18624 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1202_
timestamp 1678805552
transform 1 0 16416 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1203_
timestamp 1678805552
transform 1 0 9024 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1204_
timestamp 1678805552
transform 1 0 6912 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1205_
timestamp 1678805552
transform 1 0 12768 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1206_
timestamp 1678805552
transform 1 0 10752 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1207_
timestamp 1678805552
transform 1 0 18336 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1208_
timestamp 1678805552
transform 1 0 16416 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1209_
timestamp 1678805552
transform 1 0 18720 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1210_
timestamp 1678805552
transform 1 0 17472 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1211_
timestamp 1678805552
transform 1 0 8640 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1212_
timestamp 1678805552
transform 1 0 6912 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1213_
timestamp 1678805552
transform 1 0 13056 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1214_
timestamp 1678805552
transform 1 0 10944 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1215_
timestamp 1678805552
transform 1 0 18336 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1216_
timestamp 1678805552
transform 1 0 16992 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1217_
timestamp 1678805552
transform 1 0 2112 0 1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1218_
timestamp 1678805552
transform 1 0 1152 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1219_
timestamp 1678805552
transform 1 0 1152 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1220_
timestamp 1678805552
transform 1 0 1152 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1221_
timestamp 1678805552
transform 1 0 17856 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1222_
timestamp 1678805552
transform -1 0 11040 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1223_
timestamp 1678805552
transform -1 0 11232 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1224_
timestamp 1678805552
transform 1 0 5184 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1225_
timestamp 1678805552
transform 1 0 6336 0 -1 44604
box -50 -56 1692 834
use sg13g2_dlhq_1  _1226_
timestamp 1678805552
transform 1 0 5184 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1227_
timestamp 1678805552
transform 1 0 5184 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1228_
timestamp 1678805552
transform 1 0 4992 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1229_
timestamp 1678805552
transform 1 0 15840 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1230_
timestamp 1678805552
transform 1 0 14112 0 -1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1231_
timestamp 1678805552
transform 1 0 12576 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1232_
timestamp 1678805552
transform 1 0 10752 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1233_
timestamp 1678805552
transform 1 0 17856 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1234_
timestamp 1678805552
transform 1 0 16512 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1235_
timestamp 1678805552
transform 1 0 18720 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1236_
timestamp 1678805552
transform 1 0 16896 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1237_
timestamp 1678805552
transform 1 0 18144 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1238_
timestamp 1678805552
transform 1 0 16224 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1239_
timestamp 1678805552
transform 1 0 9600 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1240_
timestamp 1678805552
transform 1 0 7680 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1241_
timestamp 1678805552
transform -1 0 17184 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1242_
timestamp 1678805552
transform -1 0 15552 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1243_
timestamp 1678805552
transform 1 0 18240 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1244_
timestamp 1678805552
transform 1 0 14304 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1245_
timestamp 1678805552
transform 1 0 15648 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1246_
timestamp 1678805552
transform 1 0 13920 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1247_
timestamp 1678805552
transform 1 0 13344 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1248_
timestamp 1678805552
transform 1 0 10464 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1249_
timestamp 1678805552
transform 1 0 18720 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1250_
timestamp 1678805552
transform 1 0 17184 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1251_
timestamp 1678805552
transform 1 0 18432 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1252_
timestamp 1678805552
transform 1 0 16704 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1253_
timestamp 1678805552
transform 1 0 18432 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1254_
timestamp 1678805552
transform 1 0 17376 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1255_
timestamp 1678805552
transform 1 0 9120 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1256_
timestamp 1678805552
transform 1 0 7488 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1257_
timestamp 1678805552
transform 1 0 14976 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1258_
timestamp 1678805552
transform 1 0 12864 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1259_
timestamp 1678805552
transform 1 0 18624 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1260_
timestamp 1678805552
transform 1 0 16608 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1261_
timestamp 1678805552
transform 1 0 15552 0 -1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1262_
timestamp 1678805552
transform 1 0 14976 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1263_
timestamp 1678805552
transform 1 0 12288 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1264_
timestamp 1678805552
transform 1 0 11328 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1265_
timestamp 1678805552
transform 1 0 15936 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1266_
timestamp 1678805552
transform 1 0 16608 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1267_
timestamp 1678805552
transform 1 0 18528 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1268_
timestamp 1678805552
transform 1 0 16608 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1269_
timestamp 1678805552
transform 1 0 18432 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1270_
timestamp 1678805552
transform 1 0 16800 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1271_
timestamp 1678805552
transform 1 0 9792 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1272_
timestamp 1678805552
transform 1 0 8160 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1273_
timestamp 1678805552
transform 1 0 15168 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1274_
timestamp 1678805552
transform 1 0 13536 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1275_
timestamp 1678805552
transform 1 0 16704 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1276_
timestamp 1678805552
transform 1 0 15936 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1277_
timestamp 1678805552
transform 1 0 15840 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1278_
timestamp 1678805552
transform 1 0 14208 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1279_
timestamp 1678805552
transform 1 0 12576 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1280_
timestamp 1678805552
transform 1 0 10656 0 -1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1281_
timestamp 1678805552
transform 1 0 18720 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1282_
timestamp 1678805552
transform 1 0 16800 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1283_
timestamp 1678805552
transform 1 0 17088 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1284_
timestamp 1678805552
transform 1 0 16704 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1285_
timestamp 1678805552
transform 1 0 18720 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1286_
timestamp 1678805552
transform 1 0 16704 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1287_
timestamp 1678805552
transform 1 0 9312 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1288_
timestamp 1678805552
transform 1 0 7488 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1289_
timestamp 1678805552
transform 1 0 15072 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1290_
timestamp 1678805552
transform 1 0 13056 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1291_
timestamp 1678805552
transform 1 0 16416 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1292_
timestamp 1678805552
transform 1 0 15456 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1293_
timestamp 1678805552
transform 1 0 7776 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1294_
timestamp 1678805552
transform 1 0 7008 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1295_
timestamp 1678805552
transform 1 0 9888 0 1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1296_
timestamp 1678805552
transform 1 0 9216 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1297_
timestamp 1678805552
transform 1 0 4608 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1298_
timestamp 1678805552
transform 1 0 4416 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1299_
timestamp 1678805552
transform 1 0 4224 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1300_
timestamp 1678805552
transform 1 0 4128 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1301_
timestamp 1678805552
transform 1 0 10368 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1302_
timestamp 1678805552
transform 1 0 9984 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1303_
timestamp 1678805552
transform 1 0 14592 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1304_
timestamp 1678805552
transform 1 0 15648 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1305_
timestamp 1678805552
transform 1 0 4608 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1306_
timestamp 1678805552
transform 1 0 6720 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1307_
timestamp 1678805552
transform 1 0 1152 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1308_
timestamp 1678805552
transform 1 0 1152 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1309_
timestamp 1678805552
transform 1 0 11424 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1310_
timestamp 1678805552
transform 1 0 13056 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1311_
timestamp 1678805552
transform -1 0 17856 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1312_
timestamp 1678805552
transform -1 0 16704 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1313_
timestamp 1678805552
transform 1 0 5568 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1314_
timestamp 1678805552
transform 1 0 4032 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1315_
timestamp 1678805552
transform 1 0 4320 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1316_
timestamp 1678805552
transform 1 0 5280 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1317_
timestamp 1678805552
transform 1 0 8640 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1318_
timestamp 1678805552
transform 1 0 10464 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1319_
timestamp 1678805552
transform 1 0 16224 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1320_
timestamp 1678805552
transform 1 0 14496 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1321_
timestamp 1678805552
transform 1 0 8448 0 -1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1322_
timestamp 1678805552
transform 1 0 7200 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1323_
timestamp 1678805552
transform 1 0 10464 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1324_
timestamp 1678805552
transform 1 0 8736 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1325_
timestamp 1678805552
transform 1 0 12384 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1326_
timestamp 1678805552
transform 1 0 10560 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1327_
timestamp 1678805552
transform 1 0 14688 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1328_
timestamp 1678805552
transform 1 0 12960 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1329_
timestamp 1678805552
transform 1 0 5568 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1330_
timestamp 1678805552
transform 1 0 4128 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1331_
timestamp 1678805552
transform 1 0 3456 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1332_
timestamp 1678805552
transform 1 0 1152 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1333_
timestamp 1678805552
transform 1 0 12576 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1334_
timestamp 1678805552
transform 1 0 11232 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1335_
timestamp 1678805552
transform 1 0 15264 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1336_
timestamp 1678805552
transform 1 0 13632 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1337_
timestamp 1678805552
transform 1 0 5760 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1338_
timestamp 1678805552
transform 1 0 2784 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1339_
timestamp 1678805552
transform 1 0 3648 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1340_
timestamp 1678805552
transform 1 0 1152 0 1 11340
box -50 -56 1692 834
use sg13g2_dlhq_1  _1341_
timestamp 1678805552
transform -1 0 13440 0 -1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1342_
timestamp 1678805552
transform 1 0 8160 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1343_
timestamp 1678805552
transform -1 0 17280 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1344_
timestamp 1678805552
transform 1 0 14016 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1345_
timestamp 1678805552
transform 1 0 4992 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1346_
timestamp 1678805552
transform 1 0 3072 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1347_
timestamp 1678805552
transform 1 0 5280 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1348_
timestamp 1678805552
transform 1 0 3648 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1349_
timestamp 1678805552
transform 1 0 10176 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1350_
timestamp 1678805552
transform 1 0 9216 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1351_
timestamp 1678805552
transform 1 0 14208 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1352_
timestamp 1678805552
transform 1 0 12480 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1353_
timestamp 1678805552
transform 1 0 7584 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1354_
timestamp 1678805552
transform 1 0 5952 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1355_
timestamp 1678805552
transform 1 0 5952 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1356_
timestamp 1678805552
transform 1 0 4128 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1357_
timestamp 1678805552
transform 1 0 12192 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1358_
timestamp 1678805552
transform 1 0 10752 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1359_
timestamp 1678805552
transform 1 0 14784 0 -1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1360_
timestamp 1678805552
transform 1 0 12768 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1361_
timestamp 1678805552
transform 1 0 3456 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1362_
timestamp 1678805552
transform -1 0 13632 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1363_
timestamp 1678805552
transform 1 0 1440 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1364_
timestamp 1678805552
transform 1 0 1152 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1365_
timestamp 1678805552
transform 1 0 7104 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1366_
timestamp 1678805552
transform 1 0 5184 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1367_
timestamp 1678805552
transform 1 0 11424 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1368_
timestamp 1678805552
transform 1 0 9792 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1369_
timestamp 1678805552
transform 1 0 2304 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1370_
timestamp 1678805552
transform 1 0 1152 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1371_
timestamp 1678805552
transform 1 0 1920 0 1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1372_
timestamp 1678805552
transform 1 0 1152 0 -1 14364
box -50 -56 1692 834
use sg13g2_dlhq_1  _1373_
timestamp 1678805552
transform 1 0 8736 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1374_
timestamp 1678805552
transform 1 0 5184 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1375_
timestamp 1678805552
transform 1 0 14688 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1376_
timestamp 1678805552
transform 1 0 13056 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1377_
timestamp 1678805552
transform 1 0 2208 0 -1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1378_
timestamp 1678805552
transform 1 0 1248 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1379_
timestamp 1678805552
transform 1 0 1152 0 1 9828
box -50 -56 1692 834
use sg13g2_dlhq_1  _1380_
timestamp 1678805552
transform 1 0 1152 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1381_
timestamp 1678805552
transform 1 0 5088 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1382_
timestamp 1678805552
transform 1 0 5280 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1383_
timestamp 1678805552
transform 1 0 11808 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1384_
timestamp 1678805552
transform 1 0 9984 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1385_
timestamp 1678805552
transform 1 0 2784 0 -1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1386_
timestamp 1678805552
transform 1 0 1152 0 -1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1387_
timestamp 1678805552
transform 1 0 2688 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1388_
timestamp 1678805552
transform 1 0 1152 0 -1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1389_
timestamp 1678805552
transform 1 0 6912 0 1 3780
box -50 -56 1692 834
use sg13g2_dlhq_1  _1390_
timestamp 1678805552
transform 1 0 7104 0 1 756
box -50 -56 1692 834
use sg13g2_dlhq_1  _1391_
timestamp 1678805552
transform 1 0 16800 0 1 8316
box -50 -56 1692 834
use sg13g2_dlhq_1  _1392_
timestamp 1678805552
transform 1 0 18528 0 1 6804
box -50 -56 1692 834
use sg13g2_dlhq_1  _1393_
timestamp 1678805552
transform 1 0 7392 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1394_
timestamp 1678805552
transform 1 0 8736 0 -1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1395_
timestamp 1678805552
transform 1 0 9408 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1396_
timestamp 1678805552
transform 1 0 11040 0 1 12852
box -50 -56 1692 834
use sg13g2_dlhq_1  _1397_
timestamp 1678805552
transform 1 0 18624 0 1 5292
box -50 -56 1692 834
use sg13g2_dlhq_1  _1398_
timestamp 1678805552
transform 1 0 18720 0 1 2268
box -50 -56 1692 834
use sg13g2_dlhq_1  _1399_
timestamp 1678805552
transform 1 0 15360 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1400_
timestamp 1678805552
transform 1 0 14976 0 -1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1401_
timestamp 1678805552
transform 1 0 14784 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1402_
timestamp 1678805552
transform 1 0 4800 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1403_
timestamp 1678805552
transform 1 0 4224 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1404_
timestamp 1678805552
transform 1 0 2592 0 1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1405_
timestamp 1678805552
transform 1 0 11520 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1406_
timestamp 1678805552
transform 1 0 11232 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1407_
timestamp 1678805552
transform 1 0 11424 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1408_
timestamp 1678805552
transform 1 0 18048 0 -1 15876
box -50 -56 1692 834
use sg13g2_dlhq_1  _1409_
timestamp 1678805552
transform 1 0 17856 0 1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1410_
timestamp 1678805552
transform 1 0 17280 0 -1 17388
box -50 -56 1692 834
use sg13g2_dlhq_1  _1411_
timestamp 1678805552
transform 1 0 9408 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1412_
timestamp 1678805552
transform 1 0 10752 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1413_
timestamp 1678805552
transform 1 0 4704 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1414_
timestamp 1678805552
transform 1 0 3648 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1415_
timestamp 1678805552
transform 1 0 5280 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1416_
timestamp 1678805552
transform 1 0 3936 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1417_
timestamp 1678805552
transform 1 0 6240 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1418_
timestamp 1678805552
transform 1 0 7776 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1419_
timestamp 1678805552
transform 1 0 6048 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1420_
timestamp 1678805552
transform -1 0 10272 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1421_
timestamp 1678805552
transform 1 0 1152 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1422_
timestamp 1678805552
transform 1 0 1632 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1423_
timestamp 1678805552
transform -1 0 5856 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1424_
timestamp 1678805552
transform -1 0 4416 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1425_
timestamp 1678805552
transform 1 0 2784 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1426_
timestamp 1678805552
transform 1 0 1152 0 1 18900
box -50 -56 1692 834
use sg13g2_dlhq_1  _1427_
timestamp 1678805552
transform 1 0 12672 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1428_
timestamp 1678805552
transform 1 0 10752 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1429_
timestamp 1678805552
transform 1 0 7488 0 1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1430_
timestamp 1678805552
transform 1 0 5952 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1431_
timestamp 1678805552
transform 1 0 8928 0 1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1432_
timestamp 1678805552
transform 1 0 7392 0 -1 27972
box -50 -56 1692 834
use sg13g2_dlhq_1  _1433_
timestamp 1678805552
transform 1 0 12192 0 -1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1434_
timestamp 1678805552
transform 1 0 10464 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1435_
timestamp 1678805552
transform 1 0 11232 0 1 41580
box -50 -56 1692 834
use sg13g2_dlhq_1  _1436_
timestamp 1678805552
transform 1 0 11424 0 1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1437_
timestamp 1678805552
transform 1 0 11232 0 -1 40068
box -50 -56 1692 834
use sg13g2_dlhq_1  _1438_
timestamp 1678805552
transform 1 0 4416 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1439_
timestamp 1678805552
transform 1 0 3936 0 1 35532
box -50 -56 1692 834
use sg13g2_dlhq_1  _1440_
timestamp 1678805552
transform 1 0 2784 0 -1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1441_
timestamp 1678805552
transform 1 0 4224 0 -1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1442_
timestamp 1678805552
transform 1 0 4128 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1443_
timestamp 1678805552
transform 1 0 3936 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1444_
timestamp 1678805552
transform 1 0 14592 0 -1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1445_
timestamp 1678805552
transform -1 0 16608 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1446_
timestamp 1678805552
transform -1 0 16704 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1447_
timestamp 1678805552
transform 1 0 8352 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1448_
timestamp 1678805552
transform 1 0 6432 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1449_
timestamp 1678805552
transform 1 0 1152 0 1 24948
box -50 -56 1692 834
use sg13g2_dlhq_1  _1450_
timestamp 1678805552
transform 1 0 3744 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1451_
timestamp 1678805552
transform 1 0 1152 0 -1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1452_
timestamp 1678805552
transform -1 0 5856 0 -1 29484
box -50 -56 1692 834
use sg13g2_dlhq_1  _1453_
timestamp 1678805552
transform 1 0 5472 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1454_
timestamp 1678805552
transform 1 0 3840 0 -1 38556
box -50 -56 1692 834
use sg13g2_dlhq_1  _1455_
timestamp 1678805552
transform 1 0 1152 0 1 21924
box -50 -56 1692 834
use sg13g2_dlhq_1  _1456_
timestamp 1678805552
transform 1 0 2976 0 -1 26460
box -50 -56 1692 834
use sg13g2_dlhq_1  _1457_
timestamp 1678805552
transform 1 0 1152 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1458_
timestamp 1678805552
transform 1 0 1728 0 1 34020
box -50 -56 1692 834
use sg13g2_dlhq_1  _1459_
timestamp 1678805552
transform 1 0 1536 0 1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1460_
timestamp 1678805552
transform 1 0 1152 0 -1 30996
box -50 -56 1692 834
use sg13g2_dlhq_1  _1461_
timestamp 1678805552
transform 1 0 1152 0 1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1462_
timestamp 1678805552
transform 1 0 1152 0 -1 20412
box -50 -56 1692 834
use sg13g2_dlhq_1  _1463_
timestamp 1678805552
transform 1 0 11424 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1464_
timestamp 1678805552
transform 1 0 13056 0 -1 43092
box -50 -56 1692 834
use sg13g2_dlhq_1  _1465_
timestamp 1678805552
transform 1 0 6624 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1466_
timestamp 1678805552
transform 1 0 8256 0 1 37044
box -50 -56 1692 834
use sg13g2_dlhq_1  _1467_
timestamp 1678805552
transform 1 0 9312 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1468_
timestamp 1678805552
transform 1 0 10944 0 1 32508
box -50 -56 1692 834
use sg13g2_dlhq_1  _1469_
timestamp 1678805552
transform 1 0 10848 0 1 23436
box -50 -56 1692 834
use sg13g2_dlhq_1  _1470_
timestamp 1678805552
transform 1 0 12864 0 -1 23436
box -50 -56 1692 834
use sg13g2_tiehi  _1471_
timestamp 1680000651
transform 1 0 19680 0 -1 50652
box -48 -56 432 834
use sg13g2_tielo  _1472_
timestamp 1680000637
transform 1 0 19872 0 1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1473_
timestamp 1676381911
transform 1 0 19296 0 -1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1474_
timestamp 1676381911
transform 1 0 19296 0 -1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1475_
timestamp 1676381911
transform 1 0 19680 0 -1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1476_
timestamp 1676381911
transform 1 0 19296 0 1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1477_
timestamp 1676381911
transform 1 0 19680 0 1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1478_
timestamp 1676381911
transform 1 0 19872 0 -1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1479_
timestamp 1676381911
transform 1 0 19584 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1480_
timestamp 1676381911
transform 1 0 19680 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1481_
timestamp 1676381911
transform 1 0 19296 0 1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1482_
timestamp 1676381911
transform 1 0 19968 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1483_
timestamp 1676381911
transform 1 0 17568 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1484_
timestamp 1676381911
transform 1 0 19680 0 1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1485_
timestamp 1676381911
transform 1 0 19680 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1486_
timestamp 1676381911
transform 1 0 19680 0 1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1487_
timestamp 1676381911
transform 1 0 19968 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1488_
timestamp 1676381911
transform 1 0 19680 0 -1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1489_
timestamp 1676381911
transform 1 0 19680 0 1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1490_
timestamp 1676381911
transform 1 0 19584 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1491_
timestamp 1676381911
transform 1 0 19968 0 -1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1492_
timestamp 1676381911
transform 1 0 19680 0 1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1493_
timestamp 1676381911
transform 1 0 17568 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1494_
timestamp 1676381911
transform 1 0 19776 0 -1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1495_
timestamp 1676381911
transform 1 0 17184 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1496_
timestamp 1676381911
transform 1 0 19776 0 1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1497_
timestamp 1676381911
transform 1 0 17280 0 -1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1498_
timestamp 1676381911
transform 1 0 16896 0 -1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1499_
timestamp 1676381911
transform 1 0 19680 0 -1 64260
box -48 -56 432 834
use sg13g2_buf_1  _1500_
timestamp 1676381911
transform 1 0 16512 0 1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1501_
timestamp 1676381911
transform 1 0 17280 0 1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1502_
timestamp 1676381911
transform 1 0 16896 0 1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1503_
timestamp 1676381911
transform 1 0 19776 0 1 64260
box -48 -56 432 834
use sg13g2_buf_1  _1504_
timestamp 1676381911
transform 1 0 14784 0 1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1505_
timestamp 1676381911
transform 1 0 15840 0 1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1506_
timestamp 1676381911
transform -1 0 20352 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1507_
timestamp 1676381911
transform -1 0 19872 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1508_
timestamp 1676381911
transform -1 0 17568 0 1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1509_
timestamp 1676381911
transform -1 0 17952 0 1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1510_
timestamp 1676381911
transform -1 0 18240 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1511_
timestamp 1676381911
transform 1 0 16416 0 -1 65772
box -48 -56 432 834
use sg13g2_buf_1  _1512_
timestamp 1676381911
transform 1 0 16608 0 -1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1513_
timestamp 1676381911
transform -1 0 17856 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1514_
timestamp 1676381911
transform -1 0 18240 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1515_
timestamp 1676381911
transform 1 0 17088 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1516_
timestamp 1676381911
transform -1 0 19200 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1517_
timestamp 1676381911
transform -1 0 19584 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1518_
timestamp 1676381911
transform -1 0 20352 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1519_
timestamp 1676381911
transform -1 0 19968 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1520_
timestamp 1676381911
transform -1 0 20256 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1521_
timestamp 1676381911
transform -1 0 20352 0 -1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1522_
timestamp 1676381911
transform 1 0 16320 0 1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1523_
timestamp 1676381911
transform 1 0 18240 0 1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1524_
timestamp 1676381911
transform 1 0 12864 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1525_
timestamp 1676381911
transform 1 0 12096 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1526_
timestamp 1676381911
transform 1 0 1152 0 -1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1527_
timestamp 1676381911
transform -1 0 2496 0 1 74844
box -48 -56 432 834
use sg13g2_buf_1  _1528_
timestamp 1676381911
transform 1 0 1248 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1529_
timestamp 1676381911
transform -1 0 8352 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1530_
timestamp 1676381911
transform 1 0 1632 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1531_
timestamp 1676381911
transform 1 0 1248 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1532_
timestamp 1676381911
transform -1 0 4896 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1533_
timestamp 1676381911
transform 1 0 2784 0 -1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1534_
timestamp 1676381911
transform -1 0 7488 0 -1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1535_
timestamp 1676381911
transform 1 0 2784 0 -1 79380
box -48 -56 432 834
use sg13g2_buf_1  _1536_
timestamp 1676381911
transform -1 0 4896 0 1 76356
box -48 -56 432 834
use sg13g2_buf_1  _1537_
timestamp 1676381911
transform 1 0 1632 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1538_
timestamp 1676381911
transform 1 0 1344 0 1 74844
box -48 -56 432 834
use sg13g2_buf_1  _1539_
timestamp 1676381911
transform 1 0 3360 0 -1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1540_
timestamp 1676381911
transform -1 0 5664 0 1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1541_
timestamp 1676381911
transform -1 0 5280 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1542_
timestamp 1676381911
transform 1 0 4128 0 -1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1543_
timestamp 1676381911
transform 1 0 1248 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1544_
timestamp 1676381911
transform 1 0 2976 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1545_
timestamp 1676381911
transform 1 0 3744 0 -1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1546_
timestamp 1676381911
transform -1 0 11904 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1547_
timestamp 1676381911
transform 1 0 4128 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1548_
timestamp 1676381911
transform 1 0 3936 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1549_
timestamp 1676381911
transform -1 0 7104 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1550_
timestamp 1676381911
transform 1 0 1824 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1551_
timestamp 1676381911
transform -1 0 7488 0 -1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1552_
timestamp 1676381911
transform -1 0 9888 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1553_
timestamp 1676381911
transform 1 0 3168 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1554_
timestamp 1676381911
transform -1 0 18816 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1555_
timestamp 1676381911
transform 1 0 7008 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1556_
timestamp 1676381911
transform 1 0 5376 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1557_
timestamp 1676381911
transform -1 0 12864 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1558_
timestamp 1676381911
transform 1 0 5760 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1559_
timestamp 1676381911
transform 1 0 6144 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1560_
timestamp 1676381911
transform -1 0 9312 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1561_
timestamp 1676381911
transform 1 0 7584 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1562_
timestamp 1676381911
transform -1 0 16032 0 1 80892
box -48 -56 432 834
use sg13g2_buf_1  _1563_
timestamp 1676381911
transform -1 0 12000 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1564_
timestamp 1676381911
transform -1 0 13440 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1565_
timestamp 1676381911
transform -1 0 1920 0 -1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1566_
timestamp 1676381911
transform -1 0 15264 0 -1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1567_
timestamp 1676381911
transform -1 0 1536 0 1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1568_
timestamp 1676381911
transform -1 0 1920 0 1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1569_
timestamp 1676381911
transform -1 0 1824 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1570_
timestamp 1676381911
transform -1 0 2976 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1571_
timestamp 1676381911
transform -1 0 3168 0 1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1572_
timestamp 1676381911
transform -1 0 1824 0 -1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1573_
timestamp 1676381911
transform -1 0 3552 0 1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1574_
timestamp 1676381911
transform -1 0 2592 0 1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1575_
timestamp 1676381911
transform -1 0 1824 0 1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1576_
timestamp 1676381911
transform -1 0 2208 0 1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1577_
timestamp 1676381911
transform -1 0 1824 0 -1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1578_
timestamp 1676381911
transform -1 0 5280 0 -1 59724
box -48 -56 432 834
use sg13g2_buf_1  _1579_
timestamp 1676381911
transform -1 0 2208 0 1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1580_
timestamp 1676381911
transform -1 0 1824 0 1 47628
box -48 -56 432 834
use sg13g2_buf_1  _1581_
timestamp 1676381911
transform -1 0 2208 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1582_
timestamp 1676381911
transform -1 0 2208 0 -1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1583_
timestamp 1676381911
transform -1 0 12768 0 -1 74844
box -48 -56 432 834
use sg13g2_buf_1  _1584_
timestamp 1676381911
transform -1 0 13728 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1585_
timestamp 1676381911
transform -1 0 13728 0 1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1586_
timestamp 1676381911
transform -1 0 15360 0 -1 77868
box -48 -56 432 834
use sg13g2_buf_1  _1587_
timestamp 1676381911
transform -1 0 13056 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1588_
timestamp 1676381911
transform -1 0 2208 0 1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1589_
timestamp 1676381911
transform -1 0 1536 0 -1 56700
box -48 -56 432 834
use sg13g2_buf_1  _1590_
timestamp 1676381911
transform -1 0 1824 0 -1 61236
box -48 -56 432 834
use sg13g2_buf_1  _1591_
timestamp 1676381911
transform -1 0 13344 0 -1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1592_
timestamp 1676381911
transform -1 0 9984 0 1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1593_
timestamp 1676381911
transform -1 0 1632 0 -1 58212
box -48 -56 432 834
use sg13g2_buf_1  _1594_
timestamp 1676381911
transform -1 0 2592 0 1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1595_
timestamp 1676381911
transform -1 0 1824 0 -1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1596_
timestamp 1676381911
transform -1 0 3168 0 1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1597_
timestamp 1676381911
transform -1 0 2208 0 -1 49140
box -48 -56 432 834
use sg13g2_buf_1  _1598_
timestamp 1676381911
transform -1 0 8736 0 -1 52164
box -48 -56 432 834
use sg13g2_buf_1  _1599_
timestamp 1676381911
transform -1 0 1632 0 -1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1600_
timestamp 1676381911
transform -1 0 2592 0 -1 50652
box -48 -56 432 834
use sg13g2_buf_1  _1601_
timestamp 1676381911
transform -1 0 2016 0 -1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1602_
timestamp 1676381911
transform -1 0 2208 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1603_
timestamp 1676381911
transform -1 0 1824 0 -1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1604_
timestamp 1676381911
transform -1 0 2208 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1605_
timestamp 1676381911
transform -1 0 1824 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1606_
timestamp 1676381911
transform -1 0 3552 0 1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1607_
timestamp 1676381911
transform -1 0 11520 0 1 53676
box -48 -56 432 834
use sg13g2_buf_1  _1608_
timestamp 1676381911
transform -1 0 3168 0 1 55188
box -48 -56 432 834
use sg13g2_buf_1  _1609_
timestamp 1676381911
transform -1 0 2592 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1610_
timestamp 1676381911
transform -1 0 1824 0 1 62748
box -48 -56 432 834
use sg13g2_buf_1  _1611_
timestamp 1676381911
transform 1 0 16032 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1612_
timestamp 1676381911
transform 1 0 19680 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1613_
timestamp 1676381911
transform 1 0 17472 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1614_
timestamp 1676381911
transform 1 0 18720 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1615_
timestamp 1676381911
transform 1 0 18048 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1616_
timestamp 1676381911
transform 1 0 19488 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1617_
timestamp 1676381911
transform 1 0 17664 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1618_
timestamp 1676381911
transform 1 0 19296 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1619_
timestamp 1676381911
transform 1 0 19296 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1620_
timestamp 1676381911
transform 1 0 19680 0 -1 38556
box -48 -56 432 834
use sg13g2_buf_1  _1621_
timestamp 1676381911
transform 1 0 14880 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1622_
timestamp 1676381911
transform 1 0 17952 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1623_
timestamp 1676381911
transform 1 0 19296 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1624_
timestamp 1676381911
transform 1 0 18720 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1625_
timestamp 1676381911
transform 1 0 18048 0 1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1626_
timestamp 1676381911
transform 1 0 17664 0 -1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1627_
timestamp 1676381911
transform 1 0 17088 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1628_
timestamp 1676381911
transform 1 0 19104 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1629_
timestamp 1676381911
transform 1 0 17472 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1630_
timestamp 1676381911
transform 1 0 18912 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1631_
timestamp 1676381911
transform 1 0 18048 0 -1 44604
box -48 -56 432 834
use sg13g2_buf_1  _1632_
timestamp 1676381911
transform 1 0 19680 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1633_
timestamp 1676381911
transform 1 0 17856 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1634_
timestamp 1676381911
transform 1 0 18336 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1635_
timestamp 1676381911
transform 1 0 17568 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1636_
timestamp 1676381911
transform 1 0 19968 0 -1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1637_
timestamp 1676381911
transform 1 0 14880 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1638_
timestamp 1676381911
transform 1 0 16512 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1639_
timestamp 1676381911
transform 1 0 19872 0 1 41580
box -48 -56 432 834
use sg13g2_buf_1  _1640_
timestamp 1676381911
transform 1 0 19296 0 -1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1641_
timestamp 1676381911
transform 1 0 18528 0 1 43092
box -48 -56 432 834
use sg13g2_buf_1  _1642_
timestamp 1676381911
transform 1 0 19680 0 -1 46116
box -48 -56 432 834
use sg13g2_buf_1  _1643_
timestamp 1676381911
transform -1 0 14304 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1644_
timestamp 1676381911
transform 1 0 7680 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1645_
timestamp 1676381911
transform 1 0 8832 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1646_
timestamp 1676381911
transform -1 0 14688 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1647_
timestamp 1676381911
transform 1 0 4608 0 1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1648_
timestamp 1676381911
transform 1 0 5280 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1649_
timestamp 1676381911
transform 1 0 3744 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1650_
timestamp 1676381911
transform -1 0 10944 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1651_
timestamp 1676381911
transform 1 0 8832 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1652_
timestamp 1676381911
transform 1 0 8064 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1653_
timestamp 1676381911
transform 1 0 9216 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1654_
timestamp 1676381911
transform -1 0 11616 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1655_
timestamp 1676381911
transform 1 0 4896 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1656_
timestamp 1676381911
transform 1 0 4800 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1657_
timestamp 1676381911
transform 1 0 8736 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1658_
timestamp 1676381911
transform 1 0 9600 0 1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1659_
timestamp 1676381911
transform 1 0 10464 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1660_
timestamp 1676381911
transform 1 0 9024 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1661_
timestamp 1676381911
transform 1 0 10848 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1662_
timestamp 1676381911
transform 1 0 9408 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1663_
timestamp 1676381911
transform -1 0 13536 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1664_
timestamp 1676381911
transform -1 0 13920 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1665_
timestamp 1676381911
transform -1 0 13632 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1666_
timestamp 1676381911
transform 1 0 12192 0 1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1667_
timestamp 1676381911
transform -1 0 13728 0 1 82404
box -48 -56 432 834
use sg13g2_buf_1  _1668_
timestamp 1676381911
transform -1 0 15936 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1669_
timestamp 1676381911
transform -1 0 16320 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1670_
timestamp 1676381911
transform -1 0 18432 0 -1 83916
box -48 -56 432 834
use sg13g2_buf_1  _1671_
timestamp 1676381911
transform 1 0 13632 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1672_
timestamp 1676381911
transform -1 0 17664 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1673_
timestamp 1676381911
transform -1 0 17088 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1674_
timestamp 1676381911
transform -1 0 20352 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1675_
timestamp 1676381911
transform -1 0 18336 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1676_
timestamp 1676381911
transform -1 0 16704 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1677_
timestamp 1676381911
transform -1 0 17280 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1678_
timestamp 1676381911
transform -1 0 17472 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1679_
timestamp 1676381911
transform -1 0 4800 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1680_
timestamp 1676381911
transform -1 0 11712 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1681_
timestamp 1676381911
transform -1 0 1728 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1682_
timestamp 1676381911
transform -1 0 8160 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1683_
timestamp 1676381911
transform -1 0 7776 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1684_
timestamp 1676381911
transform -1 0 5472 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1685_
timestamp 1676381911
transform -1 0 3936 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1686_
timestamp 1676381911
transform -1 0 11328 0 1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1687_
timestamp 1676381911
transform -1 0 3552 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1688_
timestamp 1676381911
transform -1 0 2592 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1689_
timestamp 1676381911
transform -1 0 4896 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1690_
timestamp 1676381911
transform -1 0 1824 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1691_
timestamp 1676381911
transform -1 0 5280 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1692_
timestamp 1676381911
transform -1 0 1536 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1693_
timestamp 1676381911
transform -1 0 7584 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1694_
timestamp 1676381911
transform -1 0 3168 0 1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1695_
timestamp 1676381911
transform -1 0 9504 0 1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1696_
timestamp 1676381911
transform -1 0 5280 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1697_
timestamp 1676381911
transform -1 0 4704 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1698_
timestamp 1676381911
transform -1 0 11232 0 -1 6804
box -48 -56 432 834
use sg13g2_buf_1  _1699_
timestamp 1676381911
transform -1 0 13824 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1700_
timestamp 1676381911
transform -1 0 11424 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1701_
timestamp 1676381911
transform -1 0 10752 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1702_
timestamp 1676381911
transform -1 0 18240 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1703_
timestamp 1676381911
transform -1 0 12480 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1704_
timestamp 1676381911
transform -1 0 3936 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1705_
timestamp 1676381911
transform -1 0 2112 0 1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1706_
timestamp 1676381911
transform -1 0 17376 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1707_
timestamp 1676381911
transform -1 0 14304 0 -1 12852
box -48 -56 432 834
use sg13g2_buf_1  _1708_
timestamp 1676381911
transform -1 0 2208 0 -1 21924
box -48 -56 432 834
use sg13g2_buf_1  _1709_
timestamp 1676381911
transform -1 0 3168 0 -1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1710_
timestamp 1676381911
transform -1 0 17760 0 1 15876
box -48 -56 432 834
use sg13g2_buf_1  _1711_
timestamp 1676381911
transform -1 0 1824 0 1 14364
box -48 -56 432 834
use sg13g2_buf_1  _1712_
timestamp 1676381911
transform -1 0 3264 0 1 756
box -48 -56 432 834
use sg13g2_buf_1  _1713_
timestamp 1676381911
transform -1 0 1824 0 -1 3780
box -48 -56 432 834
use sg13g2_buf_1  _1714_
timestamp 1676381911
transform -1 0 3168 0 -1 2268
box -48 -56 432 834
use sg13g2_buf_1  _1715_
timestamp 1676381911
transform -1 0 2112 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1716_
timestamp 1676381911
transform -1 0 1824 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1717_
timestamp 1676381911
transform -1 0 3552 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1718_
timestamp 1676381911
transform -1 0 2208 0 1 5292
box -48 -56 432 834
use sg13g2_buf_1  _1719_
timestamp 1676381911
transform -1 0 3168 0 -1 8316
box -48 -56 432 834
use sg13g2_buf_1  _1720_
timestamp 1676381911
transform -1 0 1728 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1721_
timestamp 1676381911
transform -1 0 1824 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1722_
timestamp 1676381911
transform -1 0 2496 0 -1 9828
box -48 -56 432 834
use sg13g2_buf_1  _1723_
timestamp 1676381911
transform -1 0 14784 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1724_
timestamp 1676381911
transform -1 0 2208 0 -1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1725_
timestamp 1676381911
transform -1 0 3168 0 1 11340
box -48 -56 432 834
use sg13g2_buf_1  _1726_
timestamp 1676381911
transform -1 0 2208 0 -1 12852
box -48 -56 432 834
use sg13g2_antennanp  ANTENNA_1
timestamp 1679999689
transform 1 0 7008 0 -1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_2
timestamp 1679999689
transform 1 0 3264 0 -1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_3
timestamp 1679999689
transform 1 0 9216 0 1 40068
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_4
timestamp 1679999689
transform -1 0 2880 0 1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_5
timestamp 1679999689
transform 1 0 2976 0 1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_6
timestamp 1679999689
transform 1 0 6912 0 -1 43092
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_7
timestamp 1679999689
transform 1 0 4224 0 1 41580
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_8
timestamp 1679999689
transform -1 0 7104 0 1 756
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_9
timestamp 1679999689
transform 1 0 7296 0 1 79380
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_10
timestamp 1679999689
transform -1 0 7104 0 -1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_11
timestamp 1679999689
transform 1 0 7296 0 1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_12
timestamp 1679999689
transform 1 0 6816 0 -1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_13
timestamp 1679999689
transform -1 0 4704 0 -1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_14
timestamp 1679999689
transform 1 0 4992 0 1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_15
timestamp 1679999689
transform -1 0 17184 0 1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_16
timestamp 1679999689
transform 1 0 17952 0 1 77868
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_17
timestamp 1679999689
transform 1 0 18432 0 1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_18
timestamp 1679999689
transform 1 0 19584 0 -1 76356
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_19
timestamp 1679999689
transform -1 0 18624 0 -1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_20
timestamp 1679999689
transform 1 0 16032 0 1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_21
timestamp 1679999689
transform -1 0 15648 0 1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_22
timestamp 1679999689
transform -1 0 16608 0 -1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_23
timestamp 1679999689
transform 1 0 18240 0 -1 77868
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_24
timestamp 1679999689
transform 1 0 12864 0 -1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_25
timestamp 1679999689
transform -1 0 12864 0 1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_26
timestamp 1679999689
transform 1 0 12864 0 1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_27
timestamp 1679999689
transform 1 0 12096 0 1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_28
timestamp 1679999689
transform -1 0 1440 0 -1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_29
timestamp 1679999689
transform 1 0 2784 0 1 3780
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_30
timestamp 1679999689
transform 1 0 5664 0 -1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_31
timestamp 1679999689
transform -1 0 3168 0 -1 38556
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_32
timestamp 1679999689
transform 1 0 7008 0 -1 80892
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_33
timestamp 1679999689
transform 1 0 8736 0 -1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_34
timestamp 1679999689
transform 1 0 7296 0 -1 79380
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_35
timestamp 1679999689
transform 1 0 4704 0 1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_36
timestamp 1679999689
transform -1 0 5664 0 1 79380
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_37
timestamp 1679999689
transform 1 0 9216 0 1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_38
timestamp 1679999689
transform -1 0 9888 0 -1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_39
timestamp 1679999689
transform 1 0 11904 0 1 5292
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_40
timestamp 1679999689
transform -1 0 9600 0 -1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_41
timestamp 1679999689
transform -1 0 13920 0 1 2268
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_42
timestamp 1679999689
transform -1 0 5664 0 -1 30996
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_43
timestamp 1679999689
transform 1 0 6528 0 -1 82404
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_44
timestamp 1679999689
transform -1 0 5664 0 -1 32508
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_45
timestamp 1679999689
transform 1 0 6528 0 -1 83916
box -48 -56 336 834
use sg13g2_antennanp  ANTENNA_46
timestamp 1679999689
transform 1 0 19968 0 1 74844
box -48 -56 336 834
use sg13g2_buf_8  clkbuf_0_Tile_X0Y1_UserCLK
timestamp 1676451365
transform 1 0 16512 0 -1 67284
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_0__f_Tile_X0Y1_UserCLK
timestamp 1676451365
transform 1 0 18912 0 -1 58212
box -48 -56 1296 834
use sg13g2_buf_8  clkbuf_1_1__f_Tile_X0Y1_UserCLK
timestamp 1676451365
transform -1 0 16704 0 -1 74844
box -48 -56 1296 834
use sg13g2_fill_1  FILLER_0_0
timestamp 1677579658
transform 1 0 1152 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_22
timestamp 1677580104
transform 1 0 3264 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_41
timestamp 1677579658
transform 1 0 5088 0 1 756
box -48 -56 144 834
use sg13g2_fill_2  FILLER_0_172
timestamp 1677580104
transform 1 0 17664 0 1 756
box -48 -56 240 834
use sg13g2_fill_1  FILLER_0_174
timestamp 1677579658
transform 1 0 17856 0 1 756
box -48 -56 144 834
use sg13g2_decap_4  FILLER_0_196
timestamp 1679577901
transform 1 0 19968 0 1 756
box -48 -56 432 834
use sg13g2_fill_1  FILLER_1_158
timestamp 1677579658
transform 1 0 16320 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_1_176
timestamp 1677580104
transform 1 0 18048 0 -1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_1_178
timestamp 1677579658
transform 1 0 18240 0 -1 2268
box -48 -56 144 834
use sg13g2_fill_2  FILLER_2_0
timestamp 1677580104
transform 1 0 1152 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_19
timestamp 1677580104
transform 1 0 2976 0 1 2268
box -48 -56 240 834
use sg13g2_fill_2  FILLER_2_141
timestamp 1677580104
transform 1 0 14688 0 1 2268
box -48 -56 240 834
use sg13g2_fill_1  FILLER_2_143
timestamp 1677579658
transform 1 0 14880 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_2_182
timestamp 1677579658
transform 1 0 18624 0 1 2268
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_28
timestamp 1677579658
transform 1 0 3840 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_1  FILLER_3_67
timestamp 1677579658
transform 1 0 7584 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_134
timestamp 1677580104
transform 1 0 14016 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_136
timestamp 1677579658
transform 1 0 14208 0 -1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_3_170
timestamp 1677580104
transform 1 0 17472 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_3_172
timestamp 1677579658
transform 1 0 17664 0 -1 3780
box -48 -56 144 834
use sg13g2_decap_4  FILLER_3_194
timestamp 1679577901
transform 1 0 19776 0 -1 3780
box -48 -56 432 834
use sg13g2_fill_2  FILLER_3_198
timestamp 1677580104
transform 1 0 20160 0 -1 3780
box -48 -56 240 834
use sg13g2_fill_2  FILLER_4_37
timestamp 1677580104
transform 1 0 4704 0 1 3780
box -48 -56 240 834
use sg13g2_fill_1  FILLER_4_110
timestamp 1677579658
transform 1 0 11712 0 1 3780
box -48 -56 144 834
use sg13g2_fill_2  FILLER_4_128
timestamp 1677580104
transform 1 0 13440 0 1 3780
box -48 -56 240 834
use sg13g2_decap_8  FILLER_4_164
timestamp 1679581782
transform 1 0 16896 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_4_171
timestamp 1677579658
transform 1 0 17568 0 1 3780
box -48 -56 144 834
use sg13g2_decap_8  FILLER_4_193
timestamp 1679581782
transform 1 0 19680 0 1 3780
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_117
timestamp 1677579658
transform 1 0 12384 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_135
timestamp 1677579658
transform 1 0 14112 0 -1 5292
box -48 -56 144 834
use sg13g2_decap_8  FILLER_5_170
timestamp 1679581782
transform 1 0 17472 0 -1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_5_177
timestamp 1677579658
transform 1 0 18144 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_5_199
timestamp 1677579658
transform 1 0 20256 0 -1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_0
timestamp 1677580104
transform 1 0 1152 0 1 5292
box -48 -56 240 834
use sg13g2_fill_1  FILLER_6_2
timestamp 1677579658
transform 1 0 1344 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_11
timestamp 1677579658
transform 1 0 2208 0 1 5292
box -48 -56 144 834
use sg13g2_fill_2  FILLER_6_78
timestamp 1677580104
transform 1 0 8640 0 1 5292
box -48 -56 240 834
use sg13g2_decap_8  FILLER_6_153
timestamp 1679581782
transform 1 0 15840 0 1 5292
box -48 -56 720 834
use sg13g2_fill_1  FILLER_6_160
timestamp 1677579658
transform 1 0 16512 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_6_199
timestamp 1677579658
transform 1 0 20256 0 1 5292
box -48 -56 144 834
use sg13g2_fill_1  FILLER_7_17
timestamp 1677579658
transform 1 0 2784 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_7_47
timestamp 1677580104
transform 1 0 5664 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_49
timestamp 1677579658
transform 1 0 5856 0 -1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_7_105
timestamp 1679581782
transform 1 0 11232 0 -1 6804
box -48 -56 720 834
use sg13g2_decap_8  FILLER_7_133
timestamp 1679581782
transform 1 0 13920 0 -1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_7_140
timestamp 1677580104
transform 1 0 14592 0 -1 6804
box -48 -56 240 834
use sg13g2_decap_4  FILLER_7_176
timestamp 1679577901
transform 1 0 18048 0 -1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_7_197
timestamp 1677580104
transform 1 0 20064 0 -1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_7_199
timestamp 1677579658
transform 1 0 20256 0 -1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_0
timestamp 1677580104
transform 1 0 1152 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_2
timestamp 1677579658
transform 1 0 1344 0 1 6804
box -48 -56 144 834
use sg13g2_fill_2  FILLER_8_91
timestamp 1677580104
transform 1 0 9888 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_93
timestamp 1677579658
transform 1 0 10080 0 1 6804
box -48 -56 144 834
use sg13g2_decap_8  FILLER_8_111
timestamp 1679581782
transform 1 0 11808 0 1 6804
box -48 -56 720 834
use sg13g2_fill_2  FILLER_8_118
timestamp 1677580104
transform 1 0 12480 0 1 6804
box -48 -56 240 834
use sg13g2_fill_1  FILLER_8_120
timestamp 1677579658
transform 1 0 12672 0 1 6804
box -48 -56 144 834
use sg13g2_fill_1  FILLER_8_159
timestamp 1677579658
transform 1 0 16416 0 1 6804
box -48 -56 144 834
use sg13g2_decap_4  FILLER_8_177
timestamp 1679577901
transform 1 0 18144 0 1 6804
box -48 -56 432 834
use sg13g2_fill_2  FILLER_8_198
timestamp 1677580104
transform 1 0 20160 0 1 6804
box -48 -56 240 834
use sg13g2_fill_2  FILLER_9_25
timestamp 1677580104
transform 1 0 3552 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_111
timestamp 1679577901
transform 1 0 11808 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_115
timestamp 1677580104
transform 1 0 12192 0 -1 8316
box -48 -56 240 834
use sg13g2_decap_4  FILLER_9_168
timestamp 1679577901
transform 1 0 17280 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_1  FILLER_9_172
timestamp 1677579658
transform 1 0 17664 0 -1 8316
box -48 -56 144 834
use sg13g2_decap_4  FILLER_9_194
timestamp 1679577901
transform 1 0 19776 0 -1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_9_198
timestamp 1677580104
transform 1 0 20160 0 -1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_34
timestamp 1677580104
transform 1 0 4416 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_61
timestamp 1677580104
transform 1 0 7008 0 1 8316
box -48 -56 240 834
use sg13g2_decap_8  FILLER_10_84
timestamp 1679581782
transform 1 0 9216 0 1 8316
box -48 -56 720 834
use sg13g2_decap_8  FILLER_10_91
timestamp 1679581782
transform 1 0 9888 0 1 8316
box -48 -56 720 834
use sg13g2_decap_4  FILLER_10_136
timestamp 1679577901
transform 1 0 14208 0 1 8316
box -48 -56 432 834
use sg13g2_fill_2  FILLER_10_140
timestamp 1677580104
transform 1 0 14592 0 1 8316
box -48 -56 240 834
use sg13g2_fill_2  FILLER_10_180
timestamp 1677580104
transform 1 0 18432 0 1 8316
box -48 -56 240 834
use sg13g2_fill_1  FILLER_10_199
timestamp 1677579658
transform 1 0 20256 0 1 8316
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_0
timestamp 1677580104
transform 1 0 1152 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_2  FILLER_11_43
timestamp 1677580104
transform 1 0 5280 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_45
timestamp 1677579658
transform 1 0 5472 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_11_80
timestamp 1679581782
transform 1 0 8832 0 -1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_11_87
timestamp 1677580104
transform 1 0 9504 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_89
timestamp 1677579658
transform 1 0 9696 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_132
timestamp 1679577901
transform 1 0 13824 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_136
timestamp 1677579658
transform 1 0 14208 0 -1 9828
box -48 -56 144 834
use sg13g2_decap_4  FILLER_11_154
timestamp 1679577901
transform 1 0 15936 0 -1 9828
box -48 -56 432 834
use sg13g2_fill_1  FILLER_11_158
timestamp 1677579658
transform 1 0 16320 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_11_197
timestamp 1677580104
transform 1 0 20064 0 -1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_11_199
timestamp 1677579658
transform 1 0 20256 0 -1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_21
timestamp 1677580104
transform 1 0 3168 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_23
timestamp 1677579658
transform 1 0 3360 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_45
timestamp 1677579658
transform 1 0 5472 0 1 9828
box -48 -56 144 834
use sg13g2_decap_8  FILLER_12_67
timestamp 1679581782
transform 1 0 7584 0 1 9828
box -48 -56 720 834
use sg13g2_decap_4  FILLER_12_74
timestamp 1679577901
transform 1 0 8256 0 1 9828
box -48 -56 432 834
use sg13g2_decap_8  FILLER_12_95
timestamp 1679581782
transform 1 0 10272 0 1 9828
box -48 -56 720 834
use sg13g2_fill_2  FILLER_12_102
timestamp 1677580104
transform 1 0 10944 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_104
timestamp 1677579658
transform 1 0 11136 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_122
timestamp 1677579658
transform 1 0 12864 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_140
timestamp 1677579658
transform 1 0 14592 0 1 9828
box -48 -56 144 834
use sg13g2_fill_1  FILLER_12_175
timestamp 1677579658
transform 1 0 17952 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_12_197
timestamp 1677580104
transform 1 0 20064 0 1 9828
box -48 -56 240 834
use sg13g2_fill_1  FILLER_12_199
timestamp 1677579658
transform 1 0 20256 0 1 9828
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_0
timestamp 1677580104
transform 1 0 1152 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_2
timestamp 1677579658
transform 1 0 1344 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_11
timestamp 1677580104
transform 1 0 2208 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_42
timestamp 1677579658
transform 1 0 5184 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_64
timestamp 1679581782
transform 1 0 7296 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_71
timestamp 1679577901
transform 1 0 7968 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_75
timestamp 1677579658
transform 1 0 8352 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_13_114
timestamp 1677580104
transform 1 0 12096 0 -1 11340
box -48 -56 240 834
use sg13g2_fill_1  FILLER_13_116
timestamp 1677579658
transform 1 0 12288 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_142
timestamp 1679581782
transform 1 0 14784 0 -1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_13_149
timestamp 1677579658
transform 1 0 15456 0 -1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_13_171
timestamp 1679581782
transform 1 0 17568 0 -1 11340
box -48 -56 720 834
use sg13g2_decap_4  FILLER_13_178
timestamp 1679577901
transform 1 0 18240 0 -1 11340
box -48 -56 432 834
use sg13g2_fill_1  FILLER_13_199
timestamp 1677579658
transform 1 0 20256 0 -1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_29
timestamp 1677579658
transform 1 0 3936 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_68
timestamp 1679581782
transform 1 0 7680 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_96
timestamp 1677579658
transform 1 0 10368 0 1 11340
box -48 -56 144 834
use sg13g2_fill_1  FILLER_14_118
timestamp 1677579658
transform 1 0 12480 0 1 11340
box -48 -56 144 834
use sg13g2_fill_2  FILLER_14_136
timestamp 1677580104
transform 1 0 14208 0 1 11340
box -48 -56 240 834
use sg13g2_decap_8  FILLER_14_159
timestamp 1679581782
transform 1 0 16416 0 1 11340
box -48 -56 720 834
use sg13g2_fill_1  FILLER_14_166
timestamp 1677579658
transform 1 0 17088 0 1 11340
box -48 -56 144 834
use sg13g2_decap_8  FILLER_14_184
timestamp 1679581782
transform 1 0 18816 0 1 11340
box -48 -56 720 834
use sg13g2_decap_8  FILLER_14_191
timestamp 1679581782
transform 1 0 19488 0 1 11340
box -48 -56 720 834
use sg13g2_fill_2  FILLER_14_198
timestamp 1677580104
transform 1 0 20160 0 1 11340
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_0
timestamp 1677580104
transform 1 0 1152 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_2
timestamp 1677579658
transform 1 0 1344 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_15_15
timestamp 1677579658
transform 1 0 2592 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_33
timestamp 1677580104
transform 1 0 4320 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_35
timestamp 1677579658
transform 1 0 4512 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_53
timestamp 1679577901
transform 1 0 6240 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_15_57
timestamp 1677579658
transform 1 0 6624 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_15_75
timestamp 1679577901
transform 1 0 8352 0 -1 12852
box -48 -56 432 834
use sg13g2_fill_2  FILLER_15_100
timestamp 1677580104
transform 1 0 10752 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_102
timestamp 1677579658
transform 1 0 10944 0 -1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_15_124
timestamp 1679581782
transform 1 0 13056 0 -1 12852
box -48 -56 720 834
use sg13g2_fill_2  FILLER_15_131
timestamp 1677580104
transform 1 0 13728 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_15_137
timestamp 1677580104
transform 1 0 14304 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_156
timestamp 1677579658
transform 1 0 16128 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_174
timestamp 1677580104
transform 1 0 17856 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_1  FILLER_15_176
timestamp 1677579658
transform 1 0 18048 0 -1 12852
box -48 -56 144 834
use sg13g2_fill_2  FILLER_15_198
timestamp 1677580104
transform 1 0 20160 0 -1 12852
box -48 -56 240 834
use sg13g2_fill_2  FILLER_16_0
timestamp 1677580104
transform 1 0 1152 0 1 12852
box -48 -56 240 834
use sg13g2_decap_8  FILLER_16_35
timestamp 1679581782
transform 1 0 4512 0 1 12852
box -48 -56 720 834
use sg13g2_fill_1  FILLER_16_42
timestamp 1677579658
transform 1 0 5184 0 1 12852
box -48 -56 144 834
use sg13g2_fill_1  FILLER_16_64
timestamp 1677579658
transform 1 0 7296 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_82
timestamp 1679577901
transform 1 0 9024 0 1 12852
box -48 -56 432 834
use sg13g2_decap_4  FILLER_16_120
timestamp 1679577901
transform 1 0 12672 0 1 12852
box -48 -56 432 834
use sg13g2_decap_8  FILLER_16_141
timestamp 1679581782
transform 1 0 14688 0 1 12852
box -48 -56 720 834
use sg13g2_decap_4  FILLER_16_148
timestamp 1679577901
transform 1 0 15360 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_152
timestamp 1677579658
transform 1 0 15744 0 1 12852
box -48 -56 144 834
use sg13g2_decap_4  FILLER_16_178
timestamp 1679577901
transform 1 0 18240 0 1 12852
box -48 -56 432 834
use sg13g2_fill_1  FILLER_16_182
timestamp 1677579658
transform 1 0 18624 0 1 12852
box -48 -56 144 834
use sg13g2_decap_8  FILLER_17_38
timestamp 1679581782
transform 1 0 4800 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_4  FILLER_17_45
timestamp 1679577901
transform 1 0 5472 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_49
timestamp 1677580104
transform 1 0 5856 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_4  FILLER_17_72
timestamp 1679577901
transform 1 0 8064 0 -1 14364
box -48 -56 432 834
use sg13g2_decap_4  FILLER_17_97
timestamp 1679577901
transform 1 0 10464 0 -1 14364
box -48 -56 432 834
use sg13g2_fill_2  FILLER_17_101
timestamp 1677580104
transform 1 0 10848 0 -1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_17_162
timestamp 1679581782
transform 1 0 16704 0 -1 14364
box -48 -56 720 834
use sg13g2_decap_8  FILLER_17_169
timestamp 1679581782
transform 1 0 17376 0 -1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_17_176
timestamp 1677580104
transform 1 0 18048 0 -1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_17_199
timestamp 1677579658
transform 1 0 20256 0 -1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_0
timestamp 1677580104
transform 1 0 1152 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_2
timestamp 1677579658
transform 1 0 1344 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_7
timestamp 1677579658
transform 1 0 1824 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_29
timestamp 1677580104
transform 1 0 3936 0 1 14364
box -48 -56 240 834
use sg13g2_fill_2  FILLER_18_48
timestamp 1677580104
transform 1 0 5760 0 1 14364
box -48 -56 240 834
use sg13g2_decap_8  FILLER_18_67
timestamp 1679581782
transform 1 0 7584 0 1 14364
box -48 -56 720 834
use sg13g2_fill_1  FILLER_18_74
timestamp 1677579658
transform 1 0 8256 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_92
timestamp 1679577901
transform 1 0 9984 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_96
timestamp 1677579658
transform 1 0 10368 0 1 14364
box -48 -56 144 834
use sg13g2_decap_8  FILLER_18_114
timestamp 1679581782
transform 1 0 12096 0 1 14364
box -48 -56 720 834
use sg13g2_fill_2  FILLER_18_121
timestamp 1677580104
transform 1 0 12768 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_123
timestamp 1677579658
transform 1 0 12960 0 1 14364
box -48 -56 144 834
use sg13g2_fill_2  FILLER_18_141
timestamp 1677580104
transform 1 0 14688 0 1 14364
box -48 -56 240 834
use sg13g2_fill_1  FILLER_18_143
timestamp 1677579658
transform 1 0 14880 0 1 14364
box -48 -56 144 834
use sg13g2_fill_1  FILLER_18_169
timestamp 1677579658
transform 1 0 17376 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_18_195
timestamp 1679577901
transform 1 0 19872 0 1 14364
box -48 -56 432 834
use sg13g2_fill_1  FILLER_18_199
timestamp 1677579658
transform 1 0 20256 0 1 14364
box -48 -56 144 834
use sg13g2_decap_4  FILLER_19_21
timestamp 1679577901
transform 1 0 3168 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_19_25
timestamp 1677579658
transform 1 0 3552 0 -1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_19_77
timestamp 1677580104
transform 1 0 8544 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_19_96
timestamp 1679577901
transform 1 0 10368 0 -1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_19_100
timestamp 1677580104
transform 1 0 10752 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_174
timestamp 1677580104
transform 1 0 17856 0 -1 15876
box -48 -56 240 834
use sg13g2_fill_2  FILLER_19_198
timestamp 1677580104
transform 1 0 20160 0 -1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_20_4
timestamp 1679581782
transform 1 0 1536 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_11
timestamp 1677580104
transform 1 0 2208 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_13
timestamp 1677579658
transform 1 0 2400 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_35
timestamp 1679581782
transform 1 0 4512 0 1 15876
box -48 -56 720 834
use sg13g2_fill_2  FILLER_20_42
timestamp 1677580104
transform 1 0 5184 0 1 15876
box -48 -56 240 834
use sg13g2_fill_1  FILLER_20_44
timestamp 1677579658
transform 1 0 5376 0 1 15876
box -48 -56 144 834
use sg13g2_decap_4  FILLER_20_66
timestamp 1679577901
transform 1 0 7488 0 1 15876
box -48 -56 432 834
use sg13g2_fill_2  FILLER_20_70
timestamp 1677580104
transform 1 0 7872 0 1 15876
box -48 -56 240 834
use sg13g2_decap_4  FILLER_20_114
timestamp 1679577901
transform 1 0 12096 0 1 15876
box -48 -56 432 834
use sg13g2_fill_1  FILLER_20_118
timestamp 1677579658
transform 1 0 12480 0 1 15876
box -48 -56 144 834
use sg13g2_decap_8  FILLER_20_140
timestamp 1679581782
transform 1 0 14592 0 1 15876
box -48 -56 720 834
use sg13g2_fill_1  FILLER_20_147
timestamp 1677579658
transform 1 0 15264 0 1 15876
box -48 -56 144 834
use sg13g2_fill_2  FILLER_20_198
timestamp 1677580104
transform 1 0 20160 0 1 15876
box -48 -56 240 834
use sg13g2_decap_8  FILLER_21_0
timestamp 1679581782
transform 1 0 1152 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_7
timestamp 1677580104
transform 1 0 1824 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_9
timestamp 1677579658
transform 1 0 2016 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_21_31
timestamp 1679581782
transform 1 0 4128 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_21_38
timestamp 1677580104
transform 1 0 4800 0 -1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_21_40
timestamp 1677579658
transform 1 0 4992 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_21_79
timestamp 1679577901
transform 1 0 8736 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_4  FILLER_21_100
timestamp 1679577901
transform 1 0 10752 0 -1 17388
box -48 -56 432 834
use sg13g2_fill_1  FILLER_21_104
timestamp 1677579658
transform 1 0 11136 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_4  FILLER_21_122
timestamp 1679577901
transform 1 0 12864 0 -1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_21_143
timestamp 1679581782
transform 1 0 14880 0 -1 17388
box -48 -56 720 834
use sg13g2_fill_1  FILLER_21_150
timestamp 1677579658
transform 1 0 15552 0 -1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_22_17
timestamp 1679581782
transform 1 0 2784 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_24
timestamp 1679581782
transform 1 0 3456 0 1 17388
box -48 -56 720 834
use sg13g2_fill_2  FILLER_22_31
timestamp 1677580104
transform 1 0 4128 0 1 17388
box -48 -56 240 834
use sg13g2_decap_8  FILLER_22_50
timestamp 1679581782
transform 1 0 5952 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_57
timestamp 1679577901
transform 1 0 6624 0 1 17388
box -48 -56 432 834
use sg13g2_decap_8  FILLER_22_99
timestamp 1679581782
transform 1 0 10656 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_106
timestamp 1679581782
transform 1 0 11328 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_113
timestamp 1679581782
transform 1 0 12000 0 1 17388
box -48 -56 720 834
use sg13g2_decap_8  FILLER_22_120
timestamp 1679581782
transform 1 0 12672 0 1 17388
box -48 -56 720 834
use sg13g2_decap_4  FILLER_22_144
timestamp 1679577901
transform 1 0 14976 0 1 17388
box -48 -56 432 834
use sg13g2_decap_4  FILLER_22_165
timestamp 1679577901
transform 1 0 16992 0 1 17388
box -48 -56 432 834
use sg13g2_fill_2  FILLER_22_169
timestamp 1677580104
transform 1 0 17376 0 1 17388
box -48 -56 240 834
use sg13g2_fill_1  FILLER_22_199
timestamp 1677579658
transform 1 0 20256 0 1 17388
box -48 -56 144 834
use sg13g2_decap_8  FILLER_23_0
timestamp 1679581782
transform 1 0 1152 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_7
timestamp 1679577901
transform 1 0 1824 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_2  FILLER_23_11
timestamp 1677580104
transform 1 0 2208 0 -1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_23_34
timestamp 1679581782
transform 1 0 4416 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_4  FILLER_23_41
timestamp 1679577901
transform 1 0 5088 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_8  FILLER_23_66
timestamp 1679581782
transform 1 0 7488 0 -1 18900
box -48 -56 720 834
use sg13g2_decap_8  FILLER_23_73
timestamp 1679581782
transform 1 0 8160 0 -1 18900
box -48 -56 720 834
use sg13g2_fill_2  FILLER_23_80
timestamp 1677580104
transform 1 0 8832 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_23_99
timestamp 1677580104
transform 1 0 10656 0 -1 18900
box -48 -56 240 834
use sg13g2_fill_1  FILLER_23_101
timestamp 1677579658
transform 1 0 10848 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_23_140
timestamp 1679577901
transform 1 0 14592 0 -1 18900
box -48 -56 432 834
use sg13g2_decap_4  FILLER_23_174
timestamp 1679577901
transform 1 0 17856 0 -1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_23_178
timestamp 1677579658
transform 1 0 18240 0 -1 18900
box -48 -56 144 834
use sg13g2_decap_4  FILLER_24_38
timestamp 1679577901
transform 1 0 4800 0 1 18900
box -48 -56 432 834
use sg13g2_fill_1  FILLER_24_42
timestamp 1677579658
transform 1 0 5184 0 1 18900
box -48 -56 144 834
use sg13g2_fill_2  FILLER_24_98
timestamp 1677580104
transform 1 0 10560 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_138
timestamp 1677580104
transform 1 0 14400 0 1 18900
box -48 -56 240 834
use sg13g2_fill_2  FILLER_24_198
timestamp 1677580104
transform 1 0 20160 0 1 18900
box -48 -56 240 834
use sg13g2_decap_8  FILLER_25_17
timestamp 1679581782
transform 1 0 2784 0 -1 20412
box -48 -56 720 834
use sg13g2_fill_2  FILLER_25_24
timestamp 1677580104
transform 1 0 3456 0 -1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_25_77
timestamp 1677579658
transform 1 0 8544 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_95
timestamp 1679577901
transform 1 0 10272 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_25_99
timestamp 1677579658
transform 1 0 10656 0 -1 20412
box -48 -56 144 834
use sg13g2_decap_4  FILLER_25_117
timestamp 1679577901
transform 1 0 12384 0 -1 20412
box -48 -56 432 834
use sg13g2_decap_4  FILLER_25_138
timestamp 1679577901
transform 1 0 14400 0 -1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_25_177
timestamp 1677580104
transform 1 0 18144 0 -1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_17
timestamp 1679581782
transform 1 0 2784 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_24
timestamp 1679577901
transform 1 0 3456 0 1 20412
box -48 -56 432 834
use sg13g2_fill_1  FILLER_26_28
timestamp 1677579658
transform 1 0 3840 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_67
timestamp 1679581782
transform 1 0 7584 0 1 20412
box -48 -56 720 834
use sg13g2_fill_1  FILLER_26_74
timestamp 1677579658
transform 1 0 8256 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_26_117
timestamp 1679581782
transform 1 0 12384 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_124
timestamp 1679577901
transform 1 0 13056 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_128
timestamp 1677580104
transform 1 0 13440 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_152
timestamp 1677580104
transform 1 0 15744 0 1 20412
box -48 -56 240 834
use sg13g2_decap_8  FILLER_26_167
timestamp 1679581782
transform 1 0 17184 0 1 20412
box -48 -56 720 834
use sg13g2_decap_4  FILLER_26_174
timestamp 1679577901
transform 1 0 17856 0 1 20412
box -48 -56 432 834
use sg13g2_fill_2  FILLER_26_178
timestamp 1677580104
transform 1 0 18240 0 1 20412
box -48 -56 240 834
use sg13g2_fill_2  FILLER_26_197
timestamp 1677580104
transform 1 0 20064 0 1 20412
box -48 -56 240 834
use sg13g2_fill_1  FILLER_26_199
timestamp 1677579658
transform 1 0 20256 0 1 20412
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_0
timestamp 1679581782
transform 1 0 1152 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_27_11
timestamp 1677580104
transform 1 0 2208 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_27_34
timestamp 1677580104
transform 1 0 4416 0 -1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_27_36
timestamp 1677579658
transform 1 0 4608 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_54
timestamp 1679581782
transform 1 0 6336 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_8  FILLER_27_61
timestamp 1679581782
transform 1 0 7008 0 -1 21924
box -48 -56 720 834
use sg13g2_fill_1  FILLER_27_68
timestamp 1677579658
transform 1 0 7680 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_27_103
timestamp 1679581782
transform 1 0 11040 0 -1 21924
box -48 -56 720 834
use sg13g2_decap_4  FILLER_27_110
timestamp 1679577901
transform 1 0 11712 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_114
timestamp 1677579658
transform 1 0 12096 0 -1 21924
box -48 -56 144 834
use sg13g2_decap_4  FILLER_27_157
timestamp 1679577901
transform 1 0 16224 0 -1 21924
box -48 -56 432 834
use sg13g2_fill_1  FILLER_27_199
timestamp 1677579658
transform 1 0 20256 0 -1 21924
box -48 -56 144 834
use sg13g2_fill_2  FILLER_28_34
timestamp 1677580104
transform 1 0 4416 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_28_57
timestamp 1679581782
transform 1 0 6624 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_64
timestamp 1677580104
transform 1 0 7296 0 1 21924
box -48 -56 240 834
use sg13g2_fill_1  FILLER_28_66
timestamp 1677579658
transform 1 0 7488 0 1 21924
box -48 -56 144 834
use sg13g2_decap_8  FILLER_28_88
timestamp 1679581782
transform 1 0 9600 0 1 21924
box -48 -56 720 834
use sg13g2_fill_2  FILLER_28_95
timestamp 1677580104
transform 1 0 10272 0 1 21924
box -48 -56 240 834
use sg13g2_fill_2  FILLER_28_135
timestamp 1677580104
transform 1 0 14112 0 1 21924
box -48 -56 240 834
use sg13g2_decap_8  FILLER_29_17
timestamp 1679581782
transform 1 0 2784 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_24
timestamp 1677580104
transform 1 0 3456 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_70
timestamp 1679577901
transform 1 0 7872 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_74
timestamp 1677579658
transform 1 0 8256 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_109
timestamp 1677579658
transform 1 0 11616 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_29_115
timestamp 1679581782
transform 1 0 12192 0 -1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_29_139
timestamp 1677580104
transform 1 0 14496 0 -1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_29_177
timestamp 1679577901
transform 1 0 18144 0 -1 23436
box -48 -56 432 834
use sg13g2_fill_1  FILLER_29_181
timestamp 1677579658
transform 1 0 18528 0 -1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_29_199
timestamp 1677579658
transform 1 0 20256 0 -1 23436
box -48 -56 144 834
use sg13g2_decap_8  FILLER_30_0
timestamp 1679581782
transform 1 0 1152 0 1 23436
box -48 -56 720 834
use sg13g2_fill_2  FILLER_30_7
timestamp 1677580104
transform 1 0 1824 0 1 23436
box -48 -56 240 834
use sg13g2_fill_1  FILLER_30_9
timestamp 1677579658
transform 1 0 2016 0 1 23436
box -48 -56 144 834
use sg13g2_fill_1  FILLER_30_72
timestamp 1677579658
transform 1 0 8064 0 1 23436
box -48 -56 144 834
use sg13g2_fill_2  FILLER_30_94
timestamp 1677580104
transform 1 0 10176 0 1 23436
box -48 -56 240 834
use sg13g2_fill_2  FILLER_30_164
timestamp 1677580104
transform 1 0 16896 0 1 23436
box -48 -56 240 834
use sg13g2_decap_4  FILLER_31_0
timestamp 1679577901
transform 1 0 1152 0 -1 24948
box -48 -56 432 834
use sg13g2_fill_2  FILLER_31_30
timestamp 1677580104
transform 1 0 4032 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_49
timestamp 1677580104
transform 1 0 5856 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_89
timestamp 1677580104
transform 1 0 9696 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_2  FILLER_31_137
timestamp 1677580104
transform 1 0 14304 0 -1 24948
box -48 -56 240 834
use sg13g2_fill_1  FILLER_31_139
timestamp 1677579658
transform 1 0 14496 0 -1 24948
box -48 -56 144 834
use sg13g2_decap_4  FILLER_32_95
timestamp 1679577901
transform 1 0 10272 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_99
timestamp 1677579658
transform 1 0 10656 0 1 24948
box -48 -56 144 834
use sg13g2_decap_8  FILLER_32_138
timestamp 1679581782
transform 1 0 14400 0 1 24948
box -48 -56 720 834
use sg13g2_fill_2  FILLER_32_159
timestamp 1677580104
transform 1 0 16416 0 1 24948
box -48 -56 240 834
use sg13g2_decap_4  FILLER_32_195
timestamp 1679577901
transform 1 0 19872 0 1 24948
box -48 -56 432 834
use sg13g2_fill_1  FILLER_32_199
timestamp 1677579658
transform 1 0 20256 0 1 24948
box -48 -56 144 834
use sg13g2_fill_2  FILLER_33_17
timestamp 1677580104
transform 1 0 2784 0 -1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_33_60
timestamp 1679577901
transform 1 0 6912 0 -1 26460
box -48 -56 432 834
use sg13g2_decap_8  FILLER_33_115
timestamp 1679581782
transform 1 0 12192 0 -1 26460
box -48 -56 720 834
use sg13g2_decap_8  FILLER_33_122
timestamp 1679581782
transform 1 0 12864 0 -1 26460
box -48 -56 720 834
use sg13g2_fill_2  FILLER_33_197
timestamp 1677580104
transform 1 0 20064 0 -1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_33_199
timestamp 1677579658
transform 1 0 20256 0 -1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_0
timestamp 1679581782
transform 1 0 1152 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_7
timestamp 1679577901
transform 1 0 1824 0 1 26460
box -48 -56 432 834
use sg13g2_fill_1  FILLER_34_54
timestamp 1677579658
transform 1 0 6336 0 1 26460
box -48 -56 144 834
use sg13g2_decap_4  FILLER_34_70
timestamp 1679577901
transform 1 0 7872 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_74
timestamp 1677580104
transform 1 0 8256 0 1 26460
box -48 -56 240 834
use sg13g2_decap_4  FILLER_34_120
timestamp 1679577901
transform 1 0 12672 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_124
timestamp 1677580104
transform 1 0 13056 0 1 26460
box -48 -56 240 834
use sg13g2_fill_1  FILLER_34_148
timestamp 1677579658
transform 1 0 15360 0 1 26460
box -48 -56 144 834
use sg13g2_decap_8  FILLER_34_187
timestamp 1679581782
transform 1 0 19104 0 1 26460
box -48 -56 720 834
use sg13g2_decap_4  FILLER_34_194
timestamp 1679577901
transform 1 0 19776 0 1 26460
box -48 -56 432 834
use sg13g2_fill_2  FILLER_34_198
timestamp 1677580104
transform 1 0 20160 0 1 26460
box -48 -56 240 834
use sg13g2_decap_8  FILLER_35_0
timestamp 1679581782
transform 1 0 1152 0 -1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_35_7
timestamp 1679581782
transform 1 0 1824 0 -1 27972
box -48 -56 720 834
use sg13g2_fill_2  FILLER_35_14
timestamp 1677580104
transform 1 0 2496 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_1  FILLER_35_37
timestamp 1677579658
transform 1 0 4704 0 -1 27972
box -48 -56 144 834
use sg13g2_fill_1  FILLER_35_64
timestamp 1677579658
transform 1 0 7296 0 -1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_35_103
timestamp 1679577901
transform 1 0 11040 0 -1 27972
box -48 -56 432 834
use sg13g2_fill_2  FILLER_35_123
timestamp 1677580104
transform 1 0 12960 0 -1 27972
box -48 -56 240 834
use sg13g2_fill_2  FILLER_35_135
timestamp 1677580104
transform 1 0 14112 0 -1 27972
box -48 -56 240 834
use sg13g2_decap_4  FILLER_35_179
timestamp 1679577901
transform 1 0 18336 0 -1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_0
timestamp 1679581782
transform 1 0 1152 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_7
timestamp 1679581782
transform 1 0 1824 0 1 27972
box -48 -56 720 834
use sg13g2_fill_1  FILLER_36_14
timestamp 1677579658
transform 1 0 2496 0 1 27972
box -48 -56 144 834
use sg13g2_decap_4  FILLER_36_49
timestamp 1679577901
transform 1 0 5856 0 1 27972
box -48 -56 432 834
use sg13g2_decap_8  FILLER_36_73
timestamp 1679581782
transform 1 0 8160 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_36_80
timestamp 1679577901
transform 1 0 8832 0 1 27972
box -48 -56 432 834
use sg13g2_fill_1  FILLER_36_84
timestamp 1677579658
transform 1 0 9216 0 1 27972
box -48 -56 144 834
use sg13g2_decap_8  FILLER_36_102
timestamp 1679581782
transform 1 0 10944 0 1 27972
box -48 -56 720 834
use sg13g2_decap_8  FILLER_36_109
timestamp 1679581782
transform 1 0 11616 0 1 27972
box -48 -56 720 834
use sg13g2_decap_4  FILLER_37_0
timestamp 1679577901
transform 1 0 1152 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_1  FILLER_37_4
timestamp 1677579658
transform 1 0 1536 0 -1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_37_22
timestamp 1679581782
transform 1 0 3264 0 -1 29484
box -48 -56 720 834
use sg13g2_fill_2  FILLER_37_29
timestamp 1677580104
transform 1 0 3936 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_31
timestamp 1677579658
transform 1 0 4128 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_49
timestamp 1677579658
transform 1 0 5856 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_37_104
timestamp 1677579658
transform 1 0 11136 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_151
timestamp 1677580104
transform 1 0 15648 0 -1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_37_153
timestamp 1677579658
transform 1 0 15840 0 -1 29484
box -48 -56 144 834
use sg13g2_fill_2  FILLER_37_171
timestamp 1677580104
transform 1 0 17568 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_4  FILLER_37_194
timestamp 1679577901
transform 1 0 19776 0 -1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_37_198
timestamp 1677580104
transform 1 0 20160 0 -1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_0
timestamp 1679581782
transform 1 0 1152 0 1 29484
box -48 -56 720 834
use sg13g2_decap_4  FILLER_38_7
timestamp 1679577901
transform 1 0 1824 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_49
timestamp 1677580104
transform 1 0 5856 0 1 29484
box -48 -56 240 834
use sg13g2_fill_1  FILLER_38_51
timestamp 1677579658
transform 1 0 6048 0 1 29484
box -48 -56 144 834
use sg13g2_decap_4  FILLER_38_60
timestamp 1679577901
transform 1 0 6912 0 1 29484
box -48 -56 432 834
use sg13g2_fill_2  FILLER_38_64
timestamp 1677580104
transform 1 0 7296 0 1 29484
box -48 -56 240 834
use sg13g2_decap_8  FILLER_38_83
timestamp 1679581782
transform 1 0 9120 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_90
timestamp 1679581782
transform 1 0 9792 0 1 29484
box -48 -56 720 834
use sg13g2_decap_8  FILLER_38_97
timestamp 1679581782
transform 1 0 10464 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_104
timestamp 1677579658
transform 1 0 11136 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_125
timestamp 1677579658
transform 1 0 13152 0 1 29484
box -48 -56 144 834
use sg13g2_fill_1  FILLER_38_136
timestamp 1677579658
transform 1 0 14208 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_38_192
timestamp 1679581782
transform 1 0 19584 0 1 29484
box -48 -56 720 834
use sg13g2_fill_1  FILLER_38_199
timestamp 1677579658
transform 1 0 20256 0 1 29484
box -48 -56 144 834
use sg13g2_decap_8  FILLER_39_17
timestamp 1679581782
transform 1 0 2784 0 -1 30996
box -48 -56 720 834
use sg13g2_fill_2  FILLER_39_24
timestamp 1677580104
transform 1 0 3456 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_26
timestamp 1677579658
transform 1 0 3648 0 -1 30996
box -48 -56 144 834
use sg13g2_fill_2  FILLER_39_47
timestamp 1677580104
transform 1 0 5664 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_49
timestamp 1677579658
transform 1 0 5856 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_39_67
timestamp 1679577901
transform 1 0 7584 0 -1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_39_71
timestamp 1677580104
transform 1 0 7968 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_2  FILLER_39_180
timestamp 1677580104
transform 1 0 18432 0 -1 30996
box -48 -56 240 834
use sg13g2_fill_1  FILLER_39_182
timestamp 1677579658
transform 1 0 18624 0 -1 30996
box -48 -56 144 834
use sg13g2_decap_4  FILLER_40_0
timestamp 1679577901
transform 1 0 1152 0 1 30996
box -48 -56 432 834
use sg13g2_fill_2  FILLER_40_42
timestamp 1677580104
transform 1 0 5184 0 1 30996
box -48 -56 240 834
use sg13g2_decap_8  FILLER_40_107
timestamp 1679581782
transform 1 0 11424 0 1 30996
box -48 -56 720 834
use sg13g2_decap_4  FILLER_40_114
timestamp 1679577901
transform 1 0 12096 0 1 30996
box -48 -56 432 834
use sg13g2_fill_1  FILLER_40_118
timestamp 1677579658
transform 1 0 12480 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_139
timestamp 1677579658
transform 1 0 14496 0 1 30996
box -48 -56 144 834
use sg13g2_fill_1  FILLER_40_199
timestamp 1677579658
transform 1 0 20256 0 1 30996
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_0
timestamp 1679581782
transform 1 0 1152 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_28
timestamp 1679581782
transform 1 0 3840 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_35
timestamp 1679581782
transform 1 0 4512 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_42
timestamp 1677580104
transform 1 0 5184 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_2  FILLER_41_64
timestamp 1677580104
transform 1 0 7296 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_66
timestamp 1677579658
transform 1 0 7488 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_4  FILLER_41_95
timestamp 1679577901
transform 1 0 10272 0 -1 32508
box -48 -56 432 834
use sg13g2_decap_8  FILLER_41_137
timestamp 1679581782
transform 1 0 14304 0 -1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_41_161
timestamp 1679581782
transform 1 0 16608 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_41_168
timestamp 1677580104
transform 1 0 17280 0 -1 32508
box -48 -56 240 834
use sg13g2_fill_1  FILLER_41_170
timestamp 1677579658
transform 1 0 17472 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_41_192
timestamp 1679581782
transform 1 0 19584 0 -1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_41_199
timestamp 1677579658
transform 1 0 20256 0 -1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_17
timestamp 1679581782
transform 1 0 2784 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_24
timestamp 1679581782
transform 1 0 3456 0 1 32508
box -48 -56 720 834
use sg13g2_fill_1  FILLER_42_67
timestamp 1677579658
transform 1 0 7584 0 1 32508
box -48 -56 144 834
use sg13g2_decap_8  FILLER_42_119
timestamp 1679581782
transform 1 0 12576 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_126
timestamp 1679581782
transform 1 0 13248 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_133
timestamp 1679581782
transform 1 0 13920 0 1 32508
box -48 -56 720 834
use sg13g2_decap_8  FILLER_42_161
timestamp 1679581782
transform 1 0 16608 0 1 32508
box -48 -56 720 834
use sg13g2_decap_4  FILLER_42_168
timestamp 1679577901
transform 1 0 17280 0 1 32508
box -48 -56 432 834
use sg13g2_fill_2  FILLER_42_172
timestamp 1677580104
transform 1 0 17664 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_42_191
timestamp 1679581782
transform 1 0 19488 0 1 32508
box -48 -56 720 834
use sg13g2_fill_2  FILLER_42_198
timestamp 1677580104
transform 1 0 20160 0 1 32508
box -48 -56 240 834
use sg13g2_decap_8  FILLER_43_0
timestamp 1679581782
transform 1 0 1152 0 -1 34020
box -48 -56 720 834
use sg13g2_fill_2  FILLER_43_7
timestamp 1677580104
transform 1 0 1824 0 -1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_43_9
timestamp 1677579658
transform 1 0 2016 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_31
timestamp 1677579658
transform 1 0 4128 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_72
timestamp 1677579658
transform 1 0 8064 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_43_121
timestamp 1677579658
transform 1 0 12768 0 -1 34020
box -48 -56 144 834
use sg13g2_fill_2  FILLER_43_177
timestamp 1677580104
transform 1 0 18144 0 -1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_0
timestamp 1679577901
transform 1 0 1152 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_4
timestamp 1677580104
transform 1 0 1536 0 1 34020
box -48 -56 240 834
use sg13g2_decap_4  FILLER_44_23
timestamp 1679577901
transform 1 0 3360 0 1 34020
box -48 -56 432 834
use sg13g2_fill_2  FILLER_44_27
timestamp 1677580104
transform 1 0 3744 0 1 34020
box -48 -56 240 834
use sg13g2_fill_1  FILLER_44_46
timestamp 1677579658
transform 1 0 5568 0 1 34020
box -48 -56 144 834
use sg13g2_fill_1  FILLER_44_65
timestamp 1677579658
transform 1 0 7392 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_104
timestamp 1679581782
transform 1 0 11136 0 1 34020
box -48 -56 720 834
use sg13g2_decap_4  FILLER_44_111
timestamp 1679577901
transform 1 0 11808 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_115
timestamp 1677579658
transform 1 0 12192 0 1 34020
box -48 -56 144 834
use sg13g2_decap_4  FILLER_44_167
timestamp 1679577901
transform 1 0 17184 0 1 34020
box -48 -56 432 834
use sg13g2_fill_1  FILLER_44_171
timestamp 1677579658
transform 1 0 17568 0 1 34020
box -48 -56 144 834
use sg13g2_decap_8  FILLER_44_193
timestamp 1679581782
transform 1 0 19680 0 1 34020
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_0
timestamp 1679581782
transform 1 0 1152 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_28
timestamp 1679581782
transform 1 0 3840 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_35
timestamp 1679581782
transform 1 0 4512 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_65
timestamp 1679581782
transform 1 0 7392 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_72
timestamp 1679581782
transform 1 0 8064 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_79
timestamp 1679581782
transform 1 0 8736 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_86
timestamp 1677580104
transform 1 0 9408 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_105
timestamp 1679581782
transform 1 0 11232 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_112
timestamp 1677580104
transform 1 0 11904 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_45_135
timestamp 1679581782
transform 1 0 14112 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_142
timestamp 1679581782
transform 1 0 14784 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_1  FILLER_45_149
timestamp 1677579658
transform 1 0 15456 0 -1 35532
box -48 -56 144 834
use sg13g2_decap_8  FILLER_45_184
timestamp 1679581782
transform 1 0 18816 0 -1 35532
box -48 -56 720 834
use sg13g2_decap_8  FILLER_45_191
timestamp 1679581782
transform 1 0 19488 0 -1 35532
box -48 -56 720 834
use sg13g2_fill_2  FILLER_45_198
timestamp 1677580104
transform 1 0 20160 0 -1 35532
box -48 -56 240 834
use sg13g2_decap_8  FILLER_46_17
timestamp 1679581782
transform 1 0 2784 0 1 35532
box -48 -56 720 834
use sg13g2_decap_4  FILLER_46_24
timestamp 1679577901
transform 1 0 3456 0 1 35532
box -48 -56 432 834
use sg13g2_fill_1  FILLER_46_28
timestamp 1677579658
transform 1 0 3840 0 1 35532
box -48 -56 144 834
use sg13g2_fill_1  FILLER_46_46
timestamp 1677579658
transform 1 0 5568 0 1 35532
box -48 -56 144 834
use sg13g2_decap_4  FILLER_46_123
timestamp 1679577901
transform 1 0 12960 0 1 35532
box -48 -56 432 834
use sg13g2_fill_2  FILLER_46_161
timestamp 1677580104
transform 1 0 16608 0 1 35532
box -48 -56 240 834
use sg13g2_fill_2  FILLER_46_197
timestamp 1677580104
transform 1 0 20064 0 1 35532
box -48 -56 240 834
use sg13g2_fill_1  FILLER_46_199
timestamp 1677579658
transform 1 0 20256 0 1 35532
box -48 -56 144 834
use sg13g2_fill_2  FILLER_47_70
timestamp 1677580104
transform 1 0 7872 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_47_72
timestamp 1677579658
transform 1 0 8064 0 -1 37044
box -48 -56 144 834
use sg13g2_decap_4  FILLER_47_94
timestamp 1679577901
transform 1 0 10176 0 -1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_47_98
timestamp 1677580104
transform 1 0 10560 0 -1 37044
box -48 -56 240 834
use sg13g2_fill_2  FILLER_47_117
timestamp 1677580104
transform 1 0 12384 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_140
timestamp 1679581782
transform 1 0 14592 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_147
timestamp 1677580104
transform 1 0 15264 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_8  FILLER_47_170
timestamp 1679581782
transform 1 0 17472 0 -1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_47_198
timestamp 1677580104
transform 1 0 20160 0 -1 37044
box -48 -56 240 834
use sg13g2_decap_4  FILLER_48_38
timestamp 1679577901
transform 1 0 4800 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_42
timestamp 1677580104
transform 1 0 5184 0 1 37044
box -48 -56 240 834
use sg13g2_decap_4  FILLER_48_91
timestamp 1679577901
transform 1 0 9888 0 1 37044
box -48 -56 432 834
use sg13g2_fill_2  FILLER_48_95
timestamp 1677580104
transform 1 0 10272 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_135
timestamp 1677579658
transform 1 0 14112 0 1 37044
box -48 -56 144 834
use sg13g2_decap_8  FILLER_48_170
timestamp 1679581782
transform 1 0 17472 0 1 37044
box -48 -56 720 834
use sg13g2_fill_2  FILLER_48_177
timestamp 1677580104
transform 1 0 18144 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_179
timestamp 1677579658
transform 1 0 18336 0 1 37044
box -48 -56 144 834
use sg13g2_fill_2  FILLER_48_197
timestamp 1677580104
transform 1 0 20064 0 1 37044
box -48 -56 240 834
use sg13g2_fill_1  FILLER_48_199
timestamp 1677579658
transform 1 0 20256 0 1 37044
box -48 -56 144 834
use sg13g2_fill_1  FILLER_49_17
timestamp 1677579658
transform 1 0 2784 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_49_21
timestamp 1679581782
transform 1 0 3168 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_62
timestamp 1679581782
transform 1 0 7104 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_69
timestamp 1679581782
transform 1 0 7776 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_49_76
timestamp 1679581782
transform 1 0 8448 0 -1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_49_83
timestamp 1677579658
transform 1 0 9120 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_101
timestamp 1677580104
transform 1 0 10848 0 -1 38556
box -48 -56 240 834
use sg13g2_decap_8  FILLER_49_108
timestamp 1679581782
transform 1 0 11520 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_115
timestamp 1679577901
transform 1 0 12192 0 -1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_49_136
timestamp 1679581782
transform 1 0 14208 0 -1 38556
box -48 -56 720 834
use sg13g2_decap_4  FILLER_49_143
timestamp 1679577901
transform 1 0 14880 0 -1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_49_147
timestamp 1677579658
transform 1 0 15264 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_186
timestamp 1677580104
transform 1 0 19008 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_188
timestamp 1677579658
transform 1 0 19200 0 -1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_49_197
timestamp 1677580104
transform 1 0 20064 0 -1 38556
box -48 -56 240 834
use sg13g2_fill_1  FILLER_49_199
timestamp 1677579658
transform 1 0 20256 0 -1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_50_0
timestamp 1679581782
transform 1 0 1152 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_7
timestamp 1679581782
transform 1 0 1824 0 1 38556
box -48 -56 720 834
use sg13g2_fill_1  FILLER_50_14
timestamp 1677579658
transform 1 0 2496 0 1 38556
box -48 -56 144 834
use sg13g2_fill_2  FILLER_50_39
timestamp 1677580104
transform 1 0 4896 0 1 38556
box -48 -56 240 834
use sg13g2_decap_4  FILLER_50_83
timestamp 1679577901
transform 1 0 9120 0 1 38556
box -48 -56 432 834
use sg13g2_decap_8  FILLER_50_141
timestamp 1679581782
transform 1 0 14688 0 1 38556
box -48 -56 720 834
use sg13g2_decap_8  FILLER_50_148
timestamp 1679581782
transform 1 0 15360 0 1 38556
box -48 -56 720 834
use sg13g2_fill_2  FILLER_50_155
timestamp 1677580104
transform 1 0 16032 0 1 38556
box -48 -56 240 834
use sg13g2_decap_4  FILLER_50_174
timestamp 1679577901
transform 1 0 17856 0 1 38556
box -48 -56 432 834
use sg13g2_fill_1  FILLER_50_199
timestamp 1677579658
transform 1 0 20256 0 1 38556
box -48 -56 144 834
use sg13g2_decap_8  FILLER_51_0
timestamp 1679581782
transform 1 0 1152 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_4  FILLER_51_7
timestamp 1679577901
transform 1 0 1824 0 -1 40068
box -48 -56 432 834
use sg13g2_fill_2  FILLER_51_11
timestamp 1677580104
transform 1 0 2208 0 -1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_51_83
timestamp 1677579658
transform 1 0 9120 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_94
timestamp 1677579658
transform 1 0 10176 0 -1 40068
box -48 -56 144 834
use sg13g2_decap_4  FILLER_51_100
timestamp 1679577901
transform 1 0 10752 0 -1 40068
box -48 -56 432 834
use sg13g2_fill_1  FILLER_51_104
timestamp 1677579658
transform 1 0 11136 0 -1 40068
box -48 -56 144 834
use sg13g2_fill_1  FILLER_51_150
timestamp 1677579658
transform 1 0 15552 0 -1 40068
box -48 -56 144 834
use sg13g2_decap_8  FILLER_51_168
timestamp 1679581782
transform 1 0 17280 0 -1 40068
box -48 -56 720 834
use sg13g2_decap_4  FILLER_51_196
timestamp 1679577901
transform 1 0 19968 0 -1 40068
box -48 -56 432 834
use sg13g2_decap_8  FILLER_52_0
timestamp 1679581782
transform 1 0 1152 0 1 40068
box -48 -56 720 834
use sg13g2_fill_1  FILLER_52_7
timestamp 1677579658
transform 1 0 1824 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_44
timestamp 1677580104
transform 1 0 5376 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_46
timestamp 1677579658
transform 1 0 5568 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_67
timestamp 1677580104
transform 1 0 7584 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_79
timestamp 1677579658
transform 1 0 8736 0 1 40068
box -48 -56 144 834
use sg13g2_decap_4  FILLER_52_102
timestamp 1679577901
transform 1 0 10944 0 1 40068
box -48 -56 432 834
use sg13g2_fill_1  FILLER_52_106
timestamp 1677579658
transform 1 0 11328 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_52_124
timestamp 1677580104
transform 1 0 13056 0 1 40068
box -48 -56 240 834
use sg13g2_fill_2  FILLER_52_131
timestamp 1677580104
transform 1 0 13728 0 1 40068
box -48 -56 240 834
use sg13g2_decap_4  FILLER_52_171
timestamp 1679577901
transform 1 0 17568 0 1 40068
box -48 -56 432 834
use sg13g2_fill_2  FILLER_52_175
timestamp 1677580104
transform 1 0 17952 0 1 40068
box -48 -56 240 834
use sg13g2_fill_1  FILLER_52_199
timestamp 1677579658
transform 1 0 20256 0 1 40068
box -48 -56 144 834
use sg13g2_fill_2  FILLER_53_66
timestamp 1677580104
transform 1 0 7488 0 -1 41580
box -48 -56 240 834
use sg13g2_decap_8  FILLER_53_106
timestamp 1679581782
transform 1 0 11328 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_8  FILLER_53_113
timestamp 1679581782
transform 1 0 12000 0 -1 41580
box -48 -56 720 834
use sg13g2_decap_4  FILLER_53_120
timestamp 1679577901
transform 1 0 12672 0 -1 41580
box -48 -56 432 834
use sg13g2_fill_1  FILLER_53_124
timestamp 1677579658
transform 1 0 13056 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_1  FILLER_53_134
timestamp 1677579658
transform 1 0 14016 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_1  FILLER_53_152
timestamp 1677579658
transform 1 0 15744 0 -1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_54_40
timestamp 1677580104
transform 1 0 4992 0 1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_82
timestamp 1677579658
transform 1 0 9024 0 1 41580
box -48 -56 144 834
use sg13g2_fill_2  FILLER_54_147
timestamp 1677580104
transform 1 0 15264 0 1 41580
box -48 -56 240 834
use sg13g2_fill_1  FILLER_54_149
timestamp 1677579658
transform 1 0 15456 0 1 41580
box -48 -56 144 834
use sg13g2_fill_1  FILLER_54_199
timestamp 1677579658
transform 1 0 20256 0 1 41580
box -48 -56 144 834
use sg13g2_decap_8  FILLER_55_0
timestamp 1679581782
transform 1 0 1152 0 -1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_55_7
timestamp 1679581782
transform 1 0 1824 0 -1 43092
box -48 -56 720 834
use sg13g2_fill_2  FILLER_55_14
timestamp 1677580104
transform 1 0 2496 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_40
timestamp 1677580104
transform 1 0 4992 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_59
timestamp 1677579658
transform 1 0 6816 0 -1 43092
box -48 -56 144 834
use sg13g2_decap_4  FILLER_55_103
timestamp 1679577901
transform 1 0 11040 0 -1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_55_141
timestamp 1677580104
transform 1 0 14688 0 -1 43092
box -48 -56 240 834
use sg13g2_decap_8  FILLER_55_147
timestamp 1679581782
transform 1 0 15264 0 -1 43092
box -48 -56 720 834
use sg13g2_fill_1  FILLER_55_154
timestamp 1677579658
transform 1 0 15936 0 -1 43092
box -48 -56 144 834
use sg13g2_fill_1  FILLER_55_159
timestamp 1677579658
transform 1 0 16416 0 -1 43092
box -48 -56 144 834
use sg13g2_fill_2  FILLER_55_164
timestamp 1677580104
transform 1 0 16896 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_170
timestamp 1677580104
transform 1 0 17472 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_180
timestamp 1677580104
transform 1 0 18432 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_182
timestamp 1677579658
transform 1 0 18624 0 -1 43092
box -48 -56 144 834
use sg13g2_fill_2  FILLER_55_187
timestamp 1677580104
transform 1 0 19104 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_2  FILLER_55_197
timestamp 1677580104
transform 1 0 20064 0 -1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_55_199
timestamp 1677579658
transform 1 0 20256 0 -1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_0
timestamp 1679581782
transform 1 0 1152 0 1 43092
box -48 -56 720 834
use sg13g2_fill_2  FILLER_56_7
timestamp 1677580104
transform 1 0 1824 0 1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_9
timestamp 1677579658
transform 1 0 2016 0 1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_32
timestamp 1679581782
transform 1 0 4224 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_39
timestamp 1679581782
transform 1 0 4896 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_46
timestamp 1679581782
transform 1 0 5568 0 1 43092
box -48 -56 720 834
use sg13g2_fill_1  FILLER_56_53
timestamp 1677579658
transform 1 0 6240 0 1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_76
timestamp 1679581782
transform 1 0 8448 0 1 43092
box -48 -56 720 834
use sg13g2_fill_1  FILLER_56_83
timestamp 1677579658
transform 1 0 9120 0 1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_87
timestamp 1679581782
transform 1 0 9504 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_94
timestamp 1679581782
transform 1 0 10176 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_101
timestamp 1679581782
transform 1 0 10848 0 1 43092
box -48 -56 720 834
use sg13g2_fill_1  FILLER_56_108
timestamp 1677579658
transform 1 0 11520 0 1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_113
timestamp 1679581782
transform 1 0 12000 0 1 43092
box -48 -56 720 834
use sg13g2_decap_4  FILLER_56_120
timestamp 1679577901
transform 1 0 12672 0 1 43092
box -48 -56 432 834
use sg13g2_fill_2  FILLER_56_128
timestamp 1677580104
transform 1 0 13440 0 1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_130
timestamp 1677579658
transform 1 0 13632 0 1 43092
box -48 -56 144 834
use sg13g2_decap_8  FILLER_56_148
timestamp 1679581782
transform 1 0 15360 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_155
timestamp 1679581782
transform 1 0 16032 0 1 43092
box -48 -56 720 834
use sg13g2_decap_8  FILLER_56_162
timestamp 1679581782
transform 1 0 16704 0 1 43092
box -48 -56 720 834
use sg13g2_fill_1  FILLER_56_169
timestamp 1677579658
transform 1 0 17376 0 1 43092
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_178
timestamp 1677580104
transform 1 0 18240 0 1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_180
timestamp 1677579658
transform 1 0 18432 0 1 43092
box -48 -56 144 834
use sg13g2_fill_2  FILLER_56_197
timestamp 1677580104
transform 1 0 20064 0 1 43092
box -48 -56 240 834
use sg13g2_fill_1  FILLER_56_199
timestamp 1677579658
transform 1 0 20256 0 1 43092
box -48 -56 144 834
use sg13g2_decap_4  FILLER_57_0
timestamp 1679577901
transform 1 0 1152 0 -1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_57_25
timestamp 1677579658
transform 1 0 3552 0 -1 44604
box -48 -56 144 834
use sg13g2_decap_8  FILLER_57_47
timestamp 1679581782
transform 1 0 5664 0 -1 44604
box -48 -56 720 834
use sg13g2_fill_1  FILLER_57_71
timestamp 1677579658
transform 1 0 7968 0 -1 44604
box -48 -56 144 834
use sg13g2_decap_4  FILLER_57_89
timestamp 1679577901
transform 1 0 9696 0 -1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_57_93
timestamp 1677579658
transform 1 0 10080 0 -1 44604
box -48 -56 144 834
use sg13g2_decap_8  FILLER_57_132
timestamp 1679581782
transform 1 0 13824 0 -1 44604
box -48 -56 720 834
use sg13g2_decap_4  FILLER_57_139
timestamp 1679577901
transform 1 0 14496 0 -1 44604
box -48 -56 432 834
use sg13g2_decap_4  FILLER_57_168
timestamp 1679577901
transform 1 0 17280 0 -1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_57_180
timestamp 1677579658
transform 1 0 18432 0 -1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_57_198
timestamp 1677580104
transform 1 0 20160 0 -1 44604
box -48 -56 240 834
use sg13g2_decap_4  FILLER_58_46
timestamp 1679577901
transform 1 0 5568 0 1 44604
box -48 -56 432 834
use sg13g2_fill_1  FILLER_58_50
timestamp 1677579658
transform 1 0 5952 0 1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_58_89
timestamp 1677580104
transform 1 0 9696 0 1 44604
box -48 -56 240 834
use sg13g2_fill_1  FILLER_58_91
timestamp 1677579658
transform 1 0 9888 0 1 44604
box -48 -56 144 834
use sg13g2_fill_1  FILLER_58_113
timestamp 1677579658
transform 1 0 12000 0 1 44604
box -48 -56 144 834
use sg13g2_decap_8  FILLER_58_131
timestamp 1679581782
transform 1 0 13728 0 1 44604
box -48 -56 720 834
use sg13g2_decap_8  FILLER_58_138
timestamp 1679581782
transform 1 0 14400 0 1 44604
box -48 -56 720 834
use sg13g2_fill_2  FILLER_58_145
timestamp 1677580104
transform 1 0 15072 0 1 44604
box -48 -56 240 834
use sg13g2_decap_8  FILLER_58_168
timestamp 1679581782
transform 1 0 17280 0 1 44604
box -48 -56 720 834
use sg13g2_fill_1  FILLER_58_175
timestamp 1677579658
transform 1 0 17952 0 1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_58_197
timestamp 1677580104
transform 1 0 20064 0 1 44604
box -48 -56 240 834
use sg13g2_fill_1  FILLER_58_199
timestamp 1677579658
transform 1 0 20256 0 1 44604
box -48 -56 144 834
use sg13g2_fill_2  FILLER_59_0
timestamp 1677580104
transform 1 0 1152 0 -1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_2
timestamp 1677579658
transform 1 0 1344 0 -1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_59_19
timestamp 1679581782
transform 1 0 2976 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_26
timestamp 1679581782
transform 1 0 3648 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_50
timestamp 1679581782
transform 1 0 5952 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_57
timestamp 1679581782
transform 1 0 6624 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_64
timestamp 1679581782
transform 1 0 7296 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_71
timestamp 1679581782
transform 1 0 7968 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_112
timestamp 1679581782
transform 1 0 11904 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_59_119
timestamp 1679581782
transform 1 0 12576 0 -1 46116
box -48 -56 720 834
use sg13g2_decap_4  FILLER_59_126
timestamp 1679577901
transform 1 0 13248 0 -1 46116
box -48 -56 432 834
use sg13g2_decap_4  FILLER_59_147
timestamp 1679577901
transform 1 0 15264 0 -1 46116
box -48 -56 432 834
use sg13g2_fill_1  FILLER_59_151
timestamp 1677579658
transform 1 0 15648 0 -1 46116
box -48 -56 144 834
use sg13g2_fill_2  FILLER_59_186
timestamp 1677580104
transform 1 0 19008 0 -1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_188
timestamp 1677579658
transform 1 0 19200 0 -1 46116
box -48 -56 144 834
use sg13g2_fill_2  FILLER_59_197
timestamp 1677580104
transform 1 0 20064 0 -1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_59_199
timestamp 1677579658
transform 1 0 20256 0 -1 46116
box -48 -56 144 834
use sg13g2_decap_4  FILLER_60_25
timestamp 1679577901
transform 1 0 3552 0 1 46116
box -48 -56 432 834
use sg13g2_fill_1  FILLER_60_29
timestamp 1677579658
transform 1 0 3936 0 1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_60_47
timestamp 1679581782
transform 1 0 5664 0 1 46116
box -48 -56 720 834
use sg13g2_decap_8  FILLER_60_92
timestamp 1679581782
transform 1 0 9984 0 1 46116
box -48 -56 720 834
use sg13g2_fill_2  FILLER_60_99
timestamp 1677580104
transform 1 0 10656 0 1 46116
box -48 -56 240 834
use sg13g2_decap_8  FILLER_60_139
timestamp 1679581782
transform 1 0 14496 0 1 46116
box -48 -56 720 834
use sg13g2_decap_4  FILLER_60_146
timestamp 1679577901
transform 1 0 15168 0 1 46116
box -48 -56 432 834
use sg13g2_fill_1  FILLER_60_150
timestamp 1677579658
transform 1 0 15552 0 1 46116
box -48 -56 144 834
use sg13g2_decap_8  FILLER_60_168
timestamp 1679581782
transform 1 0 17280 0 1 46116
box -48 -56 720 834
use sg13g2_fill_2  FILLER_60_175
timestamp 1677580104
transform 1 0 17952 0 1 46116
box -48 -56 240 834
use sg13g2_fill_1  FILLER_60_177
timestamp 1677579658
transform 1 0 18144 0 1 46116
box -48 -56 144 834
use sg13g2_fill_1  FILLER_60_199
timestamp 1677579658
transform 1 0 20256 0 1 46116
box -48 -56 144 834
use sg13g2_fill_2  FILLER_61_0
timestamp 1677580104
transform 1 0 1152 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_1  FILLER_61_2
timestamp 1677579658
transform 1 0 1344 0 -1 47628
box -48 -56 144 834
use sg13g2_fill_2  FILLER_61_24
timestamp 1677580104
transform 1 0 3456 0 -1 47628
box -48 -56 240 834
use sg13g2_decap_4  FILLER_61_47
timestamp 1679577901
transform 1 0 5664 0 -1 47628
box -48 -56 432 834
use sg13g2_decap_4  FILLER_61_72
timestamp 1679577901
transform 1 0 8064 0 -1 47628
box -48 -56 432 834
use sg13g2_fill_1  FILLER_61_93
timestamp 1677579658
transform 1 0 10080 0 -1 47628
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_115
timestamp 1679581782
transform 1 0 12192 0 -1 47628
box -48 -56 720 834
use sg13g2_decap_8  FILLER_61_139
timestamp 1679581782
transform 1 0 14496 0 -1 47628
box -48 -56 720 834
use sg13g2_fill_1  FILLER_61_146
timestamp 1677579658
transform 1 0 15168 0 -1 47628
box -48 -56 144 834
use sg13g2_decap_8  FILLER_61_168
timestamp 1679581782
transform 1 0 17280 0 -1 47628
box -48 -56 720 834
use sg13g2_fill_2  FILLER_61_175
timestamp 1677580104
transform 1 0 17952 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_2  FILLER_61_198
timestamp 1677580104
transform 1 0 20160 0 -1 47628
box -48 -56 240 834
use sg13g2_fill_2  FILLER_62_0
timestamp 1677580104
transform 1 0 1152 0 1 47628
box -48 -56 240 834
use sg13g2_fill_1  FILLER_62_2
timestamp 1677579658
transform 1 0 1344 0 1 47628
box -48 -56 144 834
use sg13g2_fill_1  FILLER_62_36
timestamp 1677579658
transform 1 0 4608 0 1 47628
box -48 -56 144 834
use sg13g2_decap_4  FILLER_62_71
timestamp 1679577901
transform 1 0 7968 0 1 47628
box -48 -56 432 834
use sg13g2_fill_2  FILLER_62_75
timestamp 1677580104
transform 1 0 8352 0 1 47628
box -48 -56 240 834
use sg13g2_decap_4  FILLER_62_98
timestamp 1679577901
transform 1 0 10560 0 1 47628
box -48 -56 432 834
use sg13g2_decap_8  FILLER_62_191
timestamp 1679581782
transform 1 0 19488 0 1 47628
box -48 -56 720 834
use sg13g2_fill_2  FILLER_62_198
timestamp 1677580104
transform 1 0 20160 0 1 47628
box -48 -56 240 834
use sg13g2_fill_2  FILLER_63_0
timestamp 1677580104
transform 1 0 1152 0 -1 49140
box -48 -56 240 834
use sg13g2_fill_1  FILLER_63_2
timestamp 1677579658
transform 1 0 1344 0 -1 49140
box -48 -56 144 834
use sg13g2_fill_2  FILLER_63_11
timestamp 1677580104
transform 1 0 2208 0 -1 49140
box -48 -56 240 834
use sg13g2_fill_1  FILLER_63_13
timestamp 1677579658
transform 1 0 2400 0 -1 49140
box -48 -56 144 834
use sg13g2_fill_1  FILLER_63_69
timestamp 1677579658
transform 1 0 7776 0 -1 49140
box -48 -56 144 834
use sg13g2_fill_1  FILLER_63_97
timestamp 1677579658
transform 1 0 10464 0 -1 49140
box -48 -56 144 834
use sg13g2_decap_8  FILLER_63_115
timestamp 1679581782
transform 1 0 12192 0 -1 49140
box -48 -56 720 834
use sg13g2_fill_2  FILLER_63_122
timestamp 1677580104
transform 1 0 12864 0 -1 49140
box -48 -56 240 834
use sg13g2_decap_8  FILLER_63_141
timestamp 1679581782
transform 1 0 14688 0 -1 49140
box -48 -56 720 834
use sg13g2_decap_4  FILLER_63_169
timestamp 1679577901
transform 1 0 17376 0 -1 49140
box -48 -56 432 834
use sg13g2_fill_1  FILLER_63_173
timestamp 1677579658
transform 1 0 17760 0 -1 49140
box -48 -56 144 834
use sg13g2_decap_4  FILLER_63_195
timestamp 1679577901
transform 1 0 19872 0 -1 49140
box -48 -56 432 834
use sg13g2_fill_1  FILLER_63_199
timestamp 1677579658
transform 1 0 20256 0 -1 49140
box -48 -56 144 834
use sg13g2_decap_8  FILLER_64_0
timestamp 1679581782
transform 1 0 1152 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_7
timestamp 1679581782
transform 1 0 1824 0 1 49140
box -48 -56 720 834
use sg13g2_fill_1  FILLER_64_14
timestamp 1677579658
transform 1 0 2496 0 1 49140
box -48 -56 144 834
use sg13g2_decap_4  FILLER_64_53
timestamp 1679577901
transform 1 0 6240 0 1 49140
box -48 -56 432 834
use sg13g2_decap_8  FILLER_64_159
timestamp 1679581782
transform 1 0 16416 0 1 49140
box -48 -56 720 834
use sg13g2_decap_8  FILLER_64_166
timestamp 1679581782
transform 1 0 17088 0 1 49140
box -48 -56 720 834
use sg13g2_fill_1  FILLER_64_173
timestamp 1677579658
transform 1 0 17760 0 1 49140
box -48 -56 144 834
use sg13g2_decap_4  FILLER_64_195
timestamp 1679577901
transform 1 0 19872 0 1 49140
box -48 -56 432 834
use sg13g2_fill_1  FILLER_64_199
timestamp 1677579658
transform 1 0 20256 0 1 49140
box -48 -56 144 834
use sg13g2_fill_2  FILLER_65_0
timestamp 1677580104
transform 1 0 1152 0 -1 50652
box -48 -56 240 834
use sg13g2_fill_1  FILLER_65_2
timestamp 1677579658
transform 1 0 1344 0 -1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_65_66
timestamp 1677580104
transform 1 0 7488 0 -1 50652
box -48 -56 240 834
use sg13g2_fill_2  FILLER_65_98
timestamp 1677580104
transform 1 0 10560 0 -1 50652
box -48 -56 240 834
use sg13g2_fill_2  FILLER_65_197
timestamp 1677580104
transform 1 0 20064 0 -1 50652
box -48 -56 240 834
use sg13g2_fill_1  FILLER_65_199
timestamp 1677579658
transform 1 0 20256 0 -1 50652
box -48 -56 144 834
use sg13g2_decap_8  FILLER_66_21
timestamp 1679581782
transform 1 0 3168 0 1 50652
box -48 -56 720 834
use sg13g2_decap_4  FILLER_66_49
timestamp 1679577901
transform 1 0 5856 0 1 50652
box -48 -56 432 834
use sg13g2_fill_2  FILLER_66_53
timestamp 1677580104
transform 1 0 6240 0 1 50652
box -48 -56 240 834
use sg13g2_decap_4  FILLER_66_72
timestamp 1679577901
transform 1 0 8064 0 1 50652
box -48 -56 432 834
use sg13g2_fill_2  FILLER_66_93
timestamp 1677580104
transform 1 0 10080 0 1 50652
box -48 -56 240 834
use sg13g2_decap_8  FILLER_66_112
timestamp 1679581782
transform 1 0 11904 0 1 50652
box -48 -56 720 834
use sg13g2_fill_1  FILLER_66_119
timestamp 1677579658
transform 1 0 12576 0 1 50652
box -48 -56 144 834
use sg13g2_fill_1  FILLER_66_137
timestamp 1677579658
transform 1 0 14304 0 1 50652
box -48 -56 144 834
use sg13g2_decap_4  FILLER_66_153
timestamp 1679577901
transform 1 0 15840 0 1 50652
box -48 -56 432 834
use sg13g2_decap_4  FILLER_66_174
timestamp 1679577901
transform 1 0 17856 0 1 50652
box -48 -56 432 834
use sg13g2_fill_1  FILLER_66_199
timestamp 1677579658
transform 1 0 20256 0 1 50652
box -48 -56 144 834
use sg13g2_fill_2  FILLER_67_0
timestamp 1677580104
transform 1 0 1152 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_2
timestamp 1677579658
transform 1 0 1344 0 -1 52164
box -48 -56 144 834
use sg13g2_decap_4  FILLER_67_79
timestamp 1679577901
transform 1 0 8736 0 -1 52164
box -48 -56 432 834
use sg13g2_fill_1  FILLER_67_83
timestamp 1677579658
transform 1 0 9120 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_1  FILLER_67_89
timestamp 1677579658
transform 1 0 9696 0 -1 52164
box -48 -56 144 834
use sg13g2_decap_4  FILLER_67_111
timestamp 1679577901
transform 1 0 11808 0 -1 52164
box -48 -56 432 834
use sg13g2_fill_2  FILLER_67_132
timestamp 1677580104
transform 1 0 13824 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_67_164
timestamp 1677580104
transform 1 0 16896 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_166
timestamp 1677579658
transform 1 0 17088 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_1  FILLER_67_188
timestamp 1677579658
transform 1 0 19200 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_67_197
timestamp 1677580104
transform 1 0 20064 0 -1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_67_199
timestamp 1677579658
transform 1 0 20256 0 -1 52164
box -48 -56 144 834
use sg13g2_fill_2  FILLER_68_0
timestamp 1677580104
transform 1 0 1152 0 1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_2
timestamp 1677579658
transform 1 0 1344 0 1 52164
box -48 -56 144 834
use sg13g2_decap_8  FILLER_68_41
timestamp 1679581782
transform 1 0 5088 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_48
timestamp 1679581782
transform 1 0 5760 0 1 52164
box -48 -56 720 834
use sg13g2_fill_1  FILLER_68_55
timestamp 1677579658
transform 1 0 6432 0 1 52164
box -48 -56 144 834
use sg13g2_decap_8  FILLER_68_94
timestamp 1679581782
transform 1 0 10176 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_101
timestamp 1679581782
transform 1 0 10848 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_108
timestamp 1679581782
transform 1 0 11520 0 1 52164
box -48 -56 720 834
use sg13g2_decap_8  FILLER_68_115
timestamp 1679581782
transform 1 0 12192 0 1 52164
box -48 -56 720 834
use sg13g2_fill_2  FILLER_68_139
timestamp 1677580104
transform 1 0 14496 0 1 52164
box -48 -56 240 834
use sg13g2_fill_2  FILLER_68_197
timestamp 1677580104
transform 1 0 20064 0 1 52164
box -48 -56 240 834
use sg13g2_fill_1  FILLER_68_199
timestamp 1677579658
transform 1 0 20256 0 1 52164
box -48 -56 144 834
use sg13g2_fill_1  FILLER_69_0
timestamp 1677579658
transform 1 0 1152 0 -1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_69_26
timestamp 1677580104
transform 1 0 3648 0 -1 53676
box -48 -56 240 834
use sg13g2_decap_8  FILLER_69_49
timestamp 1679581782
transform 1 0 5856 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_56
timestamp 1679581782
transform 1 0 6528 0 -1 53676
box -48 -56 720 834
use sg13g2_decap_8  FILLER_69_63
timestamp 1679581782
transform 1 0 7200 0 -1 53676
box -48 -56 720 834
use sg13g2_fill_2  FILLER_69_70
timestamp 1677580104
transform 1 0 7872 0 -1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_69_72
timestamp 1677579658
transform 1 0 8064 0 -1 53676
box -48 -56 144 834
use sg13g2_fill_1  FILLER_69_128
timestamp 1677579658
transform 1 0 13440 0 -1 53676
box -48 -56 144 834
use sg13g2_decap_8  FILLER_69_170
timestamp 1679581782
transform 1 0 17472 0 -1 53676
box -48 -56 720 834
use sg13g2_fill_1  FILLER_69_177
timestamp 1677579658
transform 1 0 18144 0 -1 53676
box -48 -56 144 834
use sg13g2_fill_1  FILLER_69_199
timestamp 1677579658
transform 1 0 20256 0 -1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_0
timestamp 1677580104
transform 1 0 1152 0 1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_2
timestamp 1677579658
transform 1 0 1344 0 1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_11
timestamp 1677580104
transform 1 0 2208 0 1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_13
timestamp 1677579658
transform 1 0 2400 0 1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_70_31
timestamp 1677580104
transform 1 0 4128 0 1 53676
box -48 -56 240 834
use sg13g2_fill_2  FILLER_70_50
timestamp 1677580104
transform 1 0 5952 0 1 53676
box -48 -56 240 834
use sg13g2_fill_1  FILLER_70_52
timestamp 1677579658
transform 1 0 6144 0 1 53676
box -48 -56 144 834
use sg13g2_decap_8  FILLER_70_91
timestamp 1679581782
transform 1 0 9888 0 1 53676
box -48 -56 720 834
use sg13g2_decap_4  FILLER_70_98
timestamp 1679577901
transform 1 0 10560 0 1 53676
box -48 -56 432 834
use sg13g2_fill_2  FILLER_70_102
timestamp 1677580104
transform 1 0 10944 0 1 53676
box -48 -56 240 834
use sg13g2_decap_8  FILLER_70_159
timestamp 1679581782
transform 1 0 16416 0 1 53676
box -48 -56 720 834
use sg13g2_decap_4  FILLER_70_166
timestamp 1679577901
transform 1 0 17088 0 1 53676
box -48 -56 432 834
use sg13g2_fill_1  FILLER_70_170
timestamp 1677579658
transform 1 0 17472 0 1 53676
box -48 -56 144 834
use sg13g2_fill_2  FILLER_71_0
timestamp 1677580104
transform 1 0 1152 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_2
timestamp 1677579658
transform 1 0 1344 0 -1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_71_11
timestamp 1677580104
transform 1 0 2208 0 -1 55188
box -48 -56 240 834
use sg13g2_decap_8  FILLER_71_34
timestamp 1679581782
transform 1 0 4416 0 -1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_71_41
timestamp 1679581782
transform 1 0 5088 0 -1 55188
box -48 -56 720 834
use sg13g2_fill_1  FILLER_71_48
timestamp 1677579658
transform 1 0 5760 0 -1 55188
box -48 -56 144 834
use sg13g2_decap_4  FILLER_71_70
timestamp 1679577901
transform 1 0 7872 0 -1 55188
box -48 -56 432 834
use sg13g2_fill_1  FILLER_71_74
timestamp 1677579658
transform 1 0 8256 0 -1 55188
box -48 -56 144 834
use sg13g2_fill_1  FILLER_71_109
timestamp 1677579658
transform 1 0 11616 0 -1 55188
box -48 -56 144 834
use sg13g2_decap_4  FILLER_71_131
timestamp 1679577901
transform 1 0 13728 0 -1 55188
box -48 -56 432 834
use sg13g2_fill_1  FILLER_71_135
timestamp 1677579658
transform 1 0 14112 0 -1 55188
box -48 -56 144 834
use sg13g2_decap_4  FILLER_71_167
timestamp 1679577901
transform 1 0 17184 0 -1 55188
box -48 -56 432 834
use sg13g2_fill_1  FILLER_71_171
timestamp 1677579658
transform 1 0 17568 0 -1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_71_197
timestamp 1677580104
transform 1 0 20064 0 -1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_71_199
timestamp 1677579658
transform 1 0 20256 0 -1 55188
box -48 -56 144 834
use sg13g2_decap_8  FILLER_72_25
timestamp 1679581782
transform 1 0 3552 0 1 55188
box -48 -56 720 834
use sg13g2_decap_4  FILLER_72_32
timestamp 1679577901
transform 1 0 4224 0 1 55188
box -48 -56 432 834
use sg13g2_fill_2  FILLER_72_53
timestamp 1677580104
transform 1 0 6240 0 1 55188
box -48 -56 240 834
use sg13g2_decap_8  FILLER_72_93
timestamp 1679581782
transform 1 0 10080 0 1 55188
box -48 -56 720 834
use sg13g2_decap_4  FILLER_72_100
timestamp 1679577901
transform 1 0 10752 0 1 55188
box -48 -56 432 834
use sg13g2_fill_2  FILLER_72_104
timestamp 1677580104
transform 1 0 11136 0 1 55188
box -48 -56 240 834
use sg13g2_decap_8  FILLER_72_131
timestamp 1679581782
transform 1 0 13728 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_138
timestamp 1679581782
transform 1 0 14400 0 1 55188
box -48 -56 720 834
use sg13g2_decap_8  FILLER_72_145
timestamp 1679581782
transform 1 0 15072 0 1 55188
box -48 -56 720 834
use sg13g2_fill_2  FILLER_72_186
timestamp 1677580104
transform 1 0 19008 0 1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_188
timestamp 1677579658
transform 1 0 19200 0 1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_72_197
timestamp 1677580104
transform 1 0 20064 0 1 55188
box -48 -56 240 834
use sg13g2_fill_1  FILLER_72_199
timestamp 1677579658
transform 1 0 20256 0 1 55188
box -48 -56 144 834
use sg13g2_fill_2  FILLER_73_21
timestamp 1677580104
transform 1 0 3168 0 -1 56700
box -48 -56 240 834
use sg13g2_fill_1  FILLER_73_23
timestamp 1677579658
transform 1 0 3360 0 -1 56700
box -48 -56 144 834
use sg13g2_decap_4  FILLER_73_45
timestamp 1679577901
transform 1 0 5472 0 -1 56700
box -48 -56 432 834
use sg13g2_fill_1  FILLER_73_49
timestamp 1677579658
transform 1 0 5856 0 -1 56700
box -48 -56 144 834
use sg13g2_decap_8  FILLER_73_67
timestamp 1679581782
transform 1 0 7584 0 -1 56700
box -48 -56 720 834
use sg13g2_fill_2  FILLER_73_74
timestamp 1677580104
transform 1 0 8256 0 -1 56700
box -48 -56 240 834
use sg13g2_fill_2  FILLER_73_114
timestamp 1677580104
transform 1 0 12096 0 -1 56700
box -48 -56 240 834
use sg13g2_decap_8  FILLER_73_133
timestamp 1679581782
transform 1 0 13920 0 -1 56700
box -48 -56 720 834
use sg13g2_decap_4  FILLER_73_140
timestamp 1679577901
transform 1 0 14592 0 -1 56700
box -48 -56 432 834
use sg13g2_fill_1  FILLER_73_144
timestamp 1677579658
transform 1 0 14976 0 -1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_73_175
timestamp 1677579658
transform 1 0 17952 0 -1 56700
box -48 -56 144 834
use sg13g2_fill_2  FILLER_73_197
timestamp 1677580104
transform 1 0 20064 0 -1 56700
box -48 -56 240 834
use sg13g2_fill_1  FILLER_73_199
timestamp 1677579658
transform 1 0 20256 0 -1 56700
box -48 -56 144 834
use sg13g2_fill_2  FILLER_74_0
timestamp 1677580104
transform 1 0 1152 0 1 56700
box -48 -56 240 834
use sg13g2_fill_1  FILLER_74_2
timestamp 1677579658
transform 1 0 1344 0 1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_74_11
timestamp 1677579658
transform 1 0 2208 0 1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_74_50
timestamp 1677579658
transform 1 0 5952 0 1 56700
box -48 -56 144 834
use sg13g2_fill_2  FILLER_74_148
timestamp 1677580104
transform 1 0 15360 0 1 56700
box -48 -56 240 834
use sg13g2_fill_2  FILLER_74_197
timestamp 1677580104
transform 1 0 20064 0 1 56700
box -48 -56 240 834
use sg13g2_fill_1  FILLER_74_199
timestamp 1677579658
transform 1 0 20256 0 1 56700
box -48 -56 144 834
use sg13g2_fill_1  FILLER_75_0
timestamp 1677579658
transform 1 0 1152 0 -1 58212
box -48 -56 144 834
use sg13g2_fill_1  FILLER_75_22
timestamp 1677579658
transform 1 0 3264 0 -1 58212
box -48 -56 144 834
use sg13g2_decap_8  FILLER_75_44
timestamp 1679581782
transform 1 0 5376 0 -1 58212
box -48 -56 720 834
use sg13g2_fill_1  FILLER_75_51
timestamp 1677579658
transform 1 0 6048 0 -1 58212
box -48 -56 144 834
use sg13g2_fill_2  FILLER_75_90
timestamp 1677580104
transform 1 0 9792 0 -1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_75_92
timestamp 1677579658
transform 1 0 9984 0 -1 58212
box -48 -56 144 834
use sg13g2_fill_1  FILLER_75_110
timestamp 1677579658
transform 1 0 11712 0 -1 58212
box -48 -56 144 834
use sg13g2_decap_4  FILLER_75_128
timestamp 1679577901
transform 1 0 13440 0 -1 58212
box -48 -56 432 834
use sg13g2_fill_2  FILLER_75_132
timestamp 1677580104
transform 1 0 13824 0 -1 58212
box -48 -56 240 834
use sg13g2_fill_2  FILLER_75_198
timestamp 1677580104
transform 1 0 20160 0 -1 58212
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_0
timestamp 1677580104
transform 1 0 1152 0 1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_76_70
timestamp 1677579658
transform 1 0 7872 0 1 58212
box -48 -56 144 834
use sg13g2_decap_8  FILLER_76_109
timestamp 1679581782
transform 1 0 11616 0 1 58212
box -48 -56 720 834
use sg13g2_decap_4  FILLER_76_116
timestamp 1679577901
transform 1 0 12288 0 1 58212
box -48 -56 432 834
use sg13g2_decap_4  FILLER_76_124
timestamp 1679577901
transform 1 0 13056 0 1 58212
box -48 -56 432 834
use sg13g2_fill_2  FILLER_76_128
timestamp 1677580104
transform 1 0 13440 0 1 58212
box -48 -56 240 834
use sg13g2_fill_2  FILLER_76_164
timestamp 1677580104
transform 1 0 16896 0 1 58212
box -48 -56 240 834
use sg13g2_fill_1  FILLER_76_166
timestamp 1677579658
transform 1 0 17088 0 1 58212
box -48 -56 144 834
use sg13g2_fill_1  FILLER_77_17
timestamp 1677579658
transform 1 0 2784 0 -1 59724
box -48 -56 144 834
use sg13g2_decap_8  FILLER_77_43
timestamp 1679581782
transform 1 0 5280 0 -1 59724
box -48 -56 720 834
use sg13g2_fill_2  FILLER_77_50
timestamp 1677580104
transform 1 0 5952 0 -1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_73
timestamp 1677579658
transform 1 0 8160 0 -1 59724
box -48 -56 144 834
use sg13g2_decap_4  FILLER_77_112
timestamp 1679577901
transform 1 0 11904 0 -1 59724
box -48 -56 432 834
use sg13g2_fill_2  FILLER_77_116
timestamp 1677580104
transform 1 0 12288 0 -1 59724
box -48 -56 240 834
use sg13g2_decap_4  FILLER_77_160
timestamp 1679577901
transform 1 0 16512 0 -1 59724
box -48 -56 432 834
use sg13g2_fill_2  FILLER_77_197
timestamp 1677580104
transform 1 0 20064 0 -1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_77_199
timestamp 1677579658
transform 1 0 20256 0 -1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_78_0
timestamp 1677580104
transform 1 0 1152 0 1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_78_2
timestamp 1677579658
transform 1 0 1344 0 1 59724
box -48 -56 144 834
use sg13g2_decap_8  FILLER_78_41
timestamp 1679581782
transform 1 0 5088 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_48
timestamp 1679581782
transform 1 0 5760 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_76
timestamp 1679581782
transform 1 0 8448 0 1 59724
box -48 -56 720 834
use sg13g2_decap_8  FILLER_78_83
timestamp 1679581782
transform 1 0 9120 0 1 59724
box -48 -56 720 834
use sg13g2_decap_4  FILLER_78_90
timestamp 1679577901
transform 1 0 9792 0 1 59724
box -48 -56 432 834
use sg13g2_fill_2  FILLER_78_94
timestamp 1677580104
transform 1 0 10176 0 1 59724
box -48 -56 240 834
use sg13g2_fill_2  FILLER_78_117
timestamp 1677580104
transform 1 0 12384 0 1 59724
box -48 -56 240 834
use sg13g2_fill_2  FILLER_78_157
timestamp 1677580104
transform 1 0 16224 0 1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_78_159
timestamp 1677579658
transform 1 0 16416 0 1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_78_197
timestamp 1677580104
transform 1 0 20064 0 1 59724
box -48 -56 240 834
use sg13g2_fill_1  FILLER_78_199
timestamp 1677579658
transform 1 0 20256 0 1 59724
box -48 -56 144 834
use sg13g2_fill_2  FILLER_79_0
timestamp 1677580104
transform 1 0 1152 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_2
timestamp 1677579658
transform 1 0 1344 0 -1 61236
box -48 -56 144 834
use sg13g2_fill_1  FILLER_79_58
timestamp 1677579658
transform 1 0 6720 0 -1 61236
box -48 -56 144 834
use sg13g2_fill_2  FILLER_79_76
timestamp 1677580104
transform 1 0 8448 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_78
timestamp 1677579658
transform 1 0 8640 0 -1 61236
box -48 -56 144 834
use sg13g2_decap_4  FILLER_79_117
timestamp 1679577901
transform 1 0 12384 0 -1 61236
box -48 -56 432 834
use sg13g2_decap_4  FILLER_79_151
timestamp 1679577901
transform 1 0 15648 0 -1 61236
box -48 -56 432 834
use sg13g2_fill_2  FILLER_79_155
timestamp 1677580104
transform 1 0 16032 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_2  FILLER_79_174
timestamp 1677580104
transform 1 0 17856 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_2  FILLER_79_193
timestamp 1677580104
transform 1 0 19680 0 -1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_79_195
timestamp 1677579658
transform 1 0 19872 0 -1 61236
box -48 -56 144 834
use sg13g2_fill_1  FILLER_80_0
timestamp 1677579658
transform 1 0 1152 0 1 61236
box -48 -56 144 834
use sg13g2_decap_8  FILLER_80_39
timestamp 1679581782
transform 1 0 4896 0 1 61236
box -48 -56 720 834
use sg13g2_decap_8  FILLER_80_46
timestamp 1679581782
transform 1 0 5568 0 1 61236
box -48 -56 720 834
use sg13g2_fill_2  FILLER_80_53
timestamp 1677580104
transform 1 0 6240 0 1 61236
box -48 -56 240 834
use sg13g2_decap_8  FILLER_80_72
timestamp 1679581782
transform 1 0 8064 0 1 61236
box -48 -56 720 834
use sg13g2_fill_1  FILLER_80_79
timestamp 1677579658
transform 1 0 8736 0 1 61236
box -48 -56 144 834
use sg13g2_decap_4  FILLER_80_97
timestamp 1679577901
transform 1 0 10464 0 1 61236
box -48 -56 432 834
use sg13g2_fill_1  FILLER_80_101
timestamp 1677579658
transform 1 0 10848 0 1 61236
box -48 -56 144 834
use sg13g2_decap_4  FILLER_80_119
timestamp 1679577901
transform 1 0 12576 0 1 61236
box -48 -56 432 834
use sg13g2_fill_2  FILLER_80_123
timestamp 1677580104
transform 1 0 12960 0 1 61236
box -48 -56 240 834
use sg13g2_decap_8  FILLER_80_146
timestamp 1679581782
transform 1 0 15168 0 1 61236
box -48 -56 720 834
use sg13g2_fill_2  FILLER_80_174
timestamp 1677580104
transform 1 0 17856 0 1 61236
box -48 -56 240 834
use sg13g2_fill_2  FILLER_80_197
timestamp 1677580104
transform 1 0 20064 0 1 61236
box -48 -56 240 834
use sg13g2_fill_1  FILLER_80_199
timestamp 1677579658
transform 1 0 20256 0 1 61236
box -48 -56 144 834
use sg13g2_fill_1  FILLER_81_0
timestamp 1677579658
transform 1 0 1152 0 -1 62748
box -48 -56 144 834
use sg13g2_fill_2  FILLER_81_18
timestamp 1677580104
transform 1 0 2880 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_81_20
timestamp 1677579658
transform 1 0 3072 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_42
timestamp 1679581782
transform 1 0 5184 0 -1 62748
box -48 -56 720 834
use sg13g2_decap_4  FILLER_81_49
timestamp 1679577901
transform 1 0 5856 0 -1 62748
box -48 -56 432 834
use sg13g2_fill_2  FILLER_81_53
timestamp 1677580104
transform 1 0 6240 0 -1 62748
box -48 -56 240 834
use sg13g2_decap_8  FILLER_81_93
timestamp 1679581782
transform 1 0 10080 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_81_100
timestamp 1677580104
transform 1 0 10752 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_81_102
timestamp 1677579658
transform 1 0 10944 0 -1 62748
box -48 -56 144 834
use sg13g2_fill_2  FILLER_81_120
timestamp 1677580104
transform 1 0 12672 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_81_122
timestamp 1677579658
transform 1 0 12864 0 -1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_81_127
timestamp 1679581782
transform 1 0 13344 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_81_134
timestamp 1677580104
transform 1 0 14016 0 -1 62748
box -48 -56 240 834
use sg13g2_decap_4  FILLER_81_157
timestamp 1679577901
transform 1 0 16224 0 -1 62748
box -48 -56 432 834
use sg13g2_decap_8  FILLER_81_165
timestamp 1679581782
transform 1 0 16992 0 -1 62748
box -48 -56 720 834
use sg13g2_fill_1  FILLER_81_172
timestamp 1677579658
transform 1 0 17664 0 -1 62748
box -48 -56 144 834
use sg13g2_fill_2  FILLER_81_198
timestamp 1677580104
transform 1 0 20160 0 -1 62748
box -48 -56 240 834
use sg13g2_fill_2  FILLER_82_0
timestamp 1677580104
transform 1 0 1152 0 1 62748
box -48 -56 240 834
use sg13g2_fill_1  FILLER_82_2
timestamp 1677579658
transform 1 0 1344 0 1 62748
box -48 -56 144 834
use sg13g2_fill_1  FILLER_82_70
timestamp 1677579658
transform 1 0 7872 0 1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_82_130
timestamp 1679581782
transform 1 0 13632 0 1 62748
box -48 -56 720 834
use sg13g2_decap_4  FILLER_82_137
timestamp 1679577901
transform 1 0 14304 0 1 62748
box -48 -56 432 834
use sg13g2_fill_1  FILLER_82_141
timestamp 1677579658
transform 1 0 14688 0 1 62748
box -48 -56 144 834
use sg13g2_decap_8  FILLER_82_159
timestamp 1679581782
transform 1 0 16416 0 1 62748
box -48 -56 720 834
use sg13g2_decap_8  FILLER_82_166
timestamp 1679581782
transform 1 0 17088 0 1 62748
box -48 -56 720 834
use sg13g2_fill_2  FILLER_82_198
timestamp 1677580104
transform 1 0 20160 0 1 62748
box -48 -56 240 834
use sg13g2_fill_2  FILLER_83_0
timestamp 1677580104
transform 1 0 1152 0 -1 64260
box -48 -56 240 834
use sg13g2_decap_8  FILLER_83_19
timestamp 1679581782
transform 1 0 2976 0 -1 64260
box -48 -56 720 834
use sg13g2_fill_1  FILLER_83_26
timestamp 1677579658
transform 1 0 3648 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_4  FILLER_83_44
timestamp 1679577901
transform 1 0 5376 0 -1 64260
box -48 -56 432 834
use sg13g2_fill_2  FILLER_83_48
timestamp 1677580104
transform 1 0 5760 0 -1 64260
box -48 -56 240 834
use sg13g2_decap_4  FILLER_83_67
timestamp 1679577901
transform 1 0 7584 0 -1 64260
box -48 -56 432 834
use sg13g2_fill_2  FILLER_83_71
timestamp 1677580104
transform 1 0 7968 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_2  FILLER_83_112
timestamp 1677580104
transform 1 0 11904 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_114
timestamp 1677579658
transform 1 0 12096 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_4  FILLER_83_153
timestamp 1679577901
transform 1 0 15840 0 -1 64260
box -48 -56 432 834
use sg13g2_fill_2  FILLER_83_191
timestamp 1677580104
transform 1 0 19488 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_2  FILLER_83_197
timestamp 1677580104
transform 1 0 20064 0 -1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_83_199
timestamp 1677579658
transform 1 0 20256 0 -1 64260
box -48 -56 144 834
use sg13g2_decap_8  FILLER_84_0
timestamp 1679581782
transform 1 0 1152 0 1 64260
box -48 -56 720 834
use sg13g2_fill_1  FILLER_84_7
timestamp 1677579658
transform 1 0 1824 0 1 64260
box -48 -56 144 834
use sg13g2_fill_2  FILLER_84_67
timestamp 1677580104
transform 1 0 7584 0 1 64260
box -48 -56 240 834
use sg13g2_fill_1  FILLER_84_97
timestamp 1677579658
transform 1 0 10464 0 1 64260
box -48 -56 144 834
use sg13g2_decap_4  FILLER_84_115
timestamp 1679577901
transform 1 0 12192 0 1 64260
box -48 -56 432 834
use sg13g2_fill_2  FILLER_84_136
timestamp 1677580104
transform 1 0 14208 0 1 64260
box -48 -56 240 834
use sg13g2_decap_8  FILLER_84_155
timestamp 1679581782
transform 1 0 16032 0 1 64260
box -48 -56 720 834
use sg13g2_decap_8  FILLER_84_162
timestamp 1679581782
transform 1 0 16704 0 1 64260
box -48 -56 720 834
use sg13g2_decap_4  FILLER_84_190
timestamp 1679577901
transform 1 0 19392 0 1 64260
box -48 -56 432 834
use sg13g2_fill_2  FILLER_84_198
timestamp 1677580104
transform 1 0 20160 0 1 64260
box -48 -56 240 834
use sg13g2_decap_8  FILLER_85_0
timestamp 1679581782
transform 1 0 1152 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_85_7
timestamp 1679581782
transform 1 0 1824 0 -1 65772
box -48 -56 720 834
use sg13g2_fill_2  FILLER_85_14
timestamp 1677580104
transform 1 0 2496 0 -1 65772
box -48 -56 240 834
use sg13g2_decap_8  FILLER_85_37
timestamp 1679581782
transform 1 0 4704 0 -1 65772
box -48 -56 720 834
use sg13g2_fill_2  FILLER_85_44
timestamp 1677580104
transform 1 0 5376 0 -1 65772
box -48 -56 240 834
use sg13g2_decap_8  FILLER_85_123
timestamp 1679581782
transform 1 0 12960 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_4  FILLER_85_130
timestamp 1679577901
transform 1 0 13632 0 -1 65772
box -48 -56 432 834
use sg13g2_fill_1  FILLER_85_134
timestamp 1677579658
transform 1 0 14016 0 -1 65772
box -48 -56 144 834
use sg13g2_fill_2  FILLER_85_156
timestamp 1677580104
transform 1 0 16128 0 -1 65772
box -48 -56 240 834
use sg13g2_fill_1  FILLER_85_158
timestamp 1677579658
transform 1 0 16320 0 -1 65772
box -48 -56 144 834
use sg13g2_decap_4  FILLER_85_163
timestamp 1679577901
transform 1 0 16800 0 -1 65772
box -48 -56 432 834
use sg13g2_fill_1  FILLER_85_167
timestamp 1677579658
transform 1 0 17184 0 -1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_85_189
timestamp 1679581782
transform 1 0 19296 0 -1 65772
box -48 -56 720 834
use sg13g2_decap_4  FILLER_85_196
timestamp 1679577901
transform 1 0 19968 0 -1 65772
box -48 -56 432 834
use sg13g2_fill_2  FILLER_86_0
timestamp 1677580104
transform 1 0 1152 0 1 65772
box -48 -56 240 834
use sg13g2_fill_2  FILLER_86_19
timestamp 1677580104
transform 1 0 2976 0 1 65772
box -48 -56 240 834
use sg13g2_fill_1  FILLER_86_21
timestamp 1677579658
transform 1 0 3168 0 1 65772
box -48 -56 144 834
use sg13g2_fill_1  FILLER_86_39
timestamp 1677579658
transform 1 0 4896 0 1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_86_70
timestamp 1679581782
transform 1 0 7872 0 1 65772
box -48 -56 720 834
use sg13g2_fill_1  FILLER_86_77
timestamp 1677579658
transform 1 0 8544 0 1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_86_86
timestamp 1679581782
transform 1 0 9408 0 1 65772
box -48 -56 720 834
use sg13g2_decap_8  FILLER_86_93
timestamp 1679581782
transform 1 0 10080 0 1 65772
box -48 -56 720 834
use sg13g2_decap_4  FILLER_86_100
timestamp 1679577901
transform 1 0 10752 0 1 65772
box -48 -56 432 834
use sg13g2_decap_4  FILLER_86_155
timestamp 1679577901
transform 1 0 16032 0 1 65772
box -48 -56 432 834
use sg13g2_fill_2  FILLER_86_159
timestamp 1677580104
transform 1 0 16416 0 1 65772
box -48 -56 240 834
use sg13g2_decap_4  FILLER_86_195
timestamp 1679577901
transform 1 0 19872 0 1 65772
box -48 -56 432 834
use sg13g2_fill_1  FILLER_86_199
timestamp 1677579658
transform 1 0 20256 0 1 65772
box -48 -56 144 834
use sg13g2_decap_8  FILLER_87_0
timestamp 1679581782
transform 1 0 1152 0 -1 67284
box -48 -56 720 834
use sg13g2_decap_4  FILLER_87_7
timestamp 1679577901
transform 1 0 1824 0 -1 67284
box -48 -56 432 834
use sg13g2_fill_1  FILLER_87_11
timestamp 1677579658
transform 1 0 2208 0 -1 67284
box -48 -56 144 834
use sg13g2_decap_8  FILLER_87_33
timestamp 1679581782
transform 1 0 4320 0 -1 67284
box -48 -56 720 834
use sg13g2_fill_1  FILLER_87_40
timestamp 1677579658
transform 1 0 4992 0 -1 67284
box -48 -56 144 834
use sg13g2_fill_1  FILLER_87_58
timestamp 1677579658
transform 1 0 6720 0 -1 67284
box -48 -56 144 834
use sg13g2_decap_8  FILLER_87_127
timestamp 1679581782
transform 1 0 13344 0 -1 67284
box -48 -56 720 834
use sg13g2_fill_2  FILLER_87_134
timestamp 1677580104
transform 1 0 14016 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_2  FILLER_87_157
timestamp 1677580104
transform 1 0 16224 0 -1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_87_159
timestamp 1677579658
transform 1 0 16416 0 -1 67284
box -48 -56 144 834
use sg13g2_decap_4  FILLER_87_194
timestamp 1679577901
transform 1 0 19776 0 -1 67284
box -48 -56 432 834
use sg13g2_fill_2  FILLER_87_198
timestamp 1677580104
transform 1 0 20160 0 -1 67284
box -48 -56 240 834
use sg13g2_decap_4  FILLER_88_0
timestamp 1679577901
transform 1 0 1152 0 1 67284
box -48 -56 432 834
use sg13g2_fill_2  FILLER_88_4
timestamp 1677580104
transform 1 0 1536 0 1 67284
box -48 -56 240 834
use sg13g2_decap_8  FILLER_88_23
timestamp 1679581782
transform 1 0 3360 0 1 67284
box -48 -56 720 834
use sg13g2_decap_4  FILLER_88_30
timestamp 1679577901
transform 1 0 4032 0 1 67284
box -48 -56 432 834
use sg13g2_fill_1  FILLER_88_34
timestamp 1677579658
transform 1 0 4416 0 1 67284
box -48 -56 144 834
use sg13g2_decap_8  FILLER_88_56
timestamp 1679581782
transform 1 0 6528 0 1 67284
box -48 -56 720 834
use sg13g2_fill_1  FILLER_88_63
timestamp 1677579658
transform 1 0 7200 0 1 67284
box -48 -56 144 834
use sg13g2_decap_4  FILLER_88_100
timestamp 1679577901
transform 1 0 10752 0 1 67284
box -48 -56 432 834
use sg13g2_fill_2  FILLER_88_104
timestamp 1677580104
transform 1 0 11136 0 1 67284
box -48 -56 240 834
use sg13g2_decap_8  FILLER_88_144
timestamp 1679581782
transform 1 0 14976 0 1 67284
box -48 -56 720 834
use sg13g2_fill_2  FILLER_88_151
timestamp 1677580104
transform 1 0 15648 0 1 67284
box -48 -56 240 834
use sg13g2_fill_2  FILLER_88_170
timestamp 1677580104
transform 1 0 17472 0 1 67284
box -48 -56 240 834
use sg13g2_fill_1  FILLER_88_172
timestamp 1677579658
transform 1 0 17664 0 1 67284
box -48 -56 144 834
use sg13g2_decap_4  FILLER_88_194
timestamp 1679577901
transform 1 0 19776 0 1 67284
box -48 -56 432 834
use sg13g2_fill_2  FILLER_88_198
timestamp 1677580104
transform 1 0 20160 0 1 67284
box -48 -56 240 834
use sg13g2_decap_4  FILLER_89_0
timestamp 1679577901
transform 1 0 1152 0 -1 68796
box -48 -56 432 834
use sg13g2_decap_8  FILLER_89_25
timestamp 1679581782
transform 1 0 3552 0 -1 68796
box -48 -56 720 834
use sg13g2_decap_4  FILLER_89_32
timestamp 1679577901
transform 1 0 4224 0 -1 68796
box -48 -56 432 834
use sg13g2_fill_1  FILLER_89_36
timestamp 1677579658
transform 1 0 4608 0 -1 68796
box -48 -56 144 834
use sg13g2_fill_1  FILLER_89_54
timestamp 1677579658
transform 1 0 6336 0 -1 68796
box -48 -56 144 834
use sg13g2_decap_4  FILLER_89_110
timestamp 1679577901
transform 1 0 11712 0 -1 68796
box -48 -56 432 834
use sg13g2_fill_2  FILLER_89_114
timestamp 1677580104
transform 1 0 12096 0 -1 68796
box -48 -56 240 834
use sg13g2_fill_2  FILLER_89_150
timestamp 1677580104
transform 1 0 15552 0 -1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_89_152
timestamp 1677579658
transform 1 0 15744 0 -1 68796
box -48 -56 144 834
use sg13g2_decap_8  FILLER_89_170
timestamp 1679581782
transform 1 0 17472 0 -1 68796
box -48 -56 720 834
use sg13g2_fill_2  FILLER_89_177
timestamp 1677580104
transform 1 0 18144 0 -1 68796
box -48 -56 240 834
use sg13g2_decap_4  FILLER_89_196
timestamp 1679577901
transform 1 0 19968 0 -1 68796
box -48 -56 432 834
use sg13g2_fill_1  FILLER_90_51
timestamp 1677579658
transform 1 0 6048 0 1 68796
box -48 -56 144 834
use sg13g2_decap_4  FILLER_90_69
timestamp 1679577901
transform 1 0 7776 0 1 68796
box -48 -56 432 834
use sg13g2_fill_2  FILLER_90_73
timestamp 1677580104
transform 1 0 8160 0 1 68796
box -48 -56 240 834
use sg13g2_fill_2  FILLER_90_84
timestamp 1677580104
transform 1 0 9216 0 1 68796
box -48 -56 240 834
use sg13g2_fill_1  FILLER_90_86
timestamp 1677579658
transform 1 0 9408 0 1 68796
box -48 -56 144 834
use sg13g2_decap_4  FILLER_90_121
timestamp 1679577901
transform 1 0 12768 0 1 68796
box -48 -56 432 834
use sg13g2_decap_8  FILLER_90_163
timestamp 1679581782
transform 1 0 16800 0 1 68796
box -48 -56 720 834
use sg13g2_decap_8  FILLER_90_170
timestamp 1679581782
transform 1 0 17472 0 1 68796
box -48 -56 720 834
use sg13g2_fill_2  FILLER_90_198
timestamp 1677580104
transform 1 0 20160 0 1 68796
box -48 -56 240 834
use sg13g2_decap_4  FILLER_91_17
timestamp 1679577901
transform 1 0 2784 0 -1 70308
box -48 -56 432 834
use sg13g2_fill_1  FILLER_91_21
timestamp 1677579658
transform 1 0 3168 0 -1 70308
box -48 -56 144 834
use sg13g2_decap_8  FILLER_91_43
timestamp 1679581782
transform 1 0 5280 0 -1 70308
box -48 -56 720 834
use sg13g2_fill_1  FILLER_91_50
timestamp 1677579658
transform 1 0 5952 0 -1 70308
box -48 -56 144 834
use sg13g2_decap_4  FILLER_91_72
timestamp 1679577901
transform 1 0 8064 0 -1 70308
box -48 -56 432 834
use sg13g2_fill_2  FILLER_91_76
timestamp 1677580104
transform 1 0 8448 0 -1 70308
box -48 -56 240 834
use sg13g2_decap_8  FILLER_91_95
timestamp 1679581782
transform 1 0 10272 0 -1 70308
box -48 -56 720 834
use sg13g2_fill_2  FILLER_91_123
timestamp 1677580104
transform 1 0 12960 0 -1 70308
box -48 -56 240 834
use sg13g2_decap_8  FILLER_91_163
timestamp 1679581782
transform 1 0 16800 0 -1 70308
box -48 -56 720 834
use sg13g2_decap_4  FILLER_91_170
timestamp 1679577901
transform 1 0 17472 0 -1 70308
box -48 -56 432 834
use sg13g2_fill_2  FILLER_91_174
timestamp 1677580104
transform 1 0 17856 0 -1 70308
box -48 -56 240 834
use sg13g2_fill_2  FILLER_91_197
timestamp 1677580104
transform 1 0 20064 0 -1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_91_199
timestamp 1677579658
transform 1 0 20256 0 -1 70308
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_17
timestamp 1677580104
transform 1 0 2784 0 1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_19
timestamp 1677579658
transform 1 0 2976 0 1 70308
box -48 -56 144 834
use sg13g2_fill_2  FILLER_92_54
timestamp 1677580104
transform 1 0 6336 0 1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_94
timestamp 1677579658
transform 1 0 10176 0 1 70308
box -48 -56 144 834
use sg13g2_decap_4  FILLER_92_106
timestamp 1679577901
transform 1 0 11328 0 1 70308
box -48 -56 432 834
use sg13g2_fill_2  FILLER_92_110
timestamp 1677580104
transform 1 0 11712 0 1 70308
box -48 -56 240 834
use sg13g2_decap_8  FILLER_92_148
timestamp 1679581782
transform 1 0 15360 0 1 70308
box -48 -56 720 834
use sg13g2_fill_1  FILLER_92_155
timestamp 1677579658
transform 1 0 16032 0 1 70308
box -48 -56 144 834
use sg13g2_decap_8  FILLER_92_173
timestamp 1679581782
transform 1 0 17760 0 1 70308
box -48 -56 720 834
use sg13g2_fill_2  FILLER_92_197
timestamp 1677580104
transform 1 0 20064 0 1 70308
box -48 -56 240 834
use sg13g2_fill_1  FILLER_92_199
timestamp 1677579658
transform 1 0 20256 0 1 70308
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_0
timestamp 1677580104
transform 1 0 1152 0 -1 71820
box -48 -56 240 834
use sg13g2_decap_8  FILLER_93_23
timestamp 1679581782
transform 1 0 3360 0 -1 71820
box -48 -56 720 834
use sg13g2_fill_1  FILLER_93_30
timestamp 1677579658
transform 1 0 4032 0 -1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_93_112
timestamp 1677580104
transform 1 0 11904 0 -1 71820
box -48 -56 240 834
use sg13g2_decap_4  FILLER_93_173
timestamp 1679577901
transform 1 0 17760 0 -1 71820
box -48 -56 432 834
use sg13g2_fill_1  FILLER_93_177
timestamp 1677579658
transform 1 0 18144 0 -1 71820
box -48 -56 144 834
use sg13g2_decap_4  FILLER_93_195
timestamp 1679577901
transform 1 0 19872 0 -1 71820
box -48 -56 432 834
use sg13g2_fill_1  FILLER_93_199
timestamp 1677579658
transform 1 0 20256 0 -1 71820
box -48 -56 144 834
use sg13g2_decap_4  FILLER_94_0
timestamp 1679577901
transform 1 0 1152 0 1 71820
box -48 -56 432 834
use sg13g2_fill_1  FILLER_94_4
timestamp 1677579658
transform 1 0 1536 0 1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_94_22
timestamp 1679581782
transform 1 0 3264 0 1 71820
box -48 -56 720 834
use sg13g2_fill_2  FILLER_94_29
timestamp 1677580104
transform 1 0 3936 0 1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_94_31
timestamp 1677579658
transform 1 0 4128 0 1 71820
box -48 -56 144 834
use sg13g2_fill_2  FILLER_94_66
timestamp 1677580104
transform 1 0 7488 0 1 71820
box -48 -56 240 834
use sg13g2_fill_1  FILLER_94_107
timestamp 1677579658
transform 1 0 11424 0 1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_94_171
timestamp 1679581782
transform 1 0 17568 0 1 71820
box -48 -56 720 834
use sg13g2_fill_1  FILLER_94_178
timestamp 1677579658
transform 1 0 18240 0 1 71820
box -48 -56 144 834
use sg13g2_decap_8  FILLER_95_17
timestamp 1679581782
transform 1 0 2784 0 -1 73332
box -48 -56 720 834
use sg13g2_fill_1  FILLER_95_24
timestamp 1677579658
transform 1 0 3456 0 -1 73332
box -48 -56 144 834
use sg13g2_decap_4  FILLER_95_46
timestamp 1679577901
transform 1 0 5568 0 -1 73332
box -48 -56 432 834
use sg13g2_fill_2  FILLER_95_72
timestamp 1677580104
transform 1 0 8064 0 -1 73332
box -48 -56 240 834
use sg13g2_decap_8  FILLER_95_99
timestamp 1679581782
transform 1 0 10656 0 -1 73332
box -48 -56 720 834
use sg13g2_fill_2  FILLER_95_106
timestamp 1677580104
transform 1 0 11328 0 -1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_95_108
timestamp 1677579658
transform 1 0 11520 0 -1 73332
box -48 -56 144 834
use sg13g2_fill_2  FILLER_95_131
timestamp 1677580104
transform 1 0 13728 0 -1 73332
box -48 -56 240 834
use sg13g2_decap_8  FILLER_95_171
timestamp 1679581782
transform 1 0 17568 0 -1 73332
box -48 -56 720 834
use sg13g2_fill_1  FILLER_95_178
timestamp 1677579658
transform 1 0 18240 0 -1 73332
box -48 -56 144 834
use sg13g2_decap_4  FILLER_95_196
timestamp 1679577901
transform 1 0 19968 0 -1 73332
box -48 -56 432 834
use sg13g2_fill_2  FILLER_96_0
timestamp 1677580104
transform 1 0 1152 0 1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_2
timestamp 1677579658
transform 1 0 1344 0 1 73332
box -48 -56 144 834
use sg13g2_fill_1  FILLER_96_74
timestamp 1677579658
transform 1 0 8256 0 1 73332
box -48 -56 144 834
use sg13g2_fill_2  FILLER_96_134
timestamp 1677580104
transform 1 0 14016 0 1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_153
timestamp 1677579658
transform 1 0 15840 0 1 73332
box -48 -56 144 834
use sg13g2_decap_4  FILLER_96_157
timestamp 1679577901
transform 1 0 16224 0 1 73332
box -48 -56 432 834
use sg13g2_fill_2  FILLER_96_161
timestamp 1677580104
transform 1 0 16608 0 1 73332
box -48 -56 240 834
use sg13g2_fill_2  FILLER_96_197
timestamp 1677580104
transform 1 0 20064 0 1 73332
box -48 -56 240 834
use sg13g2_fill_1  FILLER_96_199
timestamp 1677579658
transform 1 0 20256 0 1 73332
box -48 -56 144 834
use sg13g2_decap_8  FILLER_97_0
timestamp 1679581782
transform 1 0 1152 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_4  FILLER_97_24
timestamp 1679577901
transform 1 0 3456 0 -1 74844
box -48 -56 432 834
use sg13g2_fill_1  FILLER_97_28
timestamp 1677579658
transform 1 0 3840 0 -1 74844
box -48 -56 144 834
use sg13g2_fill_2  FILLER_97_46
timestamp 1677580104
transform 1 0 5568 0 -1 74844
box -48 -56 240 834
use sg13g2_fill_1  FILLER_97_48
timestamp 1677579658
transform 1 0 5760 0 -1 74844
box -48 -56 144 834
use sg13g2_decap_8  FILLER_97_70
timestamp 1679581782
transform 1 0 7872 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_97_77
timestamp 1679581782
transform 1 0 8544 0 -1 74844
box -48 -56 720 834
use sg13g2_decap_4  FILLER_97_84
timestamp 1679577901
transform 1 0 9216 0 -1 74844
box -48 -56 432 834
use sg13g2_fill_2  FILLER_97_114
timestamp 1677580104
transform 1 0 12096 0 -1 74844
box -48 -56 240 834
use sg13g2_fill_1  FILLER_97_116
timestamp 1677579658
transform 1 0 12288 0 -1 74844
box -48 -56 144 834
use sg13g2_fill_2  FILLER_97_147
timestamp 1677580104
transform 1 0 15264 0 -1 74844
box -48 -56 240 834
use sg13g2_fill_2  FILLER_98_0
timestamp 1677580104
transform 1 0 1152 0 1 74844
box -48 -56 240 834
use sg13g2_decap_4  FILLER_98_6
timestamp 1679577901
transform 1 0 1728 0 1 74844
box -48 -56 432 834
use sg13g2_fill_1  FILLER_98_127
timestamp 1677579658
transform 1 0 13344 0 1 74844
box -48 -56 144 834
use sg13g2_fill_1  FILLER_98_145
timestamp 1677579658
transform 1 0 15072 0 1 74844
box -48 -56 144 834
use sg13g2_fill_1  FILLER_98_159
timestamp 1677579658
transform 1 0 16416 0 1 74844
box -48 -56 144 834
use sg13g2_decap_8  FILLER_98_181
timestamp 1679581782
transform 1 0 18528 0 1 74844
box -48 -56 720 834
use sg13g2_decap_8  FILLER_98_188
timestamp 1679581782
transform 1 0 19200 0 1 74844
box -48 -56 720 834
use sg13g2_fill_1  FILLER_98_195
timestamp 1677579658
transform 1 0 19872 0 1 74844
box -48 -56 144 834
use sg13g2_fill_1  FILLER_98_199
timestamp 1677579658
transform 1 0 20256 0 1 74844
box -48 -56 144 834
use sg13g2_fill_1  FILLER_99_38
timestamp 1677579658
transform 1 0 4800 0 -1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_99_74
timestamp 1679581782
transform 1 0 8256 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_99_81
timestamp 1679581782
transform 1 0 8928 0 -1 76356
box -48 -56 720 834
use sg13g2_decap_4  FILLER_99_88
timestamp 1679577901
transform 1 0 9600 0 -1 76356
box -48 -56 432 834
use sg13g2_fill_1  FILLER_99_92
timestamp 1677579658
transform 1 0 9984 0 -1 76356
box -48 -56 144 834
use sg13g2_decap_4  FILLER_99_110
timestamp 1679577901
transform 1 0 11712 0 -1 76356
box -48 -56 432 834
use sg13g2_fill_2  FILLER_99_131
timestamp 1677580104
transform 1 0 13728 0 -1 76356
box -48 -56 240 834
use sg13g2_fill_1  FILLER_99_155
timestamp 1677579658
transform 1 0 16032 0 -1 76356
box -48 -56 144 834
use sg13g2_fill_2  FILLER_99_190
timestamp 1677580104
transform 1 0 19392 0 -1 76356
box -48 -56 240 834
use sg13g2_fill_1  FILLER_99_195
timestamp 1677579658
transform 1 0 19872 0 -1 76356
box -48 -56 144 834
use sg13g2_fill_1  FILLER_100_0
timestamp 1677579658
transform 1 0 1152 0 1 76356
box -48 -56 144 834
use sg13g2_fill_1  FILLER_100_39
timestamp 1677579658
transform 1 0 4896 0 1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_100_95
timestamp 1679581782
transform 1 0 10272 0 1 76356
box -48 -56 720 834
use sg13g2_fill_1  FILLER_100_102
timestamp 1677579658
transform 1 0 10944 0 1 76356
box -48 -56 144 834
use sg13g2_decap_8  FILLER_100_120
timestamp 1679581782
transform 1 0 12672 0 1 76356
box -48 -56 720 834
use sg13g2_decap_8  FILLER_100_127
timestamp 1679581782
transform 1 0 13344 0 1 76356
box -48 -56 720 834
use sg13g2_decap_4  FILLER_100_134
timestamp 1679577901
transform 1 0 14016 0 1 76356
box -48 -56 432 834
use sg13g2_fill_1  FILLER_100_138
timestamp 1677579658
transform 1 0 14400 0 1 76356
box -48 -56 144 834
use sg13g2_fill_1  FILLER_100_173
timestamp 1677579658
transform 1 0 17760 0 1 76356
box -48 -56 144 834
use sg13g2_fill_1  FILLER_100_199
timestamp 1677579658
transform 1 0 20256 0 1 76356
box -48 -56 144 834
use sg13g2_fill_1  FILLER_101_17
timestamp 1677579658
transform 1 0 2784 0 -1 77868
box -48 -56 144 834
use sg13g2_decap_8  FILLER_101_43
timestamp 1679581782
transform 1 0 5280 0 -1 77868
box -48 -56 720 834
use sg13g2_fill_2  FILLER_101_79
timestamp 1677580104
transform 1 0 8736 0 -1 77868
box -48 -56 240 834
use sg13g2_decap_8  FILLER_101_119
timestamp 1679581782
transform 1 0 12576 0 -1 77868
box -48 -56 720 834
use sg13g2_fill_1  FILLER_101_126
timestamp 1677579658
transform 1 0 13248 0 -1 77868
box -48 -56 144 834
use sg13g2_fill_1  FILLER_101_148
timestamp 1677579658
transform 1 0 15360 0 -1 77868
box -48 -56 144 834
use sg13g2_fill_2  FILLER_101_198
timestamp 1677580104
transform 1 0 20160 0 -1 77868
box -48 -56 240 834
use sg13g2_fill_2  FILLER_102_73
timestamp 1677580104
transform 1 0 8160 0 1 77868
box -48 -56 240 834
use sg13g2_decap_4  FILLER_102_92
timestamp 1679577901
transform 1 0 9984 0 1 77868
box -48 -56 432 834
use sg13g2_decap_8  FILLER_102_117
timestamp 1679581782
transform 1 0 12384 0 1 77868
box -48 -56 720 834
use sg13g2_fill_1  FILLER_102_124
timestamp 1677579658
transform 1 0 13056 0 1 77868
box -48 -56 144 834
use sg13g2_fill_1  FILLER_102_199
timestamp 1677579658
transform 1 0 20256 0 1 77868
box -48 -56 144 834
use sg13g2_fill_1  FILLER_103_38
timestamp 1677579658
transform 1 0 4800 0 -1 79380
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_56
timestamp 1677580104
transform 1 0 6528 0 -1 79380
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_58
timestamp 1677579658
transform 1 0 6720 0 -1 79380
box -48 -56 144 834
use sg13g2_fill_1  FILLER_103_67
timestamp 1677579658
transform 1 0 7584 0 -1 79380
box -48 -56 144 834
use sg13g2_fill_2  FILLER_103_77
timestamp 1677580104
transform 1 0 8544 0 -1 79380
box -48 -56 240 834
use sg13g2_fill_1  FILLER_103_96
timestamp 1677579658
transform 1 0 10368 0 -1 79380
box -48 -56 144 834
use sg13g2_fill_1  FILLER_103_152
timestamp 1677579658
transform 1 0 15744 0 -1 79380
box -48 -56 144 834
use sg13g2_fill_1  FILLER_103_199
timestamp 1677579658
transform 1 0 20256 0 -1 79380
box -48 -56 144 834
use sg13g2_fill_1  FILLER_104_0
timestamp 1677579658
transform 1 0 1152 0 1 79380
box -48 -56 144 834
use sg13g2_fill_1  FILLER_104_26
timestamp 1677579658
transform 1 0 3648 0 1 79380
box -48 -56 144 834
use sg13g2_fill_2  FILLER_104_67
timestamp 1677580104
transform 1 0 7584 0 1 79380
box -48 -56 240 834
use sg13g2_decap_8  FILLER_104_120
timestamp 1679581782
transform 1 0 12672 0 1 79380
box -48 -56 720 834
use sg13g2_fill_2  FILLER_104_127
timestamp 1677580104
transform 1 0 13344 0 1 79380
box -48 -56 240 834
use sg13g2_fill_1  FILLER_104_129
timestamp 1677579658
transform 1 0 13536 0 1 79380
box -48 -56 144 834
use sg13g2_fill_2  FILLER_104_198
timestamp 1677580104
transform 1 0 20160 0 1 79380
box -48 -56 240 834
use sg13g2_fill_1  FILLER_105_21
timestamp 1677579658
transform 1 0 3168 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_1  FILLER_105_25
timestamp 1677579658
transform 1 0 3552 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_2  FILLER_105_54
timestamp 1677580104
transform 1 0 6336 0 -1 80892
box -48 -56 240 834
use sg13g2_fill_2  FILLER_105_85
timestamp 1677580104
transform 1 0 9312 0 -1 80892
box -48 -56 240 834
use sg13g2_fill_1  FILLER_105_87
timestamp 1677579658
transform 1 0 9504 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_1  FILLER_105_109
timestamp 1677579658
transform 1 0 11616 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_1  FILLER_105_151
timestamp 1677579658
transform 1 0 15648 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_1  FILLER_105_178
timestamp 1677579658
transform 1 0 18240 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_1  FILLER_105_199
timestamp 1677579658
transform 1 0 20256 0 -1 80892
box -48 -56 144 834
use sg13g2_fill_2  FILLER_106_17
timestamp 1677580104
transform 1 0 2784 0 1 80892
box -48 -56 240 834
use sg13g2_fill_2  FILLER_106_101
timestamp 1677580104
transform 1 0 10848 0 1 80892
box -48 -56 240 834
use sg13g2_fill_1  FILLER_106_103
timestamp 1677579658
transform 1 0 11040 0 1 80892
box -48 -56 144 834
use sg13g2_fill_1  FILLER_106_179
timestamp 1677579658
transform 1 0 18336 0 1 80892
box -48 -56 144 834
use sg13g2_fill_2  FILLER_107_21
timestamp 1677580104
transform 1 0 3168 0 -1 82404
box -48 -56 240 834
use sg13g2_fill_1  FILLER_107_136
timestamp 1677579658
transform 1 0 14208 0 -1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_107_161
timestamp 1677579658
transform 1 0 16608 0 -1 82404
box -48 -56 144 834
use sg13g2_fill_2  FILLER_107_179
timestamp 1677580104
transform 1 0 18336 0 -1 82404
box -48 -56 240 834
use sg13g2_fill_2  FILLER_107_198
timestamp 1677580104
transform 1 0 20160 0 -1 82404
box -48 -56 240 834
use sg13g2_fill_1  FILLER_108_0
timestamp 1677579658
transform 1 0 1152 0 1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_108_18
timestamp 1677579658
transform 1 0 2880 0 1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_108_43
timestamp 1677579658
transform 1 0 5280 0 1 82404
box -48 -56 144 834
use sg13g2_fill_1  FILLER_108_77
timestamp 1677579658
transform 1 0 8544 0 1 82404
box -48 -56 144 834
use sg13g2_fill_2  FILLER_108_112
timestamp 1677580104
transform 1 0 11904 0 1 82404
box -48 -56 240 834
use sg13g2_fill_2  FILLER_108_125
timestamp 1677580104
transform 1 0 13152 0 1 82404
box -48 -56 240 834
use sg13g2_fill_1  FILLER_109_0
timestamp 1677579658
transform 1 0 1152 0 -1 83916
box -48 -56 144 834
use sg13g2_fill_2  FILLER_109_59
timestamp 1677580104
transform 1 0 6816 0 -1 83916
box -48 -56 240 834
use sg13g2_fill_2  FILLER_109_112
timestamp 1677580104
transform 1 0 11904 0 -1 83916
box -48 -56 240 834
use sg13g2_fill_1  FILLER_109_158
timestamp 1677579658
transform 1 0 16320 0 -1 83916
box -48 -56 144 834
use sg13g2_fill_2  FILLER_109_184
timestamp 1677580104
transform 1 0 18816 0 -1 83916
box -48 -56 240 834
use sg13g2_fill_1  FILLER_109_199
timestamp 1677579658
transform 1 0 20256 0 -1 83916
box -48 -56 144 834
use sg13g2_fill_1  FILLER_110_0
timestamp 1677579658
transform 1 0 1152 0 1 83916
box -48 -56 144 834
use sg13g2_fill_1  FILLER_110_60
timestamp 1677579658
transform 1 0 6912 0 1 83916
box -48 -56 144 834
use sg13g2_fill_2  FILLER_110_65
timestamp 1677580104
transform 1 0 7392 0 1 83916
box -48 -56 240 834
use sg13g2_fill_2  FILLER_110_113
timestamp 1677580104
transform 1 0 12000 0 1 83916
box -48 -56 240 834
<< labels >>
flabel metal3 s 21424 24404 21504 24484 0 FreeSans 320 0 0 0 ADDR_SRAM0
port 0 nsew signal output
flabel metal3 s 21424 24740 21504 24820 0 FreeSans 320 0 0 0 ADDR_SRAM1
port 1 nsew signal output
flabel metal3 s 21424 25076 21504 25156 0 FreeSans 320 0 0 0 ADDR_SRAM2
port 2 nsew signal output
flabel metal3 s 21424 25412 21504 25492 0 FreeSans 320 0 0 0 ADDR_SRAM3
port 3 nsew signal output
flabel metal3 s 21424 25748 21504 25828 0 FreeSans 320 0 0 0 ADDR_SRAM4
port 4 nsew signal output
flabel metal3 s 21424 26084 21504 26164 0 FreeSans 320 0 0 0 ADDR_SRAM5
port 5 nsew signal output
flabel metal3 s 21424 26420 21504 26500 0 FreeSans 320 0 0 0 ADDR_SRAM6
port 6 nsew signal output
flabel metal3 s 21424 26756 21504 26836 0 FreeSans 320 0 0 0 ADDR_SRAM7
port 7 nsew signal output
flabel metal3 s 21424 27092 21504 27172 0 FreeSans 320 0 0 0 ADDR_SRAM8
port 8 nsew signal output
flabel metal3 s 21424 27428 21504 27508 0 FreeSans 320 0 0 0 ADDR_SRAM9
port 9 nsew signal output
flabel metal3 s 21424 38516 21504 38596 0 FreeSans 320 0 0 0 BM_SRAM0
port 10 nsew signal output
flabel metal3 s 21424 38852 21504 38932 0 FreeSans 320 0 0 0 BM_SRAM1
port 11 nsew signal output
flabel metal3 s 21424 41876 21504 41956 0 FreeSans 320 0 0 0 BM_SRAM10
port 12 nsew signal output
flabel metal3 s 21424 42212 21504 42292 0 FreeSans 320 0 0 0 BM_SRAM11
port 13 nsew signal output
flabel metal3 s 21424 42548 21504 42628 0 FreeSans 320 0 0 0 BM_SRAM12
port 14 nsew signal output
flabel metal3 s 21424 42884 21504 42964 0 FreeSans 320 0 0 0 BM_SRAM13
port 15 nsew signal output
flabel metal3 s 21424 43220 21504 43300 0 FreeSans 320 0 0 0 BM_SRAM14
port 16 nsew signal output
flabel metal3 s 21424 43556 21504 43636 0 FreeSans 320 0 0 0 BM_SRAM15
port 17 nsew signal output
flabel metal3 s 21424 43892 21504 43972 0 FreeSans 320 0 0 0 BM_SRAM16
port 18 nsew signal output
flabel metal3 s 21424 44228 21504 44308 0 FreeSans 320 0 0 0 BM_SRAM17
port 19 nsew signal output
flabel metal3 s 21424 44564 21504 44644 0 FreeSans 320 0 0 0 BM_SRAM18
port 20 nsew signal output
flabel metal3 s 21424 44900 21504 44980 0 FreeSans 320 0 0 0 BM_SRAM19
port 21 nsew signal output
flabel metal3 s 21424 39188 21504 39268 0 FreeSans 320 0 0 0 BM_SRAM2
port 22 nsew signal output
flabel metal3 s 21424 45236 21504 45316 0 FreeSans 320 0 0 0 BM_SRAM20
port 23 nsew signal output
flabel metal3 s 21424 45572 21504 45652 0 FreeSans 320 0 0 0 BM_SRAM21
port 24 nsew signal output
flabel metal3 s 21424 45908 21504 45988 0 FreeSans 320 0 0 0 BM_SRAM22
port 25 nsew signal output
flabel metal3 s 21424 46244 21504 46324 0 FreeSans 320 0 0 0 BM_SRAM23
port 26 nsew signal output
flabel metal3 s 21424 46580 21504 46660 0 FreeSans 320 0 0 0 BM_SRAM24
port 27 nsew signal output
flabel metal3 s 21424 46916 21504 46996 0 FreeSans 320 0 0 0 BM_SRAM25
port 28 nsew signal output
flabel metal3 s 21424 47252 21504 47332 0 FreeSans 320 0 0 0 BM_SRAM26
port 29 nsew signal output
flabel metal3 s 21424 47588 21504 47668 0 FreeSans 320 0 0 0 BM_SRAM27
port 30 nsew signal output
flabel metal3 s 21424 47924 21504 48004 0 FreeSans 320 0 0 0 BM_SRAM28
port 31 nsew signal output
flabel metal3 s 21424 48260 21504 48340 0 FreeSans 320 0 0 0 BM_SRAM29
port 32 nsew signal output
flabel metal3 s 21424 39524 21504 39604 0 FreeSans 320 0 0 0 BM_SRAM3
port 33 nsew signal output
flabel metal3 s 21424 48596 21504 48676 0 FreeSans 320 0 0 0 BM_SRAM30
port 34 nsew signal output
flabel metal3 s 21424 48932 21504 49012 0 FreeSans 320 0 0 0 BM_SRAM31
port 35 nsew signal output
flabel metal3 s 21424 39860 21504 39940 0 FreeSans 320 0 0 0 BM_SRAM4
port 36 nsew signal output
flabel metal3 s 21424 40196 21504 40276 0 FreeSans 320 0 0 0 BM_SRAM5
port 37 nsew signal output
flabel metal3 s 21424 40532 21504 40612 0 FreeSans 320 0 0 0 BM_SRAM6
port 38 nsew signal output
flabel metal3 s 21424 40868 21504 40948 0 FreeSans 320 0 0 0 BM_SRAM7
port 39 nsew signal output
flabel metal3 s 21424 41204 21504 41284 0 FreeSans 320 0 0 0 BM_SRAM8
port 40 nsew signal output
flabel metal3 s 21424 41540 21504 41620 0 FreeSans 320 0 0 0 BM_SRAM9
port 41 nsew signal output
flabel metal3 s 21424 50276 21504 50356 0 FreeSans 320 0 0 0 CLK_SRAM
port 42 nsew signal output
flabel metal3 s 21424 24068 21504 24148 0 FreeSans 320 0 0 0 CONFIGURED_top
port 43 nsew signal input
flabel metal3 s 21424 27764 21504 27844 0 FreeSans 320 0 0 0 DIN_SRAM0
port 44 nsew signal output
flabel metal3 s 21424 28100 21504 28180 0 FreeSans 320 0 0 0 DIN_SRAM1
port 45 nsew signal output
flabel metal3 s 21424 31124 21504 31204 0 FreeSans 320 0 0 0 DIN_SRAM10
port 46 nsew signal output
flabel metal3 s 21424 31460 21504 31540 0 FreeSans 320 0 0 0 DIN_SRAM11
port 47 nsew signal output
flabel metal3 s 21424 31796 21504 31876 0 FreeSans 320 0 0 0 DIN_SRAM12
port 48 nsew signal output
flabel metal3 s 21424 32132 21504 32212 0 FreeSans 320 0 0 0 DIN_SRAM13
port 49 nsew signal output
flabel metal3 s 21424 32468 21504 32548 0 FreeSans 320 0 0 0 DIN_SRAM14
port 50 nsew signal output
flabel metal3 s 21424 32804 21504 32884 0 FreeSans 320 0 0 0 DIN_SRAM15
port 51 nsew signal output
flabel metal3 s 21424 33140 21504 33220 0 FreeSans 320 0 0 0 DIN_SRAM16
port 52 nsew signal output
flabel metal3 s 21424 33476 21504 33556 0 FreeSans 320 0 0 0 DIN_SRAM17
port 53 nsew signal output
flabel metal3 s 21424 33812 21504 33892 0 FreeSans 320 0 0 0 DIN_SRAM18
port 54 nsew signal output
flabel metal3 s 21424 34148 21504 34228 0 FreeSans 320 0 0 0 DIN_SRAM19
port 55 nsew signal output
flabel metal3 s 21424 28436 21504 28516 0 FreeSans 320 0 0 0 DIN_SRAM2
port 56 nsew signal output
flabel metal3 s 21424 34484 21504 34564 0 FreeSans 320 0 0 0 DIN_SRAM20
port 57 nsew signal output
flabel metal3 s 21424 34820 21504 34900 0 FreeSans 320 0 0 0 DIN_SRAM21
port 58 nsew signal output
flabel metal3 s 21424 35156 21504 35236 0 FreeSans 320 0 0 0 DIN_SRAM22
port 59 nsew signal output
flabel metal3 s 21424 35492 21504 35572 0 FreeSans 320 0 0 0 DIN_SRAM23
port 60 nsew signal output
flabel metal3 s 21424 35828 21504 35908 0 FreeSans 320 0 0 0 DIN_SRAM24
port 61 nsew signal output
flabel metal3 s 21424 36164 21504 36244 0 FreeSans 320 0 0 0 DIN_SRAM25
port 62 nsew signal output
flabel metal3 s 21424 36500 21504 36580 0 FreeSans 320 0 0 0 DIN_SRAM26
port 63 nsew signal output
flabel metal3 s 21424 36836 21504 36916 0 FreeSans 320 0 0 0 DIN_SRAM27
port 64 nsew signal output
flabel metal3 s 21424 37172 21504 37252 0 FreeSans 320 0 0 0 DIN_SRAM28
port 65 nsew signal output
flabel metal3 s 21424 37508 21504 37588 0 FreeSans 320 0 0 0 DIN_SRAM29
port 66 nsew signal output
flabel metal3 s 21424 28772 21504 28852 0 FreeSans 320 0 0 0 DIN_SRAM3
port 67 nsew signal output
flabel metal3 s 21424 37844 21504 37924 0 FreeSans 320 0 0 0 DIN_SRAM30
port 68 nsew signal output
flabel metal3 s 21424 38180 21504 38260 0 FreeSans 320 0 0 0 DIN_SRAM31
port 69 nsew signal output
flabel metal3 s 21424 29108 21504 29188 0 FreeSans 320 0 0 0 DIN_SRAM4
port 70 nsew signal output
flabel metal3 s 21424 29444 21504 29524 0 FreeSans 320 0 0 0 DIN_SRAM5
port 71 nsew signal output
flabel metal3 s 21424 29780 21504 29860 0 FreeSans 320 0 0 0 DIN_SRAM6
port 72 nsew signal output
flabel metal3 s 21424 30116 21504 30196 0 FreeSans 320 0 0 0 DIN_SRAM7
port 73 nsew signal output
flabel metal3 s 21424 30452 21504 30532 0 FreeSans 320 0 0 0 DIN_SRAM8
port 74 nsew signal output
flabel metal3 s 21424 30788 21504 30868 0 FreeSans 320 0 0 0 DIN_SRAM9
port 75 nsew signal output
flabel metal3 s 21424 13316 21504 13396 0 FreeSans 320 0 0 0 DOUT_SRAM0
port 76 nsew signal input
flabel metal3 s 21424 13652 21504 13732 0 FreeSans 320 0 0 0 DOUT_SRAM1
port 77 nsew signal input
flabel metal3 s 21424 16676 21504 16756 0 FreeSans 320 0 0 0 DOUT_SRAM10
port 78 nsew signal input
flabel metal3 s 21424 17012 21504 17092 0 FreeSans 320 0 0 0 DOUT_SRAM11
port 79 nsew signal input
flabel metal3 s 21424 17348 21504 17428 0 FreeSans 320 0 0 0 DOUT_SRAM12
port 80 nsew signal input
flabel metal3 s 21424 17684 21504 17764 0 FreeSans 320 0 0 0 DOUT_SRAM13
port 81 nsew signal input
flabel metal3 s 21424 18020 21504 18100 0 FreeSans 320 0 0 0 DOUT_SRAM14
port 82 nsew signal input
flabel metal3 s 21424 18356 21504 18436 0 FreeSans 320 0 0 0 DOUT_SRAM15
port 83 nsew signal input
flabel metal3 s 21424 18692 21504 18772 0 FreeSans 320 0 0 0 DOUT_SRAM16
port 84 nsew signal input
flabel metal3 s 21424 19028 21504 19108 0 FreeSans 320 0 0 0 DOUT_SRAM17
port 85 nsew signal input
flabel metal3 s 21424 19364 21504 19444 0 FreeSans 320 0 0 0 DOUT_SRAM18
port 86 nsew signal input
flabel metal3 s 21424 19700 21504 19780 0 FreeSans 320 0 0 0 DOUT_SRAM19
port 87 nsew signal input
flabel metal3 s 21424 13988 21504 14068 0 FreeSans 320 0 0 0 DOUT_SRAM2
port 88 nsew signal input
flabel metal3 s 21424 20036 21504 20116 0 FreeSans 320 0 0 0 DOUT_SRAM20
port 89 nsew signal input
flabel metal3 s 21424 20372 21504 20452 0 FreeSans 320 0 0 0 DOUT_SRAM21
port 90 nsew signal input
flabel metal3 s 21424 20708 21504 20788 0 FreeSans 320 0 0 0 DOUT_SRAM22
port 91 nsew signal input
flabel metal3 s 21424 21044 21504 21124 0 FreeSans 320 0 0 0 DOUT_SRAM23
port 92 nsew signal input
flabel metal3 s 21424 21380 21504 21460 0 FreeSans 320 0 0 0 DOUT_SRAM24
port 93 nsew signal input
flabel metal3 s 21424 21716 21504 21796 0 FreeSans 320 0 0 0 DOUT_SRAM25
port 94 nsew signal input
flabel metal3 s 21424 22052 21504 22132 0 FreeSans 320 0 0 0 DOUT_SRAM26
port 95 nsew signal input
flabel metal3 s 21424 22388 21504 22468 0 FreeSans 320 0 0 0 DOUT_SRAM27
port 96 nsew signal input
flabel metal3 s 21424 22724 21504 22804 0 FreeSans 320 0 0 0 DOUT_SRAM28
port 97 nsew signal input
flabel metal3 s 21424 23060 21504 23140 0 FreeSans 320 0 0 0 DOUT_SRAM29
port 98 nsew signal input
flabel metal3 s 21424 14324 21504 14404 0 FreeSans 320 0 0 0 DOUT_SRAM3
port 99 nsew signal input
flabel metal3 s 21424 23396 21504 23476 0 FreeSans 320 0 0 0 DOUT_SRAM30
port 100 nsew signal input
flabel metal3 s 21424 23732 21504 23812 0 FreeSans 320 0 0 0 DOUT_SRAM31
port 101 nsew signal input
flabel metal3 s 21424 14660 21504 14740 0 FreeSans 320 0 0 0 DOUT_SRAM4
port 102 nsew signal input
flabel metal3 s 21424 14996 21504 15076 0 FreeSans 320 0 0 0 DOUT_SRAM5
port 103 nsew signal input
flabel metal3 s 21424 15332 21504 15412 0 FreeSans 320 0 0 0 DOUT_SRAM6
port 104 nsew signal input
flabel metal3 s 21424 15668 21504 15748 0 FreeSans 320 0 0 0 DOUT_SRAM7
port 105 nsew signal input
flabel metal3 s 21424 16004 21504 16084 0 FreeSans 320 0 0 0 DOUT_SRAM8
port 106 nsew signal input
flabel metal3 s 21424 16340 21504 16420 0 FreeSans 320 0 0 0 DOUT_SRAM9
port 107 nsew signal input
flabel metal3 s 21424 49604 21504 49684 0 FreeSans 320 0 0 0 MEN_SRAM
port 108 nsew signal output
flabel metal3 s 21424 49940 21504 50020 0 FreeSans 320 0 0 0 REN_SRAM
port 109 nsew signal output
flabel metal3 s 21424 50612 21504 50692 0 FreeSans 320 0 0 0 TIE_HIGH_SRAM
port 110 nsew signal output
flabel metal3 s 21424 50948 21504 51028 0 FreeSans 320 0 0 0 TIE_LOW_SRAM
port 111 nsew signal output
flabel metal3 s 0 59180 80 59260 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[0]
port 112 nsew signal input
flabel metal3 s 0 59516 80 59596 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[1]
port 113 nsew signal input
flabel metal3 s 0 59852 80 59932 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[2]
port 114 nsew signal input
flabel metal3 s 0 60188 80 60268 0 FreeSans 320 0 0 0 Tile_X0Y0_E1END[3]
port 115 nsew signal input
flabel metal3 s 0 63212 80 63292 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[0]
port 116 nsew signal input
flabel metal3 s 0 63548 80 63628 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[1]
port 117 nsew signal input
flabel metal3 s 0 63884 80 63964 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[2]
port 118 nsew signal input
flabel metal3 s 0 64220 80 64300 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[3]
port 119 nsew signal input
flabel metal3 s 0 64556 80 64636 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[4]
port 120 nsew signal input
flabel metal3 s 0 64892 80 64972 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[5]
port 121 nsew signal input
flabel metal3 s 0 65228 80 65308 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[6]
port 122 nsew signal input
flabel metal3 s 0 65564 80 65644 0 FreeSans 320 0 0 0 Tile_X0Y0_E2END[7]
port 123 nsew signal input
flabel metal3 s 0 60524 80 60604 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[0]
port 124 nsew signal input
flabel metal3 s 0 60860 80 60940 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[1]
port 125 nsew signal input
flabel metal3 s 0 61196 80 61276 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[2]
port 126 nsew signal input
flabel metal3 s 0 61532 80 61612 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[3]
port 127 nsew signal input
flabel metal3 s 0 61868 80 61948 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[4]
port 128 nsew signal input
flabel metal3 s 0 62204 80 62284 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[5]
port 129 nsew signal input
flabel metal3 s 0 62540 80 62620 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[6]
port 130 nsew signal input
flabel metal3 s 0 62876 80 62956 0 FreeSans 320 0 0 0 Tile_X0Y0_E2MID[7]
port 131 nsew signal input
flabel metal3 s 0 71276 80 71356 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[0]
port 132 nsew signal input
flabel metal3 s 0 74636 80 74716 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[10]
port 133 nsew signal input
flabel metal3 s 0 74972 80 75052 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[11]
port 134 nsew signal input
flabel metal3 s 0 71612 80 71692 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[1]
port 135 nsew signal input
flabel metal3 s 0 71948 80 72028 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[2]
port 136 nsew signal input
flabel metal3 s 0 72284 80 72364 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[3]
port 137 nsew signal input
flabel metal3 s 0 72620 80 72700 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[4]
port 138 nsew signal input
flabel metal3 s 0 72956 80 73036 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[5]
port 139 nsew signal input
flabel metal3 s 0 73292 80 73372 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[6]
port 140 nsew signal input
flabel metal3 s 0 73628 80 73708 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[7]
port 141 nsew signal input
flabel metal3 s 0 73964 80 74044 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[8]
port 142 nsew signal input
flabel metal3 s 0 74300 80 74380 0 FreeSans 320 0 0 0 Tile_X0Y0_E6END[9]
port 143 nsew signal input
flabel metal3 s 0 65900 80 65980 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[0]
port 144 nsew signal input
flabel metal3 s 0 69260 80 69340 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[10]
port 145 nsew signal input
flabel metal3 s 0 69596 80 69676 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[11]
port 146 nsew signal input
flabel metal3 s 0 69932 80 70012 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[12]
port 147 nsew signal input
flabel metal3 s 0 70268 80 70348 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[13]
port 148 nsew signal input
flabel metal3 s 0 70604 80 70684 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[14]
port 149 nsew signal input
flabel metal3 s 0 70940 80 71020 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[15]
port 150 nsew signal input
flabel metal3 s 0 66236 80 66316 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[1]
port 151 nsew signal input
flabel metal3 s 0 66572 80 66652 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[2]
port 152 nsew signal input
flabel metal3 s 0 66908 80 66988 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[3]
port 153 nsew signal input
flabel metal3 s 0 67244 80 67324 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[4]
port 154 nsew signal input
flabel metal3 s 0 67580 80 67660 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[5]
port 155 nsew signal input
flabel metal3 s 0 67916 80 67996 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[6]
port 156 nsew signal input
flabel metal3 s 0 68252 80 68332 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[7]
port 157 nsew signal input
flabel metal3 s 0 68588 80 68668 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[8]
port 158 nsew signal input
flabel metal3 s 0 68924 80 69004 0 FreeSans 320 0 0 0 Tile_X0Y0_EE4END[9]
port 159 nsew signal input
flabel metal3 s 0 75308 80 75388 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[0]
port 160 nsew signal input
flabel metal3 s 0 78668 80 78748 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[10]
port 161 nsew signal input
flabel metal3 s 0 79004 80 79084 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[11]
port 162 nsew signal input
flabel metal3 s 0 79340 80 79420 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[12]
port 163 nsew signal input
flabel metal3 s 0 79676 80 79756 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[13]
port 164 nsew signal input
flabel metal3 s 0 80012 80 80092 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[14]
port 165 nsew signal input
flabel metal3 s 0 80348 80 80428 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[15]
port 166 nsew signal input
flabel metal3 s 0 80684 80 80764 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[16]
port 167 nsew signal input
flabel metal3 s 0 81020 80 81100 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[17]
port 168 nsew signal input
flabel metal3 s 0 81356 80 81436 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[18]
port 169 nsew signal input
flabel metal3 s 0 81692 80 81772 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[19]
port 170 nsew signal input
flabel metal3 s 0 75644 80 75724 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[1]
port 171 nsew signal input
flabel metal3 s 0 82028 80 82108 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[20]
port 172 nsew signal input
flabel metal3 s 0 82364 80 82444 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[21]
port 173 nsew signal input
flabel metal3 s 0 82700 80 82780 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[22]
port 174 nsew signal input
flabel metal3 s 0 83036 80 83116 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[23]
port 175 nsew signal input
flabel metal3 s 0 83372 80 83452 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[24]
port 176 nsew signal input
flabel metal3 s 0 83708 80 83788 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[25]
port 177 nsew signal input
flabel metal3 s 0 84044 80 84124 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[26]
port 178 nsew signal input
flabel metal3 s 0 84380 80 84460 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[27]
port 179 nsew signal input
flabel metal3 s 0 84716 80 84796 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[28]
port 180 nsew signal input
flabel metal3 s 0 85052 80 85132 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[29]
port 181 nsew signal input
flabel metal3 s 0 75980 80 76060 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[2]
port 182 nsew signal input
flabel metal3 s 0 85388 80 85468 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[30]
port 183 nsew signal input
flabel metal3 s 0 85724 80 85804 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[31]
port 184 nsew signal input
flabel metal3 s 0 76316 80 76396 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[3]
port 185 nsew signal input
flabel metal3 s 0 76652 80 76732 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[4]
port 186 nsew signal input
flabel metal3 s 0 76988 80 77068 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[5]
port 187 nsew signal input
flabel metal3 s 0 77324 80 77404 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[6]
port 188 nsew signal input
flabel metal3 s 0 77660 80 77740 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[7]
port 189 nsew signal input
flabel metal3 s 0 77996 80 78076 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[8]
port 190 nsew signal input
flabel metal3 s 0 78332 80 78412 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData[9]
port 191 nsew signal input
flabel metal3 s 21424 51284 21504 51364 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[0]
port 192 nsew signal output
flabel metal3 s 21424 54644 21504 54724 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[10]
port 193 nsew signal output
flabel metal3 s 21424 54980 21504 55060 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[11]
port 194 nsew signal output
flabel metal3 s 21424 55316 21504 55396 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[12]
port 195 nsew signal output
flabel metal3 s 21424 55652 21504 55732 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[13]
port 196 nsew signal output
flabel metal3 s 21424 55988 21504 56068 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[14]
port 197 nsew signal output
flabel metal3 s 21424 56324 21504 56404 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[15]
port 198 nsew signal output
flabel metal3 s 21424 56660 21504 56740 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[16]
port 199 nsew signal output
flabel metal3 s 21424 56996 21504 57076 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[17]
port 200 nsew signal output
flabel metal3 s 21424 57332 21504 57412 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[18]
port 201 nsew signal output
flabel metal3 s 21424 57668 21504 57748 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[19]
port 202 nsew signal output
flabel metal3 s 21424 51620 21504 51700 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[1]
port 203 nsew signal output
flabel metal3 s 21424 58004 21504 58084 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[20]
port 204 nsew signal output
flabel metal3 s 21424 58340 21504 58420 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[21]
port 205 nsew signal output
flabel metal3 s 21424 58676 21504 58756 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[22]
port 206 nsew signal output
flabel metal3 s 21424 59012 21504 59092 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[23]
port 207 nsew signal output
flabel metal3 s 21424 59348 21504 59428 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[24]
port 208 nsew signal output
flabel metal3 s 21424 59684 21504 59764 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[25]
port 209 nsew signal output
flabel metal3 s 21424 60020 21504 60100 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[26]
port 210 nsew signal output
flabel metal3 s 21424 60356 21504 60436 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[27]
port 211 nsew signal output
flabel metal3 s 21424 60692 21504 60772 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[28]
port 212 nsew signal output
flabel metal3 s 21424 61028 21504 61108 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[29]
port 213 nsew signal output
flabel metal3 s 21424 51956 21504 52036 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[2]
port 214 nsew signal output
flabel metal3 s 21424 61364 21504 61444 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[30]
port 215 nsew signal output
flabel metal3 s 21424 61700 21504 61780 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[31]
port 216 nsew signal output
flabel metal3 s 21424 52292 21504 52372 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[3]
port 217 nsew signal output
flabel metal3 s 21424 52628 21504 52708 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[4]
port 218 nsew signal output
flabel metal3 s 21424 52964 21504 53044 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[5]
port 219 nsew signal output
flabel metal3 s 21424 53300 21504 53380 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[6]
port 220 nsew signal output
flabel metal3 s 21424 53636 21504 53716 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[7]
port 221 nsew signal output
flabel metal3 s 21424 53972 21504 54052 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[8]
port 222 nsew signal output
flabel metal3 s 21424 54308 21504 54388 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameData_O[9]
port 223 nsew signal output
flabel metal2 s 15800 85936 15880 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[0]
port 224 nsew signal output
flabel metal2 s 17720 85936 17800 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[10]
port 225 nsew signal output
flabel metal2 s 17912 85936 17992 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[11]
port 226 nsew signal output
flabel metal2 s 18104 85936 18184 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[12]
port 227 nsew signal output
flabel metal2 s 18296 85936 18376 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[13]
port 228 nsew signal output
flabel metal2 s 18488 85936 18568 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[14]
port 229 nsew signal output
flabel metal2 s 18680 85936 18760 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[15]
port 230 nsew signal output
flabel metal2 s 18872 85936 18952 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[16]
port 231 nsew signal output
flabel metal2 s 19064 85936 19144 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[17]
port 232 nsew signal output
flabel metal2 s 19256 85936 19336 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[18]
port 233 nsew signal output
flabel metal2 s 19448 85936 19528 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[19]
port 234 nsew signal output
flabel metal2 s 15992 85936 16072 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[1]
port 235 nsew signal output
flabel metal2 s 16184 85936 16264 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[2]
port 236 nsew signal output
flabel metal2 s 16376 85936 16456 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[3]
port 237 nsew signal output
flabel metal2 s 16568 85936 16648 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[4]
port 238 nsew signal output
flabel metal2 s 16760 85936 16840 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[5]
port 239 nsew signal output
flabel metal2 s 16952 85936 17032 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[6]
port 240 nsew signal output
flabel metal2 s 17144 85936 17224 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[7]
port 241 nsew signal output
flabel metal2 s 17336 85936 17416 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[8]
port 242 nsew signal output
flabel metal2 s 17528 85936 17608 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_FrameStrobe_O[9]
port 243 nsew signal output
flabel metal2 s 1784 85936 1864 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[0]
port 244 nsew signal output
flabel metal2 s 1976 85936 2056 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[1]
port 245 nsew signal output
flabel metal2 s 2168 85936 2248 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[2]
port 246 nsew signal output
flabel metal2 s 2360 85936 2440 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N1BEG[3]
port 247 nsew signal output
flabel metal2 s 2552 85936 2632 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[0]
port 248 nsew signal output
flabel metal2 s 2744 85936 2824 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[1]
port 249 nsew signal output
flabel metal2 s 2936 85936 3016 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[2]
port 250 nsew signal output
flabel metal2 s 3128 85936 3208 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[3]
port 251 nsew signal output
flabel metal2 s 3320 85936 3400 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[4]
port 252 nsew signal output
flabel metal2 s 3512 85936 3592 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[5]
port 253 nsew signal output
flabel metal2 s 3704 85936 3784 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[6]
port 254 nsew signal output
flabel metal2 s 3896 85936 3976 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEG[7]
port 255 nsew signal output
flabel metal2 s 4088 85936 4168 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[0]
port 256 nsew signal output
flabel metal2 s 4280 85936 4360 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[1]
port 257 nsew signal output
flabel metal2 s 4472 85936 4552 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[2]
port 258 nsew signal output
flabel metal2 s 4664 85936 4744 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[3]
port 259 nsew signal output
flabel metal2 s 4856 85936 4936 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[4]
port 260 nsew signal output
flabel metal2 s 5048 85936 5128 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[5]
port 261 nsew signal output
flabel metal2 s 5240 85936 5320 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[6]
port 262 nsew signal output
flabel metal2 s 5432 85936 5512 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N2BEGb[7]
port 263 nsew signal output
flabel metal2 s 5624 85936 5704 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[0]
port 264 nsew signal output
flabel metal2 s 7544 85936 7624 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[10]
port 265 nsew signal output
flabel metal2 s 7736 85936 7816 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[11]
port 266 nsew signal output
flabel metal2 s 7928 85936 8008 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[12]
port 267 nsew signal output
flabel metal2 s 8120 85936 8200 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[13]
port 268 nsew signal output
flabel metal2 s 8312 85936 8392 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[14]
port 269 nsew signal output
flabel metal2 s 8504 85936 8584 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[15]
port 270 nsew signal output
flabel metal2 s 5816 85936 5896 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[1]
port 271 nsew signal output
flabel metal2 s 6008 85936 6088 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[2]
port 272 nsew signal output
flabel metal2 s 6200 85936 6280 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[3]
port 273 nsew signal output
flabel metal2 s 6392 85936 6472 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[4]
port 274 nsew signal output
flabel metal2 s 6584 85936 6664 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[5]
port 275 nsew signal output
flabel metal2 s 6776 85936 6856 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[6]
port 276 nsew signal output
flabel metal2 s 6968 85936 7048 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[7]
port 277 nsew signal output
flabel metal2 s 7160 85936 7240 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[8]
port 278 nsew signal output
flabel metal2 s 7352 85936 7432 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_N4BEG[9]
port 279 nsew signal output
flabel metal2 s 8696 85936 8776 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[0]
port 280 nsew signal input
flabel metal2 s 8888 85936 8968 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[1]
port 281 nsew signal input
flabel metal2 s 9080 85936 9160 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[2]
port 282 nsew signal input
flabel metal2 s 9272 85936 9352 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S1END[3]
port 283 nsew signal input
flabel metal2 s 11000 85936 11080 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[0]
port 284 nsew signal input
flabel metal2 s 11192 85936 11272 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[1]
port 285 nsew signal input
flabel metal2 s 11384 85936 11464 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[2]
port 286 nsew signal input
flabel metal2 s 11576 85936 11656 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[3]
port 287 nsew signal input
flabel metal2 s 11768 85936 11848 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[4]
port 288 nsew signal input
flabel metal2 s 11960 85936 12040 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[5]
port 289 nsew signal input
flabel metal2 s 12152 85936 12232 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[6]
port 290 nsew signal input
flabel metal2 s 12344 85936 12424 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2END[7]
port 291 nsew signal input
flabel metal2 s 9464 85936 9544 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[0]
port 292 nsew signal input
flabel metal2 s 9656 85936 9736 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[1]
port 293 nsew signal input
flabel metal2 s 9848 85936 9928 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[2]
port 294 nsew signal input
flabel metal2 s 10040 85936 10120 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[3]
port 295 nsew signal input
flabel metal2 s 10232 85936 10312 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[4]
port 296 nsew signal input
flabel metal2 s 10424 85936 10504 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[5]
port 297 nsew signal input
flabel metal2 s 10616 85936 10696 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[6]
port 298 nsew signal input
flabel metal2 s 10808 85936 10888 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S2MID[7]
port 299 nsew signal input
flabel metal2 s 12536 85936 12616 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[0]
port 300 nsew signal input
flabel metal2 s 14456 85936 14536 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[10]
port 301 nsew signal input
flabel metal2 s 14648 85936 14728 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[11]
port 302 nsew signal input
flabel metal2 s 14840 85936 14920 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[12]
port 303 nsew signal input
flabel metal2 s 15032 85936 15112 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[13]
port 304 nsew signal input
flabel metal2 s 15224 85936 15304 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[14]
port 305 nsew signal input
flabel metal2 s 15416 85936 15496 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[15]
port 306 nsew signal input
flabel metal2 s 12728 85936 12808 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[1]
port 307 nsew signal input
flabel metal2 s 12920 85936 13000 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[2]
port 308 nsew signal input
flabel metal2 s 13112 85936 13192 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[3]
port 309 nsew signal input
flabel metal2 s 13304 85936 13384 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[4]
port 310 nsew signal input
flabel metal2 s 13496 85936 13576 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[5]
port 311 nsew signal input
flabel metal2 s 13688 85936 13768 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[6]
port 312 nsew signal input
flabel metal2 s 13880 85936 13960 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[7]
port 313 nsew signal input
flabel metal2 s 14072 85936 14152 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[8]
port 314 nsew signal input
flabel metal2 s 14264 85936 14344 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_S4END[9]
port 315 nsew signal input
flabel metal2 s 15608 85936 15688 86016 0 FreeSans 320 0 0 0 Tile_X0Y0_UserCLKo
port 316 nsew signal output
flabel metal3 s 0 43052 80 43132 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[0]
port 317 nsew signal output
flabel metal3 s 0 43388 80 43468 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[1]
port 318 nsew signal output
flabel metal3 s 0 43724 80 43804 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[2]
port 319 nsew signal output
flabel metal3 s 0 44060 80 44140 0 FreeSans 320 0 0 0 Tile_X0Y0_W1BEG[3]
port 320 nsew signal output
flabel metal3 s 0 44396 80 44476 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[0]
port 321 nsew signal output
flabel metal3 s 0 44732 80 44812 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[1]
port 322 nsew signal output
flabel metal3 s 0 45068 80 45148 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[2]
port 323 nsew signal output
flabel metal3 s 0 45404 80 45484 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[3]
port 324 nsew signal output
flabel metal3 s 0 45740 80 45820 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[4]
port 325 nsew signal output
flabel metal3 s 0 46076 80 46156 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[5]
port 326 nsew signal output
flabel metal3 s 0 46412 80 46492 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[6]
port 327 nsew signal output
flabel metal3 s 0 46748 80 46828 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEG[7]
port 328 nsew signal output
flabel metal3 s 0 47084 80 47164 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[0]
port 329 nsew signal output
flabel metal3 s 0 47420 80 47500 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[1]
port 330 nsew signal output
flabel metal3 s 0 47756 80 47836 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[2]
port 331 nsew signal output
flabel metal3 s 0 48092 80 48172 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[3]
port 332 nsew signal output
flabel metal3 s 0 48428 80 48508 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[4]
port 333 nsew signal output
flabel metal3 s 0 48764 80 48844 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[5]
port 334 nsew signal output
flabel metal3 s 0 49100 80 49180 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[6]
port 335 nsew signal output
flabel metal3 s 0 49436 80 49516 0 FreeSans 320 0 0 0 Tile_X0Y0_W2BEGb[7]
port 336 nsew signal output
flabel metal3 s 0 55148 80 55228 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[0]
port 337 nsew signal output
flabel metal3 s 0 58508 80 58588 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[10]
port 338 nsew signal output
flabel metal3 s 0 58844 80 58924 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[11]
port 339 nsew signal output
flabel metal3 s 0 55484 80 55564 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[1]
port 340 nsew signal output
flabel metal3 s 0 55820 80 55900 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[2]
port 341 nsew signal output
flabel metal3 s 0 56156 80 56236 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[3]
port 342 nsew signal output
flabel metal3 s 0 56492 80 56572 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[4]
port 343 nsew signal output
flabel metal3 s 0 56828 80 56908 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[5]
port 344 nsew signal output
flabel metal3 s 0 57164 80 57244 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[6]
port 345 nsew signal output
flabel metal3 s 0 57500 80 57580 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[7]
port 346 nsew signal output
flabel metal3 s 0 57836 80 57916 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[8]
port 347 nsew signal output
flabel metal3 s 0 58172 80 58252 0 FreeSans 320 0 0 0 Tile_X0Y0_W6BEG[9]
port 348 nsew signal output
flabel metal3 s 0 49772 80 49852 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[0]
port 349 nsew signal output
flabel metal3 s 0 53132 80 53212 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[10]
port 350 nsew signal output
flabel metal3 s 0 53468 80 53548 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[11]
port 351 nsew signal output
flabel metal3 s 0 53804 80 53884 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[12]
port 352 nsew signal output
flabel metal3 s 0 54140 80 54220 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[13]
port 353 nsew signal output
flabel metal3 s 0 54476 80 54556 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[14]
port 354 nsew signal output
flabel metal3 s 0 54812 80 54892 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[15]
port 355 nsew signal output
flabel metal3 s 0 50108 80 50188 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[1]
port 356 nsew signal output
flabel metal3 s 0 50444 80 50524 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[2]
port 357 nsew signal output
flabel metal3 s 0 50780 80 50860 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[3]
port 358 nsew signal output
flabel metal3 s 0 51116 80 51196 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[4]
port 359 nsew signal output
flabel metal3 s 0 51452 80 51532 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[5]
port 360 nsew signal output
flabel metal3 s 0 51788 80 51868 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[6]
port 361 nsew signal output
flabel metal3 s 0 52124 80 52204 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[7]
port 362 nsew signal output
flabel metal3 s 0 52460 80 52540 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[8]
port 363 nsew signal output
flabel metal3 s 0 52796 80 52876 0 FreeSans 320 0 0 0 Tile_X0Y0_WW4BEG[9]
port 364 nsew signal output
flabel metal3 s 0 16172 80 16252 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[0]
port 365 nsew signal input
flabel metal3 s 0 16508 80 16588 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[1]
port 366 nsew signal input
flabel metal3 s 0 16844 80 16924 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[2]
port 367 nsew signal input
flabel metal3 s 0 17180 80 17260 0 FreeSans 320 0 0 0 Tile_X0Y1_E1END[3]
port 368 nsew signal input
flabel metal3 s 0 20204 80 20284 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[0]
port 369 nsew signal input
flabel metal3 s 0 20540 80 20620 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[1]
port 370 nsew signal input
flabel metal3 s 0 20876 80 20956 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[2]
port 371 nsew signal input
flabel metal3 s 0 21212 80 21292 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[3]
port 372 nsew signal input
flabel metal3 s 0 21548 80 21628 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[4]
port 373 nsew signal input
flabel metal3 s 0 21884 80 21964 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[5]
port 374 nsew signal input
flabel metal3 s 0 22220 80 22300 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[6]
port 375 nsew signal input
flabel metal3 s 0 22556 80 22636 0 FreeSans 320 0 0 0 Tile_X0Y1_E2END[7]
port 376 nsew signal input
flabel metal3 s 0 17516 80 17596 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[0]
port 377 nsew signal input
flabel metal3 s 0 17852 80 17932 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[1]
port 378 nsew signal input
flabel metal3 s 0 18188 80 18268 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[2]
port 379 nsew signal input
flabel metal3 s 0 18524 80 18604 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[3]
port 380 nsew signal input
flabel metal3 s 0 18860 80 18940 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[4]
port 381 nsew signal input
flabel metal3 s 0 19196 80 19276 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[5]
port 382 nsew signal input
flabel metal3 s 0 19532 80 19612 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[6]
port 383 nsew signal input
flabel metal3 s 0 19868 80 19948 0 FreeSans 320 0 0 0 Tile_X0Y1_E2MID[7]
port 384 nsew signal input
flabel metal3 s 0 28268 80 28348 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[0]
port 385 nsew signal input
flabel metal3 s 0 31628 80 31708 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[10]
port 386 nsew signal input
flabel metal3 s 0 31964 80 32044 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[11]
port 387 nsew signal input
flabel metal3 s 0 28604 80 28684 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[1]
port 388 nsew signal input
flabel metal3 s 0 28940 80 29020 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[2]
port 389 nsew signal input
flabel metal3 s 0 29276 80 29356 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[3]
port 390 nsew signal input
flabel metal3 s 0 29612 80 29692 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[4]
port 391 nsew signal input
flabel metal3 s 0 29948 80 30028 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[5]
port 392 nsew signal input
flabel metal3 s 0 30284 80 30364 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[6]
port 393 nsew signal input
flabel metal3 s 0 30620 80 30700 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[7]
port 394 nsew signal input
flabel metal3 s 0 30956 80 31036 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[8]
port 395 nsew signal input
flabel metal3 s 0 31292 80 31372 0 FreeSans 320 0 0 0 Tile_X0Y1_E6END[9]
port 396 nsew signal input
flabel metal3 s 0 22892 80 22972 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[0]
port 397 nsew signal input
flabel metal3 s 0 26252 80 26332 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[10]
port 398 nsew signal input
flabel metal3 s 0 26588 80 26668 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[11]
port 399 nsew signal input
flabel metal3 s 0 26924 80 27004 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[12]
port 400 nsew signal input
flabel metal3 s 0 27260 80 27340 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[13]
port 401 nsew signal input
flabel metal3 s 0 27596 80 27676 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[14]
port 402 nsew signal input
flabel metal3 s 0 27932 80 28012 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[15]
port 403 nsew signal input
flabel metal3 s 0 23228 80 23308 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[1]
port 404 nsew signal input
flabel metal3 s 0 23564 80 23644 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[2]
port 405 nsew signal input
flabel metal3 s 0 23900 80 23980 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[3]
port 406 nsew signal input
flabel metal3 s 0 24236 80 24316 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[4]
port 407 nsew signal input
flabel metal3 s 0 24572 80 24652 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[5]
port 408 nsew signal input
flabel metal3 s 0 24908 80 24988 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[6]
port 409 nsew signal input
flabel metal3 s 0 25244 80 25324 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[7]
port 410 nsew signal input
flabel metal3 s 0 25580 80 25660 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[8]
port 411 nsew signal input
flabel metal3 s 0 25916 80 25996 0 FreeSans 320 0 0 0 Tile_X0Y1_EE4END[9]
port 412 nsew signal input
flabel metal3 s 0 32300 80 32380 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[0]
port 413 nsew signal input
flabel metal3 s 0 35660 80 35740 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[10]
port 414 nsew signal input
flabel metal3 s 0 35996 80 36076 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[11]
port 415 nsew signal input
flabel metal3 s 0 36332 80 36412 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[12]
port 416 nsew signal input
flabel metal3 s 0 36668 80 36748 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[13]
port 417 nsew signal input
flabel metal3 s 0 37004 80 37084 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[14]
port 418 nsew signal input
flabel metal3 s 0 37340 80 37420 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[15]
port 419 nsew signal input
flabel metal3 s 0 37676 80 37756 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[16]
port 420 nsew signal input
flabel metal3 s 0 38012 80 38092 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[17]
port 421 nsew signal input
flabel metal3 s 0 38348 80 38428 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[18]
port 422 nsew signal input
flabel metal3 s 0 38684 80 38764 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[19]
port 423 nsew signal input
flabel metal3 s 0 32636 80 32716 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[1]
port 424 nsew signal input
flabel metal3 s 0 39020 80 39100 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[20]
port 425 nsew signal input
flabel metal3 s 0 39356 80 39436 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[21]
port 426 nsew signal input
flabel metal3 s 0 39692 80 39772 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[22]
port 427 nsew signal input
flabel metal3 s 0 40028 80 40108 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[23]
port 428 nsew signal input
flabel metal3 s 0 40364 80 40444 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[24]
port 429 nsew signal input
flabel metal3 s 0 40700 80 40780 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[25]
port 430 nsew signal input
flabel metal3 s 0 41036 80 41116 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[26]
port 431 nsew signal input
flabel metal3 s 0 41372 80 41452 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[27]
port 432 nsew signal input
flabel metal3 s 0 41708 80 41788 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[28]
port 433 nsew signal input
flabel metal3 s 0 42044 80 42124 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[29]
port 434 nsew signal input
flabel metal3 s 0 32972 80 33052 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[2]
port 435 nsew signal input
flabel metal3 s 0 42380 80 42460 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[30]
port 436 nsew signal input
flabel metal3 s 0 42716 80 42796 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[31]
port 437 nsew signal input
flabel metal3 s 0 33308 80 33388 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[3]
port 438 nsew signal input
flabel metal3 s 0 33644 80 33724 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[4]
port 439 nsew signal input
flabel metal3 s 0 33980 80 34060 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[5]
port 440 nsew signal input
flabel metal3 s 0 34316 80 34396 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[6]
port 441 nsew signal input
flabel metal3 s 0 34652 80 34732 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[7]
port 442 nsew signal input
flabel metal3 s 0 34988 80 35068 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[8]
port 443 nsew signal input
flabel metal3 s 0 35324 80 35404 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData[9]
port 444 nsew signal input
flabel metal3 s 21424 62036 21504 62116 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[0]
port 445 nsew signal output
flabel metal3 s 21424 65396 21504 65476 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[10]
port 446 nsew signal output
flabel metal3 s 21424 65732 21504 65812 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[11]
port 447 nsew signal output
flabel metal3 s 21424 66068 21504 66148 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[12]
port 448 nsew signal output
flabel metal3 s 21424 66404 21504 66484 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[13]
port 449 nsew signal output
flabel metal3 s 21424 66740 21504 66820 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[14]
port 450 nsew signal output
flabel metal3 s 21424 67076 21504 67156 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[15]
port 451 nsew signal output
flabel metal3 s 21424 67412 21504 67492 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[16]
port 452 nsew signal output
flabel metal3 s 21424 67748 21504 67828 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[17]
port 453 nsew signal output
flabel metal3 s 21424 68084 21504 68164 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[18]
port 454 nsew signal output
flabel metal3 s 21424 68420 21504 68500 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[19]
port 455 nsew signal output
flabel metal3 s 21424 62372 21504 62452 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[1]
port 456 nsew signal output
flabel metal3 s 21424 68756 21504 68836 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[20]
port 457 nsew signal output
flabel metal3 s 21424 69092 21504 69172 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[21]
port 458 nsew signal output
flabel metal3 s 21424 69428 21504 69508 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[22]
port 459 nsew signal output
flabel metal3 s 21424 69764 21504 69844 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[23]
port 460 nsew signal output
flabel metal3 s 21424 70100 21504 70180 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[24]
port 461 nsew signal output
flabel metal3 s 21424 70436 21504 70516 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[25]
port 462 nsew signal output
flabel metal3 s 21424 70772 21504 70852 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[26]
port 463 nsew signal output
flabel metal3 s 21424 71108 21504 71188 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[27]
port 464 nsew signal output
flabel metal3 s 21424 71444 21504 71524 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[28]
port 465 nsew signal output
flabel metal3 s 21424 71780 21504 71860 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[29]
port 466 nsew signal output
flabel metal3 s 21424 62708 21504 62788 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[2]
port 467 nsew signal output
flabel metal3 s 21424 72116 21504 72196 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[30]
port 468 nsew signal output
flabel metal3 s 21424 72452 21504 72532 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[31]
port 469 nsew signal output
flabel metal3 s 21424 63044 21504 63124 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[3]
port 470 nsew signal output
flabel metal3 s 21424 63380 21504 63460 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[4]
port 471 nsew signal output
flabel metal3 s 21424 63716 21504 63796 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[5]
port 472 nsew signal output
flabel metal3 s 21424 64052 21504 64132 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[6]
port 473 nsew signal output
flabel metal3 s 21424 64388 21504 64468 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[7]
port 474 nsew signal output
flabel metal3 s 21424 64724 21504 64804 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[8]
port 475 nsew signal output
flabel metal3 s 21424 65060 21504 65140 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameData_O[9]
port 476 nsew signal output
flabel metal2 s 15800 0 15880 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[0]
port 477 nsew signal input
flabel metal2 s 17720 0 17800 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[10]
port 478 nsew signal input
flabel metal2 s 17912 0 17992 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[11]
port 479 nsew signal input
flabel metal2 s 18104 0 18184 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[12]
port 480 nsew signal input
flabel metal2 s 18296 0 18376 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[13]
port 481 nsew signal input
flabel metal2 s 18488 0 18568 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[14]
port 482 nsew signal input
flabel metal2 s 18680 0 18760 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[15]
port 483 nsew signal input
flabel metal2 s 18872 0 18952 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[16]
port 484 nsew signal input
flabel metal2 s 19064 0 19144 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[17]
port 485 nsew signal input
flabel metal2 s 19256 0 19336 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[18]
port 486 nsew signal input
flabel metal2 s 19448 0 19528 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[19]
port 487 nsew signal input
flabel metal2 s 15992 0 16072 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[1]
port 488 nsew signal input
flabel metal2 s 16184 0 16264 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[2]
port 489 nsew signal input
flabel metal2 s 16376 0 16456 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[3]
port 490 nsew signal input
flabel metal2 s 16568 0 16648 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[4]
port 491 nsew signal input
flabel metal2 s 16760 0 16840 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[5]
port 492 nsew signal input
flabel metal2 s 16952 0 17032 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[6]
port 493 nsew signal input
flabel metal2 s 17144 0 17224 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[7]
port 494 nsew signal input
flabel metal2 s 17336 0 17416 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[8]
port 495 nsew signal input
flabel metal2 s 17528 0 17608 80 0 FreeSans 320 0 0 0 Tile_X0Y1_FrameStrobe[9]
port 496 nsew signal input
flabel metal2 s 1784 0 1864 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[0]
port 497 nsew signal input
flabel metal2 s 1976 0 2056 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[1]
port 498 nsew signal input
flabel metal2 s 2168 0 2248 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[2]
port 499 nsew signal input
flabel metal2 s 2360 0 2440 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N1END[3]
port 500 nsew signal input
flabel metal2 s 4088 0 4168 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[0]
port 501 nsew signal input
flabel metal2 s 4280 0 4360 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[1]
port 502 nsew signal input
flabel metal2 s 4472 0 4552 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[2]
port 503 nsew signal input
flabel metal2 s 4664 0 4744 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[3]
port 504 nsew signal input
flabel metal2 s 4856 0 4936 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[4]
port 505 nsew signal input
flabel metal2 s 5048 0 5128 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[5]
port 506 nsew signal input
flabel metal2 s 5240 0 5320 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[6]
port 507 nsew signal input
flabel metal2 s 5432 0 5512 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2END[7]
port 508 nsew signal input
flabel metal2 s 2552 0 2632 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[0]
port 509 nsew signal input
flabel metal2 s 2744 0 2824 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[1]
port 510 nsew signal input
flabel metal2 s 2936 0 3016 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[2]
port 511 nsew signal input
flabel metal2 s 3128 0 3208 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[3]
port 512 nsew signal input
flabel metal2 s 3320 0 3400 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[4]
port 513 nsew signal input
flabel metal2 s 3512 0 3592 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[5]
port 514 nsew signal input
flabel metal2 s 3704 0 3784 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[6]
port 515 nsew signal input
flabel metal2 s 3896 0 3976 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N2MID[7]
port 516 nsew signal input
flabel metal2 s 5624 0 5704 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[0]
port 517 nsew signal input
flabel metal2 s 7544 0 7624 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[10]
port 518 nsew signal input
flabel metal2 s 7736 0 7816 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[11]
port 519 nsew signal input
flabel metal2 s 7928 0 8008 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[12]
port 520 nsew signal input
flabel metal2 s 8120 0 8200 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[13]
port 521 nsew signal input
flabel metal2 s 8312 0 8392 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[14]
port 522 nsew signal input
flabel metal2 s 8504 0 8584 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[15]
port 523 nsew signal input
flabel metal2 s 5816 0 5896 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[1]
port 524 nsew signal input
flabel metal2 s 6008 0 6088 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[2]
port 525 nsew signal input
flabel metal2 s 6200 0 6280 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[3]
port 526 nsew signal input
flabel metal2 s 6392 0 6472 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[4]
port 527 nsew signal input
flabel metal2 s 6584 0 6664 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[5]
port 528 nsew signal input
flabel metal2 s 6776 0 6856 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[6]
port 529 nsew signal input
flabel metal2 s 6968 0 7048 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[7]
port 530 nsew signal input
flabel metal2 s 7160 0 7240 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[8]
port 531 nsew signal input
flabel metal2 s 7352 0 7432 80 0 FreeSans 320 0 0 0 Tile_X0Y1_N4END[9]
port 532 nsew signal input
flabel metal2 s 8696 0 8776 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[0]
port 533 nsew signal output
flabel metal2 s 8888 0 8968 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[1]
port 534 nsew signal output
flabel metal2 s 9080 0 9160 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[2]
port 535 nsew signal output
flabel metal2 s 9272 0 9352 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S1BEG[3]
port 536 nsew signal output
flabel metal2 s 9464 0 9544 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[0]
port 537 nsew signal output
flabel metal2 s 9656 0 9736 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[1]
port 538 nsew signal output
flabel metal2 s 9848 0 9928 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[2]
port 539 nsew signal output
flabel metal2 s 10040 0 10120 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[3]
port 540 nsew signal output
flabel metal2 s 10232 0 10312 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[4]
port 541 nsew signal output
flabel metal2 s 10424 0 10504 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[5]
port 542 nsew signal output
flabel metal2 s 10616 0 10696 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[6]
port 543 nsew signal output
flabel metal2 s 10808 0 10888 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEG[7]
port 544 nsew signal output
flabel metal2 s 11000 0 11080 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[0]
port 545 nsew signal output
flabel metal2 s 11192 0 11272 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[1]
port 546 nsew signal output
flabel metal2 s 11384 0 11464 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[2]
port 547 nsew signal output
flabel metal2 s 11576 0 11656 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[3]
port 548 nsew signal output
flabel metal2 s 11768 0 11848 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[4]
port 549 nsew signal output
flabel metal2 s 11960 0 12040 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[5]
port 550 nsew signal output
flabel metal2 s 12152 0 12232 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[6]
port 551 nsew signal output
flabel metal2 s 12344 0 12424 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S2BEGb[7]
port 552 nsew signal output
flabel metal2 s 12536 0 12616 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[0]
port 553 nsew signal output
flabel metal2 s 14456 0 14536 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[10]
port 554 nsew signal output
flabel metal2 s 14648 0 14728 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[11]
port 555 nsew signal output
flabel metal2 s 14840 0 14920 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[12]
port 556 nsew signal output
flabel metal2 s 15032 0 15112 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[13]
port 557 nsew signal output
flabel metal2 s 15224 0 15304 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[14]
port 558 nsew signal output
flabel metal2 s 15416 0 15496 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[15]
port 559 nsew signal output
flabel metal2 s 12728 0 12808 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[1]
port 560 nsew signal output
flabel metal2 s 12920 0 13000 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[2]
port 561 nsew signal output
flabel metal2 s 13112 0 13192 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[3]
port 562 nsew signal output
flabel metal2 s 13304 0 13384 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[4]
port 563 nsew signal output
flabel metal2 s 13496 0 13576 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[5]
port 564 nsew signal output
flabel metal2 s 13688 0 13768 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[6]
port 565 nsew signal output
flabel metal2 s 13880 0 13960 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[7]
port 566 nsew signal output
flabel metal2 s 14072 0 14152 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[8]
port 567 nsew signal output
flabel metal2 s 14264 0 14344 80 0 FreeSans 320 0 0 0 Tile_X0Y1_S4BEG[9]
port 568 nsew signal output
flabel metal2 s 15608 0 15688 80 0 FreeSans 320 0 0 0 Tile_X0Y1_UserCLK
port 569 nsew signal input
flabel metal3 s 0 44 80 124 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[0]
port 570 nsew signal output
flabel metal3 s 0 380 80 460 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[1]
port 571 nsew signal output
flabel metal3 s 0 716 80 796 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[2]
port 572 nsew signal output
flabel metal3 s 0 1052 80 1132 0 FreeSans 320 0 0 0 Tile_X0Y1_W1BEG[3]
port 573 nsew signal output
flabel metal3 s 0 1388 80 1468 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[0]
port 574 nsew signal output
flabel metal3 s 0 1724 80 1804 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[1]
port 575 nsew signal output
flabel metal3 s 0 2060 80 2140 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[2]
port 576 nsew signal output
flabel metal3 s 0 2396 80 2476 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[3]
port 577 nsew signal output
flabel metal3 s 0 2732 80 2812 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[4]
port 578 nsew signal output
flabel metal3 s 0 3068 80 3148 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[5]
port 579 nsew signal output
flabel metal3 s 0 3404 80 3484 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[6]
port 580 nsew signal output
flabel metal3 s 0 3740 80 3820 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEG[7]
port 581 nsew signal output
flabel metal3 s 0 4076 80 4156 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[0]
port 582 nsew signal output
flabel metal3 s 0 4412 80 4492 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[1]
port 583 nsew signal output
flabel metal3 s 0 4748 80 4828 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[2]
port 584 nsew signal output
flabel metal3 s 0 5084 80 5164 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[3]
port 585 nsew signal output
flabel metal3 s 0 5420 80 5500 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[4]
port 586 nsew signal output
flabel metal3 s 0 5756 80 5836 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[5]
port 587 nsew signal output
flabel metal3 s 0 6092 80 6172 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[6]
port 588 nsew signal output
flabel metal3 s 0 6428 80 6508 0 FreeSans 320 0 0 0 Tile_X0Y1_W2BEGb[7]
port 589 nsew signal output
flabel metal3 s 0 12140 80 12220 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[0]
port 590 nsew signal output
flabel metal3 s 0 15500 80 15580 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[10]
port 591 nsew signal output
flabel metal3 s 0 15836 80 15916 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[11]
port 592 nsew signal output
flabel metal3 s 0 12476 80 12556 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[1]
port 593 nsew signal output
flabel metal3 s 0 12812 80 12892 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[2]
port 594 nsew signal output
flabel metal3 s 0 13148 80 13228 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[3]
port 595 nsew signal output
flabel metal3 s 0 13484 80 13564 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[4]
port 596 nsew signal output
flabel metal3 s 0 13820 80 13900 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[5]
port 597 nsew signal output
flabel metal3 s 0 14156 80 14236 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[6]
port 598 nsew signal output
flabel metal3 s 0 14492 80 14572 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[7]
port 599 nsew signal output
flabel metal3 s 0 14828 80 14908 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[8]
port 600 nsew signal output
flabel metal3 s 0 15164 80 15244 0 FreeSans 320 0 0 0 Tile_X0Y1_W6BEG[9]
port 601 nsew signal output
flabel metal3 s 0 6764 80 6844 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[0]
port 602 nsew signal output
flabel metal3 s 0 10124 80 10204 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[10]
port 603 nsew signal output
flabel metal3 s 0 10460 80 10540 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[11]
port 604 nsew signal output
flabel metal3 s 0 10796 80 10876 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[12]
port 605 nsew signal output
flabel metal3 s 0 11132 80 11212 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[13]
port 606 nsew signal output
flabel metal3 s 0 11468 80 11548 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[14]
port 607 nsew signal output
flabel metal3 s 0 11804 80 11884 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[15]
port 608 nsew signal output
flabel metal3 s 0 7100 80 7180 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[1]
port 609 nsew signal output
flabel metal3 s 0 7436 80 7516 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[2]
port 610 nsew signal output
flabel metal3 s 0 7772 80 7852 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[3]
port 611 nsew signal output
flabel metal3 s 0 8108 80 8188 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[4]
port 612 nsew signal output
flabel metal3 s 0 8444 80 8524 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[5]
port 613 nsew signal output
flabel metal3 s 0 8780 80 8860 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[6]
port 614 nsew signal output
flabel metal3 s 0 9116 80 9196 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[7]
port 615 nsew signal output
flabel metal3 s 0 9452 80 9532 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[8]
port 616 nsew signal output
flabel metal3 s 0 9788 80 9868 0 FreeSans 320 0 0 0 Tile_X0Y1_WW4BEG[9]
port 617 nsew signal output
flabel metal6 s 4892 0 5332 86016 0 FreeSans 2624 90 0 0 VGND
port 618 nsew ground bidirectional
flabel metal6 s 4892 0 5332 328 0 FreeSans 2624 0 0 0 VGND
port 618 nsew ground bidirectional
flabel metal6 s 4892 85688 5332 86016 0 FreeSans 2624 0 0 0 VGND
port 618 nsew ground bidirectional
flabel metal6 s 20012 0 20452 86016 0 FreeSans 2624 90 0 0 VGND
port 618 nsew ground bidirectional
flabel metal6 s 20012 0 20452 328 0 FreeSans 2624 0 0 0 VGND
port 618 nsew ground bidirectional
flabel metal6 s 20012 85688 20452 86016 0 FreeSans 2624 0 0 0 VGND
port 618 nsew ground bidirectional
flabel metal6 s 3652 0 4092 86016 0 FreeSans 2624 90 0 0 VPWR
port 619 nsew power bidirectional
flabel metal6 s 3652 0 4092 328 0 FreeSans 2624 0 0 0 VPWR
port 619 nsew power bidirectional
flabel metal6 s 3652 85688 4092 86016 0 FreeSans 2624 0 0 0 VPWR
port 619 nsew power bidirectional
flabel metal6 s 18772 0 19212 86016 0 FreeSans 2624 90 0 0 VPWR
port 619 nsew power bidirectional
flabel metal6 s 18772 0 19212 328 0 FreeSans 2624 0 0 0 VPWR
port 619 nsew power bidirectional
flabel metal6 s 18772 85688 19212 86016 0 FreeSans 2624 0 0 0 VPWR
port 619 nsew power bidirectional
flabel metal3 s 21424 49268 21504 49348 0 FreeSans 320 0 0 0 WEN_SRAM
port 620 nsew signal output
rlabel metal1 10802 83916 10802 83916 0 VGND
rlabel metal1 10752 84672 10752 84672 0 VPWR
rlabel metal2 12096 23604 12096 23604 0 ADDR_SRAM0
rlabel metal3 8208 23268 8208 23268 0 ADDR_SRAM1
rlabel metal3 14178 25116 14178 25116 0 ADDR_SRAM2
rlabel metal3 14208 36288 14208 36288 0 ADDR_SRAM3
rlabel metal3 20802 25788 20802 25788 0 ADDR_SRAM4
rlabel metal3 21426 26124 21426 26124 0 ADDR_SRAM5
rlabel metal3 21042 26460 21042 26460 0 ADDR_SRAM6
rlabel metal4 17088 31416 17088 31416 0 ADDR_SRAM7
rlabel metal3 21282 27132 21282 27132 0 ADDR_SRAM8
rlabel metal3 21186 27468 21186 27468 0 ADDR_SRAM9
rlabel metal3 21042 38556 21042 38556 0 BM_SRAM0
rlabel metal2 16560 35877 16560 35877 0 BM_SRAM1
rlabel metal3 21426 41916 21426 41916 0 BM_SRAM10
rlabel metal3 21234 42252 21234 42252 0 BM_SRAM11
rlabel metal3 20640 20160 20640 20160 0 BM_SRAM12
rlabel metal3 21186 42924 21186 42924 0 BM_SRAM13
rlabel metal4 20832 39942 20832 39942 0 BM_SRAM14
rlabel metal3 21426 43596 21426 43596 0 BM_SRAM15
rlabel metal3 15984 53004 15984 53004 0 BM_SRAM16
rlabel metal3 20994 44268 20994 44268 0 BM_SRAM17
rlabel metal3 21090 44604 21090 44604 0 BM_SRAM18
rlabel metal3 20784 74592 20784 74592 0 BM_SRAM19
rlabel metal3 21090 39228 21090 39228 0 BM_SRAM2
rlabel metal3 18192 65184 18192 65184 0 BM_SRAM20
rlabel metal2 17280 44436 17280 44436 0 BM_SRAM21
rlabel metal3 21138 45948 21138 45948 0 BM_SRAM22
rlabel metal4 19968 69342 19968 69342 0 BM_SRAM23
rlabel metal3 20802 46620 20802 46620 0 BM_SRAM24
rlabel metal2 19968 48006 19968 48006 0 BM_SRAM25
rlabel metal3 21186 47292 21186 47292 0 BM_SRAM26
rlabel metal3 20994 47628 20994 47628 0 BM_SRAM27
rlabel metal3 21378 47964 21378 47964 0 BM_SRAM28
rlabel metal2 17280 48594 17280 48594 0 BM_SRAM29
rlabel metal3 20802 39564 20802 39564 0 BM_SRAM3
rlabel metal3 21186 48636 21186 48636 0 BM_SRAM30
rlabel metal3 20928 54180 20928 54180 0 BM_SRAM31
rlabel metal2 20448 22176 20448 22176 0 BM_SRAM4
rlabel metal2 20400 33852 20400 33852 0 BM_SRAM5
rlabel metal3 21042 40572 21042 40572 0 BM_SRAM6
rlabel metal3 18144 40782 18144 40782 0 BM_SRAM7
rlabel metal3 21330 41244 21330 41244 0 BM_SRAM8
rlabel metal3 21282 41580 21282 41580 0 BM_SRAM9
rlabel metal2 19584 50232 19584 50232 0 CLK_SRAM
rlabel via3 21426 24108 21426 24108 0 CONFIGURED_top
rlabel metal2 19296 27258 19296 27258 0 DIN_SRAM0
rlabel metal3 19026 28140 19026 28140 0 DIN_SRAM1
rlabel metal3 21186 31164 21186 31164 0 DIN_SRAM10
rlabel metal3 21042 31500 21042 31500 0 DIN_SRAM11
rlabel metal2 20544 21882 20544 21882 0 DIN_SRAM12
rlabel metal3 20802 32172 20802 32172 0 DIN_SRAM13
rlabel metal3 21042 32508 21042 32508 0 DIN_SRAM14
rlabel metal3 21282 32844 21282 32844 0 DIN_SRAM15
rlabel metal2 16752 68964 16752 68964 0 DIN_SRAM16
rlabel metal3 21378 33516 21378 33516 0 DIN_SRAM17
rlabel metal3 21138 33852 21138 33852 0 DIN_SRAM18
rlabel metal2 20544 71106 20544 71106 0 DIN_SRAM19
rlabel metal2 11040 28854 11040 28854 0 DIN_SRAM2
rlabel metal3 21090 34524 21090 34524 0 DIN_SRAM20
rlabel metal3 20898 34860 20898 34860 0 DIN_SRAM21
rlabel metal3 21378 35196 21378 35196 0 DIN_SRAM22
rlabel metal3 21378 35532 21378 35532 0 DIN_SRAM23
rlabel metal3 19458 35868 19458 35868 0 DIN_SRAM24
rlabel metal3 21138 36204 21138 36204 0 DIN_SRAM25
rlabel metal3 21378 36540 21378 36540 0 DIN_SRAM26
rlabel metal3 21378 36876 21378 36876 0 DIN_SRAM27
rlabel metal3 20802 37212 20802 37212 0 DIN_SRAM28
rlabel metal3 19074 37548 19074 37548 0 DIN_SRAM29
rlabel metal3 20850 28812 20850 28812 0 DIN_SRAM3
rlabel metal2 19104 43680 19104 43680 0 DIN_SRAM30
rlabel metal3 19632 54180 19632 54180 0 DIN_SRAM31
rlabel metal3 20496 24696 20496 24696 0 DIN_SRAM4
rlabel metal3 21090 29484 21090 29484 0 DIN_SRAM5
rlabel metal3 20802 29820 20802 29820 0 DIN_SRAM6
rlabel metal3 19122 30156 19122 30156 0 DIN_SRAM7
rlabel metal2 19488 30114 19488 30114 0 DIN_SRAM8
rlabel metal2 16512 30996 16512 30996 0 DIN_SRAM9
rlabel metal2 13344 13692 13344 13692 0 DOUT_SRAM0
rlabel metal3 18240 12936 18240 12936 0 DOUT_SRAM1
rlabel metal3 18930 16716 18930 16716 0 DOUT_SRAM10
rlabel via3 21426 17052 21426 17052 0 DOUT_SRAM11
rlabel metal3 21042 17388 21042 17388 0 DOUT_SRAM12
rlabel metal2 6096 16296 6096 16296 0 DOUT_SRAM13
rlabel metal2 7776 13020 7776 13020 0 DOUT_SRAM14
rlabel metal4 18240 16926 18240 16926 0 DOUT_SRAM15
rlabel metal3 19170 18732 19170 18732 0 DOUT_SRAM16
rlabel metal3 20802 19068 20802 19068 0 DOUT_SRAM17
rlabel metal3 21138 19404 21138 19404 0 DOUT_SRAM18
rlabel metal3 21042 19740 21042 19740 0 DOUT_SRAM19
rlabel metal3 20850 14028 20850 14028 0 DOUT_SRAM2
rlabel metal3 15744 19992 15744 19992 0 DOUT_SRAM20
rlabel metal3 20994 20412 20994 20412 0 DOUT_SRAM21
rlabel metal3 21426 20748 21426 20748 0 DOUT_SRAM22
rlabel metal4 12048 28980 12048 28980 0 DOUT_SRAM23
rlabel metal3 15120 32760 15120 32760 0 DOUT_SRAM24
rlabel metal3 20802 21756 20802 21756 0 DOUT_SRAM25
rlabel metal3 20802 22092 20802 22092 0 DOUT_SRAM26
rlabel metal3 20802 22428 20802 22428 0 DOUT_SRAM27
rlabel metal3 15504 30240 15504 30240 0 DOUT_SRAM28
rlabel metal3 21234 23100 21234 23100 0 DOUT_SRAM29
rlabel metal3 20994 14364 20994 14364 0 DOUT_SRAM3
rlabel metal3 20994 23436 20994 23436 0 DOUT_SRAM30
rlabel metal4 576 39144 576 39144 0 DOUT_SRAM31
rlabel metal2 19824 13020 19824 13020 0 DOUT_SRAM4
rlabel metal2 2304 13986 2304 13986 0 DOUT_SRAM5
rlabel metal3 20802 15372 20802 15372 0 DOUT_SRAM6
rlabel metal2 15264 14742 15264 14742 0 DOUT_SRAM7
rlabel metal3 20994 16044 20994 16044 0 DOUT_SRAM8
rlabel metal3 16392 16380 16392 16380 0 DOUT_SRAM9
rlabel metal3 21090 49644 21090 49644 0 MEN_SRAM
rlabel metal3 20802 49980 20802 49980 0 REN_SRAM
rlabel metal3 21090 50652 21090 50652 0 TIE_HIGH_SRAM
rlabel metal3 20802 50988 20802 50988 0 TIE_LOW_SRAM
rlabel metal2 14400 65352 14400 65352 0 Tile_X0Y0_E1END[0]
rlabel metal2 15456 55104 15456 55104 0 Tile_X0Y0_E1END[1]
rlabel metal2 13824 53130 13824 53130 0 Tile_X0Y0_E1END[2]
rlabel metal3 17760 67620 17760 67620 0 Tile_X0Y0_E1END[3]
rlabel metal3 270 63252 270 63252 0 Tile_X0Y0_E2END[0]
rlabel metal2 4416 65268 4416 65268 0 Tile_X0Y0_E2END[1]
rlabel metal3 1290 63924 1290 63924 0 Tile_X0Y0_E2END[2]
rlabel metal3 270 64260 270 64260 0 Tile_X0Y0_E2END[3]
rlabel metal3 1134 64596 1134 64596 0 Tile_X0Y0_E2END[4]
rlabel metal2 2208 66654 2208 66654 0 Tile_X0Y0_E2END[5]
rlabel metal3 3360 65310 3360 65310 0 Tile_X0Y0_E2END[6]
rlabel metal3 798 65604 798 65604 0 Tile_X0Y0_E2END[7]
rlabel metal3 174 60564 174 60564 0 Tile_X0Y0_E2MID[0]
rlabel metal3 126 60900 126 60900 0 Tile_X0Y0_E2MID[1]
rlabel metal2 1536 62034 1536 62034 0 Tile_X0Y0_E2MID[2]
rlabel metal3 1422 61572 1422 61572 0 Tile_X0Y0_E2MID[3]
rlabel metal3 126 61908 126 61908 0 Tile_X0Y0_E2MID[4]
rlabel metal2 1824 68418 1824 68418 0 Tile_X0Y0_E2MID[5]
rlabel metal3 654 62580 654 62580 0 Tile_X0Y0_E2MID[6]
rlabel metal2 1680 68628 1680 68628 0 Tile_X0Y0_E2MID[7]
rlabel metal3 702 71316 702 71316 0 Tile_X0Y0_E6END[0]
rlabel metal2 2304 68082 2304 68082 0 Tile_X0Y0_E6END[10]
rlabel metal3 654 75012 654 75012 0 Tile_X0Y0_E6END[11]
rlabel metal3 702 71652 702 71652 0 Tile_X0Y0_E6END[1]
rlabel metal2 18624 66276 18624 66276 0 Tile_X0Y0_E6END[2]
rlabel metal2 19200 72240 19200 72240 0 Tile_X0Y0_E6END[3]
rlabel metal2 12912 71484 12912 71484 0 Tile_X0Y0_E6END[4]
rlabel metal2 1440 72240 1440 72240 0 Tile_X0Y0_E6END[5]
rlabel metal3 14400 54768 14400 54768 0 Tile_X0Y0_E6END[6]
rlabel metal3 18672 69972 18672 69972 0 Tile_X0Y0_E6END[7]
rlabel metal2 16320 72576 16320 72576 0 Tile_X0Y0_E6END[8]
rlabel metal3 12576 49854 12576 49854 0 Tile_X0Y0_E6END[9]
rlabel metal2 15840 71904 15840 71904 0 Tile_X0Y0_EE4END[0]
rlabel metal3 1230 69300 1230 69300 0 Tile_X0Y0_EE4END[10]
rlabel metal2 19008 72114 19008 72114 0 Tile_X0Y0_EE4END[11]
rlabel metal3 78 69972 78 69972 0 Tile_X0Y0_EE4END[12]
rlabel metal3 510 70308 510 70308 0 Tile_X0Y0_EE4END[13]
rlabel metal3 558 70644 558 70644 0 Tile_X0Y0_EE4END[14]
rlabel metal3 16800 71316 16800 71316 0 Tile_X0Y0_EE4END[15]
rlabel metal3 624 51744 624 51744 0 Tile_X0Y0_EE4END[1]
rlabel metal2 18048 63126 18048 63126 0 Tile_X0Y0_EE4END[2]
rlabel metal2 18528 78992 18528 78992 0 Tile_X0Y0_EE4END[3]
rlabel via2 78 67284 78 67284 0 Tile_X0Y0_EE4END[4]
rlabel metal3 1296 49980 1296 49980 0 Tile_X0Y0_EE4END[5]
rlabel metal3 174 67956 174 67956 0 Tile_X0Y0_EE4END[6]
rlabel metal2 18432 67956 18432 67956 0 Tile_X0Y0_EE4END[7]
rlabel metal2 16224 71904 16224 71904 0 Tile_X0Y0_EE4END[8]
rlabel metal3 126 68964 126 68964 0 Tile_X0Y0_EE4END[9]
rlabel metal3 1680 70644 1680 70644 0 Tile_X0Y0_FrameData[0]
rlabel metal2 1344 46368 1344 46368 0 Tile_X0Y0_FrameData[10]
rlabel via2 12000 49644 12000 49644 0 Tile_X0Y0_FrameData[11]
rlabel metal3 414 79380 414 79380 0 Tile_X0Y0_FrameData[12]
rlabel metal2 14880 67662 14880 67662 0 Tile_X0Y0_FrameData[13]
rlabel metal2 13968 72324 13968 72324 0 Tile_X0Y0_FrameData[14]
rlabel metal3 654 80388 654 80388 0 Tile_X0Y0_FrameData[15]
rlabel metal3 19248 50316 19248 50316 0 Tile_X0Y0_FrameData[16]
rlabel metal2 18336 50904 18336 50904 0 Tile_X0Y0_FrameData[17]
rlabel metal4 1920 48510 1920 48510 0 Tile_X0Y0_FrameData[18]
rlabel metal3 13536 72408 13536 72408 0 Tile_X0Y0_FrameData[19]
rlabel metal2 15360 76608 15360 76608 0 Tile_X0Y0_FrameData[1]
rlabel metal3 462 82068 462 82068 0 Tile_X0Y0_FrameData[20]
rlabel metal3 2496 82740 2496 82740 0 Tile_X0Y0_FrameData[21]
rlabel metal3 1230 82740 1230 82740 0 Tile_X0Y0_FrameData[22]
rlabel metal2 13248 68838 13248 68838 0 Tile_X0Y0_FrameData[23]
rlabel metal2 14448 50316 14448 50316 0 Tile_X0Y0_FrameData[24]
rlabel metal2 17760 48552 17760 48552 0 Tile_X0Y0_FrameData[25]
rlabel metal2 1488 52500 1488 52500 0 Tile_X0Y0_FrameData[26]
rlabel metal2 12720 50988 12720 50988 0 Tile_X0Y0_FrameData[27]
rlabel metal3 13440 83664 13440 83664 0 Tile_X0Y0_FrameData[28]
rlabel metal2 1440 66192 1440 66192 0 Tile_X0Y0_FrameData[29]
rlabel metal2 2016 45276 2016 45276 0 Tile_X0Y0_FrameData[2]
rlabel metal2 13440 71148 13440 71148 0 Tile_X0Y0_FrameData[30]
rlabel metal2 2112 84126 2112 84126 0 Tile_X0Y0_FrameData[31]
rlabel metal2 12960 47166 12960 47166 0 Tile_X0Y0_FrameData[3]
rlabel metal2 1248 69888 1248 69888 0 Tile_X0Y0_FrameData[4]
rlabel metal2 13248 53970 13248 53970 0 Tile_X0Y0_FrameData[5]
rlabel metal2 1392 82068 1392 82068 0 Tile_X0Y0_FrameData[6]
rlabel metal2 1344 82488 1344 82488 0 Tile_X0Y0_FrameData[7]
rlabel metal3 1824 69132 1824 69132 0 Tile_X0Y0_FrameData[8]
rlabel metal2 1872 67620 1872 67620 0 Tile_X0Y0_FrameData[9]
rlabel metal3 21282 51324 21282 51324 0 Tile_X0Y0_FrameData_O[0]
rlabel metal2 19968 55062 19968 55062 0 Tile_X0Y0_FrameData_O[10]
rlabel metal3 20706 55020 20706 55020 0 Tile_X0Y0_FrameData_O[11]
rlabel metal3 21090 55356 21090 55356 0 Tile_X0Y0_FrameData_O[12]
rlabel metal3 20994 55692 20994 55692 0 Tile_X0Y0_FrameData_O[13]
rlabel metal2 19680 56784 19680 56784 0 Tile_X0Y0_FrameData_O[14]
rlabel metal3 20802 56364 20802 56364 0 Tile_X0Y0_FrameData_O[15]
rlabel metal3 21090 56700 21090 56700 0 Tile_X0Y0_FrameData_O[16]
rlabel metal3 21090 57036 21090 57036 0 Tile_X0Y0_FrameData_O[17]
rlabel metal3 21090 57372 21090 57372 0 Tile_X0Y0_FrameData_O[18]
rlabel metal3 20802 57708 20802 57708 0 Tile_X0Y0_FrameData_O[19]
rlabel metal3 20802 51660 20802 51660 0 Tile_X0Y0_FrameData_O[1]
rlabel metal4 19872 59766 19872 59766 0 Tile_X0Y0_FrameData_O[20]
rlabel metal3 19458 58380 19458 58380 0 Tile_X0Y0_FrameData_O[21]
rlabel metal2 19872 60144 19872 60144 0 Tile_X0Y0_FrameData_O[22]
rlabel metal3 17568 59094 17568 59094 0 Tile_X0Y0_FrameData_O[23]
rlabel metal3 21378 59388 21378 59388 0 Tile_X0Y0_FrameData_O[24]
rlabel metal3 21138 59724 21138 59724 0 Tile_X0Y0_FrameData_O[25]
rlabel metal2 16800 59976 16800 59976 0 Tile_X0Y0_FrameData_O[26]
rlabel metal2 17568 60354 17568 60354 0 Tile_X0Y0_FrameData_O[27]
rlabel metal2 17184 60522 17184 60522 0 Tile_X0Y0_FrameData_O[28]
rlabel metal3 19872 64428 19872 64428 0 Tile_X0Y0_FrameData_O[29]
rlabel metal2 19584 52164 19584 52164 0 Tile_X0Y0_FrameData_O[2]
rlabel metal3 21138 61404 21138 61404 0 Tile_X0Y0_FrameData_O[30]
rlabel metal3 18786 61740 18786 61740 0 Tile_X0Y0_FrameData_O[31]
rlabel metal3 20706 52332 20706 52332 0 Tile_X0Y0_FrameData_O[3]
rlabel metal3 20802 52668 20802 52668 0 Tile_X0Y0_FrameData_O[4]
rlabel metal2 19872 53424 19872 53424 0 Tile_X0Y0_FrameData_O[5]
rlabel metal3 20802 53340 20802 53340 0 Tile_X0Y0_FrameData_O[6]
rlabel metal3 20994 53676 20994 53676 0 Tile_X0Y0_FrameData_O[7]
rlabel metal3 20850 54012 20850 54012 0 Tile_X0Y0_FrameData_O[8]
rlabel metal2 17856 54264 17856 54264 0 Tile_X0Y0_FrameData_O[9]
rlabel metal2 20064 84504 20064 84504 0 Tile_X0Y0_FrameStrobe_O[0]
rlabel metal3 18336 84504 18336 84504 0 Tile_X0Y0_FrameStrobe_O[10]
rlabel metal3 18624 84420 18624 84420 0 Tile_X0Y0_FrameStrobe_O[11]
rlabel metal2 20064 83076 20064 83076 0 Tile_X0Y0_FrameStrobe_O[12]
rlabel metal3 19008 84084 19008 84084 0 Tile_X0Y0_FrameStrobe_O[13]
rlabel metal2 19968 84000 19968 84000 0 Tile_X0Y0_FrameStrobe_O[14]
rlabel metal2 18720 85314 18720 85314 0 Tile_X0Y0_FrameStrobe_O[15]
rlabel metal2 18912 85398 18912 85398 0 Tile_X0Y0_FrameStrobe_O[16]
rlabel metal2 19104 85482 19104 85482 0 Tile_X0Y0_FrameStrobe_O[17]
rlabel metal2 13152 84798 13152 84798 0 Tile_X0Y0_FrameStrobe_O[18]
rlabel metal4 12384 84126 12384 84126 0 Tile_X0Y0_FrameStrobe_O[19]
rlabel metal2 19584 84294 19584 84294 0 Tile_X0Y0_FrameStrobe_O[1]
rlabel metal2 16224 85440 16224 85440 0 Tile_X0Y0_FrameStrobe_O[2]
rlabel metal3 17136 78456 17136 78456 0 Tile_X0Y0_FrameStrobe_O[3]
rlabel metal2 16608 85188 16608 85188 0 Tile_X0Y0_FrameStrobe_O[4]
rlabel metal3 16656 65268 16656 65268 0 Tile_X0Y0_FrameStrobe_O[5]
rlabel metal2 16992 85188 16992 85188 0 Tile_X0Y0_FrameStrobe_O[6]
rlabel metal2 17568 77952 17568 77952 0 Tile_X0Y0_FrameStrobe_O[7]
rlabel metal2 17376 84558 17376 84558 0 Tile_X0Y0_FrameStrobe_O[8]
rlabel metal2 17568 83928 17568 83928 0 Tile_X0Y0_FrameStrobe_O[9]
rlabel metal3 9936 74508 9936 74508 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 11808 74757 11808 74757 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 6240 67921 6240 67921 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit10.Q
rlabel metal2 4704 67704 4704 67704 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit11.Q
rlabel metal3 4512 71484 4512 71484 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 5856 71733 5856 71733 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 3264 83160 3264 83160 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 4896 82236 4896 82236 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 9024 80805 9024 80805 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 7488 80430 7488 80430 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit17.Q
rlabel metal2 6240 82359 6240 82359 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 4704 82110 4704 82110 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 12672 46410 12672 46410 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 8304 82803 8304 82803 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 6720 83034 6720 83034 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit21.Q
rlabel metal3 11712 82992 11712 82992 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 10032 83580 10032 83580 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 9984 73038 9984 73038 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 10128 73668 10128 73668 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 15037 60724 15037 60724 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 14112 59640 14112 59640 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 11808 71652 11808 71652 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 11616 71358 11616 71358 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 14352 47040 14352 47040 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 15936 76062 15936 76062 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 15744 76272 15744 76272 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 11088 69384 11088 69384 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 12672 69671 12672 69671 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 14928 77700 14928 77700 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit6.Q
rlabel metal2 16896 78757 16896 78757 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit7.Q
rlabel metal2 3552 80136 3552 80136 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 5472 80808 5472 80808 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame0_bit9.Q
rlabel metal3 6192 65940 6192 65940 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit0.Q
rlabel metal3 6720 66108 6720 66108 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 12816 49476 12816 49476 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit10.Q
rlabel via1 14544 49480 14544 49480 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 11520 66990 11520 66990 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit12.Q
rlabel via1 13104 66943 13104 66943 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 13824 80598 13824 80598 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 15360 80805 15360 80805 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit15.Q
rlabel metal3 9936 78204 9936 78204 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit16.Q
rlabel via2 12096 78206 12096 78206 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 12768 47922 12768 47922 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit18.Q
rlabel metal2 14304 48265 14304 48265 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 9216 65646 9216 65646 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 11520 67914 11520 67914 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 13056 67921 13056 67921 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit21.Q
rlabel metal2 13824 82740 13824 82740 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 15456 83041 15456 83041 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 10656 79128 10656 79128 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit24.Q
rlabel via1 12240 79039 12240 79039 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 12576 50274 12576 50274 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit26.Q
rlabel via1 14160 50311 14160 50311 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 11136 65478 11136 65478 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 12672 65685 12672 65685 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 9312 65310 9312 65310 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 14496 82110 14496 82110 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 16032 82611 16032 82611 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 7104 75936 7104 75936 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 6816 76272 6816 76272 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 2208 76650 2208 76650 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit6.Q
rlabel metal2 1920 77574 1920 77574 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit7.Q
rlabel metal2 10752 77574 10752 77574 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 12528 76860 12528 76860 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 18864 45948 18864 45948 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 20016 45192 20016 45192 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 17856 57330 17856 57330 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 19392 57715 19392 57715 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit11.Q
rlabel metal2 18240 71526 18240 71526 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 19920 71484 19920 71484 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit13.Q
rlabel metal2 15744 72902 15744 72902 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit14.Q
rlabel metal3 17472 72996 17472 72996 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 18048 49980 18048 49980 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 19632 49539 19632 49539 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 17808 60060 17808 60060 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 19440 60123 19440 60123 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 17952 63168 17952 63168 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit2.Q
rlabel metal3 18432 81060 18432 81060 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 19968 77371 19968 77371 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 14304 65688 14304 65688 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit22.Q
rlabel via1 15888 65431 15888 65431 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit23.Q
rlabel metal3 15744 48804 15744 48804 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit24.Q
rlabel via1 17136 48799 17136 48799 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 17376 52458 17376 52458 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 18912 52287 18912 52287 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 17952 68334 17952 68334 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit28.Q
rlabel metal3 19680 71064 19680 71064 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 19680 65940 19680 65940 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 7008 73584 7008 73584 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 7584 72996 7584 72996 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 18768 78372 18768 78372 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 20736 78162 20736 78162 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 17424 65436 17424 65436 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 19008 65811 19008 65811 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit7.Q
rlabel metal2 15456 44216 15456 44216 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit8.Q
rlabel metal2 16992 44559 16992 44559 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame2_bit9.Q
rlabel metal3 18144 47292 18144 47292 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 19968 44436 19968 44436 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 17856 55020 17856 55020 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 19392 55143 19392 55143 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit11.Q
rlabel metal3 18192 69636 18192 69636 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit12.Q
rlabel metal3 19680 69804 19680 69804 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 15696 72660 15696 72660 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 17664 75684 17664 75684 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 18000 48804 18000 48804 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit16.Q
rlabel via1 19632 48799 19632 48799 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 17760 59388 17760 59388 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit18.Q
rlabel via1 19440 59383 19440 59383 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 17856 62412 17856 62412 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 18288 81816 18288 81816 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 18720 82992 18720 82992 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 14400 67578 14400 67578 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 15936 67071 15936 67071 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 15456 47544 15456 47544 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 16992 47541 16992 47541 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit25.Q
rlabel metal2 17472 52458 17472 52458 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 19008 52591 19008 52591 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 17568 70518 17568 70518 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 19488 67239 19488 67239 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit29.Q
rlabel metal3 18768 65520 18768 65520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 14976 70014 14976 70014 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 16512 70599 16512 70599 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit31.Q
rlabel metal3 18192 73500 18192 73500 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit4.Q
rlabel metal3 19968 73164 19968 73164 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 17424 64596 17424 64596 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit6.Q
rlabel via1 19152 64600 19152 64600 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 15264 43890 15264 43890 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 17040 45003 17040 45003 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 8064 53760 8064 53760 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 9648 54075 9648 54075 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 11520 55272 11520 55272 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 13200 55020 13200 55020 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit11.Q
rlabel metal3 13680 78204 13680 78204 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 14880 78505 14880 78505 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 13104 57099 13104 57099 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 11520 57339 11520 57339 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit15.Q
rlabel via1 9840 55528 9840 55528 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit16.Q
rlabel metal3 8112 55356 8112 55356 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 4032 53382 4032 53382 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit18.Q
rlabel via1 5616 53335 5616 53335 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit19.Q
rlabel metal3 3648 44268 3648 44268 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 6624 60354 6624 60354 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 8208 60123 8208 60123 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit21.Q
rlabel metal2 13344 63385 13344 63385 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 11808 63387 11808 63387 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 9504 58125 9504 58125 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 7968 58128 7968 58128 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 5184 56403 5184 56403 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 3648 56406 3648 56406 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 4896 62493 4896 62493 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit28.Q
rlabel metal2 3360 62464 3360 62464 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit29.Q
rlabel via1 5424 44263 5424 44263 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 14976 69258 14976 69258 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 16512 69475 16512 69475 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 4704 62412 4704 62412 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 3168 62293 3168 62293 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 11520 75474 11520 75474 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 13056 75229 13056 75229 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 11424 53382 11424 53382 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 13152 53589 13152 53589 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 6240 47544 6240 47544 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit0.Q
rlabel via1 7824 47287 7824 47287 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 10368 47544 10368 47544 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit10.Q
rlabel via1 11952 47287 11952 47287 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 6048 63042 6048 63042 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 7584 63385 7584 63385 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit13.Q
rlabel metal2 9600 56616 9600 56616 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit14.Q
rlabel metal2 10368 56403 10368 56403 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 6528 51996 6528 51996 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 8016 51240 8016 51240 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit17.Q
rlabel metal2 4032 51114 4032 51114 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit18.Q
rlabel metal3 5616 50484 5616 50484 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 3600 44100 3600 44100 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 6336 60018 6336 60018 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 7872 59889 7872 59889 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 13776 56448 13776 56448 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit22.Q
rlabel via2 15071 57045 15071 57045 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 8352 52458 8352 52458 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 9888 52801 9888 52801 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 3264 52458 3264 52458 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 4608 52038 4608 52038 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 4704 60060 4704 60060 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 3168 60015 3168 60015 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit29.Q
rlabel metal2 5448 44982 5448 44982 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit3.Q
rlabel metal3 9984 63084 9984 63084 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit30.Q
rlabel metal3 10992 63084 10992 63084 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 4224 55104 4224 55104 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit4.Q
rlabel metal3 3360 54180 3360 54180 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit5.Q
rlabel metal2 14112 64344 14112 64344 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit6.Q
rlabel metal3 15744 64428 15744 64428 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 9984 51534 9984 51534 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit8.Q
rlabel metal3 11808 51282 11808 51282 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame5_bit9.Q
rlabel via1 13584 44263 13584 44263 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 12000 44310 12000 44310 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit1.Q
rlabel metal2 2784 47292 2784 47292 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 4320 48265 4320 48265 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit11.Q
rlabel metal2 3552 57918 3552 57918 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 5088 57915 5088 57915 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit13.Q
rlabel metal2 10080 59430 10080 59430 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 11568 58800 11568 58800 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit15.Q
rlabel metal2 5952 49056 5952 49056 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit16.Q
rlabel metal2 7488 49431 7488 49431 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 3840 47334 3840 47334 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit18.Q
rlabel via1 5424 47287 5424 47287 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit19.Q
rlabel metal2 11760 45003 11760 45003 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 4176 57036 4176 57036 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit20.Q
rlabel metal2 2592 57379 2592 57379 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 6192 57036 6192 57036 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 7776 57337 7776 57337 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 8160 46410 8160 46410 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit24.Q
rlabel metal3 9888 46872 9888 46872 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit25.Q
rlabel metal2 2784 50148 2784 50148 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 4320 49693 4320 49693 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 3264 60144 3264 60144 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 4800 60193 4800 60193 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 10176 45234 10176 45234 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 10512 60060 10512 60060 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 12144 60123 12144 60123 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit31.Q
rlabel metal3 16128 54264 16128 54264 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit4.Q
rlabel metal3 14544 54264 14544 54264 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 6048 55104 6048 55104 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 7584 55143 7584 55143 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 7872 44898 7872 44898 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 9552 44436 9552 44436 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 16704 75516 16704 75516 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 18240 75271 18240 75271 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit1.Q
rlabel via1 7632 74503 7632 74503 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 6048 74760 6048 74760 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 8256 62286 8256 62286 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 9792 62661 9792 62661 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 5760 64512 5760 64512 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 7296 64430 7296 64430 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 6240 70224 6240 70224 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 7728 69384 7728 69384 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit17.Q
rlabel metal3 12960 72996 12960 72996 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 13440 72492 13440 72492 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 1440 77238 1440 77238 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 13344 72450 13344 72450 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 16512 54852 16512 54852 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 15264 56280 15264 56280 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 17088 57330 17088 57330 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 14880 52584 14880 52584 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit24.Q
rlabel via2 14688 53340 14688 53340 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 16800 51744 16800 51744 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit26.Q
rlabel metal2 19776 82698 19776 82698 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 17760 82572 17760 82572 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 15264 84084 15264 84084 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 3168 73759 3168 73759 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit3.Q
rlabel metal2 12096 61527 12096 61527 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit30.Q
rlabel metal2 10560 60942 10560 60942 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 2880 65520 2880 65520 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit4.Q
rlabel via1 4464 65431 4464 65431 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit5.Q
rlabel metal2 2592 69174 2592 69174 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 3264 69633 3264 69633 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 10176 82992 10176 82992 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 4512 78505 4512 78505 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 2400 68712 2400 68712 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit0.Q
rlabel via1 4080 66943 4080 66943 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit1.Q
rlabel metal4 3456 73290 3456 73290 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit10.Q
rlabel metal2 4992 70053 4992 70053 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit11.Q
rlabel metal2 5280 73500 5280 73500 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit12.Q
rlabel metal2 3984 73668 3984 73668 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit13.Q
rlabel metal2 6480 78792 6480 78792 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit14.Q
rlabel metal2 7104 78750 7104 78750 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit15.Q
rlabel metal2 8448 79002 8448 79002 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit16.Q
rlabel metal2 9216 50484 9216 50484 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit17.Q
rlabel metal2 9504 50064 9504 50064 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit18.Q
rlabel metal3 10464 49476 10464 49476 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit19.Q
rlabel metal2 1536 72954 1536 72954 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit2.Q
rlabel metal2 9504 67711 9504 67711 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit20.Q
rlabel metal2 7968 67830 7968 67830 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit21.Q
rlabel metal2 9984 68544 9984 68544 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit22.Q
rlabel via1 11376 80551 11376 80551 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit23.Q
rlabel metal3 11616 81228 11616 81228 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 12672 82698 12672 82698 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit25.Q
rlabel metal2 14976 74757 14976 74757 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit26.Q
rlabel metal3 13680 73920 13680 73920 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 14352 60060 14352 60060 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit28.Q
rlabel metal3 16176 59556 16176 59556 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit29.Q
rlabel metal2 3072 73623 3072 73623 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit3.Q
rlabel metal3 8208 70644 8208 70644 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit30.Q
rlabel metal2 10080 70140 10080 70140 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit31.Q
rlabel metal2 2688 76902 2688 76902 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit4.Q
rlabel metal2 4224 77035 4224 77035 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit5.Q
rlabel metal2 2640 75180 2640 75180 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit6.Q
rlabel metal2 4272 75243 4272 75243 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit7.Q
rlabel metal2 2112 66402 2112 66402 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit8.Q
rlabel metal2 3648 64645 3648 64645 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame8_bit9.Q
rlabel metal2 9984 77371 9984 77371 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit22.Q
rlabel metal2 8448 76650 8448 76650 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit23.Q
rlabel metal2 14688 62202 14688 62202 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit24.Q
rlabel via1 15984 62407 15984 62407 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit25.Q
rlabel metal2 7968 71694 7968 71694 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit26.Q
rlabel metal2 9504 71733 9504 71733 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit27.Q
rlabel metal2 15840 79674 15840 79674 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit28.Q
rlabel metal2 17280 82236 17280 82236 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit29.Q
rlabel metal3 1344 80598 1344 80598 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit30.Q
rlabel metal2 2880 80889 2880 80889 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_ConfigMem.Inst_frame9_bit31.Q
rlabel metal2 12576 57204 12576 57204 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG0
rlabel via1 6899 66949 6899 66949 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG1
rlabel metal2 7584 52374 7584 52374 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG2
rlabel metal3 3984 60060 3984 60060 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG3
rlabel metal2 13536 70980 13536 70980 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG4
rlabel metal2 11760 53508 11760 53508 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG5
rlabel metal3 8304 52500 8304 52500 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG6
rlabel metal2 14928 68880 14928 68880 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS2_BEG7
rlabel metal2 16032 67956 16032 67956 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG0
rlabel metal3 16176 54432 16176 54432 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG1
rlabel metal3 14304 52500 14304 52500 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG10
rlabel metal2 11952 70896 11952 70896 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG11
rlabel metal3 14640 65436 14640 65436 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG12
rlabel metal3 16848 54432 16848 54432 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG13
rlabel metal2 14592 51324 14592 51324 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG14
rlabel metal2 19008 66906 19008 66906 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG15
rlabel metal2 14784 53592 14784 53592 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG2
rlabel metal2 12384 63210 12384 63210 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG3
rlabel metal3 12720 70644 12720 70644 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG4
rlabel metal2 16512 47040 16512 47040 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG5
rlabel metal2 15168 52416 15168 52416 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG6
rlabel metal3 17856 69132 17856 69132 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG7
rlabel metal2 12768 70749 12768 70749 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG8
rlabel metal2 19104 49140 19104 49140 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.J_NS4_BEG9
rlabel metal3 6240 75978 6240 75978 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG0
rlabel metal5 14448 64764 14448 64764 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG1
rlabel metal3 1584 71820 1584 71820 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG2
rlabel metal2 8208 84336 8208 84336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1BEG3
rlabel metal2 912 51324 912 51324 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END0
rlabel metal3 13104 33852 13104 33852 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END1
rlabel metal2 11424 70728 11424 70728 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END2
rlabel metal4 14496 52038 14496 52038 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N1END3
rlabel metal3 2124 76776 2124 76776 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG0
rlabel metal3 1440 83496 1440 83496 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG1
rlabel metal2 3264 71736 3264 71736 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG2
rlabel metal3 3504 82152 3504 82152 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG3
rlabel metal2 7440 79044 7440 79044 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG4
rlabel metal4 2496 71736 2496 71736 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG5
rlabel metal3 5280 70140 5280 70140 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG6
rlabel metal3 2016 84336 2016 84336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEG7
rlabel metal4 1440 75138 1440 75138 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb0
rlabel metal4 1056 74844 1056 74844 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb1
rlabel metal3 3648 35280 3648 35280 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb2
rlabel metal4 672 44688 672 44688 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb3
rlabel metal3 5664 82068 5664 82068 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb4
rlabel metal5 5472 29652 5472 29652 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb5
rlabel metal3 5424 31248 5424 31248 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb6
rlabel metal5 9080 82068 9080 82068 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N2BEGb7
rlabel metal2 5856 82362 5856 82362 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG0
rlabel metal5 8636 48048 8636 48048 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG1
rlabel metal2 8544 69678 8544 69678 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG2
rlabel metal3 9744 84336 9744 84336 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.N4BEG3
rlabel metal2 3984 1932 3984 1932 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG0
rlabel metal4 1056 37632 1056 37632 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG1
rlabel metal5 7920 12600 7920 12600 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG2
rlabel metal3 8352 37296 8352 37296 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG3
rlabel metal3 960 62832 960 62832 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG4
rlabel metal3 10080 33348 10080 33348 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG5
rlabel metal2 6144 31290 6144 31290 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG6
rlabel metal3 8736 70056 8736 70056 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S2BEG7
rlabel metal3 15120 70560 15120 70560 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG0
rlabel metal3 16080 31500 16080 31500 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG1
rlabel metal3 16656 51744 16656 51744 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG2
rlabel metal3 18144 1848 18144 1848 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.S4BEG3
rlabel metal3 11808 45360 11808 45360 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG0
rlabel metal2 13536 43512 13536 43512 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG1
rlabel metal2 11904 44646 11904 44646 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG2
rlabel metal3 15744 54936 15744 54936 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W1BEG3
rlabel metal2 1440 45696 1440 45696 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG0
rlabel metal2 9600 44940 9600 44940 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG1
rlabel metal2 1776 45696 1776 45696 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG2
rlabel metal2 2736 52836 2736 52836 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG3
rlabel metal4 2496 56784 2496 56784 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG4
rlabel metal2 7584 48048 7584 48048 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG5
rlabel metal3 4512 46536 4512 46536 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG6
rlabel metal2 2352 50232 2352 50232 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEG7
rlabel metal2 7968 57036 7968 57036 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb0
rlabel metal2 2112 47880 2112 47880 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb1
rlabel metal2 1728 49014 1728 49014 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb2
rlabel metal3 4992 59304 4992 59304 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb3
rlabel metal2 2112 61782 2112 61782 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb4
rlabel metal2 7968 47754 7968 47754 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb5
rlabel metal2 2112 45276 2112 45276 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb6
rlabel metal2 2160 50232 2160 50232 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W2BEGb7
rlabel metal2 12672 74718 12672 74718 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG0
rlabel metal2 13344 54138 13344 54138 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG1
rlabel metal2 5376 57162 5376 57162 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG10
rlabel metal2 2496 62874 2496 62874 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG11
rlabel metal2 13248 55524 13248 55524 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG2
rlabel metal2 15264 77784 15264 77784 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG3
rlabel metal2 12960 57792 12960 57792 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG4
rlabel metal2 2112 57330 2112 57330 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG5
rlabel metal3 1440 53886 1440 53886 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG6
rlabel metal2 1728 60690 1728 60690 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG7
rlabel metal2 13248 62622 13248 62622 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG8
rlabel metal2 9744 58044 9744 58044 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.W6BEG9
rlabel metal4 1728 56364 1728 56364 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG0
rlabel metal2 11424 51492 11424 51492 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG1
rlabel metal2 2016 53466 2016 53466 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG10
rlabel metal2 3456 55986 3456 55986 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG11
rlabel metal2 11472 56028 11472 56028 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG12
rlabel metal2 9648 53928 9648 53928 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG13
rlabel metal2 2496 45024 2496 45024 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG14
rlabel metal2 2592 62916 2592 62916 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG15
rlabel metal2 2208 48090 2208 48090 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG2
rlabel metal3 8208 53676 8208 53676 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG3
rlabel metal2 1344 54138 1344 54138 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG4
rlabel metal2 2400 51114 2400 51114 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG5
rlabel metal2 5760 52080 5760 52080 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG6
rlabel metal2 2112 54936 2112 54936 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG7
rlabel metal2 1728 55776 1728 55776 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG8
rlabel metal2 2112 54012 2112 54012 0 Tile_X0Y0_IHP_SRAM_top.Inst_IHP_SRAM_top_switch_matrix.WW4BEG9
rlabel metal3 6912 36876 6912 36876 0 Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_10.A
rlabel metal3 13776 67956 13776 67956 0 Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_11.A
rlabel metal3 16608 52080 16608 52080 0 Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_8.A
rlabel metal3 7824 66696 7824 66696 0 Tile_X0Y0_IHP_SRAM_top.N4BEG_outbuf_9.A
rlabel metal2 1824 83928 1824 83928 0 Tile_X0Y0_N1BEG[0]
rlabel metal2 2256 75432 2256 75432 0 Tile_X0Y0_N1BEG[1]
rlabel metal2 1536 76650 1536 76650 0 Tile_X0Y0_N1BEG[2]
rlabel metal2 2400 85482 2400 85482 0 Tile_X0Y0_N1BEG[3]
rlabel metal2 2592 84936 2592 84936 0 Tile_X0Y0_N2BEG[0]
rlabel metal2 1536 83790 1536 83790 0 Tile_X0Y0_N2BEG[1]
rlabel metal2 2976 84936 2976 84936 0 Tile_X0Y0_N2BEG[2]
rlabel metal2 3024 82236 3024 82236 0 Tile_X0Y0_N2BEG[3]
rlabel metal2 7104 82236 7104 82236 0 Tile_X0Y0_N2BEG[4]
rlabel metal2 3024 79212 3024 79212 0 Tile_X0Y0_N2BEG[5]
rlabel metal2 3744 85440 3744 85440 0 Tile_X0Y0_N2BEG[6]
rlabel metal2 1920 84672 1920 84672 0 Tile_X0Y0_N2BEG[7]
rlabel metal2 4128 84936 4128 84936 0 Tile_X0Y0_N2BEGb[0]
rlabel metal2 3648 82530 3648 82530 0 Tile_X0Y0_N2BEGb[1]
rlabel metal2 4512 83970 4512 83970 0 Tile_X0Y0_N2BEGb[2]
rlabel metal2 4704 84852 4704 84852 0 Tile_X0Y0_N2BEGb[3]
rlabel metal2 4416 83160 4416 83160 0 Tile_X0Y0_N2BEGb[4]
rlabel metal2 1536 84504 1536 84504 0 Tile_X0Y0_N2BEGb[5]
rlabel metal3 2976 82572 2976 82572 0 Tile_X0Y0_N2BEGb[6]
rlabel metal2 4032 82614 4032 82614 0 Tile_X0Y0_N2BEGb[7]
rlabel metal3 11952 5880 11952 5880 0 Tile_X0Y0_N4BEG[0]
rlabel metal2 5664 83748 5664 83748 0 Tile_X0Y0_N4BEG[10]
rlabel metal2 12576 83454 12576 83454 0 Tile_X0Y0_N4BEG[11]
rlabel metal2 6096 82992 6096 82992 0 Tile_X0Y0_N4BEG[12]
rlabel metal2 6432 83076 6432 83076 0 Tile_X0Y0_N4BEG[13]
rlabel metal3 8688 83748 8688 83748 0 Tile_X0Y0_N4BEG[14]
rlabel metal3 8208 84420 8208 84420 0 Tile_X0Y0_N4BEG[15]
rlabel metal2 1056 18816 1056 18816 0 Tile_X0Y0_N4BEG[1]
rlabel metal3 768 27048 768 27048 0 Tile_X0Y0_N4BEG[2]
rlabel metal5 7628 65856 7628 65856 0 Tile_X0Y0_N4BEG[3]
rlabel via5 2132 3612 2132 3612 0 Tile_X0Y0_N4BEG[4]
rlabel metal3 7248 16548 7248 16548 0 Tile_X0Y0_N4BEG[5]
rlabel metal2 6816 85776 6816 85776 0 Tile_X0Y0_N4BEG[6]
rlabel metal4 1824 34776 1824 34776 0 Tile_X0Y0_N4BEG[7]
rlabel metal2 7200 84894 7200 84894 0 Tile_X0Y0_N4BEG[8]
rlabel metal2 7344 84420 7344 84420 0 Tile_X0Y0_N4BEG[9]
rlabel metal3 10560 71568 10560 71568 0 Tile_X0Y0_S1END[0]
rlabel metal2 13584 53508 13584 53508 0 Tile_X0Y0_S1END[1]
rlabel metal2 11712 65520 11712 65520 0 Tile_X0Y0_S1END[2]
rlabel metal2 14976 54936 14976 54936 0 Tile_X0Y0_S1END[3]
rlabel metal2 11040 84558 11040 84558 0 Tile_X0Y0_S2END[0]
rlabel metal3 10272 71820 10272 71820 0 Tile_X0Y0_S2END[1]
rlabel metal2 11424 85230 11424 85230 0 Tile_X0Y0_S2END[2]
rlabel metal2 11616 84936 11616 84936 0 Tile_X0Y0_S2END[3]
rlabel metal2 11808 85482 11808 85482 0 Tile_X0Y0_S2END[4]
rlabel metal2 12000 85230 12000 85230 0 Tile_X0Y0_S2END[5]
rlabel metal2 12192 85734 12192 85734 0 Tile_X0Y0_S2END[6]
rlabel metal2 12384 85650 12384 85650 0 Tile_X0Y0_S2END[7]
rlabel metal3 2832 2352 2832 2352 0 Tile_X0Y0_S2MID[0]
rlabel metal3 960 46662 960 46662 0 Tile_X0Y0_S2MID[1]
rlabel metal2 4896 71358 4896 71358 0 Tile_X0Y0_S2MID[2]
rlabel metal2 10080 85104 10080 85104 0 Tile_X0Y0_S2MID[3]
rlabel metal2 7008 2142 7008 2142 0 Tile_X0Y0_S2MID[4]
rlabel metal2 6912 82614 6912 82614 0 Tile_X0Y0_S2MID[5]
rlabel metal2 5424 32340 5424 32340 0 Tile_X0Y0_S2MID[6]
rlabel metal5 10688 83496 10688 83496 0 Tile_X0Y0_S2MID[7]
rlabel metal2 12576 84810 12576 84810 0 Tile_X0Y0_S4END[0]
rlabel metal2 14496 85146 14496 85146 0 Tile_X0Y0_S4END[10]
rlabel metal2 14688 85566 14688 85566 0 Tile_X0Y0_S4END[11]
rlabel metal2 14880 85020 14880 85020 0 Tile_X0Y0_S4END[12]
rlabel metal2 15072 84726 15072 84726 0 Tile_X0Y0_S4END[13]
rlabel metal2 15264 85356 15264 85356 0 Tile_X0Y0_S4END[14]
rlabel metal2 15456 84936 15456 84936 0 Tile_X0Y0_S4END[15]
rlabel metal2 12096 53424 12096 53424 0 Tile_X0Y0_S4END[1]
rlabel metal2 12960 85230 12960 85230 0 Tile_X0Y0_S4END[2]
rlabel metal2 13824 78330 13824 78330 0 Tile_X0Y0_S4END[3]
rlabel metal2 13344 85356 13344 85356 0 Tile_X0Y0_S4END[4]
rlabel metal2 13824 15876 13824 15876 0 Tile_X0Y0_S4END[5]
rlabel metal2 9312 15036 9312 15036 0 Tile_X0Y0_S4END[6]
rlabel metal2 19440 12516 19440 12516 0 Tile_X0Y0_S4END[7]
rlabel metal2 14112 85104 14112 85104 0 Tile_X0Y0_S4END[8]
rlabel metal2 14304 84726 14304 84726 0 Tile_X0Y0_S4END[9]
rlabel metal2 15648 84936 15648 84936 0 Tile_X0Y0_UserCLKo
rlabel metal2 11712 43050 11712 43050 0 Tile_X0Y0_W1BEG[0]
rlabel metal3 78 43428 78 43428 0 Tile_X0Y0_W1BEG[1]
rlabel metal3 846 43764 846 43764 0 Tile_X0Y0_W1BEG[2]
rlabel metal3 7518 44100 7518 44100 0 Tile_X0Y0_W1BEG[3]
rlabel metal3 654 44436 654 44436 0 Tile_X0Y0_W2BEG[0]
rlabel metal3 846 44772 846 44772 0 Tile_X0Y0_W2BEG[1]
rlabel metal3 798 45108 798 45108 0 Tile_X0Y0_W2BEG[2]
rlabel metal3 1290 45444 1290 45444 0 Tile_X0Y0_W2BEG[3]
rlabel metal3 1290 45780 1290 45780 0 Tile_X0Y0_W2BEG[4]
rlabel metal3 798 46116 798 46116 0 Tile_X0Y0_W2BEG[5]
rlabel metal2 3264 46368 3264 46368 0 Tile_X0Y0_W2BEG[6]
rlabel metal3 1182 46788 1182 46788 0 Tile_X0Y0_W2BEG[7]
rlabel metal3 366 47124 366 47124 0 Tile_X0Y0_W2BEGb[0]
rlabel metal3 990 47460 990 47460 0 Tile_X0Y0_W2BEGb[1]
rlabel metal3 750 47796 750 47796 0 Tile_X0Y0_W2BEGb[2]
rlabel metal3 1614 48132 1614 48132 0 Tile_X0Y0_W2BEGb[3]
rlabel metal3 1038 48468 1038 48468 0 Tile_X0Y0_W2BEGb[4]
rlabel metal2 1584 48216 1584 48216 0 Tile_X0Y0_W2BEGb[5]
rlabel metal2 1776 45528 1776 45528 0 Tile_X0Y0_W2BEGb[6]
rlabel metal3 990 49476 990 49476 0 Tile_X0Y0_W2BEGb[7]
rlabel metal3 510 55188 510 55188 0 Tile_X0Y0_W6BEG[0]
rlabel metal2 1344 58128 1344 58128 0 Tile_X0Y0_W6BEG[10]
rlabel metal3 510 58884 510 58884 0 Tile_X0Y0_W6BEG[11]
rlabel metal2 13488 55020 13488 55020 0 Tile_X0Y0_W6BEG[1]
rlabel metal2 13440 55314 13440 55314 0 Tile_X0Y0_W6BEG[2]
rlabel metal5 14540 77280 14540 77280 0 Tile_X0Y0_W6BEG[3]
rlabel metal2 10080 57456 10080 57456 0 Tile_X0Y0_W6BEG[4]
rlabel metal3 990 56868 990 56868 0 Tile_X0Y0_W6BEG[5]
rlabel metal2 1248 56868 1248 56868 0 Tile_X0Y0_W6BEG[6]
rlabel metal3 750 57540 750 57540 0 Tile_X0Y0_W6BEG[7]
rlabel metal3 702 57876 702 57876 0 Tile_X0Y0_W6BEG[8]
rlabel metal3 1290 58212 1290 58212 0 Tile_X0Y0_W6BEG[9]
rlabel metal3 798 49812 798 49812 0 Tile_X0Y0_WW4BEG[0]
rlabel metal3 78 53172 78 53172 0 Tile_X0Y0_WW4BEG[10]
rlabel metal3 1662 53508 1662 53508 0 Tile_X0Y0_WW4BEG[11]
rlabel metal3 126 53844 126 53844 0 Tile_X0Y0_WW4BEG[12]
rlabel metal3 1290 54180 1290 54180 0 Tile_X0Y0_WW4BEG[13]
rlabel metal2 2304 46242 2304 46242 0 Tile_X0Y0_WW4BEG[14]
rlabel metal3 750 54852 750 54852 0 Tile_X0Y0_WW4BEG[15]
rlabel metal2 2880 50484 2880 50484 0 Tile_X0Y0_WW4BEG[1]
rlabel metal2 1872 48972 1872 48972 0 Tile_X0Y0_WW4BEG[2]
rlabel metal2 8448 51198 8448 51198 0 Tile_X0Y0_WW4BEG[3]
rlabel metal3 702 51156 702 51156 0 Tile_X0Y0_WW4BEG[4]
rlabel metal2 2160 50064 2160 50064 0 Tile_X0Y0_WW4BEG[5]
rlabel metal3 894 51828 894 51828 0 Tile_X0Y0_WW4BEG[6]
rlabel metal3 1230 52164 1230 52164 0 Tile_X0Y0_WW4BEG[7]
rlabel metal3 846 52500 846 52500 0 Tile_X0Y0_WW4BEG[8]
rlabel metal3 942 52836 942 52836 0 Tile_X0Y0_WW4BEG[9]
rlabel metal2 18672 20076 18672 20076 0 Tile_X0Y1_E1END[0]
rlabel metal2 17952 34188 17952 34188 0 Tile_X0Y1_E1END[1]
rlabel metal2 12384 36288 12384 36288 0 Tile_X0Y1_E1END[2]
rlabel metal3 13632 34482 13632 34482 0 Tile_X0Y1_E1END[3]
rlabel metal2 11040 20496 11040 20496 0 Tile_X0Y1_E2END[0]
rlabel metal2 5568 23520 5568 23520 0 Tile_X0Y1_E2END[1]
rlabel metal2 6336 20874 6336 20874 0 Tile_X0Y1_E2END[2]
rlabel metal3 8160 33180 8160 33180 0 Tile_X0Y1_E2END[3]
rlabel metal2 3168 40908 3168 40908 0 Tile_X0Y1_E2END[4]
rlabel metal3 990 21924 990 21924 0 Tile_X0Y1_E2END[5]
rlabel metal4 2880 24528 2880 24528 0 Tile_X0Y1_E2END[6]
rlabel metal2 2784 23898 2784 23898 0 Tile_X0Y1_E2END[7]
rlabel metal3 5598 17556 5598 17556 0 Tile_X0Y1_E2MID[0]
rlabel metal3 846 17892 846 17892 0 Tile_X0Y1_E2MID[1]
rlabel metal2 2448 29652 2448 29652 0 Tile_X0Y1_E2MID[2]
rlabel metal2 2208 39774 2208 39774 0 Tile_X0Y1_E2MID[3]
rlabel metal3 3120 27636 3120 27636 0 Tile_X0Y1_E2MID[4]
rlabel via2 78 19236 78 19236 0 Tile_X0Y1_E2MID[5]
rlabel metal3 942 19572 942 19572 0 Tile_X0Y1_E2MID[6]
rlabel metal3 2064 22512 2064 22512 0 Tile_X0Y1_E2MID[7]
rlabel metal2 17856 26670 17856 26670 0 Tile_X0Y1_E6END[0]
rlabel metal2 2496 31878 2496 31878 0 Tile_X0Y1_E6END[10]
rlabel metal2 18912 36960 18912 36960 0 Tile_X0Y1_E6END[11]
rlabel metal3 4272 30996 4272 30996 0 Tile_X0Y1_E6END[1]
rlabel metal3 78 28980 78 28980 0 Tile_X0Y1_E6END[2]
rlabel metal3 606 29316 606 29316 0 Tile_X0Y1_E6END[3]
rlabel metal3 654 29652 654 29652 0 Tile_X0Y1_E6END[4]
rlabel metal2 1440 31962 1440 31962 0 Tile_X0Y1_E6END[5]
rlabel metal2 13056 31542 13056 31542 0 Tile_X0Y1_E6END[6]
rlabel metal3 654 30660 654 30660 0 Tile_X0Y1_E6END[7]
rlabel metal3 222 30996 222 30996 0 Tile_X0Y1_E6END[8]
rlabel metal2 2976 33264 2976 33264 0 Tile_X0Y1_E6END[9]
rlabel metal2 18048 29484 18048 29484 0 Tile_X0Y1_EE4END[0]
rlabel metal3 894 26292 894 26292 0 Tile_X0Y1_EE4END[10]
rlabel metal3 1038 26628 1038 26628 0 Tile_X0Y1_EE4END[11]
rlabel metal3 846 26964 846 26964 0 Tile_X0Y1_EE4END[12]
rlabel metal3 606 27300 606 27300 0 Tile_X0Y1_EE4END[13]
rlabel metal3 1278 27636 1278 27636 0 Tile_X0Y1_EE4END[14]
rlabel metal3 1182 27972 1182 27972 0 Tile_X0Y1_EE4END[15]
rlabel metal3 174 23268 174 23268 0 Tile_X0Y1_EE4END[1]
rlabel metal3 78 23604 78 23604 0 Tile_X0Y1_EE4END[2]
rlabel metal4 384 23856 384 23856 0 Tile_X0Y1_EE4END[3]
rlabel metal2 18624 24444 18624 24444 0 Tile_X0Y1_EE4END[4]
rlabel metal3 1086 24612 1086 24612 0 Tile_X0Y1_EE4END[5]
rlabel metal2 12576 32130 12576 32130 0 Tile_X0Y1_EE4END[6]
rlabel metal3 318 25284 318 25284 0 Tile_X0Y1_EE4END[7]
rlabel metal3 18096 29064 18096 29064 0 Tile_X0Y1_EE4END[8]
rlabel metal2 15408 26208 15408 26208 0 Tile_X0Y1_EE4END[9]
rlabel metal2 15936 4914 15936 4914 0 Tile_X0Y1_FrameData[0]
rlabel metal2 15168 1596 15168 1596 0 Tile_X0Y1_FrameData[10]
rlabel metal2 11904 1134 11904 1134 0 Tile_X0Y1_FrameData[11]
rlabel metal2 1296 14028 1296 14028 0 Tile_X0Y1_FrameData[12]
rlabel metal2 1248 15624 1248 15624 0 Tile_X0Y1_FrameData[13]
rlabel metal2 13632 30618 13632 30618 0 Tile_X0Y1_FrameData[14]
rlabel metal2 1296 37380 1296 37380 0 Tile_X0Y1_FrameData[15]
rlabel metal2 16512 2058 16512 2058 0 Tile_X0Y1_FrameData[16]
rlabel metal2 5280 1176 5280 1176 0 Tile_X0Y1_FrameData[17]
rlabel metal2 1344 19740 1344 19740 0 Tile_X0Y1_FrameData[18]
rlabel metal2 1344 21084 1344 21084 0 Tile_X0Y1_FrameData[19]
rlabel metal4 16320 16002 16320 16002 0 Tile_X0Y1_FrameData[1]
rlabel metal2 1344 30198 1344 30198 0 Tile_X0Y1_FrameData[20]
rlabel metal3 846 39396 846 39396 0 Tile_X0Y1_FrameData[21]
rlabel metal2 1248 19194 1248 19194 0 Tile_X0Y1_FrameData[22]
rlabel metal3 894 40068 894 40068 0 Tile_X0Y1_FrameData[23]
rlabel metal3 2208 40362 2208 40362 0 Tile_X0Y1_FrameData[24]
rlabel metal2 1296 22260 1296 22260 0 Tile_X0Y1_FrameData[25]
rlabel metal2 7248 1092 7248 1092 0 Tile_X0Y1_FrameData[26]
rlabel metal4 2016 39774 2016 39774 0 Tile_X0Y1_FrameData[27]
rlabel metal3 1680 7980 1680 7980 0 Tile_X0Y1_FrameData[28]
rlabel metal2 1248 22974 1248 22974 0 Tile_X0Y1_FrameData[29]
rlabel metal3 126 33012 126 33012 0 Tile_X0Y1_FrameData[2]
rlabel metal2 13104 30240 13104 30240 0 Tile_X0Y1_FrameData[30]
rlabel metal3 1296 25284 1296 25284 0 Tile_X0Y1_FrameData[31]
rlabel metal3 13344 17094 13344 17094 0 Tile_X0Y1_FrameData[3]
rlabel metal2 1248 38262 1248 38262 0 Tile_X0Y1_FrameData[4]
rlabel metal3 1392 38472 1392 38472 0 Tile_X0Y1_FrameData[5]
rlabel metal3 1440 41244 1440 41244 0 Tile_X0Y1_FrameData[6]
rlabel metal2 2208 43386 2208 43386 0 Tile_X0Y1_FrameData[7]
rlabel metal2 16560 14028 16560 14028 0 Tile_X0Y1_FrameData[8]
rlabel metal2 18576 1932 18576 1932 0 Tile_X0Y1_FrameData[9]
rlabel metal3 13680 49224 13680 49224 0 Tile_X0Y1_FrameData_O[0]
rlabel metal3 18498 65436 18498 65436 0 Tile_X0Y1_FrameData_O[10]
rlabel metal3 21138 65772 21138 65772 0 Tile_X0Y1_FrameData_O[11]
rlabel metal3 20994 66108 20994 66108 0 Tile_X0Y1_FrameData_O[12]
rlabel metal3 17826 66444 17826 66444 0 Tile_X0Y1_FrameData_O[13]
rlabel metal3 21234 66780 21234 66780 0 Tile_X0Y1_FrameData_O[14]
rlabel metal3 21090 67116 21090 67116 0 Tile_X0Y1_FrameData_O[15]
rlabel metal3 20802 67452 20802 67452 0 Tile_X0Y1_FrameData_O[16]
rlabel metal3 21186 67788 21186 67788 0 Tile_X0Y1_FrameData_O[17]
rlabel metal3 21042 68124 21042 68124 0 Tile_X0Y1_FrameData_O[18]
rlabel metal3 21186 68460 21186 68460 0 Tile_X0Y1_FrameData_O[19]
rlabel metal3 20850 62412 20850 62412 0 Tile_X0Y1_FrameData_O[1]
rlabel metal3 20994 68796 20994 68796 0 Tile_X0Y1_FrameData_O[20]
rlabel metal3 20994 69132 20994 69132 0 Tile_X0Y1_FrameData_O[21]
rlabel metal3 21042 69468 21042 69468 0 Tile_X0Y1_FrameData_O[22]
rlabel metal3 16944 54180 16944 54180 0 Tile_X0Y1_FrameData_O[23]
rlabel metal3 19650 70140 19650 70140 0 Tile_X0Y1_FrameData_O[24]
rlabel metal3 20448 41412 20448 41412 0 Tile_X0Y1_FrameData_O[25]
rlabel metal3 18306 70812 18306 70812 0 Tile_X0Y1_FrameData_O[26]
rlabel metal3 19122 71148 19122 71148 0 Tile_X0Y1_FrameData_O[27]
rlabel metal3 21138 71484 21138 71484 0 Tile_X0Y1_FrameData_O[28]
rlabel via3 21426 71820 21426 71820 0 Tile_X0Y1_FrameData_O[29]
rlabel metal3 20994 62748 20994 62748 0 Tile_X0Y1_FrameData_O[2]
rlabel metal3 19938 72156 19938 72156 0 Tile_X0Y1_FrameData_O[30]
rlabel metal3 21282 72492 21282 72492 0 Tile_X0Y1_FrameData_O[31]
rlabel metal3 21234 63084 21234 63084 0 Tile_X0Y1_FrameData_O[3]
rlabel metal2 18336 43302 18336 43302 0 Tile_X0Y1_FrameData_O[4]
rlabel metal3 21330 63756 21330 63756 0 Tile_X0Y1_FrameData_O[5]
rlabel metal4 17952 53340 17952 53340 0 Tile_X0Y1_FrameData_O[6]
rlabel metal3 21042 64428 21042 64428 0 Tile_X0Y1_FrameData_O[7]
rlabel metal3 21234 64764 21234 64764 0 Tile_X0Y1_FrameData_O[8]
rlabel metal3 21330 65100 21330 65100 0 Tile_X0Y1_FrameData_O[9]
rlabel metal2 20640 82404 20640 82404 0 Tile_X0Y1_FrameStrobe[0]
rlabel metal2 17760 660 17760 660 0 Tile_X0Y1_FrameStrobe[10]
rlabel metal2 17952 786 17952 786 0 Tile_X0Y1_FrameStrobe[11]
rlabel metal2 18144 660 18144 660 0 Tile_X0Y1_FrameStrobe[12]
rlabel metal2 18336 618 18336 618 0 Tile_X0Y1_FrameStrobe[13]
rlabel metal2 18528 450 18528 450 0 Tile_X0Y1_FrameStrobe[14]
rlabel metal2 18720 660 18720 660 0 Tile_X0Y1_FrameStrobe[15]
rlabel metal2 18912 366 18912 366 0 Tile_X0Y1_FrameStrobe[16]
rlabel metal2 19104 534 19104 534 0 Tile_X0Y1_FrameStrobe[17]
rlabel metal2 19296 156 19296 156 0 Tile_X0Y1_FrameStrobe[18]
rlabel metal2 19488 114 19488 114 0 Tile_X0Y1_FrameStrobe[19]
rlabel metal2 2496 38892 2496 38892 0 Tile_X0Y1_FrameStrobe[1]
rlabel metal2 18240 19404 18240 19404 0 Tile_X0Y1_FrameStrobe[2]
rlabel metal3 17952 18312 17952 18312 0 Tile_X0Y1_FrameStrobe[3]
rlabel metal2 2496 16632 2496 16632 0 Tile_X0Y1_FrameStrobe[4]
rlabel metal2 2496 11760 2496 11760 0 Tile_X0Y1_FrameStrobe[5]
rlabel metal3 2016 15372 2016 15372 0 Tile_X0Y1_FrameStrobe[6]
rlabel metal2 17184 240 17184 240 0 Tile_X0Y1_FrameStrobe[7]
rlabel metal2 2304 20370 2304 20370 0 Tile_X0Y1_FrameStrobe[8]
rlabel metal2 17568 492 17568 492 0 Tile_X0Y1_FrameStrobe[9]
rlabel metal2 17376 5250 17376 5250 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit0.Q
rlabel metal2 18336 5719 18336 5719 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit1.Q
rlabel metal2 13680 1260 13680 1260 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit10.Q
rlabel metal3 8016 924 8016 924 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit11.Q
rlabel metal2 2688 37128 2688 37128 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit12.Q
rlabel metal2 2688 36330 2688 36330 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit13.Q
rlabel metal2 4608 39067 4608 39067 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit14.Q
rlabel metal2 2736 37632 2736 37632 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit15.Q
rlabel metal2 7008 2646 7008 2646 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit16.Q
rlabel metal2 6768 1260 6768 1260 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit17.Q
rlabel metal3 6240 3192 6240 3192 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit18.Q
rlabel metal2 5088 3234 5088 3234 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit19.Q
rlabel metal2 12768 16506 12768 16506 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit2.Q
rlabel metal2 5760 30366 5760 30366 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit20.Q
rlabel metal2 7104 31423 7104 31423 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit21.Q
rlabel metal3 9360 5124 9360 5124 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit22.Q
rlabel metal2 10656 4578 10656 4578 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit23.Q
rlabel metal2 15168 21210 15168 21210 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit24.Q
rlabel metal3 15168 21756 15168 21756 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit25.Q
rlabel metal2 12576 27510 12576 27510 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit26.Q
rlabel metal2 12288 26544 12288 26544 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit27.Q
rlabel metal2 8736 33222 8736 33222 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit28.Q
rlabel metal2 9600 32256 9600 32256 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit29.Q
rlabel metal2 14304 16513 14304 16513 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit3.Q
rlabel metal2 15072 26628 15072 26628 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit30.Q
rlabel metal2 14736 27048 14736 27048 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit31.Q
rlabel metal2 8832 17682 8832 17682 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit4.Q
rlabel metal2 10656 17472 10656 17472 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit5.Q
rlabel metal2 15792 9660 15792 9660 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit6.Q
rlabel metal3 17568 10416 17568 10416 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit7.Q
rlabel metal3 4512 2016 4512 2016 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit8.Q
rlabel metal2 4896 1757 4896 1757 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame0_bit9.Q
rlabel metal2 7296 40026 7296 40026 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit0.Q
rlabel metal2 8832 39312 8832 39312 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit1.Q
rlabel metal2 12768 15582 12768 15582 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit10.Q
rlabel metal2 14544 14952 14544 14952 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit11.Q
rlabel metal2 8496 20244 8496 20244 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit12.Q
rlabel metal2 10176 20496 10176 20496 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit13.Q
rlabel metal2 18432 14280 18432 14280 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit14.Q
rlabel metal2 20256 13727 20256 13727 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit15.Q
rlabel metal2 17952 2772 17952 2772 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit16.Q
rlabel metal2 19824 1260 19824 1260 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit17.Q
rlabel metal2 12576 19194 12576 19194 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit18.Q
rlabel via1 14160 19240 14160 19240 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit19.Q
rlabel metal2 9504 42798 9504 42798 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit2.Q
rlabel metal2 8736 19194 8736 19194 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit20.Q
rlabel metal2 10560 18984 10560 18984 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit21.Q
rlabel metal3 18096 9660 18096 9660 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit22.Q
rlabel metal2 20112 8904 20112 8904 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit23.Q
rlabel metal2 18000 7308 18000 7308 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit24.Q
rlabel metal3 19728 6636 19728 6636 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit25.Q
rlabel metal2 12768 18606 12768 18606 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit26.Q
rlabel metal3 14592 17976 14592 17976 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit27.Q
rlabel metal2 8352 15708 8352 15708 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit28.Q
rlabel metal2 9888 15582 9888 15582 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit29.Q
rlabel metal2 19680 41111 19680 41111 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit3.Q
rlabel metal2 18720 11970 18720 11970 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit30.Q
rlabel metal2 19944 12432 19944 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit31.Q
rlabel metal2 2304 40908 2304 40908 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit4.Q
rlabel metal2 2880 40908 2880 40908 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit5.Q
rlabel metal2 4128 40453 4128 40453 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit6.Q
rlabel metal3 3792 42756 3792 42756 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit7.Q
rlabel metal3 18192 2856 18192 2856 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit8.Q
rlabel metal2 19656 4116 19656 4116 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame1_bit9.Q
rlabel metal2 9312 34178 9312 34178 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit0.Q
rlabel metal2 10704 33852 10704 33852 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit1.Q
rlabel metal2 15744 40488 15744 40488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit10.Q
rlabel metal2 17232 39900 17232 39900 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit11.Q
rlabel metal3 16896 29148 16896 29148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit12.Q
rlabel metal2 19608 29148 19608 29148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit13.Q
rlabel metal3 14352 33684 14352 33684 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit14.Q
rlabel metal2 16224 33765 16224 33765 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit15.Q
rlabel metal2 9504 36078 9504 36078 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit16.Q
rlabel metal2 11136 35616 11136 35616 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit17.Q
rlabel metal2 17760 39480 17760 39480 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit18.Q
rlabel metal2 19680 39981 19680 39981 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit19.Q
rlabel metal2 18864 38388 18864 38388 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit2.Q
rlabel metal2 18480 19488 18480 19488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit20.Q
rlabel metal2 20400 18732 20400 18732 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit21.Q
rlabel metal2 18048 34188 18048 34188 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit22.Q
rlabel metal2 19392 33728 19392 33728 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit23.Q
rlabel metal2 12288 37128 12288 37128 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit24.Q
rlabel metal3 13968 38052 13968 38052 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit25.Q
rlabel metal2 15696 41412 15696 41412 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit26.Q
rlabel metal2 17376 41664 17376 41664 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit27.Q
rlabel metal2 6480 41412 6480 41412 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit28.Q
rlabel metal3 7440 41916 7440 41916 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit29.Q
rlabel metal2 19920 37632 19920 37632 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit3.Q
rlabel metal2 8928 41706 8928 41706 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit30.Q
rlabel metal2 7776 43722 7776 43722 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit31.Q
rlabel metal2 18528 22344 18528 22344 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit4.Q
rlabel metal2 20016 20580 20016 20580 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit5.Q
rlabel metal2 18528 34314 18528 34314 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit6.Q
rlabel metal2 20400 30828 20400 30828 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit7.Q
rlabel metal3 12384 36708 12384 36708 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit8.Q
rlabel metal3 14688 35700 14688 35700 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame2_bit9.Q
rlabel metal2 9312 29232 9312 29232 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit0.Q
rlabel metal2 10848 28847 10848 28847 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit1.Q
rlabel metal2 15744 37716 15744 37716 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit10.Q
rlabel metal2 17256 38136 17256 38136 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit11.Q
rlabel metal2 17520 29316 17520 29316 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit12.Q
rlabel metal3 18768 29400 18768 29400 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit13.Q
rlabel metal2 15072 30870 15072 30870 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit14.Q
rlabel metal2 16704 30912 16704 30912 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit15.Q
rlabel metal2 9648 30828 9648 30828 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit16.Q
rlabel metal2 11280 30828 11280 30828 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit17.Q
rlabel metal2 18336 36414 18336 36414 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit18.Q
rlabel metal2 19920 36120 19920 36120 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit19.Q
rlabel metal2 18240 28056 18240 28056 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit2.Q
rlabel metal2 18432 21630 18432 21630 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit20.Q
rlabel metal2 20016 19488 20016 19488 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit21.Q
rlabel metal2 18144 31626 18144 31626 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit22.Q
rlabel metal2 17472 30408 17472 30408 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit23.Q
rlabel metal2 12288 35448 12288 35448 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit24.Q
rlabel metal2 13824 34895 13824 34895 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit25.Q
rlabel metal3 16080 35700 16080 35700 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit26.Q
rlabel metal2 17136 34944 17136 34944 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit27.Q
rlabel metal2 18192 25536 18192 25536 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit28.Q
rlabel metal2 20064 23268 20064 23268 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit29.Q
rlabel metal2 20400 23940 20400 23940 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit3.Q
rlabel metal2 14784 32928 14784 32928 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit30.Q
rlabel metal2 16464 32340 16464 32340 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit31.Q
rlabel metal2 18528 24654 18528 24654 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit4.Q
rlabel metal3 19344 23940 19344 23940 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit5.Q
rlabel metal2 18384 30828 18384 30828 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit6.Q
rlabel metal2 20208 27720 20208 27720 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit7.Q
rlabel metal2 12480 32214 12480 32214 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit8.Q
rlabel metal2 14112 31668 14112 31668 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame3_bit9.Q
rlabel metal2 16032 12936 16032 12936 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit0.Q
rlabel metal2 17712 12600 17712 12600 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit1.Q
rlabel metal2 14592 13727 14592 13727 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit10.Q
rlabel metal2 13008 12600 13008 12600 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit11.Q
rlabel metal2 2640 17976 2640 17976 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit12.Q
rlabel metal2 2784 15708 2784 15708 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit13.Q
rlabel metal2 8256 12894 8256 12894 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit14.Q
rlabel metal2 6192 12600 6192 12600 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit15.Q
rlabel metal2 17088 16513 17088 16513 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit16.Q
rlabel metal2 16128 15582 16128 15582 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit17.Q
rlabel metal2 11520 23604 11520 23604 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit18.Q
rlabel metal2 11856 24360 11856 24360 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit19.Q
rlabel metal2 12000 11424 12000 11424 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit2.Q
rlabel metal2 1968 24612 1968 24612 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit20.Q
rlabel metal2 5856 23730 5856 23730 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit21.Q
rlabel metal3 6240 26124 6240 26124 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit22.Q
rlabel metal2 6624 25990 6624 25990 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit23.Q
rlabel metal2 10752 38640 10752 38640 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit24.Q
rlabel metal2 11424 38682 11424 38682 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit25.Q
rlabel metal2 8544 25830 8544 25830 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit26.Q
rlabel metal2 9792 26166 9792 26166 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit27.Q
rlabel metal2 17280 26880 17280 26880 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit28.Q
rlabel metal3 18336 26292 18336 26292 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit29.Q
rlabel metal2 10224 10416 10224 10416 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit3.Q
rlabel metal2 14880 28266 14880 28266 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit30.Q
rlabel metal2 16560 27804 16560 27804 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit31.Q
rlabel metal2 7200 18813 7200 18813 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit4.Q
rlabel metal2 5760 17976 5760 17976 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit5.Q
rlabel metal2 5568 12138 5568 12138 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit6.Q
rlabel metal2 7080 13188 7080 13188 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit7.Q
rlabel metal2 15168 14448 15168 14448 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit8.Q
rlabel metal2 16704 15001 16704 15001 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame4_bit9.Q
rlabel metal2 14016 5376 14016 5376 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit0.Q
rlabel metal2 15696 5124 15696 5124 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit1.Q
rlabel metal2 9696 8820 9696 8820 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit10.Q
rlabel metal2 11520 9531 11520 9531 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit11.Q
rlabel metal2 2688 12768 2688 12768 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit12.Q
rlabel metal2 4512 19537 4512 19537 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit13.Q
rlabel metal3 4896 8820 4896 8820 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit14.Q
rlabel metal3 7152 8148 7152 8148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit15.Q
rlabel metal2 15168 3276 15168 3276 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit16.Q
rlabel metal2 16704 3283 16704 3283 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit17.Q
rlabel metal3 12672 10416 12672 10416 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit18.Q
rlabel metal2 14112 11253 14112 11253 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit19.Q
rlabel metal2 11616 7308 11616 7308 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit2.Q
rlabel metal2 2688 7308 2688 7308 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit20.Q
rlabel metal2 4992 10458 4992 10458 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit21.Q
rlabel metal2 5760 8148 5760 8148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit22.Q
rlabel metal3 7248 9660 7248 9660 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit23.Q
rlabel metal2 14544 10416 14544 10416 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit24.Q
rlabel metal2 16176 10416 16176 10416 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit25.Q
rlabel metal2 12384 8610 12384 8610 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit26.Q
rlabel metal2 13920 8402 13920 8402 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit27.Q
rlabel metal2 10272 15960 10272 15960 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit28.Q
rlabel metal2 11952 14952 11952 14952 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit29.Q
rlabel metal4 10080 7686 10080 7686 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit3.Q
rlabel metal2 8544 11508 8544 11508 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit30.Q
rlabel metal2 10032 11172 10032 11172 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit31.Q
rlabel metal2 5280 15708 5280 15708 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit4.Q
rlabel metal2 6816 16373 6816 16373 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit5.Q
rlabel metal3 4992 4368 4992 4368 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit6.Q
rlabel metal2 6528 6720 6528 6720 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit7.Q
rlabel metal2 15552 8190 15552 8190 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit8.Q
rlabel metal3 15408 8148 15408 8148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame5_bit9.Q
rlabel metal2 11616 2856 11616 2856 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit0.Q
rlabel metal2 13344 3693 13344 3693 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit1.Q
rlabel metal3 7584 2100 7584 2100 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit10.Q
rlabel metal2 10272 1722 10272 1722 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit11.Q
rlabel metal3 3408 14196 3408 14196 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit12.Q
rlabel metal2 3456 15876 3456 15876 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit13.Q
rlabel metal3 2784 11004 2784 11004 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit14.Q
rlabel metal2 4128 9905 4128 9905 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit15.Q
rlabel metal3 11568 2100 11568 2100 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit16.Q
rlabel metal3 13152 2604 13152 2604 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit17.Q
rlabel metal2 6720 4242 6720 4242 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit18.Q
rlabel metal2 8640 2310 8640 2310 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit19.Q
rlabel metal3 7728 4368 7728 4368 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit2.Q
rlabel metal2 2352 12516 2352 12516 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit20.Q
rlabel metal3 2976 7434 2976 7434 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit21.Q
rlabel metal2 12384 5628 12384 5628 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit22.Q
rlabel metal2 4992 1680 4992 1680 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit23.Q
rlabel metal2 14592 7098 14592 7098 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit24.Q
rlabel metal2 16272 6636 16272 6636 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit25.Q
rlabel metal3 12288 5082 12288 5082 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit26.Q
rlabel metal2 13680 5880 13680 5880 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit27.Q
rlabel metal2 5664 15582 5664 15582 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit28.Q
rlabel metal2 7488 15120 7488 15120 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit29.Q
rlabel metal2 7008 6932 7008 6932 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit3.Q
rlabel metal2 7440 6636 7440 6636 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit30.Q
rlabel metal2 9120 7056 9120 7056 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit31.Q
rlabel metal3 2976 12096 2976 12096 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit4.Q
rlabel metal2 2064 12600 2064 12600 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit5.Q
rlabel metal2 2880 1260 2880 1260 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit6.Q
rlabel metal2 3744 3990 3744 3990 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit7.Q
rlabel metal2 14544 2100 14544 2100 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit8.Q
rlabel metal2 16176 2100 16176 2100 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame6_bit9.Q
rlabel metal2 5760 20706 5760 20706 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit0.Q
rlabel metal2 6816 20370 6816 20370 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit1.Q
rlabel metal2 14496 29536 14496 29536 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit10.Q
rlabel metal2 13056 29778 13056 29778 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit11.Q
rlabel metal2 5760 25452 5760 25452 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit12.Q
rlabel metal2 6288 29148 6288 29148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit13.Q
rlabel metal2 6288 26796 6288 26796 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit14.Q
rlabel metal2 16128 19194 16128 19194 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit15.Q
rlabel metal2 16560 18732 16560 18732 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit16.Q
rlabel metal2 17472 18564 17472 18564 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit17.Q
rlabel metal2 20256 3192 20256 3192 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit18.Q
rlabel metal2 20064 5040 20064 5040 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit19.Q
rlabel metal2 4800 22437 4800 22437 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit2.Q
rlabel metal2 12672 13440 12672 13440 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit20.Q
rlabel metal2 10944 13734 10944 13734 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit21.Q
rlabel metal2 10224 12684 10224 12684 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit22.Q
rlabel metal2 8880 13440 8880 13440 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit23.Q
rlabel metal2 20064 7770 20064 7770 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit24.Q
rlabel metal2 18288 8904 18288 8904 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit25.Q
rlabel metal2 8640 1218 8640 1218 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit26.Q
rlabel via1 8784 4120 8784 4120 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit27.Q
rlabel metal2 2736 8148 2736 8148 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit28.Q
rlabel metal2 4272 12600 4272 12600 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit29.Q
rlabel metal2 6288 21672 6288 21672 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit3.Q
rlabel metal3 3120 9072 3120 9072 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit30.Q
rlabel metal2 4320 6006 4320 6006 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit31.Q
rlabel metal2 12240 20244 12240 20244 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit4.Q
rlabel metal2 10560 21042 10560 21042 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit5.Q
rlabel metal3 18288 17220 18288 17220 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit6.Q
rlabel metal2 20160 16821 20160 16821 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit7.Q
rlabel metal2 20064 15582 20064 15582 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit8.Q
rlabel metal2 13440 29106 13440 29106 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame7_bit9.Q
rlabel metal2 8352 23730 8352 23730 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit0.Q
rlabel metal2 9888 23522 9888 23522 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit1.Q
rlabel metal2 6144 37044 6144 37044 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit10.Q
rlabel metal3 13776 39732 13776 39732 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit11.Q
rlabel metal2 12960 39984 12960 39984 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit12.Q
rlabel metal2 13680 41244 13680 41244 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit13.Q
rlabel metal2 12288 22218 12288 22218 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit14.Q
rlabel metal2 13776 21756 13776 21756 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit15.Q
rlabel metal2 9216 27678 9216 27678 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit16.Q
rlabel metal2 10464 27090 10464 27090 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit17.Q
rlabel metal2 7536 30828 7536 30828 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit18.Q
rlabel metal2 9072 30072 9072 30072 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit19.Q
rlabel metal3 16992 23772 16992 23772 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit2.Q
rlabel metal2 12576 25242 12576 25242 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit20.Q
rlabel metal2 14208 25032 14208 25032 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit21.Q
rlabel metal2 2016 20958 2016 20958 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit22.Q
rlabel metal2 4320 22722 4320 22722 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit23.Q
rlabel metal2 2400 26166 2400 26166 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit24.Q
rlabel metal2 3984 26859 3984 26859 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit25.Q
rlabel metal3 3360 29316 3360 29316 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit26.Q
rlabel metal3 2352 26292 2352 26292 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit27.Q
rlabel metal2 9408 24903 9408 24903 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit28.Q
rlabel metal2 7872 24570 7872 24570 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit29.Q
rlabel metal3 14928 23268 14928 23268 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit3.Q
rlabel metal2 9312 22010 9312 22010 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit30.Q
rlabel metal2 7776 22554 7776 22554 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit31.Q
rlabel metal3 16416 24360 16416 24360 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit4.Q
rlabel metal2 6336 34440 6336 34440 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit5.Q
rlabel metal2 6144 34776 6144 34776 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit6.Q
rlabel metal2 7680 33726 7680 33726 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit7.Q
rlabel metal2 5472 37128 5472 37128 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit8.Q
rlabel metal3 5664 36120 5664 36120 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame8_bit9.Q
rlabel metal2 14400 23310 14400 23310 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit10.Q
rlabel metal2 12672 23730 12672 23730 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit11.Q
rlabel metal2 12480 33383 12480 33383 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit12.Q
rlabel metal2 10896 33012 10896 33012 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit13.Q
rlabel metal2 9888 36957 9888 36957 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit14.Q
rlabel metal2 8352 36960 8352 36960 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit15.Q
rlabel metal2 14592 42217 14592 42217 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit16.Q
rlabel metal2 13056 42210 13056 42210 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit17.Q
rlabel metal3 2364 24612 2364 24612 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit18.Q
rlabel metal2 2688 20706 2688 20706 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit19.Q
rlabel metal2 2304 32634 2304 32634 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit20.Q
rlabel metal2 3120 31500 3120 31500 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit21.Q
rlabel metal2 3264 34650 3264 34650 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit22.Q
rlabel metal2 2688 34146 2688 34146 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit23.Q
rlabel metal2 4464 26292 4464 26292 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit24.Q
rlabel metal2 2640 22512 2640 22512 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit25.Q
rlabel metal2 5376 38556 5376 38556 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit26.Q
rlabel metal2 6960 38388 6960 38388 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit27.Q
rlabel metal2 4272 29316 4272 29316 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit28.Q
rlabel metal2 2256 29820 2256 29820 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit29.Q
rlabel metal3 5040 30828 5040 30828 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit30.Q
rlabel metal2 2736 25536 2736 25536 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_ConfigMem.Inst_frame9_bit31.Q
rlabel metal2 9984 16212 9984 16212 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG10
rlabel metal3 17952 19404 17952 19404 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG11
rlabel metal2 17088 13146 17088 13146 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG12
rlabel metal3 14304 16044 14304 16044 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG13
rlabel metal2 13344 35826 13344 35826 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG14
rlabel metal2 16800 18186 16800 18186 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG15
rlabel metal2 19200 16254 19200 16254 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG4
rlabel metal2 14304 19026 14304 19026 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG5
rlabel metal2 13536 32928 13536 32928 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG6
rlabel metal2 13728 12684 13728 12684 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG7
rlabel metal2 19296 16002 19296 16002 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG8
rlabel metal2 15792 31332 15792 31332 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.J_NS4_BEG9
rlabel metal3 14112 21084 14112 21084 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG0
rlabel metal5 8304 23940 8304 23940 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG1
rlabel metal3 9120 31164 9120 31164 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG2
rlabel metal4 14544 22596 14544 22596 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S1BEG3
rlabel metal3 4512 10080 4512 10080 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG0
rlabel metal3 5808 6636 5808 6636 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG1
rlabel metal2 1152 15372 1152 15372 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG2
rlabel metal3 10224 24696 10224 24696 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG3
rlabel metal3 8976 2688 8976 2688 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG4
rlabel metal3 7824 3780 7824 3780 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG5
rlabel metal3 7104 6048 7104 6048 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG6
rlabel metal3 11856 16044 11856 16044 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S2BEG7
rlabel metal2 18192 15708 18192 15708 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG0
rlabel metal3 16272 18900 16272 18900 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG1
rlabel metal4 17184 10668 17184 10668 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG2
rlabel metal3 16032 17640 16032 17640 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.S4BEG3
rlabel metal2 18336 5124 18336 5124 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG0
rlabel metal2 11808 12684 11808 12684 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG1
rlabel metal2 10368 13692 10368 13692 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG2
rlabel metal2 19392 8736 19392 8736 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W1BEG3
rlabel metal2 7728 7896 7728 7896 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG0
rlabel metal2 5424 11844 5424 11844 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG1
rlabel metal2 4416 10122 4416 10122 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG2
rlabel metal2 13536 3906 13536 3906 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG3
rlabel metal3 6576 6972 6576 6972 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG4
rlabel metal3 2352 12012 2352 12012 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG5
rlabel metal2 4800 8778 4800 8778 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG6
rlabel metal3 1728 12390 1728 12390 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEG7
rlabel metal3 7776 8904 7776 8904 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb0
rlabel metal2 1440 17472 1440 17472 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb1
rlabel metal2 7488 10584 7488 10584 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb2
rlabel metal2 13488 2520 13488 2520 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb3
rlabel metal2 9408 7098 9408 7098 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb4
rlabel metal3 5424 12768 5424 12768 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb5
rlabel metal2 4656 5712 4656 5712 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb6
rlabel metal2 11136 6678 11136 6678 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W2BEGb7
rlabel metal2 13728 8988 13728 8988 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG0
rlabel metal2 12096 14910 12096 14910 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG1
rlabel metal2 7968 14700 7968 14700 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG10
rlabel metal3 17472 16296 17472 16296 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG11
rlabel metal2 10512 12432 10512 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG2
rlabel metal3 17952 13272 17952 13272 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG3
rlabel metal3 12192 11172 12192 11172 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG4
rlabel metal3 5472 14784 5472 14784 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG5
rlabel metal2 2016 13188 2016 13188 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG6
rlabel metal3 17088 14784 17088 14784 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG7
rlabel metal2 14352 12432 14352 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG8
rlabel metal2 2112 21588 2112 21588 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.W6BEG9
rlabel metal2 1728 14616 1728 14616 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG0
rlabel metal2 3168 1512 3168 1512 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG1
rlabel metal2 1728 11004 1728 11004 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG10
rlabel metal2 2400 9198 2400 9198 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG11
rlabel metal3 14400 11508 14400 11508 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG12
rlabel metal4 2112 12432 2112 12432 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG13
rlabel metal3 5328 11760 5328 11760 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG14
rlabel metal3 16320 12390 16320 12390 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG15
rlabel metal2 1728 3906 1728 3906 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG2
rlabel metal2 15840 4746 15840 4746 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG3
rlabel metal2 9888 8736 9888 8736 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG4
rlabel metal2 1728 5964 1728 5964 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG5
rlabel metal3 5184 7896 5184 7896 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG6
rlabel metal2 2112 5544 2112 5544 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG7
rlabel metal2 11712 8988 11712 8988 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG8
rlabel metal3 2064 12264 2064 12264 0 Tile_X0Y1_IHP_SRAM_bot.Inst_IHP_SRAM_bot_switch_matrix.WW4BEG9
rlabel metal2 14832 19404 14832 19404 0 Tile_X0Y1_N1END[0]
rlabel metal2 12864 14994 12864 14994 0 Tile_X0Y1_N1END[1]
rlabel metal3 2064 4536 2064 4536 0 Tile_X0Y1_N1END[2]
rlabel metal2 18480 12516 18480 12516 0 Tile_X0Y1_N1END[3]
rlabel metal2 4128 870 4128 870 0 Tile_X0Y1_N2END[0]
rlabel metal2 4320 912 4320 912 0 Tile_X0Y1_N2END[1]
rlabel metal2 4512 450 4512 450 0 Tile_X0Y1_N2END[2]
rlabel metal2 4704 492 4704 492 0 Tile_X0Y1_N2END[3]
rlabel metal2 4896 324 4896 324 0 Tile_X0Y1_N2END[4]
rlabel metal2 5088 324 5088 324 0 Tile_X0Y1_N2END[5]
rlabel metal2 5280 240 5280 240 0 Tile_X0Y1_N2END[6]
rlabel metal3 7824 3612 7824 3612 0 Tile_X0Y1_N2END[7]
rlabel metal2 2592 492 2592 492 0 Tile_X0Y1_N2MID[0]
rlabel metal3 5616 67620 5616 67620 0 Tile_X0Y1_N2MID[1]
rlabel metal2 2976 324 2976 324 0 Tile_X0Y1_N2MID[2]
rlabel metal2 3168 534 3168 534 0 Tile_X0Y1_N2MID[3]
rlabel metal2 3360 282 3360 282 0 Tile_X0Y1_N2MID[4]
rlabel metal2 3264 1596 3264 1596 0 Tile_X0Y1_N2MID[5]
rlabel metal2 3744 660 3744 660 0 Tile_X0Y1_N2MID[6]
rlabel metal2 3936 366 3936 366 0 Tile_X0Y1_N2MID[7]
rlabel metal2 12480 8610 12480 8610 0 Tile_X0Y1_N4END[0]
rlabel metal3 5184 1050 5184 1050 0 Tile_X0Y1_N4END[10]
rlabel metal3 7440 3108 7440 3108 0 Tile_X0Y1_N4END[11]
rlabel metal3 1920 126 1920 126 0 Tile_X0Y1_N4END[12]
rlabel metal2 8112 3192 8112 3192 0 Tile_X0Y1_N4END[13]
rlabel metal2 8352 660 8352 660 0 Tile_X0Y1_N4END[14]
rlabel metal2 8544 156 8544 156 0 Tile_X0Y1_N4END[15]
rlabel metal2 13248 15876 13248 15876 0 Tile_X0Y1_N4END[1]
rlabel metal3 8400 11676 8400 11676 0 Tile_X0Y1_N4END[2]
rlabel metal2 6240 114 6240 114 0 Tile_X0Y1_N4END[3]
rlabel metal2 6432 618 6432 618 0 Tile_X0Y1_N4END[4]
rlabel metal2 6624 366 6624 366 0 Tile_X0Y1_N4END[5]
rlabel metal2 6816 576 6816 576 0 Tile_X0Y1_N4END[6]
rlabel metal2 7008 198 7008 198 0 Tile_X0Y1_N4END[7]
rlabel metal2 7200 492 7200 492 0 Tile_X0Y1_N4END[8]
rlabel metal2 7248 5460 7248 5460 0 Tile_X0Y1_N4END[9]
rlabel metal2 8736 576 8736 576 0 Tile_X0Y1_S1BEG[0]
rlabel metal2 8928 660 8928 660 0 Tile_X0Y1_S1BEG[1]
rlabel metal2 9120 870 9120 870 0 Tile_X0Y1_S1BEG[2]
rlabel metal2 9312 282 9312 282 0 Tile_X0Y1_S1BEG[3]
rlabel metal2 9504 870 9504 870 0 Tile_X0Y1_S2BEG[0]
rlabel metal2 9696 576 9696 576 0 Tile_X0Y1_S2BEG[1]
rlabel metal2 9888 912 9888 912 0 Tile_X0Y1_S2BEG[2]
rlabel metal2 10080 324 10080 324 0 Tile_X0Y1_S2BEG[3]
rlabel metal2 10272 534 10272 534 0 Tile_X0Y1_S2BEG[4]
rlabel metal2 10464 366 10464 366 0 Tile_X0Y1_S2BEG[5]
rlabel metal2 10656 492 10656 492 0 Tile_X0Y1_S2BEG[6]
rlabel metal2 10848 324 10848 324 0 Tile_X0Y1_S2BEG[7]
rlabel metal2 11040 156 11040 156 0 Tile_X0Y1_S2BEGb[0]
rlabel metal2 11232 534 11232 534 0 Tile_X0Y1_S2BEGb[1]
rlabel metal2 11424 1794 11424 1794 0 Tile_X0Y1_S2BEGb[2]
rlabel metal2 11616 1122 11616 1122 0 Tile_X0Y1_S2BEGb[3]
rlabel metal2 11808 828 11808 828 0 Tile_X0Y1_S2BEGb[4]
rlabel metal2 12000 870 12000 870 0 Tile_X0Y1_S2BEGb[5]
rlabel metal2 12192 1458 12192 1458 0 Tile_X0Y1_S2BEGb[6]
rlabel metal2 12384 660 12384 660 0 Tile_X0Y1_S2BEGb[7]
rlabel metal2 12576 492 12576 492 0 Tile_X0Y1_S4BEG[0]
rlabel metal2 14496 912 14496 912 0 Tile_X0Y1_S4BEG[10]
rlabel metal2 19968 1008 19968 1008 0 Tile_X0Y1_S4BEG[11]
rlabel metal2 18048 714 18048 714 0 Tile_X0Y1_S4BEG[12]
rlabel metal3 15744 3192 15744 3192 0 Tile_X0Y1_S4BEG[13]
rlabel metal2 15264 156 15264 156 0 Tile_X0Y1_S4BEG[14]
rlabel metal2 15456 786 15456 786 0 Tile_X0Y1_S4BEG[15]
rlabel metal2 12768 660 12768 660 0 Tile_X0Y1_S4BEG[1]
rlabel metal2 12960 492 12960 492 0 Tile_X0Y1_S4BEG[2]
rlabel metal2 13152 618 13152 618 0 Tile_X0Y1_S4BEG[3]
rlabel metal2 13344 660 13344 660 0 Tile_X0Y1_S4BEG[4]
rlabel metal2 13536 450 13536 450 0 Tile_X0Y1_S4BEG[5]
rlabel metal2 13728 408 13728 408 0 Tile_X0Y1_S4BEG[6]
rlabel metal2 13920 492 13920 492 0 Tile_X0Y1_S4BEG[7]
rlabel metal2 14016 3192 14016 3192 0 Tile_X0Y1_S4BEG[8]
rlabel metal2 14304 492 14304 492 0 Tile_X0Y1_S4BEG[9]
rlabel metal2 15648 408 15648 408 0 Tile_X0Y1_UserCLK
rlabel metal3 126 84 126 84 0 Tile_X0Y1_W1BEG[0]
rlabel metal4 8448 1176 8448 1176 0 Tile_X0Y1_W1BEG[1]
rlabel metal3 750 756 750 756 0 Tile_X0Y1_W1BEG[2]
rlabel metal3 1230 1092 1230 1092 0 Tile_X0Y1_W1BEG[3]
rlabel metal3 126 1428 126 1428 0 Tile_X0Y1_W2BEG[0]
rlabel metal3 126 1764 126 1764 0 Tile_X0Y1_W2BEG[1]
rlabel metal3 318 2100 318 2100 0 Tile_X0Y1_W2BEG[2]
rlabel metal3 4440 2436 4440 2436 0 Tile_X0Y1_W2BEG[3]
rlabel metal3 462 2772 462 2772 0 Tile_X0Y1_W2BEG[4]
rlabel metal3 1182 3108 1182 3108 0 Tile_X0Y1_W2BEG[5]
rlabel metal3 222 3444 222 3444 0 Tile_X0Y1_W2BEG[6]
rlabel metal3 990 3780 990 3780 0 Tile_X0Y1_W2BEG[7]
rlabel metal4 4128 6678 4128 6678 0 Tile_X0Y1_W2BEGb[0]
rlabel metal3 672 16044 672 16044 0 Tile_X0Y1_W2BEGb[1]
rlabel metal3 6864 9996 6864 9996 0 Tile_X0Y1_W2BEGb[2]
rlabel metal3 702 5124 702 5124 0 Tile_X0Y1_W2BEGb[3]
rlabel metal3 9216 5628 9216 5628 0 Tile_X0Y1_W2BEGb[4]
rlabel metal3 1290 5796 1290 5796 0 Tile_X0Y1_W2BEGb[5]
rlabel metal3 126 6132 126 6132 0 Tile_X0Y1_W2BEGb[6]
rlabel metal3 78 6468 78 6468 0 Tile_X0Y1_W2BEGb[7]
rlabel metal2 13536 9870 13536 9870 0 Tile_X0Y1_W6BEG[0]
rlabel metal2 2880 15456 2880 15456 0 Tile_X0Y1_W6BEG[10]
rlabel metal2 17472 15960 17472 15960 0 Tile_X0Y1_W6BEG[11]
rlabel metal2 11136 12432 11136 12432 0 Tile_X0Y1_W6BEG[1]
rlabel metal3 1038 12852 1038 12852 0 Tile_X0Y1_W6BEG[2]
rlabel metal3 414 13188 414 13188 0 Tile_X0Y1_W6BEG[3]
rlabel metal2 12192 12726 12192 12726 0 Tile_X0Y1_W6BEG[4]
rlabel metal2 3648 14196 3648 14196 0 Tile_X0Y1_W6BEG[5]
rlabel metal2 1824 13818 1824 13818 0 Tile_X0Y1_W6BEG[6]
rlabel metal3 654 14532 654 14532 0 Tile_X0Y1_W6BEG[7]
rlabel metal3 1134 14868 1134 14868 0 Tile_X0Y1_W6BEG[8]
rlabel metal3 990 15204 990 15204 0 Tile_X0Y1_W6BEG[9]
rlabel metal3 1152 13188 1152 13188 0 Tile_X0Y1_WW4BEG[0]
rlabel metal3 798 10164 798 10164 0 Tile_X0Y1_WW4BEG[10]
rlabel metal2 2208 10080 2208 10080 0 Tile_X0Y1_WW4BEG[11]
rlabel metal3 7278 10836 7278 10836 0 Tile_X0Y1_WW4BEG[12]
rlabel metal3 990 11172 990 11172 0 Tile_X0Y1_WW4BEG[13]
rlabel metal3 1470 11508 1470 11508 0 Tile_X0Y1_WW4BEG[14]
rlabel metal3 990 11844 990 11844 0 Tile_X0Y1_WW4BEG[15]
rlabel metal3 2016 924 2016 924 0 Tile_X0Y1_WW4BEG[1]
rlabel metal2 1584 3612 1584 3612 0 Tile_X0Y1_WW4BEG[2]
rlabel metal2 2880 2142 2880 2142 0 Tile_X0Y1_WW4BEG[3]
rlabel metal3 942 8148 942 8148 0 Tile_X0Y1_WW4BEG[4]
rlabel metal2 1488 5880 1488 5880 0 Tile_X0Y1_WW4BEG[5]
rlabel metal2 3264 8484 3264 8484 0 Tile_X0Y1_WW4BEG[6]
rlabel metal2 1920 7518 1920 7518 0 Tile_X0Y1_WW4BEG[7]
rlabel metal3 1566 9492 1566 9492 0 Tile_X0Y1_WW4BEG[8]
rlabel metal2 1440 9744 1440 9744 0 Tile_X0Y1_WW4BEG[9]
rlabel via2 21426 49308 21426 49308 0 WEN_SRAM
rlabel metal2 9600 39228 9600 39228 0 _0000_
rlabel metal2 2592 39942 2592 39942 0 _0001_
rlabel metal2 9120 43008 9120 43008 0 _0002_
rlabel metal2 14784 59892 14784 59892 0 _0003_
rlabel metal2 10560 70602 10560 70602 0 _0004_
rlabel metal2 16128 74550 16128 74550 0 _0005_
rlabel metal2 10464 73206 10464 73206 0 _0006_
rlabel metal3 15168 26964 15168 26964 0 _0007_
rlabel metal3 9936 32172 9936 32172 0 _0008_
rlabel metal3 11808 27636 11808 27636 0 _0009_
rlabel metal2 15936 21798 15936 21798 0 _0010_
rlabel metal2 8640 78372 8640 78372 0 _0011_
rlabel metal3 8736 48804 8736 48804 0 _0012_
rlabel metal2 9312 66444 9312 66444 0 _0013_
rlabel metal2 11904 80976 11904 80976 0 _0014_
rlabel metal3 11952 70644 11952 70644 0 _0015_
rlabel metal3 16128 57036 16128 57036 0 _0016_
rlabel metal2 15648 52038 15648 52038 0 _0017_
rlabel metal3 19248 79968 19248 79968 0 _0018_
rlabel metal2 15072 25284 15072 25284 0 _0019_
rlabel metal2 16896 24612 16896 24612 0 _0020_
rlabel metal2 7392 34356 7392 34356 0 _0021_
rlabel metal3 6672 33684 6672 33684 0 _0022_
rlabel metal2 5712 35868 5712 35868 0 _0023_
rlabel metal3 6816 36708 6816 36708 0 _0024_
rlabel metal2 13200 41244 13200 41244 0 _0025_
rlabel metal3 13728 39480 13728 39480 0 _0026_
rlabel metal2 18624 18270 18624 18270 0 _0027_
rlabel metal2 19776 14952 19776 14952 0 _0028_
rlabel metal3 12768 29148 12768 29148 0 _0029_
rlabel metal3 14112 29064 14112 29064 0 _0030_
rlabel metal2 6816 29316 6816 29316 0 _0031_
rlabel metal2 7488 28140 7488 28140 0 _0032_
rlabel metal2 14880 19194 14880 19194 0 _0033_
rlabel metal2 17664 19404 17664 19404 0 _0034_
rlabel metal2 10848 40614 10848 40614 0 _0035_
rlabel metal2 7968 43428 7968 43428 0 _0036_
rlabel metal2 2976 40824 2976 40824 0 _0037_
rlabel metal2 7949 73668 7949 73668 0 _0038_
rlabel via1 7202 66108 7202 66108 0 _0039_
rlabel metal3 10205 64596 10205 64596 0 _0040_
rlabel metal2 6336 75516 6336 75516 0 _0041_
rlabel via2 1437 79800 1437 79800 0 _0042_
rlabel metal2 5232 2100 5232 2100 0 _0043_
rlabel metal3 9840 40404 9840 40404 0 _0044_
rlabel metal2 9888 40530 9888 40530 0 _0045_
rlabel metal2 9600 41118 9600 41118 0 _0046_
rlabel metal2 11136 41338 11136 41338 0 _0047_
rlabel metal2 9408 42252 9408 42252 0 _0048_
rlabel metal2 10560 41496 10560 41496 0 _0049_
rlabel metal2 10656 41412 10656 41412 0 _0050_
rlabel metal2 11040 41202 11040 41202 0 _0051_
rlabel metal3 15408 41244 15408 41244 0 _0052_
rlabel metal2 9840 39816 9840 39816 0 _0053_
rlabel metal2 9600 39732 9600 39732 0 _0054_
rlabel metal3 15654 40404 15654 40404 0 _0055_
rlabel metal2 20160 40572 20160 40572 0 _0056_
rlabel metal3 15072 60900 15072 60900 0 _0057_
rlabel metal2 14496 60858 14496 60858 0 _0058_
rlabel metal3 15216 61068 15216 61068 0 _0059_
rlabel metal3 12528 15456 12528 15456 0 _0060_
rlabel metal2 12864 27720 12864 27720 0 _0061_
rlabel metal2 12480 27300 12480 27300 0 _0062_
rlabel metal2 11952 33684 11952 33684 0 _0063_
rlabel metal2 11040 71652 11040 71652 0 _0064_
rlabel metal2 11520 70980 11520 70980 0 _0065_
rlabel metal2 9408 70770 9408 70770 0 _0066_
rlabel metal2 8832 16170 8832 16170 0 _0067_
rlabel metal2 8544 32844 8544 32844 0 _0068_
rlabel metal2 9072 33852 9072 33852 0 _0069_
rlabel metal2 9504 33432 9504 33432 0 _0070_
rlabel metal3 15696 75012 15696 75012 0 _0071_
rlabel metal2 15744 75516 15744 75516 0 _0072_
rlabel metal3 17184 75180 17184 75180 0 _0073_
rlabel metal3 18144 14028 18144 14028 0 _0074_
rlabel metal2 15072 27300 15072 27300 0 _0075_
rlabel metal2 15504 26292 15504 26292 0 _0076_
rlabel metal3 14880 36120 14880 36120 0 _0077_
rlabel metal2 3840 7308 3840 7308 0 _0078_
rlabel metal2 2880 37086 2880 37086 0 _0079_
rlabel metal2 16224 14826 16224 14826 0 _0080_
rlabel metal2 18432 18396 18432 18396 0 _0081_
rlabel metal2 12960 29363 12960 29363 0 _0082_
rlabel metal2 7248 14028 7248 14028 0 _0083_
rlabel metal3 16080 16212 16080 16212 0 _0084_
rlabel metal2 9984 74256 9984 74256 0 _0085_
rlabel metal2 10080 73416 10080 73416 0 _0086_
rlabel metal3 14496 74550 14496 74550 0 _0087_
rlabel metal2 18528 8442 18528 8442 0 _0088_
rlabel metal3 15168 21588 15168 21588 0 _0089_
rlabel metal2 15648 21084 15648 21084 0 _0090_
rlabel metal3 14544 22260 14544 22260 0 _0091_
rlabel metal2 7296 73752 7296 73752 0 _0092_
rlabel metal3 7776 73164 7776 73164 0 _0093_
rlabel metal2 5760 66024 5760 66024 0 _0094_
rlabel metal3 7392 65940 7392 65940 0 _0095_
rlabel metal2 9504 65447 9504 65447 0 _0096_
rlabel metal2 9792 64344 9792 64344 0 _0097_
rlabel metal3 7632 76020 7632 76020 0 _0098_
rlabel metal2 6912 76104 6912 76104 0 _0099_
rlabel metal2 2064 76860 2064 76860 0 _0100_
rlabel metal3 1632 79674 1632 79674 0 _0101_
rlabel metal2 8064 78750 8064 78750 0 _0102_
rlabel metal2 8064 77448 8064 77448 0 _0103_
rlabel metal2 8160 77490 8160 77490 0 _0104_
rlabel metal2 8352 78456 8352 78456 0 _0105_
rlabel metal2 7728 78876 7728 78876 0 _0106_
rlabel metal2 8016 77700 8016 77700 0 _0107_
rlabel metal4 8256 79170 8256 79170 0 _0108_
rlabel metal2 7968 48930 7968 48930 0 _0109_
rlabel metal2 10320 49476 10320 49476 0 _0110_
rlabel metal2 10416 48972 10416 48972 0 _0111_
rlabel metal2 8256 48888 8256 48888 0 _0112_
rlabel metal3 8448 47964 8448 47964 0 _0113_
rlabel metal2 10848 49434 10848 49434 0 _0114_
rlabel metal3 9888 47964 9888 47964 0 _0115_
rlabel metal2 10656 67200 10656 67200 0 _0116_
rlabel metal3 8688 67620 8688 67620 0 _0117_
rlabel metal2 9984 67830 9984 67830 0 _0118_
rlabel metal3 10272 67620 10272 67620 0 _0119_
rlabel metal2 10368 68502 10368 68502 0 _0120_
rlabel metal2 9744 68460 9744 68460 0 _0121_
rlabel metal3 9264 68376 9264 68376 0 _0122_
rlabel metal2 12048 81228 12048 81228 0 _0123_
rlabel metal2 12480 82488 12480 82488 0 _0124_
rlabel metal2 11520 81270 11520 81270 0 _0125_
rlabel metal3 12240 81060 12240 81060 0 _0126_
rlabel metal2 11568 82236 11568 82236 0 _0127_
rlabel metal3 11904 80640 11904 80640 0 _0128_
rlabel metal2 12384 82488 12384 82488 0 _0129_
rlabel metal2 12000 70728 12000 70728 0 _0130_
rlabel metal2 13680 72240 13680 72240 0 _0131_
rlabel metal2 13344 73458 13344 73458 0 _0132_
rlabel metal2 12432 70644 12432 70644 0 _0133_
rlabel metal3 14496 70644 14496 70644 0 _0134_
rlabel metal2 14400 71526 14400 71526 0 _0135_
rlabel metal2 15072 70770 15072 70770 0 _0136_
rlabel metal3 16800 55020 16800 55020 0 _0137_
rlabel metal2 16896 57078 16896 57078 0 _0138_
rlabel metal2 17376 56532 17376 56532 0 _0139_
rlabel metal2 16992 56868 16992 56868 0 _0140_
rlabel metal3 17232 56364 17232 56364 0 _0141_
rlabel metal2 16992 56574 16992 56574 0 _0142_
rlabel metal2 17616 56364 17616 56364 0 _0143_
rlabel metal3 15648 50988 15648 50988 0 _0144_
rlabel metal3 14592 50988 14592 50988 0 _0145_
rlabel metal2 14784 51072 14784 51072 0 _0146_
rlabel metal2 15360 50988 15360 50988 0 _0147_
rlabel metal3 15840 51240 15840 51240 0 _0148_
rlabel metal2 16609 51875 16609 51875 0 _0149_
rlabel metal2 16416 51702 16416 51702 0 _0150_
rlabel metal2 19392 83286 19392 83286 0 _0151_
rlabel metal3 17040 79044 17040 79044 0 _0152_
rlabel metal2 17952 79128 17952 79128 0 _0153_
rlabel metal3 18432 83076 18432 83076 0 _0154_
rlabel metal3 17520 83412 17520 83412 0 _0155_
rlabel metal3 16656 79716 16656 79716 0 _0156_
rlabel metal2 15600 79968 15600 79968 0 _0157_
rlabel metal2 13824 13860 13824 13860 0 _0158_
rlabel metal2 10368 34692 10368 34692 0 _0159_
rlabel metal2 14352 15624 14352 15624 0 _0160_
rlabel metal2 19680 18186 19680 18186 0 _0161_
rlabel metal2 12000 23730 12000 23730 0 _0162_
rlabel metal2 10416 23772 10416 23772 0 _0163_
rlabel metal2 10560 23352 10560 23352 0 _0164_
rlabel metal2 6048 23352 6048 23352 0 _0165_
rlabel metal2 1920 23730 1920 23730 0 _0166_
rlabel metal2 5952 23184 5952 23184 0 _0167_
rlabel metal2 6816 25578 6816 25578 0 _0168_
rlabel metal2 7296 26880 7296 26880 0 _0169_
rlabel metal2 6720 25830 6720 25830 0 _0170_
rlabel metal2 11328 38346 11328 38346 0 _0171_
rlabel metal2 9792 39354 9792 39354 0 _0172_
rlabel metal3 10800 38220 10800 38220 0 _0173_
rlabel metal3 10176 26124 10176 26124 0 _0174_
rlabel metal2 7584 26460 7584 26460 0 _0175_
rlabel metal2 10272 26376 10272 26376 0 _0176_
rlabel metal2 17664 23352 17664 23352 0 _0177_
rlabel metal2 17760 23898 17760 23898 0 _0178_
rlabel metal2 16512 24948 16512 24948 0 _0179_
rlabel metal3 16416 23100 16416 23100 0 _0180_
rlabel metal2 16752 23268 16752 23268 0 _0181_
rlabel metal2 15552 25242 15552 25242 0 _0182_
rlabel metal2 17472 23310 17472 23310 0 _0183_
rlabel metal2 16320 26040 16320 26040 0 _0184_
rlabel metal2 15840 25620 15840 25620 0 _0185_
rlabel metal4 16320 25074 16320 25074 0 _0186_
rlabel metal2 5760 34440 5760 34440 0 _0187_
rlabel metal3 6480 34356 6480 34356 0 _0188_
rlabel metal2 7008 34440 7008 34440 0 _0189_
rlabel metal2 7968 33390 7968 33390 0 _0190_
rlabel metal2 7632 33516 7632 33516 0 _0191_
rlabel metal2 7200 32886 7200 32886 0 _0192_
rlabel metal2 7296 33096 7296 33096 0 _0193_
rlabel metal2 7200 33600 7200 33600 0 _0194_
rlabel metal2 7488 33012 7488 33012 0 _0195_
rlabel metal2 7392 33894 7392 33894 0 _0196_
rlabel metal3 6768 35280 6768 35280 0 _0197_
rlabel metal3 6768 35868 6768 35868 0 _0198_
rlabel metal2 6048 36078 6048 36078 0 _0199_
rlabel metal2 6432 36404 6432 36404 0 _0200_
rlabel metal2 6624 36750 6624 36750 0 _0201_
rlabel metal2 7680 36918 7680 36918 0 _0202_
rlabel metal3 6240 37380 6240 37380 0 _0203_
rlabel metal2 7392 36162 7392 36162 0 _0204_
rlabel metal2 7104 36960 7104 36960 0 _0205_
rlabel metal2 6912 36624 6912 36624 0 _0206_
rlabel metal3 12624 38892 12624 38892 0 _0207_
rlabel metal3 13824 39060 13824 39060 0 _0208_
rlabel metal2 15408 39900 15408 39900 0 _0209_
rlabel metal2 13920 40194 13920 40194 0 _0210_
rlabel metal2 13632 40572 13632 40572 0 _0211_
rlabel metal2 14688 40362 14688 40362 0 _0212_
rlabel metal2 14784 39816 14784 39816 0 _0213_
rlabel metal2 14304 39102 14304 39102 0 _0214_
rlabel metal3 14784 38892 14784 38892 0 _0215_
rlabel metal2 14496 39186 14496 39186 0 _0216_
rlabel metal2 20400 17220 20400 17220 0 _0217_
rlabel metal2 19920 17724 19920 17724 0 _0218_
rlabel metal2 17952 16884 17952 16884 0 _0219_
rlabel metal2 19728 15540 19728 15540 0 _0220_
rlabel metal3 18960 15372 18960 15372 0 _0221_
rlabel metal2 19776 16170 19776 16170 0 _0222_
rlabel metal3 19248 16212 19248 16212 0 _0223_
rlabel metal2 19488 15540 19488 15540 0 _0224_
rlabel metal2 19248 14700 19248 14700 0 _0225_
rlabel metal3 18768 14952 18768 14952 0 _0226_
rlabel metal2 11424 30240 11424 30240 0 _0227_
rlabel metal2 14976 29190 14976 29190 0 _0228_
rlabel metal3 14976 28308 14976 28308 0 _0229_
rlabel metal2 15552 29274 15552 29274 0 _0230_
rlabel metal2 13248 27678 13248 27678 0 _0231_
rlabel metal2 12960 28602 12960 28602 0 _0232_
rlabel metal2 12864 28518 12864 28518 0 _0233_
rlabel metal2 14064 29988 14064 29988 0 _0234_
rlabel metal2 13728 27888 13728 27888 0 _0235_
rlabel metal2 13584 27636 13584 27636 0 _0236_
rlabel metal2 6144 29400 6144 29400 0 _0237_
rlabel metal3 6960 29148 6960 29148 0 _0238_
rlabel metal3 7536 27636 7536 27636 0 _0239_
rlabel metal3 6288 29064 6288 29064 0 _0240_
rlabel metal3 6576 27048 6576 27048 0 _0241_
rlabel metal2 6528 27090 6528 27090 0 _0242_
rlabel metal2 6432 25620 6432 25620 0 _0243_
rlabel metal2 7584 28518 7584 28518 0 _0244_
rlabel metal2 6816 27300 6816 27300 0 _0245_
rlabel metal2 7200 27888 7200 27888 0 _0246_
rlabel metal3 17280 20412 17280 20412 0 _0247_
rlabel metal3 16848 19236 16848 19236 0 _0248_
rlabel metal2 15552 19026 15552 19026 0 _0249_
rlabel metal2 17760 19992 17760 19992 0 _0250_
rlabel metal2 15072 19530 15072 19530 0 _0251_
rlabel metal2 17184 18826 17184 18826 0 _0252_
rlabel metal2 17280 18522 17280 18522 0 _0253_
rlabel metal2 16800 20118 16800 20118 0 _0254_
rlabel metal2 17424 18732 17424 18732 0 _0255_
rlabel metal3 16176 20580 16176 20580 0 _0256_
rlabel metal2 7104 40908 7104 40908 0 _0257_
rlabel metal2 7440 42588 7440 42588 0 _0258_
rlabel metal2 7392 41160 7392 41160 0 _0259_
rlabel metal3 6768 40656 6768 40656 0 _0260_
rlabel via1 7018 41244 7018 41244 0 _0261_
rlabel metal2 10752 40152 10752 40152 0 _0262_
rlabel metal2 7776 41412 7776 41412 0 _0263_
rlabel metal2 8112 40404 8112 40404 0 _0264_
rlabel metal3 8640 40656 8640 40656 0 _0265_
rlabel metal3 8400 40404 8400 40404 0 _0266_
rlabel metal2 6192 40404 6192 40404 0 _0267_
rlabel metal2 6192 40656 6192 40656 0 _0268_
rlabel metal2 7872 40488 7872 40488 0 _0269_
rlabel metal2 8160 41118 8160 41118 0 _0270_
rlabel metal2 7200 41790 7200 41790 0 _0271_
rlabel metal2 8160 41832 8160 41832 0 _0272_
rlabel metal3 7920 41916 7920 41916 0 _0273_
rlabel metal2 8448 42000 8448 42000 0 _0274_
rlabel metal2 8640 42252 8640 42252 0 _0275_
rlabel metal2 8544 41916 8544 41916 0 _0276_
rlabel metal2 8352 43176 8352 43176 0 _0277_
rlabel metal2 8064 42966 8064 42966 0 _0278_
rlabel metal2 4320 40446 4320 40446 0 _0279_
rlabel metal3 4416 39816 4416 39816 0 _0280_
rlabel metal2 4704 39984 4704 39984 0 _0281_
rlabel metal2 4032 41370 4032 41370 0 _0282_
rlabel metal2 4800 43134 4800 43134 0 _0283_
rlabel metal2 2016 40698 2016 40698 0 _0284_
rlabel metal3 4032 41160 4032 41160 0 _0285_
rlabel metal3 4416 40404 4416 40404 0 _0286_
rlabel metal2 4512 40530 4512 40530 0 _0287_
rlabel metal2 3360 42252 3360 42252 0 _0288_
rlabel metal2 3504 41076 3504 41076 0 _0289_
rlabel metal3 4128 41916 4128 41916 0 _0290_
rlabel metal2 3552 42294 3552 42294 0 _0291_
rlabel metal2 2880 42210 2880 42210 0 _0292_
rlabel metal2 4032 41874 4032 41874 0 _0293_
rlabel metal2 4416 41454 4416 41454 0 _0294_
rlabel metal2 4128 42294 4128 42294 0 _0295_
rlabel metal2 4416 42672 4416 42672 0 _0296_
rlabel metal2 16992 65520 16992 65520 0 clknet_0_Tile_X0Y1_UserCLK
rlabel metal2 19440 54012 19440 54012 0 clknet_1_0__leaf_Tile_X0Y1_UserCLK
rlabel metal2 15840 81312 15840 81312 0 clknet_1_1__leaf_Tile_X0Y1_UserCLK
<< properties >>
string FIXED_BBOX 0 0 21504 86016
<< end >>
