VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO W_TT_IF2
  CLASS BLOCK ;
  FOREIGN W_TT_IF2 ;
  ORIGIN 0.000 0.000 ;
  SIZE 107.520 BY 430.080 ;
  PIN CLK_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 174.100 0.400 174.500 ;
    END
  END CLK_TT_PROJECT
  PIN ENA_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.632400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 170.740 0.400 171.140 ;
    END
  END ENA_TT_PROJECT
  PIN RST_N_TT_PROJECT
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.958400 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 177.460 0.400 177.860 ;
    END
  END RST_N_TT_PROJECT
  PIN Tile_X0Y0_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 295.900 107.520 296.300 ;
    END
  END Tile_X0Y0_E1BEG[0]
  PIN Tile_X0Y0_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 297.580 107.520 297.980 ;
    END
  END Tile_X0Y0_E1BEG[1]
  PIN Tile_X0Y0_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 299.260 107.520 299.660 ;
    END
  END Tile_X0Y0_E1BEG[2]
  PIN Tile_X0Y0_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 300.940 107.520 301.340 ;
    END
  END Tile_X0Y0_E1BEG[3]
  PIN Tile_X0Y0_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 302.620 107.520 303.020 ;
    END
  END Tile_X0Y0_E2BEG[0]
  PIN Tile_X0Y0_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 304.300 107.520 304.700 ;
    END
  END Tile_X0Y0_E2BEG[1]
  PIN Tile_X0Y0_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 305.980 107.520 306.380 ;
    END
  END Tile_X0Y0_E2BEG[2]
  PIN Tile_X0Y0_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 307.660 107.520 308.060 ;
    END
  END Tile_X0Y0_E2BEG[3]
  PIN Tile_X0Y0_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 309.340 107.520 309.740 ;
    END
  END Tile_X0Y0_E2BEG[4]
  PIN Tile_X0Y0_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 311.020 107.520 311.420 ;
    END
  END Tile_X0Y0_E2BEG[5]
  PIN Tile_X0Y0_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 312.700 107.520 313.100 ;
    END
  END Tile_X0Y0_E2BEG[6]
  PIN Tile_X0Y0_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 314.380 107.520 314.780 ;
    END
  END Tile_X0Y0_E2BEG[7]
  PIN Tile_X0Y0_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 316.060 107.520 316.460 ;
    END
  END Tile_X0Y0_E2BEGb[0]
  PIN Tile_X0Y0_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 317.740 107.520 318.140 ;
    END
  END Tile_X0Y0_E2BEGb[1]
  PIN Tile_X0Y0_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 319.420 107.520 319.820 ;
    END
  END Tile_X0Y0_E2BEGb[2]
  PIN Tile_X0Y0_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 321.100 107.520 321.500 ;
    END
  END Tile_X0Y0_E2BEGb[3]
  PIN Tile_X0Y0_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 322.780 107.520 323.180 ;
    END
  END Tile_X0Y0_E2BEGb[4]
  PIN Tile_X0Y0_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 324.460 107.520 324.860 ;
    END
  END Tile_X0Y0_E2BEGb[5]
  PIN Tile_X0Y0_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 326.140 107.520 326.540 ;
    END
  END Tile_X0Y0_E2BEGb[6]
  PIN Tile_X0Y0_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 327.820 107.520 328.220 ;
    END
  END Tile_X0Y0_E2BEGb[7]
  PIN Tile_X0Y0_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 356.380 107.520 356.780 ;
    END
  END Tile_X0Y0_E6BEG[0]
  PIN Tile_X0Y0_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 373.180 107.520 373.580 ;
    END
  END Tile_X0Y0_E6BEG[10]
  PIN Tile_X0Y0_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 374.860 107.520 375.260 ;
    END
  END Tile_X0Y0_E6BEG[11]
  PIN Tile_X0Y0_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 358.060 107.520 358.460 ;
    END
  END Tile_X0Y0_E6BEG[1]
  PIN Tile_X0Y0_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 359.740 107.520 360.140 ;
    END
  END Tile_X0Y0_E6BEG[2]
  PIN Tile_X0Y0_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 361.420 107.520 361.820 ;
    END
  END Tile_X0Y0_E6BEG[3]
  PIN Tile_X0Y0_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 363.100 107.520 363.500 ;
    END
  END Tile_X0Y0_E6BEG[4]
  PIN Tile_X0Y0_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 364.780 107.520 365.180 ;
    END
  END Tile_X0Y0_E6BEG[5]
  PIN Tile_X0Y0_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 366.460 107.520 366.860 ;
    END
  END Tile_X0Y0_E6BEG[6]
  PIN Tile_X0Y0_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 368.140 107.520 368.540 ;
    END
  END Tile_X0Y0_E6BEG[7]
  PIN Tile_X0Y0_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 369.820 107.520 370.220 ;
    END
  END Tile_X0Y0_E6BEG[8]
  PIN Tile_X0Y0_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 371.500 107.520 371.900 ;
    END
  END Tile_X0Y0_E6BEG[9]
  PIN Tile_X0Y0_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 329.500 107.520 329.900 ;
    END
  END Tile_X0Y0_EE4BEG[0]
  PIN Tile_X0Y0_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 346.300 107.520 346.700 ;
    END
  END Tile_X0Y0_EE4BEG[10]
  PIN Tile_X0Y0_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 347.980 107.520 348.380 ;
    END
  END Tile_X0Y0_EE4BEG[11]
  PIN Tile_X0Y0_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 349.660 107.520 350.060 ;
    END
  END Tile_X0Y0_EE4BEG[12]
  PIN Tile_X0Y0_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 351.340 107.520 351.740 ;
    END
  END Tile_X0Y0_EE4BEG[13]
  PIN Tile_X0Y0_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 353.020 107.520 353.420 ;
    END
  END Tile_X0Y0_EE4BEG[14]
  PIN Tile_X0Y0_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 354.700 107.520 355.100 ;
    END
  END Tile_X0Y0_EE4BEG[15]
  PIN Tile_X0Y0_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 331.180 107.520 331.580 ;
    END
  END Tile_X0Y0_EE4BEG[1]
  PIN Tile_X0Y0_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 332.860 107.520 333.260 ;
    END
  END Tile_X0Y0_EE4BEG[2]
  PIN Tile_X0Y0_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 334.540 107.520 334.940 ;
    END
  END Tile_X0Y0_EE4BEG[3]
  PIN Tile_X0Y0_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 336.220 107.520 336.620 ;
    END
  END Tile_X0Y0_EE4BEG[4]
  PIN Tile_X0Y0_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 337.900 107.520 338.300 ;
    END
  END Tile_X0Y0_EE4BEG[5]
  PIN Tile_X0Y0_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 339.580 107.520 339.980 ;
    END
  END Tile_X0Y0_EE4BEG[6]
  PIN Tile_X0Y0_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 341.260 107.520 341.660 ;
    END
  END Tile_X0Y0_EE4BEG[7]
  PIN Tile_X0Y0_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 342.940 107.520 343.340 ;
    END
  END Tile_X0Y0_EE4BEG[8]
  PIN Tile_X0Y0_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 344.620 107.520 345.020 ;
    END
  END Tile_X0Y0_EE4BEG[9]
  PIN Tile_X0Y0_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.445600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 180.820 0.400 181.220 ;
    END
  END Tile_X0Y0_FrameData[0]
  PIN Tile_X0Y0_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.420 0.400 214.820 ;
    END
  END Tile_X0Y0_FrameData[10]
  PIN Tile_X0Y0_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 217.780 0.400 218.180 ;
    END
  END Tile_X0Y0_FrameData[11]
  PIN Tile_X0Y0_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 221.140 0.400 221.540 ;
    END
  END Tile_X0Y0_FrameData[12]
  PIN Tile_X0Y0_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 224.500 0.400 224.900 ;
    END
  END Tile_X0Y0_FrameData[13]
  PIN Tile_X0Y0_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 227.860 0.400 228.260 ;
    END
  END Tile_X0Y0_FrameData[14]
  PIN Tile_X0Y0_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 231.220 0.400 231.620 ;
    END
  END Tile_X0Y0_FrameData[15]
  PIN Tile_X0Y0_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 234.580 0.400 234.980 ;
    END
  END Tile_X0Y0_FrameData[16]
  PIN Tile_X0Y0_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 237.940 0.400 238.340 ;
    END
  END Tile_X0Y0_FrameData[17]
  PIN Tile_X0Y0_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 241.300 0.400 241.700 ;
    END
  END Tile_X0Y0_FrameData[18]
  PIN Tile_X0Y0_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 244.660 0.400 245.060 ;
    END
  END Tile_X0Y0_FrameData[19]
  PIN Tile_X0Y0_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.445600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 184.180 0.400 184.580 ;
    END
  END Tile_X0Y0_FrameData[1]
  PIN Tile_X0Y0_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 248.020 0.400 248.420 ;
    END
  END Tile_X0Y0_FrameData[20]
  PIN Tile_X0Y0_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 251.380 0.400 251.780 ;
    END
  END Tile_X0Y0_FrameData[21]
  PIN Tile_X0Y0_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.740 0.400 255.140 ;
    END
  END Tile_X0Y0_FrameData[22]
  PIN Tile_X0Y0_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 258.100 0.400 258.500 ;
    END
  END Tile_X0Y0_FrameData[23]
  PIN Tile_X0Y0_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 261.460 0.400 261.860 ;
    END
  END Tile_X0Y0_FrameData[24]
  PIN Tile_X0Y0_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 264.820 0.400 265.220 ;
    END
  END Tile_X0Y0_FrameData[25]
  PIN Tile_X0Y0_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 268.180 0.400 268.580 ;
    END
  END Tile_X0Y0_FrameData[26]
  PIN Tile_X0Y0_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 271.540 0.400 271.940 ;
    END
  END Tile_X0Y0_FrameData[27]
  PIN Tile_X0Y0_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 274.900 0.400 275.300 ;
    END
  END Tile_X0Y0_FrameData[28]
  PIN Tile_X0Y0_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.260 0.400 278.660 ;
    END
  END Tile_X0Y0_FrameData[29]
  PIN Tile_X0Y0_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.445600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 187.540 0.400 187.940 ;
    END
  END Tile_X0Y0_FrameData[2]
  PIN Tile_X0Y0_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 281.620 0.400 282.020 ;
    END
  END Tile_X0Y0_FrameData[30]
  PIN Tile_X0Y0_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 284.980 0.400 285.380 ;
    END
  END Tile_X0Y0_FrameData[31]
  PIN Tile_X0Y0_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.445600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 190.900 0.400 191.300 ;
    END
  END Tile_X0Y0_FrameData[3]
  PIN Tile_X0Y0_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.445600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 194.260 0.400 194.660 ;
    END
  END Tile_X0Y0_FrameData[4]
  PIN Tile_X0Y0_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.445600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 197.620 0.400 198.020 ;
    END
  END Tile_X0Y0_FrameData[5]
  PIN Tile_X0Y0_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.445600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 200.980 0.400 201.380 ;
    END
  END Tile_X0Y0_FrameData[6]
  PIN Tile_X0Y0_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.445600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 204.340 0.400 204.740 ;
    END
  END Tile_X0Y0_FrameData[7]
  PIN Tile_X0Y0_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 207.700 0.400 208.100 ;
    END
  END Tile_X0Y0_FrameData[8]
  PIN Tile_X0Y0_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 211.060 0.400 211.460 ;
    END
  END Tile_X0Y0_FrameData[9]
  PIN Tile_X0Y0_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 376.540 107.520 376.940 ;
    END
  END Tile_X0Y0_FrameData_O[0]
  PIN Tile_X0Y0_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 393.340 107.520 393.740 ;
    END
  END Tile_X0Y0_FrameData_O[10]
  PIN Tile_X0Y0_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 395.020 107.520 395.420 ;
    END
  END Tile_X0Y0_FrameData_O[11]
  PIN Tile_X0Y0_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 396.700 107.520 397.100 ;
    END
  END Tile_X0Y0_FrameData_O[12]
  PIN Tile_X0Y0_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 398.380 107.520 398.780 ;
    END
  END Tile_X0Y0_FrameData_O[13]
  PIN Tile_X0Y0_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 400.060 107.520 400.460 ;
    END
  END Tile_X0Y0_FrameData_O[14]
  PIN Tile_X0Y0_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 401.740 107.520 402.140 ;
    END
  END Tile_X0Y0_FrameData_O[15]
  PIN Tile_X0Y0_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 403.420 107.520 403.820 ;
    END
  END Tile_X0Y0_FrameData_O[16]
  PIN Tile_X0Y0_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 405.100 107.520 405.500 ;
    END
  END Tile_X0Y0_FrameData_O[17]
  PIN Tile_X0Y0_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 406.780 107.520 407.180 ;
    END
  END Tile_X0Y0_FrameData_O[18]
  PIN Tile_X0Y0_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 408.460 107.520 408.860 ;
    END
  END Tile_X0Y0_FrameData_O[19]
  PIN Tile_X0Y0_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 378.220 107.520 378.620 ;
    END
  END Tile_X0Y0_FrameData_O[1]
  PIN Tile_X0Y0_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 410.140 107.520 410.540 ;
    END
  END Tile_X0Y0_FrameData_O[20]
  PIN Tile_X0Y0_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 411.820 107.520 412.220 ;
    END
  END Tile_X0Y0_FrameData_O[21]
  PIN Tile_X0Y0_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 413.500 107.520 413.900 ;
    END
  END Tile_X0Y0_FrameData_O[22]
  PIN Tile_X0Y0_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 415.180 107.520 415.580 ;
    END
  END Tile_X0Y0_FrameData_O[23]
  PIN Tile_X0Y0_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 416.860 107.520 417.260 ;
    END
  END Tile_X0Y0_FrameData_O[24]
  PIN Tile_X0Y0_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 418.540 107.520 418.940 ;
    END
  END Tile_X0Y0_FrameData_O[25]
  PIN Tile_X0Y0_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 420.220 107.520 420.620 ;
    END
  END Tile_X0Y0_FrameData_O[26]
  PIN Tile_X0Y0_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 421.900 107.520 422.300 ;
    END
  END Tile_X0Y0_FrameData_O[27]
  PIN Tile_X0Y0_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 423.580 107.520 423.980 ;
    END
  END Tile_X0Y0_FrameData_O[28]
  PIN Tile_X0Y0_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 425.260 107.520 425.660 ;
    END
  END Tile_X0Y0_FrameData_O[29]
  PIN Tile_X0Y0_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 379.900 107.520 380.300 ;
    END
  END Tile_X0Y0_FrameData_O[2]
  PIN Tile_X0Y0_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 426.940 107.520 427.340 ;
    END
  END Tile_X0Y0_FrameData_O[30]
  PIN Tile_X0Y0_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 428.620 107.520 429.020 ;
    END
  END Tile_X0Y0_FrameData_O[31]
  PIN Tile_X0Y0_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 381.580 107.520 381.980 ;
    END
  END Tile_X0Y0_FrameData_O[3]
  PIN Tile_X0Y0_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 383.260 107.520 383.660 ;
    END
  END Tile_X0Y0_FrameData_O[4]
  PIN Tile_X0Y0_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 384.940 107.520 385.340 ;
    END
  END Tile_X0Y0_FrameData_O[5]
  PIN Tile_X0Y0_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 386.620 107.520 387.020 ;
    END
  END Tile_X0Y0_FrameData_O[6]
  PIN Tile_X0Y0_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 388.300 107.520 388.700 ;
    END
  END Tile_X0Y0_FrameData_O[7]
  PIN Tile_X0Y0_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 389.980 107.520 390.380 ;
    END
  END Tile_X0Y0_FrameData_O[8]
  PIN Tile_X0Y0_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 391.660 107.520 392.060 ;
    END
  END Tile_X0Y0_FrameData_O[9]
  PIN Tile_X0Y0_FrameStrobe_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.000 429.680 79.400 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[0]
  PIN Tile_X0Y0_FrameStrobe_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 88.600 429.680 89.000 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[10]
  PIN Tile_X0Y0_FrameStrobe_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 89.560 429.680 89.960 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[11]
  PIN Tile_X0Y0_FrameStrobe_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 90.520 429.680 90.920 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[12]
  PIN Tile_X0Y0_FrameStrobe_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 91.480 429.680 91.880 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[13]
  PIN Tile_X0Y0_FrameStrobe_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 92.440 429.680 92.840 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[14]
  PIN Tile_X0Y0_FrameStrobe_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 93.400 429.680 93.800 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[15]
  PIN Tile_X0Y0_FrameStrobe_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 429.680 94.760 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[16]
  PIN Tile_X0Y0_FrameStrobe_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 95.320 429.680 95.720 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[17]
  PIN Tile_X0Y0_FrameStrobe_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 96.280 429.680 96.680 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[18]
  PIN Tile_X0Y0_FrameStrobe_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 97.240 429.680 97.640 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[19]
  PIN Tile_X0Y0_FrameStrobe_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 79.960 429.680 80.360 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[1]
  PIN Tile_X0Y0_FrameStrobe_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 429.680 81.320 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[2]
  PIN Tile_X0Y0_FrameStrobe_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 81.880 429.680 82.280 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[3]
  PIN Tile_X0Y0_FrameStrobe_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 82.840 429.680 83.240 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[4]
  PIN Tile_X0Y0_FrameStrobe_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 83.800 429.680 84.200 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[5]
  PIN Tile_X0Y0_FrameStrobe_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 84.760 429.680 85.160 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[6]
  PIN Tile_X0Y0_FrameStrobe_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 85.720 429.680 86.120 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[7]
  PIN Tile_X0Y0_FrameStrobe_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 86.680 429.680 87.080 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[8]
  PIN Tile_X0Y0_FrameStrobe_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 87.640 429.680 88.040 430.080 ;
    END
  END Tile_X0Y0_FrameStrobe_O[9]
  PIN Tile_X0Y0_N1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 8.920 429.680 9.320 430.080 ;
    END
  END Tile_X0Y0_N1BEG[0]
  PIN Tile_X0Y0_N1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 9.880 429.680 10.280 430.080 ;
    END
  END Tile_X0Y0_N1BEG[1]
  PIN Tile_X0Y0_N1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 10.840 429.680 11.240 430.080 ;
    END
  END Tile_X0Y0_N1BEG[2]
  PIN Tile_X0Y0_N1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 11.800 429.680 12.200 430.080 ;
    END
  END Tile_X0Y0_N1BEG[3]
  PIN Tile_X0Y0_N2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 12.760 429.680 13.160 430.080 ;
    END
  END Tile_X0Y0_N2BEG[0]
  PIN Tile_X0Y0_N2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 13.720 429.680 14.120 430.080 ;
    END
  END Tile_X0Y0_N2BEG[1]
  PIN Tile_X0Y0_N2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 14.680 429.680 15.080 430.080 ;
    END
  END Tile_X0Y0_N2BEG[2]
  PIN Tile_X0Y0_N2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 15.640 429.680 16.040 430.080 ;
    END
  END Tile_X0Y0_N2BEG[3]
  PIN Tile_X0Y0_N2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 16.600 429.680 17.000 430.080 ;
    END
  END Tile_X0Y0_N2BEG[4]
  PIN Tile_X0Y0_N2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 17.560 429.680 17.960 430.080 ;
    END
  END Tile_X0Y0_N2BEG[5]
  PIN Tile_X0Y0_N2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 18.520 429.680 18.920 430.080 ;
    END
  END Tile_X0Y0_N2BEG[6]
  PIN Tile_X0Y0_N2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 19.480 429.680 19.880 430.080 ;
    END
  END Tile_X0Y0_N2BEG[7]
  PIN Tile_X0Y0_N2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 429.680 20.840 430.080 ;
    END
  END Tile_X0Y0_N2BEGb[0]
  PIN Tile_X0Y0_N2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 21.400 429.680 21.800 430.080 ;
    END
  END Tile_X0Y0_N2BEGb[1]
  PIN Tile_X0Y0_N2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 22.360 429.680 22.760 430.080 ;
    END
  END Tile_X0Y0_N2BEGb[2]
  PIN Tile_X0Y0_N2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 23.320 429.680 23.720 430.080 ;
    END
  END Tile_X0Y0_N2BEGb[3]
  PIN Tile_X0Y0_N2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 24.280 429.680 24.680 430.080 ;
    END
  END Tile_X0Y0_N2BEGb[4]
  PIN Tile_X0Y0_N2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 25.240 429.680 25.640 430.080 ;
    END
  END Tile_X0Y0_N2BEGb[5]
  PIN Tile_X0Y0_N2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 26.200 429.680 26.600 430.080 ;
    END
  END Tile_X0Y0_N2BEGb[6]
  PIN Tile_X0Y0_N2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 429.680 27.560 430.080 ;
    END
  END Tile_X0Y0_N2BEGb[7]
  PIN Tile_X0Y0_N4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 28.120 429.680 28.520 430.080 ;
    END
  END Tile_X0Y0_N4BEG[0]
  PIN Tile_X0Y0_N4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 37.720 429.680 38.120 430.080 ;
    END
  END Tile_X0Y0_N4BEG[10]
  PIN Tile_X0Y0_N4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 38.680 429.680 39.080 430.080 ;
    END
  END Tile_X0Y0_N4BEG[11]
  PIN Tile_X0Y0_N4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 39.640 429.680 40.040 430.080 ;
    END
  END Tile_X0Y0_N4BEG[12]
  PIN Tile_X0Y0_N4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 429.680 41.000 430.080 ;
    END
  END Tile_X0Y0_N4BEG[13]
  PIN Tile_X0Y0_N4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 41.560 429.680 41.960 430.080 ;
    END
  END Tile_X0Y0_N4BEG[14]
  PIN Tile_X0Y0_N4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 42.520 429.680 42.920 430.080 ;
    END
  END Tile_X0Y0_N4BEG[15]
  PIN Tile_X0Y0_N4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 29.080 429.680 29.480 430.080 ;
    END
  END Tile_X0Y0_N4BEG[1]
  PIN Tile_X0Y0_N4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 30.040 429.680 30.440 430.080 ;
    END
  END Tile_X0Y0_N4BEG[2]
  PIN Tile_X0Y0_N4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.000 429.680 31.400 430.080 ;
    END
  END Tile_X0Y0_N4BEG[3]
  PIN Tile_X0Y0_N4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 31.960 429.680 32.360 430.080 ;
    END
  END Tile_X0Y0_N4BEG[4]
  PIN Tile_X0Y0_N4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 32.920 429.680 33.320 430.080 ;
    END
  END Tile_X0Y0_N4BEG[5]
  PIN Tile_X0Y0_N4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 33.880 429.680 34.280 430.080 ;
    END
  END Tile_X0Y0_N4BEG[6]
  PIN Tile_X0Y0_N4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 34.840 429.680 35.240 430.080 ;
    END
  END Tile_X0Y0_N4BEG[7]
  PIN Tile_X0Y0_N4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 35.800 429.680 36.200 430.080 ;
    END
  END Tile_X0Y0_N4BEG[8]
  PIN Tile_X0Y0_N4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 36.760 429.680 37.160 430.080 ;
    END
  END Tile_X0Y0_N4BEG[9]
  PIN Tile_X0Y0_S1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.307800 ;
    PORT
      LAYER Metal2 ;
        RECT 43.480 429.680 43.880 430.080 ;
    END
  END Tile_X0Y0_S1END[0]
  PIN Tile_X0Y0_S1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.307800 ;
    PORT
      LAYER Metal2 ;
        RECT 44.440 429.680 44.840 430.080 ;
    END
  END Tile_X0Y0_S1END[1]
  PIN Tile_X0Y0_S1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.307800 ;
    PORT
      LAYER Metal2 ;
        RECT 45.400 429.680 45.800 430.080 ;
    END
  END Tile_X0Y0_S1END[2]
  PIN Tile_X0Y0_S1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.307800 ;
    PORT
      LAYER Metal2 ;
        RECT 46.360 429.680 46.760 430.080 ;
    END
  END Tile_X0Y0_S1END[3]
  PIN Tile_X0Y0_S2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 55.000 429.680 55.400 430.080 ;
    END
  END Tile_X0Y0_S2END[0]
  PIN Tile_X0Y0_S2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 55.960 429.680 56.360 430.080 ;
    END
  END Tile_X0Y0_S2END[1]
  PIN Tile_X0Y0_S2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 56.920 429.680 57.320 430.080 ;
    END
  END Tile_X0Y0_S2END[2]
  PIN Tile_X0Y0_S2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 57.880 429.680 58.280 430.080 ;
    END
  END Tile_X0Y0_S2END[3]
  PIN Tile_X0Y0_S2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 58.840 429.680 59.240 430.080 ;
    END
  END Tile_X0Y0_S2END[4]
  PIN Tile_X0Y0_S2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 59.800 429.680 60.200 430.080 ;
    END
  END Tile_X0Y0_S2END[5]
  PIN Tile_X0Y0_S2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 429.680 61.160 430.080 ;
    END
  END Tile_X0Y0_S2END[6]
  PIN Tile_X0Y0_S2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 61.720 429.680 62.120 430.080 ;
    END
  END Tile_X0Y0_S2END[7]
  PIN Tile_X0Y0_S2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.455000 ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 429.680 47.720 430.080 ;
    END
  END Tile_X0Y0_S2MID[0]
  PIN Tile_X0Y0_S2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.455000 ;
    PORT
      LAYER Metal2 ;
        RECT 48.280 429.680 48.680 430.080 ;
    END
  END Tile_X0Y0_S2MID[1]
  PIN Tile_X0Y0_S2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.877500 ;
    PORT
      LAYER Metal2 ;
        RECT 49.240 429.680 49.640 430.080 ;
    END
  END Tile_X0Y0_S2MID[2]
  PIN Tile_X0Y0_S2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 10.657400 ;
    ANTENNADIFFAREA 32.246399 ;
    PORT
      LAYER Metal2 ;
        RECT 50.200 429.680 50.600 430.080 ;
    END
  END Tile_X0Y0_S2MID[3]
  PIN Tile_X0Y0_S2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 51.160 429.680 51.560 430.080 ;
    END
  END Tile_X0Y0_S2MID[4]
  PIN Tile_X0Y0_S2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 52.120 429.680 52.520 430.080 ;
    END
  END Tile_X0Y0_S2MID[5]
  PIN Tile_X0Y0_S2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 53.080 429.680 53.480 430.080 ;
    END
  END Tile_X0Y0_S2MID[6]
  PIN Tile_X0Y0_S2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal2 ;
        RECT 54.040 429.680 54.440 430.080 ;
    END
  END Tile_X0Y0_S2MID[7]
  PIN Tile_X0Y0_S4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 62.680 429.680 63.080 430.080 ;
    END
  END Tile_X0Y0_S4END[0]
  PIN Tile_X0Y0_S4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 72.280 429.680 72.680 430.080 ;
    END
  END Tile_X0Y0_S4END[10]
  PIN Tile_X0Y0_S4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 73.240 429.680 73.640 430.080 ;
    END
  END Tile_X0Y0_S4END[11]
  PIN Tile_X0Y0_S4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 74.200 429.680 74.600 430.080 ;
    END
  END Tile_X0Y0_S4END[12]
  PIN Tile_X0Y0_S4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 75.160 429.680 75.560 430.080 ;
    END
  END Tile_X0Y0_S4END[13]
  PIN Tile_X0Y0_S4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 76.120 429.680 76.520 430.080 ;
    END
  END Tile_X0Y0_S4END[14]
  PIN Tile_X0Y0_S4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 77.080 429.680 77.480 430.080 ;
    END
  END Tile_X0Y0_S4END[15]
  PIN Tile_X0Y0_S4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 63.640 429.680 64.040 430.080 ;
    END
  END Tile_X0Y0_S4END[1]
  PIN Tile_X0Y0_S4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 64.600 429.680 65.000 430.080 ;
    END
  END Tile_X0Y0_S4END[2]
  PIN Tile_X0Y0_S4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 65.560 429.680 65.960 430.080 ;
    END
  END Tile_X0Y0_S4END[3]
  PIN Tile_X0Y0_S4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 66.520 429.680 66.920 430.080 ;
    END
  END Tile_X0Y0_S4END[4]
  PIN Tile_X0Y0_S4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 67.480 429.680 67.880 430.080 ;
    END
  END Tile_X0Y0_S4END[5]
  PIN Tile_X0Y0_S4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.440 429.680 68.840 430.080 ;
    END
  END Tile_X0Y0_S4END[6]
  PIN Tile_X0Y0_S4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 429.680 69.800 430.080 ;
    END
  END Tile_X0Y0_S4END[7]
  PIN Tile_X0Y0_S4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.789100 ;
    ANTENNADIFFAREA 2.015400 ;
    PORT
      LAYER Metal2 ;
        RECT 70.360 429.680 70.760 430.080 ;
    END
  END Tile_X0Y0_S4END[8]
  PIN Tile_X0Y0_S4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 71.320 429.680 71.720 430.080 ;
    END
  END Tile_X0Y0_S4END[9]
  PIN Tile_X0Y0_UserCLKo
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 78.040 429.680 78.440 430.080 ;
    END
  END Tile_X0Y0_UserCLKo
  PIN Tile_X0Y0_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 215.260 107.520 215.660 ;
    END
  END Tile_X0Y0_W1END[0]
  PIN Tile_X0Y0_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 216.940 107.520 217.340 ;
    END
  END Tile_X0Y0_W1END[1]
  PIN Tile_X0Y0_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 218.620 107.520 219.020 ;
    END
  END Tile_X0Y0_W1END[2]
  PIN Tile_X0Y0_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 220.300 107.520 220.700 ;
    END
  END Tile_X0Y0_W1END[3]
  PIN Tile_X0Y0_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 235.420 107.520 235.820 ;
    END
  END Tile_X0Y0_W2END[0]
  PIN Tile_X0Y0_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 237.100 107.520 237.500 ;
    END
  END Tile_X0Y0_W2END[1]
  PIN Tile_X0Y0_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 238.780 107.520 239.180 ;
    END
  END Tile_X0Y0_W2END[2]
  PIN Tile_X0Y0_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 240.460 107.520 240.860 ;
    END
  END Tile_X0Y0_W2END[3]
  PIN Tile_X0Y0_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 242.140 107.520 242.540 ;
    END
  END Tile_X0Y0_W2END[4]
  PIN Tile_X0Y0_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 243.820 107.520 244.220 ;
    END
  END Tile_X0Y0_W2END[5]
  PIN Tile_X0Y0_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 245.500 107.520 245.900 ;
    END
  END Tile_X0Y0_W2END[6]
  PIN Tile_X0Y0_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 247.180 107.520 247.580 ;
    END
  END Tile_X0Y0_W2END[7]
  PIN Tile_X0Y0_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 221.980 107.520 222.380 ;
    END
  END Tile_X0Y0_W2MID[0]
  PIN Tile_X0Y0_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 223.660 107.520 224.060 ;
    END
  END Tile_X0Y0_W2MID[1]
  PIN Tile_X0Y0_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 225.340 107.520 225.740 ;
    END
  END Tile_X0Y0_W2MID[2]
  PIN Tile_X0Y0_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 227.020 107.520 227.420 ;
    END
  END Tile_X0Y0_W2MID[3]
  PIN Tile_X0Y0_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 228.700 107.520 229.100 ;
    END
  END Tile_X0Y0_W2MID[4]
  PIN Tile_X0Y0_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 230.380 107.520 230.780 ;
    END
  END Tile_X0Y0_W2MID[5]
  PIN Tile_X0Y0_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 232.060 107.520 232.460 ;
    END
  END Tile_X0Y0_W2MID[6]
  PIN Tile_X0Y0_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 233.740 107.520 234.140 ;
    END
  END Tile_X0Y0_W2MID[7]
  PIN Tile_X0Y0_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.734000 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 275.740 107.520 276.140 ;
    END
  END Tile_X0Y0_W6END[0]
  PIN Tile_X0Y0_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.947200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 292.540 107.520 292.940 ;
    END
  END Tile_X0Y0_W6END[10]
  PIN Tile_X0Y0_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.947200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 294.220 107.520 294.620 ;
    END
  END Tile_X0Y0_W6END[11]
  PIN Tile_X0Y0_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.734000 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 277.420 107.520 277.820 ;
    END
  END Tile_X0Y0_W6END[1]
  PIN Tile_X0Y0_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.734000 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 279.100 107.520 279.500 ;
    END
  END Tile_X0Y0_W6END[2]
  PIN Tile_X0Y0_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.734000 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 280.780 107.520 281.180 ;
    END
  END Tile_X0Y0_W6END[3]
  PIN Tile_X0Y0_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.947200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 282.460 107.520 282.860 ;
    END
  END Tile_X0Y0_W6END[4]
  PIN Tile_X0Y0_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.947200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 284.140 107.520 284.540 ;
    END
  END Tile_X0Y0_W6END[5]
  PIN Tile_X0Y0_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.947200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 285.820 107.520 286.220 ;
    END
  END Tile_X0Y0_W6END[6]
  PIN Tile_X0Y0_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.947200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 287.500 107.520 287.900 ;
    END
  END Tile_X0Y0_W6END[7]
  PIN Tile_X0Y0_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.947200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 289.180 107.520 289.580 ;
    END
  END Tile_X0Y0_W6END[8]
  PIN Tile_X0Y0_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.947200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 290.860 107.520 291.260 ;
    END
  END Tile_X0Y0_W6END[9]
  PIN Tile_X0Y0_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 248.860 107.520 249.260 ;
    END
  END Tile_X0Y0_WW4END[0]
  PIN Tile_X0Y0_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 265.660 107.520 266.060 ;
    END
  END Tile_X0Y0_WW4END[10]
  PIN Tile_X0Y0_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 267.340 107.520 267.740 ;
    END
  END Tile_X0Y0_WW4END[11]
  PIN Tile_X0Y0_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 269.020 107.520 269.420 ;
    END
  END Tile_X0Y0_WW4END[12]
  PIN Tile_X0Y0_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 270.700 107.520 271.100 ;
    END
  END Tile_X0Y0_WW4END[13]
  PIN Tile_X0Y0_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 272.380 107.520 272.780 ;
    END
  END Tile_X0Y0_WW4END[14]
  PIN Tile_X0Y0_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.492200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 274.060 107.520 274.460 ;
    END
  END Tile_X0Y0_WW4END[15]
  PIN Tile_X0Y0_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 250.540 107.520 250.940 ;
    END
  END Tile_X0Y0_WW4END[1]
  PIN Tile_X0Y0_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 252.220 107.520 252.620 ;
    END
  END Tile_X0Y0_WW4END[2]
  PIN Tile_X0Y0_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 253.900 107.520 254.300 ;
    END
  END Tile_X0Y0_WW4END[3]
  PIN Tile_X0Y0_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 255.580 107.520 255.980 ;
    END
  END Tile_X0Y0_WW4END[4]
  PIN Tile_X0Y0_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 257.260 107.520 257.660 ;
    END
  END Tile_X0Y0_WW4END[5]
  PIN Tile_X0Y0_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 258.940 107.520 259.340 ;
    END
  END Tile_X0Y0_WW4END[6]
  PIN Tile_X0Y0_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 260.620 107.520 261.020 ;
    END
  END Tile_X0Y0_WW4END[7]
  PIN Tile_X0Y0_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 262.300 107.520 262.700 ;
    END
  END Tile_X0Y0_WW4END[8]
  PIN Tile_X0Y0_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 263.980 107.520 264.380 ;
    END
  END Tile_X0Y0_WW4END[9]
  PIN Tile_X0Y1_E1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 80.860 107.520 81.260 ;
    END
  END Tile_X0Y1_E1BEG[0]
  PIN Tile_X0Y1_E1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 82.540 107.520 82.940 ;
    END
  END Tile_X0Y1_E1BEG[1]
  PIN Tile_X0Y1_E1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 84.220 107.520 84.620 ;
    END
  END Tile_X0Y1_E1BEG[2]
  PIN Tile_X0Y1_E1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 85.900 107.520 86.300 ;
    END
  END Tile_X0Y1_E1BEG[3]
  PIN Tile_X0Y1_E2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 87.580 107.520 87.980 ;
    END
  END Tile_X0Y1_E2BEG[0]
  PIN Tile_X0Y1_E2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 89.260 107.520 89.660 ;
    END
  END Tile_X0Y1_E2BEG[1]
  PIN Tile_X0Y1_E2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 90.940 107.520 91.340 ;
    END
  END Tile_X0Y1_E2BEG[2]
  PIN Tile_X0Y1_E2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 92.620 107.520 93.020 ;
    END
  END Tile_X0Y1_E2BEG[3]
  PIN Tile_X0Y1_E2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 94.300 107.520 94.700 ;
    END
  END Tile_X0Y1_E2BEG[4]
  PIN Tile_X0Y1_E2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 95.980 107.520 96.380 ;
    END
  END Tile_X0Y1_E2BEG[5]
  PIN Tile_X0Y1_E2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 97.660 107.520 98.060 ;
    END
  END Tile_X0Y1_E2BEG[6]
  PIN Tile_X0Y1_E2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 99.340 107.520 99.740 ;
    END
  END Tile_X0Y1_E2BEG[7]
  PIN Tile_X0Y1_E2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 101.020 107.520 101.420 ;
    END
  END Tile_X0Y1_E2BEGb[0]
  PIN Tile_X0Y1_E2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 102.700 107.520 103.100 ;
    END
  END Tile_X0Y1_E2BEGb[1]
  PIN Tile_X0Y1_E2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 104.380 107.520 104.780 ;
    END
  END Tile_X0Y1_E2BEGb[2]
  PIN Tile_X0Y1_E2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 106.060 107.520 106.460 ;
    END
  END Tile_X0Y1_E2BEGb[3]
  PIN Tile_X0Y1_E2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 107.740 107.520 108.140 ;
    END
  END Tile_X0Y1_E2BEGb[4]
  PIN Tile_X0Y1_E2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 109.420 107.520 109.820 ;
    END
  END Tile_X0Y1_E2BEGb[5]
  PIN Tile_X0Y1_E2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 111.100 107.520 111.500 ;
    END
  END Tile_X0Y1_E2BEGb[6]
  PIN Tile_X0Y1_E2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 112.780 107.520 113.180 ;
    END
  END Tile_X0Y1_E2BEGb[7]
  PIN Tile_X0Y1_E6BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 141.340 107.520 141.740 ;
    END
  END Tile_X0Y1_E6BEG[0]
  PIN Tile_X0Y1_E6BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 158.140 107.520 158.540 ;
    END
  END Tile_X0Y1_E6BEG[10]
  PIN Tile_X0Y1_E6BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 159.820 107.520 160.220 ;
    END
  END Tile_X0Y1_E6BEG[11]
  PIN Tile_X0Y1_E6BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 143.020 107.520 143.420 ;
    END
  END Tile_X0Y1_E6BEG[1]
  PIN Tile_X0Y1_E6BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 144.700 107.520 145.100 ;
    END
  END Tile_X0Y1_E6BEG[2]
  PIN Tile_X0Y1_E6BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 146.380 107.520 146.780 ;
    END
  END Tile_X0Y1_E6BEG[3]
  PIN Tile_X0Y1_E6BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 148.060 107.520 148.460 ;
    END
  END Tile_X0Y1_E6BEG[4]
  PIN Tile_X0Y1_E6BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 149.740 107.520 150.140 ;
    END
  END Tile_X0Y1_E6BEG[5]
  PIN Tile_X0Y1_E6BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 151.420 107.520 151.820 ;
    END
  END Tile_X0Y1_E6BEG[6]
  PIN Tile_X0Y1_E6BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 153.100 107.520 153.500 ;
    END
  END Tile_X0Y1_E6BEG[7]
  PIN Tile_X0Y1_E6BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 154.780 107.520 155.180 ;
    END
  END Tile_X0Y1_E6BEG[8]
  PIN Tile_X0Y1_E6BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 156.460 107.520 156.860 ;
    END
  END Tile_X0Y1_E6BEG[9]
  PIN Tile_X0Y1_EE4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 114.460 107.520 114.860 ;
    END
  END Tile_X0Y1_EE4BEG[0]
  PIN Tile_X0Y1_EE4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 131.260 107.520 131.660 ;
    END
  END Tile_X0Y1_EE4BEG[10]
  PIN Tile_X0Y1_EE4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 132.940 107.520 133.340 ;
    END
  END Tile_X0Y1_EE4BEG[11]
  PIN Tile_X0Y1_EE4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 134.620 107.520 135.020 ;
    END
  END Tile_X0Y1_EE4BEG[12]
  PIN Tile_X0Y1_EE4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 136.300 107.520 136.700 ;
    END
  END Tile_X0Y1_EE4BEG[13]
  PIN Tile_X0Y1_EE4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 137.980 107.520 138.380 ;
    END
  END Tile_X0Y1_EE4BEG[14]
  PIN Tile_X0Y1_EE4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 139.660 107.520 140.060 ;
    END
  END Tile_X0Y1_EE4BEG[15]
  PIN Tile_X0Y1_EE4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 116.140 107.520 116.540 ;
    END
  END Tile_X0Y1_EE4BEG[1]
  PIN Tile_X0Y1_EE4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 117.820 107.520 118.220 ;
    END
  END Tile_X0Y1_EE4BEG[2]
  PIN Tile_X0Y1_EE4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 119.500 107.520 119.900 ;
    END
  END Tile_X0Y1_EE4BEG[3]
  PIN Tile_X0Y1_EE4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 121.180 107.520 121.580 ;
    END
  END Tile_X0Y1_EE4BEG[4]
  PIN Tile_X0Y1_EE4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 122.860 107.520 123.260 ;
    END
  END Tile_X0Y1_EE4BEG[5]
  PIN Tile_X0Y1_EE4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 124.540 107.520 124.940 ;
    END
  END Tile_X0Y1_EE4BEG[6]
  PIN Tile_X0Y1_EE4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 126.220 107.520 126.620 ;
    END
  END Tile_X0Y1_EE4BEG[7]
  PIN Tile_X0Y1_EE4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 127.900 107.520 128.300 ;
    END
  END Tile_X0Y1_EE4BEG[8]
  PIN Tile_X0Y1_EE4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 129.580 107.520 129.980 ;
    END
  END Tile_X0Y1_EE4BEG[9]
  PIN Tile_X0Y1_FrameData[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 288.340 0.400 288.740 ;
    END
  END Tile_X0Y1_FrameData[0]
  PIN Tile_X0Y1_FrameData[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 321.940 0.400 322.340 ;
    END
  END Tile_X0Y1_FrameData[10]
  PIN Tile_X0Y1_FrameData[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 325.300 0.400 325.700 ;
    END
  END Tile_X0Y1_FrameData[11]
  PIN Tile_X0Y1_FrameData[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 328.660 0.400 329.060 ;
    END
  END Tile_X0Y1_FrameData[12]
  PIN Tile_X0Y1_FrameData[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 332.020 0.400 332.420 ;
    END
  END Tile_X0Y1_FrameData[13]
  PIN Tile_X0Y1_FrameData[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 335.380 0.400 335.780 ;
    END
  END Tile_X0Y1_FrameData[14]
  PIN Tile_X0Y1_FrameData[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 338.740 0.400 339.140 ;
    END
  END Tile_X0Y1_FrameData[15]
  PIN Tile_X0Y1_FrameData[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.100 0.400 342.500 ;
    END
  END Tile_X0Y1_FrameData[16]
  PIN Tile_X0Y1_FrameData[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 345.460 0.400 345.860 ;
    END
  END Tile_X0Y1_FrameData[17]
  PIN Tile_X0Y1_FrameData[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 348.820 0.400 349.220 ;
    END
  END Tile_X0Y1_FrameData[18]
  PIN Tile_X0Y1_FrameData[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 352.180 0.400 352.580 ;
    END
  END Tile_X0Y1_FrameData[19]
  PIN Tile_X0Y1_FrameData[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 291.700 0.400 292.100 ;
    END
  END Tile_X0Y1_FrameData[1]
  PIN Tile_X0Y1_FrameData[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 355.540 0.400 355.940 ;
    END
  END Tile_X0Y1_FrameData[20]
  PIN Tile_X0Y1_FrameData[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 358.900 0.400 359.300 ;
    END
  END Tile_X0Y1_FrameData[21]
  PIN Tile_X0Y1_FrameData[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 362.260 0.400 362.660 ;
    END
  END Tile_X0Y1_FrameData[22]
  PIN Tile_X0Y1_FrameData[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 50.906700 ;
    ANTENNADIFFAREA 163.247391 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 365.620 0.400 366.020 ;
    END
  END Tile_X0Y1_FrameData[23]
  PIN Tile_X0Y1_FrameData[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 368.980 0.400 369.380 ;
    END
  END Tile_X0Y1_FrameData[24]
  PIN Tile_X0Y1_FrameData[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 372.340 0.400 372.740 ;
    END
  END Tile_X0Y1_FrameData[25]
  PIN Tile_X0Y1_FrameData[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 375.700 0.400 376.100 ;
    END
  END Tile_X0Y1_FrameData[26]
  PIN Tile_X0Y1_FrameData[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 379.060 0.400 379.460 ;
    END
  END Tile_X0Y1_FrameData[27]
  PIN Tile_X0Y1_FrameData[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 382.420 0.400 382.820 ;
    END
  END Tile_X0Y1_FrameData[28]
  PIN Tile_X0Y1_FrameData[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 385.780 0.400 386.180 ;
    END
  END Tile_X0Y1_FrameData[29]
  PIN Tile_X0Y1_FrameData[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 295.060 0.400 295.460 ;
    END
  END Tile_X0Y1_FrameData[2]
  PIN Tile_X0Y1_FrameData[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 389.140 0.400 389.540 ;
    END
  END Tile_X0Y1_FrameData[30]
  PIN Tile_X0Y1_FrameData[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.101900 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 392.500 0.400 392.900 ;
    END
  END Tile_X0Y1_FrameData[31]
  PIN Tile_X0Y1_FrameData[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 298.420 0.400 298.820 ;
    END
  END Tile_X0Y1_FrameData[3]
  PIN Tile_X0Y1_FrameData[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 301.780 0.400 302.180 ;
    END
  END Tile_X0Y1_FrameData[4]
  PIN Tile_X0Y1_FrameData[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 305.140 0.400 305.540 ;
    END
  END Tile_X0Y1_FrameData[5]
  PIN Tile_X0Y1_FrameData[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 308.500 0.400 308.900 ;
    END
  END Tile_X0Y1_FrameData[6]
  PIN Tile_X0Y1_FrameData[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 311.860 0.400 312.260 ;
    END
  END Tile_X0Y1_FrameData[7]
  PIN Tile_X0Y1_FrameData[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 7.101900 ;
    ANTENNADIFFAREA 18.138599 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 315.220 0.400 315.620 ;
    END
  END Tile_X0Y1_FrameData[8]
  PIN Tile_X0Y1_FrameData[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.626300 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.580 0.400 318.980 ;
    END
  END Tile_X0Y1_FrameData[9]
  PIN Tile_X0Y1_FrameData_O[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 161.500 107.520 161.900 ;
    END
  END Tile_X0Y1_FrameData_O[0]
  PIN Tile_X0Y1_FrameData_O[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 178.300 107.520 178.700 ;
    END
  END Tile_X0Y1_FrameData_O[10]
  PIN Tile_X0Y1_FrameData_O[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 179.980 107.520 180.380 ;
    END
  END Tile_X0Y1_FrameData_O[11]
  PIN Tile_X0Y1_FrameData_O[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 181.660 107.520 182.060 ;
    END
  END Tile_X0Y1_FrameData_O[12]
  PIN Tile_X0Y1_FrameData_O[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 183.340 107.520 183.740 ;
    END
  END Tile_X0Y1_FrameData_O[13]
  PIN Tile_X0Y1_FrameData_O[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 185.020 107.520 185.420 ;
    END
  END Tile_X0Y1_FrameData_O[14]
  PIN Tile_X0Y1_FrameData_O[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 186.700 107.520 187.100 ;
    END
  END Tile_X0Y1_FrameData_O[15]
  PIN Tile_X0Y1_FrameData_O[16]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 188.380 107.520 188.780 ;
    END
  END Tile_X0Y1_FrameData_O[16]
  PIN Tile_X0Y1_FrameData_O[17]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 190.060 107.520 190.460 ;
    END
  END Tile_X0Y1_FrameData_O[17]
  PIN Tile_X0Y1_FrameData_O[18]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 191.740 107.520 192.140 ;
    END
  END Tile_X0Y1_FrameData_O[18]
  PIN Tile_X0Y1_FrameData_O[19]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 193.420 107.520 193.820 ;
    END
  END Tile_X0Y1_FrameData_O[19]
  PIN Tile_X0Y1_FrameData_O[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 163.180 107.520 163.580 ;
    END
  END Tile_X0Y1_FrameData_O[1]
  PIN Tile_X0Y1_FrameData_O[20]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 195.100 107.520 195.500 ;
    END
  END Tile_X0Y1_FrameData_O[20]
  PIN Tile_X0Y1_FrameData_O[21]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 196.780 107.520 197.180 ;
    END
  END Tile_X0Y1_FrameData_O[21]
  PIN Tile_X0Y1_FrameData_O[22]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 198.460 107.520 198.860 ;
    END
  END Tile_X0Y1_FrameData_O[22]
  PIN Tile_X0Y1_FrameData_O[23]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 200.140 107.520 200.540 ;
    END
  END Tile_X0Y1_FrameData_O[23]
  PIN Tile_X0Y1_FrameData_O[24]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 201.820 107.520 202.220 ;
    END
  END Tile_X0Y1_FrameData_O[24]
  PIN Tile_X0Y1_FrameData_O[25]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 203.500 107.520 203.900 ;
    END
  END Tile_X0Y1_FrameData_O[25]
  PIN Tile_X0Y1_FrameData_O[26]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 205.180 107.520 205.580 ;
    END
  END Tile_X0Y1_FrameData_O[26]
  PIN Tile_X0Y1_FrameData_O[27]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 206.860 107.520 207.260 ;
    END
  END Tile_X0Y1_FrameData_O[27]
  PIN Tile_X0Y1_FrameData_O[28]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 208.540 107.520 208.940 ;
    END
  END Tile_X0Y1_FrameData_O[28]
  PIN Tile_X0Y1_FrameData_O[29]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 210.220 107.520 210.620 ;
    END
  END Tile_X0Y1_FrameData_O[29]
  PIN Tile_X0Y1_FrameData_O[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 164.860 107.520 165.260 ;
    END
  END Tile_X0Y1_FrameData_O[2]
  PIN Tile_X0Y1_FrameData_O[30]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 211.900 107.520 212.300 ;
    END
  END Tile_X0Y1_FrameData_O[30]
  PIN Tile_X0Y1_FrameData_O[31]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 213.580 107.520 213.980 ;
    END
  END Tile_X0Y1_FrameData_O[31]
  PIN Tile_X0Y1_FrameData_O[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 166.540 107.520 166.940 ;
    END
  END Tile_X0Y1_FrameData_O[3]
  PIN Tile_X0Y1_FrameData_O[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 168.220 107.520 168.620 ;
    END
  END Tile_X0Y1_FrameData_O[4]
  PIN Tile_X0Y1_FrameData_O[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 169.900 107.520 170.300 ;
    END
  END Tile_X0Y1_FrameData_O[5]
  PIN Tile_X0Y1_FrameData_O[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 171.580 107.520 171.980 ;
    END
  END Tile_X0Y1_FrameData_O[6]
  PIN Tile_X0Y1_FrameData_O[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 173.260 107.520 173.660 ;
    END
  END Tile_X0Y1_FrameData_O[7]
  PIN Tile_X0Y1_FrameData_O[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 174.940 107.520 175.340 ;
    END
  END Tile_X0Y1_FrameData_O[8]
  PIN Tile_X0Y1_FrameData_O[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 176.620 107.520 177.020 ;
    END
  END Tile_X0Y1_FrameData_O[9]
  PIN Tile_X0Y1_FrameStrobe[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.326300 ;
    PORT
      LAYER Metal2 ;
        RECT 79.000 0.000 79.400 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[0]
  PIN Tile_X0Y1_FrameStrobe[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 88.600 0.000 89.000 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[10]
  PIN Tile_X0Y1_FrameStrobe[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 89.560 0.000 89.960 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[11]
  PIN Tile_X0Y1_FrameStrobe[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 90.520 0.000 90.920 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[12]
  PIN Tile_X0Y1_FrameStrobe[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 91.480 0.000 91.880 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[13]
  PIN Tile_X0Y1_FrameStrobe[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 92.440 0.000 92.840 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[14]
  PIN Tile_X0Y1_FrameStrobe[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 93.400 0.000 93.800 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[15]
  PIN Tile_X0Y1_FrameStrobe[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 94.360 0.000 94.760 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[16]
  PIN Tile_X0Y1_FrameStrobe[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 95.320 0.000 95.720 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[17]
  PIN Tile_X0Y1_FrameStrobe[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 96.280 0.000 96.680 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[18]
  PIN Tile_X0Y1_FrameStrobe[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 97.240 0.000 97.640 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[19]
  PIN Tile_X0Y1_FrameStrobe[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.326300 ;
    PORT
      LAYER Metal2 ;
        RECT 79.960 0.000 80.360 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[1]
  PIN Tile_X0Y1_FrameStrobe[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.326300 ;
    PORT
      LAYER Metal2 ;
        RECT 80.920 0.000 81.320 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[2]
  PIN Tile_X0Y1_FrameStrobe[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.326300 ;
    PORT
      LAYER Metal2 ;
        RECT 81.880 0.000 82.280 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[3]
  PIN Tile_X0Y1_FrameStrobe[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.326300 ;
    PORT
      LAYER Metal2 ;
        RECT 82.840 0.000 83.240 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[4]
  PIN Tile_X0Y1_FrameStrobe[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.326300 ;
    PORT
      LAYER Metal2 ;
        RECT 83.800 0.000 84.200 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[5]
  PIN Tile_X0Y1_FrameStrobe[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 13.326300 ;
    PORT
      LAYER Metal2 ;
        RECT 84.760 0.000 85.160 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[6]
  PIN Tile_X0Y1_FrameStrobe[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 11.683100 ;
    PORT
      LAYER Metal2 ;
        RECT 85.720 0.000 86.120 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[7]
  PIN Tile_X0Y1_FrameStrobe[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 86.680 0.000 87.080 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[8]
  PIN Tile_X0Y1_FrameStrobe[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 87.640 0.000 88.040 0.400 ;
    END
  END Tile_X0Y1_FrameStrobe[9]
  PIN Tile_X0Y1_N1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.311700 ;
    PORT
      LAYER Metal2 ;
        RECT 8.920 0.000 9.320 0.400 ;
    END
  END Tile_X0Y1_N1END[0]
  PIN Tile_X0Y1_N1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.311700 ;
    PORT
      LAYER Metal2 ;
        RECT 9.880 0.000 10.280 0.400 ;
    END
  END Tile_X0Y1_N1END[1]
  PIN Tile_X0Y1_N1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.311700 ;
    PORT
      LAYER Metal2 ;
        RECT 10.840 0.000 11.240 0.400 ;
    END
  END Tile_X0Y1_N1END[2]
  PIN Tile_X0Y1_N1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.311700 ;
    PORT
      LAYER Metal2 ;
        RECT 11.800 0.000 12.200 0.400 ;
    END
  END Tile_X0Y1_N1END[3]
  PIN Tile_X0Y1_N2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.226200 ;
    PORT
      LAYER Metal2 ;
        RECT 20.440 0.000 20.840 0.400 ;
    END
  END Tile_X0Y1_N2END[0]
  PIN Tile_X0Y1_N2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.226200 ;
    PORT
      LAYER Metal2 ;
        RECT 21.400 0.000 21.800 0.400 ;
    END
  END Tile_X0Y1_N2END[1]
  PIN Tile_X0Y1_N2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.678600 ;
    PORT
      LAYER Metal2 ;
        RECT 22.360 0.000 22.760 0.400 ;
    END
  END Tile_X0Y1_N2END[2]
  PIN Tile_X0Y1_N2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.620100 ;
    PORT
      LAYER Metal2 ;
        RECT 23.320 0.000 23.720 0.400 ;
    END
  END Tile_X0Y1_N2END[3]
  PIN Tile_X0Y1_N2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 24.280 0.000 24.680 0.400 ;
    END
  END Tile_X0Y1_N2END[4]
  PIN Tile_X0Y1_N2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 25.240 0.000 25.640 0.400 ;
    END
  END Tile_X0Y1_N2END[5]
  PIN Tile_X0Y1_N2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 26.200 0.000 26.600 0.400 ;
    END
  END Tile_X0Y1_N2END[6]
  PIN Tile_X0Y1_N2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal2 ;
        RECT 27.160 0.000 27.560 0.400 ;
    END
  END Tile_X0Y1_N2END[7]
  PIN Tile_X0Y1_N2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.439400 ;
    PORT
      LAYER Metal2 ;
        RECT 12.760 0.000 13.160 0.400 ;
    END
  END Tile_X0Y1_N2MID[0]
  PIN Tile_X0Y1_N2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.439400 ;
    PORT
      LAYER Metal2 ;
        RECT 13.720 0.000 14.120 0.400 ;
    END
  END Tile_X0Y1_N2MID[1]
  PIN Tile_X0Y1_N2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.439400 ;
    PORT
      LAYER Metal2 ;
        RECT 14.680 0.000 15.080 0.400 ;
    END
  END Tile_X0Y1_N2MID[2]
  PIN Tile_X0Y1_N2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.439400 ;
    PORT
      LAYER Metal2 ;
        RECT 15.640 0.000 16.040 0.400 ;
    END
  END Tile_X0Y1_N2MID[3]
  PIN Tile_X0Y1_N2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.643200 ;
    ANTENNADIFFAREA 4.030800 ;
    PORT
      LAYER Metal2 ;
        RECT 16.600 0.000 17.000 0.400 ;
    END
  END Tile_X0Y1_N2MID[4]
  PIN Tile_X0Y1_N2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.643200 ;
    ANTENNADIFFAREA 4.030800 ;
    PORT
      LAYER Metal2 ;
        RECT 17.560 0.000 17.960 0.400 ;
    END
  END Tile_X0Y1_N2MID[5]
  PIN Tile_X0Y1_N2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.878800 ;
    PORT
      LAYER Metal2 ;
        RECT 18.520 0.000 18.920 0.400 ;
    END
  END Tile_X0Y1_N2MID[6]
  PIN Tile_X0Y1_N2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.860000 ;
    ANTENNADIFFAREA 8.061600 ;
    PORT
      LAYER Metal2 ;
        RECT 19.480 0.000 19.880 0.400 ;
    END
  END Tile_X0Y1_N2MID[7]
  PIN Tile_X0Y1_N4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 28.120 0.000 28.520 0.400 ;
    END
  END Tile_X0Y1_N4END[0]
  PIN Tile_X0Y1_N4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 37.720 0.000 38.120 0.400 ;
    END
  END Tile_X0Y1_N4END[10]
  PIN Tile_X0Y1_N4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 38.680 0.000 39.080 0.400 ;
    END
  END Tile_X0Y1_N4END[11]
  PIN Tile_X0Y1_N4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 39.640 0.000 40.040 0.400 ;
    END
  END Tile_X0Y1_N4END[12]
  PIN Tile_X0Y1_N4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 40.600 0.000 41.000 0.400 ;
    END
  END Tile_X0Y1_N4END[13]
  PIN Tile_X0Y1_N4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 41.560 0.000 41.960 0.400 ;
    END
  END Tile_X0Y1_N4END[14]
  PIN Tile_X0Y1_N4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 42.520 0.000 42.920 0.400 ;
    END
  END Tile_X0Y1_N4END[15]
  PIN Tile_X0Y1_N4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 29.080 0.000 29.480 0.400 ;
    END
  END Tile_X0Y1_N4END[1]
  PIN Tile_X0Y1_N4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 30.040 0.000 30.440 0.400 ;
    END
  END Tile_X0Y1_N4END[2]
  PIN Tile_X0Y1_N4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.000 0.000 31.400 0.400 ;
    END
  END Tile_X0Y1_N4END[3]
  PIN Tile_X0Y1_N4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 31.960 0.000 32.360 0.400 ;
    END
  END Tile_X0Y1_N4END[4]
  PIN Tile_X0Y1_N4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 32.920 0.000 33.320 0.400 ;
    END
  END Tile_X0Y1_N4END[5]
  PIN Tile_X0Y1_N4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 33.880 0.000 34.280 0.400 ;
    END
  END Tile_X0Y1_N4END[6]
  PIN Tile_X0Y1_N4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal2 ;
        RECT 34.840 0.000 35.240 0.400 ;
    END
  END Tile_X0Y1_N4END[7]
  PIN Tile_X0Y1_N4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 35.800 0.000 36.200 0.400 ;
    END
  END Tile_X0Y1_N4END[8]
  PIN Tile_X0Y1_N4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.180700 ;
    PORT
      LAYER Metal2 ;
        RECT 36.760 0.000 37.160 0.400 ;
    END
  END Tile_X0Y1_N4END[9]
  PIN Tile_X0Y1_S1BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 43.480 0.000 43.880 0.400 ;
    END
  END Tile_X0Y1_S1BEG[0]
  PIN Tile_X0Y1_S1BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 44.440 0.000 44.840 0.400 ;
    END
  END Tile_X0Y1_S1BEG[1]
  PIN Tile_X0Y1_S1BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 45.400 0.000 45.800 0.400 ;
    END
  END Tile_X0Y1_S1BEG[2]
  PIN Tile_X0Y1_S1BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 46.360 0.000 46.760 0.400 ;
    END
  END Tile_X0Y1_S1BEG[3]
  PIN Tile_X0Y1_S2BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 47.320 0.000 47.720 0.400 ;
    END
  END Tile_X0Y1_S2BEG[0]
  PIN Tile_X0Y1_S2BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 48.280 0.000 48.680 0.400 ;
    END
  END Tile_X0Y1_S2BEG[1]
  PIN Tile_X0Y1_S2BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 49.240 0.000 49.640 0.400 ;
    END
  END Tile_X0Y1_S2BEG[2]
  PIN Tile_X0Y1_S2BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 50.200 0.000 50.600 0.400 ;
    END
  END Tile_X0Y1_S2BEG[3]
  PIN Tile_X0Y1_S2BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 51.160 0.000 51.560 0.400 ;
    END
  END Tile_X0Y1_S2BEG[4]
  PIN Tile_X0Y1_S2BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 52.120 0.000 52.520 0.400 ;
    END
  END Tile_X0Y1_S2BEG[5]
  PIN Tile_X0Y1_S2BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 53.080 0.000 53.480 0.400 ;
    END
  END Tile_X0Y1_S2BEG[6]
  PIN Tile_X0Y1_S2BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 54.040 0.000 54.440 0.400 ;
    END
  END Tile_X0Y1_S2BEG[7]
  PIN Tile_X0Y1_S2BEGb[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 55.000 0.000 55.400 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[0]
  PIN Tile_X0Y1_S2BEGb[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 55.960 0.000 56.360 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[1]
  PIN Tile_X0Y1_S2BEGb[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 56.920 0.000 57.320 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[2]
  PIN Tile_X0Y1_S2BEGb[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 57.880 0.000 58.280 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[3]
  PIN Tile_X0Y1_S2BEGb[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 58.840 0.000 59.240 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[4]
  PIN Tile_X0Y1_S2BEGb[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 59.800 0.000 60.200 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[5]
  PIN Tile_X0Y1_S2BEGb[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 60.760 0.000 61.160 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[6]
  PIN Tile_X0Y1_S2BEGb[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 61.720 0.000 62.120 0.400 ;
    END
  END Tile_X0Y1_S2BEGb[7]
  PIN Tile_X0Y1_S4BEG[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 62.680 0.000 63.080 0.400 ;
    END
  END Tile_X0Y1_S4BEG[0]
  PIN Tile_X0Y1_S4BEG[10]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 72.280 0.000 72.680 0.400 ;
    END
  END Tile_X0Y1_S4BEG[10]
  PIN Tile_X0Y1_S4BEG[11]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 73.240 0.000 73.640 0.400 ;
    END
  END Tile_X0Y1_S4BEG[11]
  PIN Tile_X0Y1_S4BEG[12]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 74.200 0.000 74.600 0.400 ;
    END
  END Tile_X0Y1_S4BEG[12]
  PIN Tile_X0Y1_S4BEG[13]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 75.160 0.000 75.560 0.400 ;
    END
  END Tile_X0Y1_S4BEG[13]
  PIN Tile_X0Y1_S4BEG[14]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 76.120 0.000 76.520 0.400 ;
    END
  END Tile_X0Y1_S4BEG[14]
  PIN Tile_X0Y1_S4BEG[15]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 77.080 0.000 77.480 0.400 ;
    END
  END Tile_X0Y1_S4BEG[15]
  PIN Tile_X0Y1_S4BEG[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 63.640 0.000 64.040 0.400 ;
    END
  END Tile_X0Y1_S4BEG[1]
  PIN Tile_X0Y1_S4BEG[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 64.600 0.000 65.000 0.400 ;
    END
  END Tile_X0Y1_S4BEG[2]
  PIN Tile_X0Y1_S4BEG[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 65.560 0.000 65.960 0.400 ;
    END
  END Tile_X0Y1_S4BEG[3]
  PIN Tile_X0Y1_S4BEG[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 66.520 0.000 66.920 0.400 ;
    END
  END Tile_X0Y1_S4BEG[4]
  PIN Tile_X0Y1_S4BEG[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 67.480 0.000 67.880 0.400 ;
    END
  END Tile_X0Y1_S4BEG[5]
  PIN Tile_X0Y1_S4BEG[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 68.440 0.000 68.840 0.400 ;
    END
  END Tile_X0Y1_S4BEG[6]
  PIN Tile_X0Y1_S4BEG[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 0.000 69.800 0.400 ;
    END
  END Tile_X0Y1_S4BEG[7]
  PIN Tile_X0Y1_S4BEG[8]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 70.360 0.000 70.760 0.400 ;
    END
  END Tile_X0Y1_S4BEG[8]
  PIN Tile_X0Y1_S4BEG[9]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.708600 ;
    PORT
      LAYER Metal2 ;
        RECT 71.320 0.000 71.720 0.400 ;
    END
  END Tile_X0Y1_S4BEG[9]
  PIN Tile_X0Y1_UserCLK
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.725400 ;
    PORT
      LAYER Metal2 ;
        RECT 78.040 0.000 78.440 0.400 ;
    END
  END Tile_X0Y1_UserCLK
  PIN Tile_X0Y1_W1END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 0.220 107.520 0.620 ;
    END
  END Tile_X0Y1_W1END[0]
  PIN Tile_X0Y1_W1END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 1.900 107.520 2.300 ;
    END
  END Tile_X0Y1_W1END[1]
  PIN Tile_X0Y1_W1END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 3.580 107.520 3.980 ;
    END
  END Tile_X0Y1_W1END[2]
  PIN Tile_X0Y1_W1END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 5.260 107.520 5.660 ;
    END
  END Tile_X0Y1_W1END[3]
  PIN Tile_X0Y1_W2END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 20.380 107.520 20.780 ;
    END
  END Tile_X0Y1_W2END[0]
  PIN Tile_X0Y1_W2END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.820300 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 22.060 107.520 22.460 ;
    END
  END Tile_X0Y1_W2END[1]
  PIN Tile_X0Y1_W2END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.881400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 23.740 107.520 24.140 ;
    END
  END Tile_X0Y1_W2END[2]
  PIN Tile_X0Y1_W2END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.917800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 25.420 107.520 25.820 ;
    END
  END Tile_X0Y1_W2END[3]
  PIN Tile_X0Y1_W2END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.898300 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 27.100 107.520 27.500 ;
    END
  END Tile_X0Y1_W2END[4]
  PIN Tile_X0Y1_W2END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.910000 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 28.780 107.520 29.180 ;
    END
  END Tile_X0Y1_W2END[5]
  PIN Tile_X0Y1_W2END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 30.460 107.520 30.860 ;
    END
  END Tile_X0Y1_W2END[6]
  PIN Tile_X0Y1_W2END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 32.140 107.520 32.540 ;
    END
  END Tile_X0Y1_W2END[7]
  PIN Tile_X0Y1_W2MID[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.881400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 6.940 107.520 7.340 ;
    END
  END Tile_X0Y1_W2MID[0]
  PIN Tile_X0Y1_W2MID[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 8.620 107.520 9.020 ;
    END
  END Tile_X0Y1_W2MID[1]
  PIN Tile_X0Y1_W2MID[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 10.300 107.520 10.700 ;
    END
  END Tile_X0Y1_W2MID[2]
  PIN Tile_X0Y1_W2MID[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.787800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 11.980 107.520 12.380 ;
    END
  END Tile_X0Y1_W2MID[3]
  PIN Tile_X0Y1_W2MID[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 13.660 107.520 14.060 ;
    END
  END Tile_X0Y1_W2MID[4]
  PIN Tile_X0Y1_W2MID[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 15.340 107.520 15.740 ;
    END
  END Tile_X0Y1_W2MID[5]
  PIN Tile_X0Y1_W2MID[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.910000 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 17.020 107.520 17.420 ;
    END
  END Tile_X0Y1_W2MID[6]
  PIN Tile_X0Y1_W2MID[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 18.700 107.520 19.100 ;
    END
  END Tile_X0Y1_W2MID[7]
  PIN Tile_X0Y1_W6END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.668200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 60.700 107.520 61.100 ;
    END
  END Tile_X0Y1_W6END[0]
  PIN Tile_X0Y1_W6END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 77.500 107.520 77.900 ;
    END
  END Tile_X0Y1_W6END[10]
  PIN Tile_X0Y1_W6END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 79.180 107.520 79.580 ;
    END
  END Tile_X0Y1_W6END[11]
  PIN Tile_X0Y1_W6END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.668200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 62.380 107.520 62.780 ;
    END
  END Tile_X0Y1_W6END[1]
  PIN Tile_X0Y1_W6END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.668200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 64.060 107.520 64.460 ;
    END
  END Tile_X0Y1_W6END[2]
  PIN Tile_X0Y1_W6END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.668200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 65.740 107.520 66.140 ;
    END
  END Tile_X0Y1_W6END[3]
  PIN Tile_X0Y1_W6END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 67.420 107.520 67.820 ;
    END
  END Tile_X0Y1_W6END[4]
  PIN Tile_X0Y1_W6END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 69.100 107.520 69.500 ;
    END
  END Tile_X0Y1_W6END[5]
  PIN Tile_X0Y1_W6END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 70.780 107.520 71.180 ;
    END
  END Tile_X0Y1_W6END[6]
  PIN Tile_X0Y1_W6END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 72.460 107.520 72.860 ;
    END
  END Tile_X0Y1_W6END[7]
  PIN Tile_X0Y1_W6END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 74.140 107.520 74.540 ;
    END
  END Tile_X0Y1_W6END[8]
  PIN Tile_X0Y1_W6END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 75.820 107.520 76.220 ;
    END
  END Tile_X0Y1_W6END[9]
  PIN Tile_X0Y1_WW4END[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 33.820 107.520 34.220 ;
    END
  END Tile_X0Y1_WW4END[0]
  PIN Tile_X0Y1_WW4END[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 50.620 107.520 51.020 ;
    END
  END Tile_X0Y1_WW4END[10]
  PIN Tile_X0Y1_WW4END[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 52.300 107.520 52.700 ;
    END
  END Tile_X0Y1_WW4END[11]
  PIN Tile_X0Y1_WW4END[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 53.980 107.520 54.380 ;
    END
  END Tile_X0Y1_WW4END[12]
  PIN Tile_X0Y1_WW4END[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 55.660 107.520 56.060 ;
    END
  END Tile_X0Y1_WW4END[13]
  PIN Tile_X0Y1_WW4END[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 57.340 107.520 57.740 ;
    END
  END Tile_X0Y1_WW4END[14]
  PIN Tile_X0Y1_WW4END[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 59.020 107.520 59.420 ;
    END
  END Tile_X0Y1_WW4END[15]
  PIN Tile_X0Y1_WW4END[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 35.500 107.520 35.900 ;
    END
  END Tile_X0Y1_WW4END[1]
  PIN Tile_X0Y1_WW4END[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 37.180 107.520 37.580 ;
    END
  END Tile_X0Y1_WW4END[2]
  PIN Tile_X0Y1_WW4END[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.426400 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 38.860 107.520 39.260 ;
    END
  END Tile_X0Y1_WW4END[3]
  PIN Tile_X0Y1_WW4END[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 40.540 107.520 40.940 ;
    END
  END Tile_X0Y1_WW4END[4]
  PIN Tile_X0Y1_WW4END[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 42.220 107.520 42.620 ;
    END
  END Tile_X0Y1_WW4END[5]
  PIN Tile_X0Y1_WW4END[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 43.900 107.520 44.300 ;
    END
  END Tile_X0Y1_WW4END[6]
  PIN Tile_X0Y1_WW4END[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 45.580 107.520 45.980 ;
    END
  END Tile_X0Y1_WW4END[7]
  PIN Tile_X0Y1_WW4END[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 47.260 107.520 47.660 ;
    END
  END Tile_X0Y1_WW4END[8]
  PIN Tile_X0Y1_WW4END[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.213200 ;
    PORT
      LAYER Metal3 ;
        RECT 107.120 48.940 107.520 49.340 ;
    END
  END Tile_X0Y1_WW4END[9]
  PIN UIO_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 143.860 0.400 144.260 ;
    END
  END UIO_IN_TT_PROJECT0
  PIN UIO_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 147.220 0.400 147.620 ;
    END
  END UIO_IN_TT_PROJECT1
  PIN UIO_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.580 0.400 150.980 ;
    END
  END UIO_IN_TT_PROJECT2
  PIN UIO_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.662000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 153.940 0.400 154.340 ;
    END
  END UIO_IN_TT_PROJECT3
  PIN UIO_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.649200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 157.300 0.400 157.700 ;
    END
  END UIO_IN_TT_PROJECT4
  PIN UIO_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.649200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 160.660 0.400 161.060 ;
    END
  END UIO_IN_TT_PROJECT5
  PIN UIO_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.649200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 164.020 0.400 164.420 ;
    END
  END UIO_IN_TT_PROJECT6
  PIN UIO_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.649200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 167.380 0.400 167.780 ;
    END
  END UIO_IN_TT_PROJECT7
  PIN UIO_OE_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.066000 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 90.100 0.400 90.500 ;
    END
  END UIO_OE_TT_PROJECT0
  PIN UIO_OE_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.639600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 93.460 0.400 93.860 ;
    END
  END UIO_OE_TT_PROJECT1
  PIN UIO_OE_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 96.820 0.400 97.220 ;
    END
  END UIO_OE_TT_PROJECT2
  PIN UIO_OE_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 100.180 0.400 100.580 ;
    END
  END UIO_OE_TT_PROJECT3
  PIN UIO_OE_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 103.540 0.400 103.940 ;
    END
  END UIO_OE_TT_PROJECT4
  PIN UIO_OE_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 106.900 0.400 107.300 ;
    END
  END UIO_OE_TT_PROJECT5
  PIN UIO_OE_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 110.260 0.400 110.660 ;
    END
  END UIO_OE_TT_PROJECT6
  PIN UIO_OE_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.852800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 113.620 0.400 114.020 ;
    END
  END UIO_OE_TT_PROJECT7
  PIN UIO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 5.538000 ;
    ANTENNADIFFAREA 14.107800 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 63.220 0.400 63.620 ;
    END
  END UIO_OUT_TT_PROJECT0
  PIN UIO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 66.580 0.400 66.980 ;
    END
  END UIO_OUT_TT_PROJECT1
  PIN UIO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 69.940 0.400 70.340 ;
    END
  END UIO_OUT_TT_PROJECT2
  PIN UIO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 73.300 0.400 73.700 ;
    END
  END UIO_OUT_TT_PROJECT3
  PIN UIO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 76.660 0.400 77.060 ;
    END
  END UIO_OUT_TT_PROJECT4
  PIN UIO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 80.020 0.400 80.420 ;
    END
  END UIO_OUT_TT_PROJECT5
  PIN UIO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 83.380 0.400 83.780 ;
    END
  END UIO_OUT_TT_PROJECT6
  PIN UIO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.279200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.740 0.400 87.140 ;
    END
  END UIO_OUT_TT_PROJECT7
  PIN UI_IN_TT_PROJECT0
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 116.980 0.400 117.380 ;
    END
  END UI_IN_TT_PROJECT0
  PIN UI_IN_TT_PROJECT1
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 120.340 0.400 120.740 ;
    END
  END UI_IN_TT_PROJECT1
  PIN UI_IN_TT_PROJECT2
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 123.700 0.400 124.100 ;
    END
  END UI_IN_TT_PROJECT2
  PIN UI_IN_TT_PROJECT3
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 1.008100 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 127.060 0.400 127.460 ;
    END
  END UI_IN_TT_PROJECT3
  PIN UI_IN_TT_PROJECT4
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 130.420 0.400 130.820 ;
    END
  END UI_IN_TT_PROJECT4
  PIN UI_IN_TT_PROJECT5
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 133.780 0.400 134.180 ;
    END
  END UI_IN_TT_PROJECT5
  PIN UI_IN_TT_PROJECT6
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 137.140 0.400 137.540 ;
    END
  END UI_IN_TT_PROJECT6
  PIN UI_IN_TT_PROJECT7
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.677200 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 140.500 0.400 140.900 ;
    END
  END UI_IN_TT_PROJECT7
  PIN UO_OUT_TT_PROJECT0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.770600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 36.340 0.400 36.740 ;
    END
  END UO_OUT_TT_PROJECT0
  PIN UO_OUT_TT_PROJECT1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.770600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 39.700 0.400 40.100 ;
    END
  END UO_OUT_TT_PROJECT1
  PIN UO_OUT_TT_PROJECT2
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.770600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 43.060 0.400 43.460 ;
    END
  END UO_OUT_TT_PROJECT2
  PIN UO_OUT_TT_PROJECT3
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.770600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 46.420 0.400 46.820 ;
    END
  END UO_OUT_TT_PROJECT3
  PIN UO_OUT_TT_PROJECT4
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.770600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 49.780 0.400 50.180 ;
    END
  END UO_OUT_TT_PROJECT4
  PIN UO_OUT_TT_PROJECT5
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.770600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 53.140 0.400 53.540 ;
    END
  END UO_OUT_TT_PROJECT5
  PIN UO_OUT_TT_PROJECT6
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.770600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 56.500 0.400 56.900 ;
    END
  END UO_OUT_TT_PROJECT6
  PIN UO_OUT_TT_PROJECT7
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.770600 ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 59.860 0.400 60.260 ;
    END
  END UO_OUT_TT_PROJECT7
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER TopMetal1 ;
        RECT 24.460 0.000 26.660 430.080 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 100.060 0.000 102.260 430.080 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER TopMetal1 ;
        RECT 18.260 0.000 20.460 430.080 ;
    END
    PORT
      LAYER TopMetal1 ;
        RECT 93.860 0.000 96.060 430.080 ;
    END
  END VPWR
  OBS
      LAYER GatPoly ;
        RECT 5.760 3.630 101.760 423.510 ;
      LAYER Metal1 ;
        RECT 5.760 3.560 102.260 423.580 ;
      LAYER Metal2 ;
        RECT 0.375 429.470 8.710 429.680 ;
        RECT 9.530 429.470 9.670 429.680 ;
        RECT 10.490 429.470 10.630 429.680 ;
        RECT 11.450 429.470 11.590 429.680 ;
        RECT 12.410 429.470 12.550 429.680 ;
        RECT 13.370 429.470 13.510 429.680 ;
        RECT 14.330 429.470 14.470 429.680 ;
        RECT 15.290 429.470 15.430 429.680 ;
        RECT 16.250 429.470 16.390 429.680 ;
        RECT 17.210 429.470 17.350 429.680 ;
        RECT 18.170 429.470 18.310 429.680 ;
        RECT 19.130 429.470 19.270 429.680 ;
        RECT 20.090 429.470 20.230 429.680 ;
        RECT 21.050 429.470 21.190 429.680 ;
        RECT 22.010 429.470 22.150 429.680 ;
        RECT 22.970 429.470 23.110 429.680 ;
        RECT 23.930 429.470 24.070 429.680 ;
        RECT 24.890 429.470 25.030 429.680 ;
        RECT 25.850 429.470 25.990 429.680 ;
        RECT 26.810 429.470 26.950 429.680 ;
        RECT 27.770 429.470 27.910 429.680 ;
        RECT 28.730 429.470 28.870 429.680 ;
        RECT 29.690 429.470 29.830 429.680 ;
        RECT 30.650 429.470 30.790 429.680 ;
        RECT 31.610 429.470 31.750 429.680 ;
        RECT 32.570 429.470 32.710 429.680 ;
        RECT 33.530 429.470 33.670 429.680 ;
        RECT 34.490 429.470 34.630 429.680 ;
        RECT 35.450 429.470 35.590 429.680 ;
        RECT 36.410 429.470 36.550 429.680 ;
        RECT 37.370 429.470 37.510 429.680 ;
        RECT 38.330 429.470 38.470 429.680 ;
        RECT 39.290 429.470 39.430 429.680 ;
        RECT 40.250 429.470 40.390 429.680 ;
        RECT 41.210 429.470 41.350 429.680 ;
        RECT 42.170 429.470 42.310 429.680 ;
        RECT 43.130 429.470 43.270 429.680 ;
        RECT 44.090 429.470 44.230 429.680 ;
        RECT 45.050 429.470 45.190 429.680 ;
        RECT 46.010 429.470 46.150 429.680 ;
        RECT 46.970 429.470 47.110 429.680 ;
        RECT 47.930 429.470 48.070 429.680 ;
        RECT 48.890 429.470 49.030 429.680 ;
        RECT 49.850 429.470 49.990 429.680 ;
        RECT 50.810 429.470 50.950 429.680 ;
        RECT 51.770 429.470 51.910 429.680 ;
        RECT 52.730 429.470 52.870 429.680 ;
        RECT 53.690 429.470 53.830 429.680 ;
        RECT 54.650 429.470 54.790 429.680 ;
        RECT 55.610 429.470 55.750 429.680 ;
        RECT 56.570 429.470 56.710 429.680 ;
        RECT 57.530 429.470 57.670 429.680 ;
        RECT 58.490 429.470 58.630 429.680 ;
        RECT 59.450 429.470 59.590 429.680 ;
        RECT 60.410 429.470 60.550 429.680 ;
        RECT 61.370 429.470 61.510 429.680 ;
        RECT 62.330 429.470 62.470 429.680 ;
        RECT 63.290 429.470 63.430 429.680 ;
        RECT 64.250 429.470 64.390 429.680 ;
        RECT 65.210 429.470 65.350 429.680 ;
        RECT 66.170 429.470 66.310 429.680 ;
        RECT 67.130 429.470 67.270 429.680 ;
        RECT 68.090 429.470 68.230 429.680 ;
        RECT 69.050 429.470 69.190 429.680 ;
        RECT 70.010 429.470 70.150 429.680 ;
        RECT 70.970 429.470 71.110 429.680 ;
        RECT 71.930 429.470 72.070 429.680 ;
        RECT 72.890 429.470 73.030 429.680 ;
        RECT 73.850 429.470 73.990 429.680 ;
        RECT 74.810 429.470 74.950 429.680 ;
        RECT 75.770 429.470 75.910 429.680 ;
        RECT 76.730 429.470 76.870 429.680 ;
        RECT 77.690 429.470 77.830 429.680 ;
        RECT 78.650 429.470 78.790 429.680 ;
        RECT 79.610 429.470 79.750 429.680 ;
        RECT 80.570 429.470 80.710 429.680 ;
        RECT 81.530 429.470 81.670 429.680 ;
        RECT 82.490 429.470 82.630 429.680 ;
        RECT 83.450 429.470 83.590 429.680 ;
        RECT 84.410 429.470 84.550 429.680 ;
        RECT 85.370 429.470 85.510 429.680 ;
        RECT 86.330 429.470 86.470 429.680 ;
        RECT 87.290 429.470 87.430 429.680 ;
        RECT 88.250 429.470 88.390 429.680 ;
        RECT 89.210 429.470 89.350 429.680 ;
        RECT 90.170 429.470 90.310 429.680 ;
        RECT 91.130 429.470 91.270 429.680 ;
        RECT 92.090 429.470 92.230 429.680 ;
        RECT 93.050 429.470 93.190 429.680 ;
        RECT 94.010 429.470 94.150 429.680 ;
        RECT 94.970 429.470 95.110 429.680 ;
        RECT 95.930 429.470 96.070 429.680 ;
        RECT 96.890 429.470 97.030 429.680 ;
        RECT 97.850 429.470 107.145 429.680 ;
        RECT 0.375 0.610 107.145 429.470 ;
        RECT 0.375 0.100 8.710 0.610 ;
        RECT 9.530 0.100 9.670 0.610 ;
        RECT 10.490 0.100 10.630 0.610 ;
        RECT 11.450 0.100 11.590 0.610 ;
        RECT 12.410 0.100 12.550 0.610 ;
        RECT 13.370 0.100 13.510 0.610 ;
        RECT 14.330 0.100 14.470 0.610 ;
        RECT 15.290 0.100 15.430 0.610 ;
        RECT 16.250 0.100 16.390 0.610 ;
        RECT 17.210 0.100 17.350 0.610 ;
        RECT 18.170 0.100 18.310 0.610 ;
        RECT 19.130 0.100 19.270 0.610 ;
        RECT 20.090 0.100 20.230 0.610 ;
        RECT 21.050 0.100 21.190 0.610 ;
        RECT 22.010 0.100 22.150 0.610 ;
        RECT 22.970 0.100 23.110 0.610 ;
        RECT 23.930 0.100 24.070 0.610 ;
        RECT 24.890 0.100 25.030 0.610 ;
        RECT 25.850 0.100 25.990 0.610 ;
        RECT 26.810 0.100 26.950 0.610 ;
        RECT 27.770 0.100 27.910 0.610 ;
        RECT 28.730 0.100 28.870 0.610 ;
        RECT 29.690 0.100 29.830 0.610 ;
        RECT 30.650 0.100 30.790 0.610 ;
        RECT 31.610 0.100 31.750 0.610 ;
        RECT 32.570 0.100 32.710 0.610 ;
        RECT 33.530 0.100 33.670 0.610 ;
        RECT 34.490 0.100 34.630 0.610 ;
        RECT 35.450 0.100 35.590 0.610 ;
        RECT 36.410 0.100 36.550 0.610 ;
        RECT 37.370 0.100 37.510 0.610 ;
        RECT 38.330 0.100 38.470 0.610 ;
        RECT 39.290 0.100 39.430 0.610 ;
        RECT 40.250 0.100 40.390 0.610 ;
        RECT 41.210 0.100 41.350 0.610 ;
        RECT 42.170 0.100 42.310 0.610 ;
        RECT 43.130 0.100 43.270 0.610 ;
        RECT 44.090 0.100 44.230 0.610 ;
        RECT 45.050 0.100 45.190 0.610 ;
        RECT 46.010 0.100 46.150 0.610 ;
        RECT 46.970 0.100 47.110 0.610 ;
        RECT 47.930 0.100 48.070 0.610 ;
        RECT 48.890 0.100 49.030 0.610 ;
        RECT 49.850 0.100 49.990 0.610 ;
        RECT 50.810 0.100 50.950 0.610 ;
        RECT 51.770 0.100 51.910 0.610 ;
        RECT 52.730 0.100 52.870 0.610 ;
        RECT 53.690 0.100 53.830 0.610 ;
        RECT 54.650 0.100 54.790 0.610 ;
        RECT 55.610 0.100 55.750 0.610 ;
        RECT 56.570 0.100 56.710 0.610 ;
        RECT 57.530 0.100 57.670 0.610 ;
        RECT 58.490 0.100 58.630 0.610 ;
        RECT 59.450 0.100 59.590 0.610 ;
        RECT 60.410 0.100 60.550 0.610 ;
        RECT 61.370 0.100 61.510 0.610 ;
        RECT 62.330 0.100 62.470 0.610 ;
        RECT 63.290 0.100 63.430 0.610 ;
        RECT 64.250 0.100 64.390 0.610 ;
        RECT 65.210 0.100 65.350 0.610 ;
        RECT 66.170 0.100 66.310 0.610 ;
        RECT 67.130 0.100 67.270 0.610 ;
        RECT 68.090 0.100 68.230 0.610 ;
        RECT 69.050 0.100 69.190 0.610 ;
        RECT 70.010 0.100 70.150 0.610 ;
        RECT 70.970 0.100 71.110 0.610 ;
        RECT 71.930 0.100 72.070 0.610 ;
        RECT 72.890 0.100 73.030 0.610 ;
        RECT 73.850 0.100 73.990 0.610 ;
        RECT 74.810 0.100 74.950 0.610 ;
        RECT 75.770 0.100 75.910 0.610 ;
        RECT 76.730 0.100 76.870 0.610 ;
        RECT 77.690 0.100 77.830 0.610 ;
        RECT 78.650 0.100 78.790 0.610 ;
        RECT 79.610 0.100 79.750 0.610 ;
        RECT 80.570 0.100 80.710 0.610 ;
        RECT 81.530 0.100 81.670 0.610 ;
        RECT 82.490 0.100 82.630 0.610 ;
        RECT 83.450 0.100 83.590 0.610 ;
        RECT 84.410 0.100 84.550 0.610 ;
        RECT 85.370 0.100 85.510 0.610 ;
        RECT 86.330 0.100 86.470 0.610 ;
        RECT 87.290 0.100 87.430 0.610 ;
        RECT 88.250 0.100 88.390 0.610 ;
        RECT 89.210 0.100 89.350 0.610 ;
        RECT 90.170 0.100 90.310 0.610 ;
        RECT 91.130 0.100 91.270 0.610 ;
        RECT 92.090 0.100 92.230 0.610 ;
        RECT 93.050 0.100 93.190 0.610 ;
        RECT 94.010 0.100 94.150 0.610 ;
        RECT 94.970 0.100 95.110 0.610 ;
        RECT 95.930 0.100 96.070 0.610 ;
        RECT 96.890 0.100 97.030 0.610 ;
        RECT 97.850 0.100 107.145 0.610 ;
      LAYER Metal3 ;
        RECT 0.100 429.230 107.185 429.765 ;
        RECT 0.100 428.410 106.910 429.230 ;
        RECT 0.100 427.550 107.185 428.410 ;
        RECT 0.100 426.730 106.910 427.550 ;
        RECT 0.100 425.870 107.185 426.730 ;
        RECT 0.100 425.050 106.910 425.870 ;
        RECT 0.100 424.190 107.185 425.050 ;
        RECT 0.100 423.370 106.910 424.190 ;
        RECT 0.100 422.510 107.185 423.370 ;
        RECT 0.100 421.690 106.910 422.510 ;
        RECT 0.100 420.830 107.185 421.690 ;
        RECT 0.100 420.010 106.910 420.830 ;
        RECT 0.100 419.150 107.185 420.010 ;
        RECT 0.100 418.330 106.910 419.150 ;
        RECT 0.100 417.470 107.185 418.330 ;
        RECT 0.100 416.650 106.910 417.470 ;
        RECT 0.100 415.790 107.185 416.650 ;
        RECT 0.100 414.970 106.910 415.790 ;
        RECT 0.100 414.110 107.185 414.970 ;
        RECT 0.100 413.290 106.910 414.110 ;
        RECT 0.100 412.430 107.185 413.290 ;
        RECT 0.100 411.610 106.910 412.430 ;
        RECT 0.100 410.750 107.185 411.610 ;
        RECT 0.100 409.930 106.910 410.750 ;
        RECT 0.100 409.070 107.185 409.930 ;
        RECT 0.100 408.250 106.910 409.070 ;
        RECT 0.100 407.390 107.185 408.250 ;
        RECT 0.100 406.570 106.910 407.390 ;
        RECT 0.100 405.710 107.185 406.570 ;
        RECT 0.100 404.890 106.910 405.710 ;
        RECT 0.100 404.030 107.185 404.890 ;
        RECT 0.100 403.210 106.910 404.030 ;
        RECT 0.100 402.350 107.185 403.210 ;
        RECT 0.100 401.530 106.910 402.350 ;
        RECT 0.100 400.670 107.185 401.530 ;
        RECT 0.100 399.850 106.910 400.670 ;
        RECT 0.100 398.990 107.185 399.850 ;
        RECT 0.100 398.170 106.910 398.990 ;
        RECT 0.100 397.310 107.185 398.170 ;
        RECT 0.100 396.490 106.910 397.310 ;
        RECT 0.100 395.630 107.185 396.490 ;
        RECT 0.100 394.810 106.910 395.630 ;
        RECT 0.100 393.950 107.185 394.810 ;
        RECT 0.100 393.130 106.910 393.950 ;
        RECT 0.100 393.110 107.185 393.130 ;
        RECT 0.610 392.290 107.185 393.110 ;
        RECT 0.100 392.270 107.185 392.290 ;
        RECT 0.100 391.450 106.910 392.270 ;
        RECT 0.100 390.590 107.185 391.450 ;
        RECT 0.100 389.770 106.910 390.590 ;
        RECT 0.100 389.750 107.185 389.770 ;
        RECT 0.610 388.930 107.185 389.750 ;
        RECT 0.100 388.910 107.185 388.930 ;
        RECT 0.100 388.090 106.910 388.910 ;
        RECT 0.100 387.230 107.185 388.090 ;
        RECT 0.100 386.410 106.910 387.230 ;
        RECT 0.100 386.390 107.185 386.410 ;
        RECT 0.610 385.570 107.185 386.390 ;
        RECT 0.100 385.550 107.185 385.570 ;
        RECT 0.100 384.730 106.910 385.550 ;
        RECT 0.100 383.870 107.185 384.730 ;
        RECT 0.100 383.050 106.910 383.870 ;
        RECT 0.100 383.030 107.185 383.050 ;
        RECT 0.610 382.210 107.185 383.030 ;
        RECT 0.100 382.190 107.185 382.210 ;
        RECT 0.100 381.370 106.910 382.190 ;
        RECT 0.100 380.510 107.185 381.370 ;
        RECT 0.100 379.690 106.910 380.510 ;
        RECT 0.100 379.670 107.185 379.690 ;
        RECT 0.610 378.850 107.185 379.670 ;
        RECT 0.100 378.830 107.185 378.850 ;
        RECT 0.100 378.010 106.910 378.830 ;
        RECT 0.100 377.150 107.185 378.010 ;
        RECT 0.100 376.330 106.910 377.150 ;
        RECT 0.100 376.310 107.185 376.330 ;
        RECT 0.610 375.490 107.185 376.310 ;
        RECT 0.100 375.470 107.185 375.490 ;
        RECT 0.100 374.650 106.910 375.470 ;
        RECT 0.100 373.790 107.185 374.650 ;
        RECT 0.100 372.970 106.910 373.790 ;
        RECT 0.100 372.950 107.185 372.970 ;
        RECT 0.610 372.130 107.185 372.950 ;
        RECT 0.100 372.110 107.185 372.130 ;
        RECT 0.100 371.290 106.910 372.110 ;
        RECT 0.100 370.430 107.185 371.290 ;
        RECT 0.100 369.610 106.910 370.430 ;
        RECT 0.100 369.590 107.185 369.610 ;
        RECT 0.610 368.770 107.185 369.590 ;
        RECT 0.100 368.750 107.185 368.770 ;
        RECT 0.100 367.930 106.910 368.750 ;
        RECT 0.100 367.070 107.185 367.930 ;
        RECT 0.100 366.250 106.910 367.070 ;
        RECT 0.100 366.230 107.185 366.250 ;
        RECT 0.610 365.410 107.185 366.230 ;
        RECT 0.100 365.390 107.185 365.410 ;
        RECT 0.100 364.570 106.910 365.390 ;
        RECT 0.100 363.710 107.185 364.570 ;
        RECT 0.100 362.890 106.910 363.710 ;
        RECT 0.100 362.870 107.185 362.890 ;
        RECT 0.610 362.050 107.185 362.870 ;
        RECT 0.100 362.030 107.185 362.050 ;
        RECT 0.100 361.210 106.910 362.030 ;
        RECT 0.100 360.350 107.185 361.210 ;
        RECT 0.100 359.530 106.910 360.350 ;
        RECT 0.100 359.510 107.185 359.530 ;
        RECT 0.610 358.690 107.185 359.510 ;
        RECT 0.100 358.670 107.185 358.690 ;
        RECT 0.100 357.850 106.910 358.670 ;
        RECT 0.100 356.990 107.185 357.850 ;
        RECT 0.100 356.170 106.910 356.990 ;
        RECT 0.100 356.150 107.185 356.170 ;
        RECT 0.610 355.330 107.185 356.150 ;
        RECT 0.100 355.310 107.185 355.330 ;
        RECT 0.100 354.490 106.910 355.310 ;
        RECT 0.100 353.630 107.185 354.490 ;
        RECT 0.100 352.810 106.910 353.630 ;
        RECT 0.100 352.790 107.185 352.810 ;
        RECT 0.610 351.970 107.185 352.790 ;
        RECT 0.100 351.950 107.185 351.970 ;
        RECT 0.100 351.130 106.910 351.950 ;
        RECT 0.100 350.270 107.185 351.130 ;
        RECT 0.100 349.450 106.910 350.270 ;
        RECT 0.100 349.430 107.185 349.450 ;
        RECT 0.610 348.610 107.185 349.430 ;
        RECT 0.100 348.590 107.185 348.610 ;
        RECT 0.100 347.770 106.910 348.590 ;
        RECT 0.100 346.910 107.185 347.770 ;
        RECT 0.100 346.090 106.910 346.910 ;
        RECT 0.100 346.070 107.185 346.090 ;
        RECT 0.610 345.250 107.185 346.070 ;
        RECT 0.100 345.230 107.185 345.250 ;
        RECT 0.100 344.410 106.910 345.230 ;
        RECT 0.100 343.550 107.185 344.410 ;
        RECT 0.100 342.730 106.910 343.550 ;
        RECT 0.100 342.710 107.185 342.730 ;
        RECT 0.610 341.890 107.185 342.710 ;
        RECT 0.100 341.870 107.185 341.890 ;
        RECT 0.100 341.050 106.910 341.870 ;
        RECT 0.100 340.190 107.185 341.050 ;
        RECT 0.100 339.370 106.910 340.190 ;
        RECT 0.100 339.350 107.185 339.370 ;
        RECT 0.610 338.530 107.185 339.350 ;
        RECT 0.100 338.510 107.185 338.530 ;
        RECT 0.100 337.690 106.910 338.510 ;
        RECT 0.100 336.830 107.185 337.690 ;
        RECT 0.100 336.010 106.910 336.830 ;
        RECT 0.100 335.990 107.185 336.010 ;
        RECT 0.610 335.170 107.185 335.990 ;
        RECT 0.100 335.150 107.185 335.170 ;
        RECT 0.100 334.330 106.910 335.150 ;
        RECT 0.100 333.470 107.185 334.330 ;
        RECT 0.100 332.650 106.910 333.470 ;
        RECT 0.100 332.630 107.185 332.650 ;
        RECT 0.610 331.810 107.185 332.630 ;
        RECT 0.100 331.790 107.185 331.810 ;
        RECT 0.100 330.970 106.910 331.790 ;
        RECT 0.100 330.110 107.185 330.970 ;
        RECT 0.100 329.290 106.910 330.110 ;
        RECT 0.100 329.270 107.185 329.290 ;
        RECT 0.610 328.450 107.185 329.270 ;
        RECT 0.100 328.430 107.185 328.450 ;
        RECT 0.100 327.610 106.910 328.430 ;
        RECT 0.100 326.750 107.185 327.610 ;
        RECT 0.100 325.930 106.910 326.750 ;
        RECT 0.100 325.910 107.185 325.930 ;
        RECT 0.610 325.090 107.185 325.910 ;
        RECT 0.100 325.070 107.185 325.090 ;
        RECT 0.100 324.250 106.910 325.070 ;
        RECT 0.100 323.390 107.185 324.250 ;
        RECT 0.100 322.570 106.910 323.390 ;
        RECT 0.100 322.550 107.185 322.570 ;
        RECT 0.610 321.730 107.185 322.550 ;
        RECT 0.100 321.710 107.185 321.730 ;
        RECT 0.100 320.890 106.910 321.710 ;
        RECT 0.100 320.030 107.185 320.890 ;
        RECT 0.100 319.210 106.910 320.030 ;
        RECT 0.100 319.190 107.185 319.210 ;
        RECT 0.610 318.370 107.185 319.190 ;
        RECT 0.100 318.350 107.185 318.370 ;
        RECT 0.100 317.530 106.910 318.350 ;
        RECT 0.100 316.670 107.185 317.530 ;
        RECT 0.100 315.850 106.910 316.670 ;
        RECT 0.100 315.830 107.185 315.850 ;
        RECT 0.610 315.010 107.185 315.830 ;
        RECT 0.100 314.990 107.185 315.010 ;
        RECT 0.100 314.170 106.910 314.990 ;
        RECT 0.100 313.310 107.185 314.170 ;
        RECT 0.100 312.490 106.910 313.310 ;
        RECT 0.100 312.470 107.185 312.490 ;
        RECT 0.610 311.650 107.185 312.470 ;
        RECT 0.100 311.630 107.185 311.650 ;
        RECT 0.100 310.810 106.910 311.630 ;
        RECT 0.100 309.950 107.185 310.810 ;
        RECT 0.100 309.130 106.910 309.950 ;
        RECT 0.100 309.110 107.185 309.130 ;
        RECT 0.610 308.290 107.185 309.110 ;
        RECT 0.100 308.270 107.185 308.290 ;
        RECT 0.100 307.450 106.910 308.270 ;
        RECT 0.100 306.590 107.185 307.450 ;
        RECT 0.100 305.770 106.910 306.590 ;
        RECT 0.100 305.750 107.185 305.770 ;
        RECT 0.610 304.930 107.185 305.750 ;
        RECT 0.100 304.910 107.185 304.930 ;
        RECT 0.100 304.090 106.910 304.910 ;
        RECT 0.100 303.230 107.185 304.090 ;
        RECT 0.100 302.410 106.910 303.230 ;
        RECT 0.100 302.390 107.185 302.410 ;
        RECT 0.610 301.570 107.185 302.390 ;
        RECT 0.100 301.550 107.185 301.570 ;
        RECT 0.100 300.730 106.910 301.550 ;
        RECT 0.100 299.870 107.185 300.730 ;
        RECT 0.100 299.050 106.910 299.870 ;
        RECT 0.100 299.030 107.185 299.050 ;
        RECT 0.610 298.210 107.185 299.030 ;
        RECT 0.100 298.190 107.185 298.210 ;
        RECT 0.100 297.370 106.910 298.190 ;
        RECT 0.100 296.510 107.185 297.370 ;
        RECT 0.100 295.690 106.910 296.510 ;
        RECT 0.100 295.670 107.185 295.690 ;
        RECT 0.610 294.850 107.185 295.670 ;
        RECT 0.100 294.830 107.185 294.850 ;
        RECT 0.100 294.010 106.910 294.830 ;
        RECT 0.100 293.150 107.185 294.010 ;
        RECT 0.100 292.330 106.910 293.150 ;
        RECT 0.100 292.310 107.185 292.330 ;
        RECT 0.610 291.490 107.185 292.310 ;
        RECT 0.100 291.470 107.185 291.490 ;
        RECT 0.100 290.650 106.910 291.470 ;
        RECT 0.100 289.790 107.185 290.650 ;
        RECT 0.100 288.970 106.910 289.790 ;
        RECT 0.100 288.950 107.185 288.970 ;
        RECT 0.610 288.130 107.185 288.950 ;
        RECT 0.100 288.110 107.185 288.130 ;
        RECT 0.100 287.290 106.910 288.110 ;
        RECT 0.100 286.430 107.185 287.290 ;
        RECT 0.100 285.610 106.910 286.430 ;
        RECT 0.100 285.590 107.185 285.610 ;
        RECT 0.610 284.770 107.185 285.590 ;
        RECT 0.100 284.750 107.185 284.770 ;
        RECT 0.100 283.930 106.910 284.750 ;
        RECT 0.100 283.070 107.185 283.930 ;
        RECT 0.100 282.250 106.910 283.070 ;
        RECT 0.100 282.230 107.185 282.250 ;
        RECT 0.610 281.410 107.185 282.230 ;
        RECT 0.100 281.390 107.185 281.410 ;
        RECT 0.100 280.570 106.910 281.390 ;
        RECT 0.100 279.710 107.185 280.570 ;
        RECT 0.100 278.890 106.910 279.710 ;
        RECT 0.100 278.870 107.185 278.890 ;
        RECT 0.610 278.050 107.185 278.870 ;
        RECT 0.100 278.030 107.185 278.050 ;
        RECT 0.100 277.210 106.910 278.030 ;
        RECT 0.100 276.350 107.185 277.210 ;
        RECT 0.100 275.530 106.910 276.350 ;
        RECT 0.100 275.510 107.185 275.530 ;
        RECT 0.610 274.690 107.185 275.510 ;
        RECT 0.100 274.670 107.185 274.690 ;
        RECT 0.100 273.850 106.910 274.670 ;
        RECT 0.100 272.990 107.185 273.850 ;
        RECT 0.100 272.170 106.910 272.990 ;
        RECT 0.100 272.150 107.185 272.170 ;
        RECT 0.610 271.330 107.185 272.150 ;
        RECT 0.100 271.310 107.185 271.330 ;
        RECT 0.100 270.490 106.910 271.310 ;
        RECT 0.100 269.630 107.185 270.490 ;
        RECT 0.100 268.810 106.910 269.630 ;
        RECT 0.100 268.790 107.185 268.810 ;
        RECT 0.610 267.970 107.185 268.790 ;
        RECT 0.100 267.950 107.185 267.970 ;
        RECT 0.100 267.130 106.910 267.950 ;
        RECT 0.100 266.270 107.185 267.130 ;
        RECT 0.100 265.450 106.910 266.270 ;
        RECT 0.100 265.430 107.185 265.450 ;
        RECT 0.610 264.610 107.185 265.430 ;
        RECT 0.100 264.590 107.185 264.610 ;
        RECT 0.100 263.770 106.910 264.590 ;
        RECT 0.100 262.910 107.185 263.770 ;
        RECT 0.100 262.090 106.910 262.910 ;
        RECT 0.100 262.070 107.185 262.090 ;
        RECT 0.610 261.250 107.185 262.070 ;
        RECT 0.100 261.230 107.185 261.250 ;
        RECT 0.100 260.410 106.910 261.230 ;
        RECT 0.100 259.550 107.185 260.410 ;
        RECT 0.100 258.730 106.910 259.550 ;
        RECT 0.100 258.710 107.185 258.730 ;
        RECT 0.610 257.890 107.185 258.710 ;
        RECT 0.100 257.870 107.185 257.890 ;
        RECT 0.100 257.050 106.910 257.870 ;
        RECT 0.100 256.190 107.185 257.050 ;
        RECT 0.100 255.370 106.910 256.190 ;
        RECT 0.100 255.350 107.185 255.370 ;
        RECT 0.610 254.530 107.185 255.350 ;
        RECT 0.100 254.510 107.185 254.530 ;
        RECT 0.100 253.690 106.910 254.510 ;
        RECT 0.100 252.830 107.185 253.690 ;
        RECT 0.100 252.010 106.910 252.830 ;
        RECT 0.100 251.990 107.185 252.010 ;
        RECT 0.610 251.170 107.185 251.990 ;
        RECT 0.100 251.150 107.185 251.170 ;
        RECT 0.100 250.330 106.910 251.150 ;
        RECT 0.100 249.470 107.185 250.330 ;
        RECT 0.100 248.650 106.910 249.470 ;
        RECT 0.100 248.630 107.185 248.650 ;
        RECT 0.610 247.810 107.185 248.630 ;
        RECT 0.100 247.790 107.185 247.810 ;
        RECT 0.100 246.970 106.910 247.790 ;
        RECT 0.100 246.110 107.185 246.970 ;
        RECT 0.100 245.290 106.910 246.110 ;
        RECT 0.100 245.270 107.185 245.290 ;
        RECT 0.610 244.450 107.185 245.270 ;
        RECT 0.100 244.430 107.185 244.450 ;
        RECT 0.100 243.610 106.910 244.430 ;
        RECT 0.100 242.750 107.185 243.610 ;
        RECT 0.100 241.930 106.910 242.750 ;
        RECT 0.100 241.910 107.185 241.930 ;
        RECT 0.610 241.090 107.185 241.910 ;
        RECT 0.100 241.070 107.185 241.090 ;
        RECT 0.100 240.250 106.910 241.070 ;
        RECT 0.100 239.390 107.185 240.250 ;
        RECT 0.100 238.570 106.910 239.390 ;
        RECT 0.100 238.550 107.185 238.570 ;
        RECT 0.610 237.730 107.185 238.550 ;
        RECT 0.100 237.710 107.185 237.730 ;
        RECT 0.100 236.890 106.910 237.710 ;
        RECT 0.100 236.030 107.185 236.890 ;
        RECT 0.100 235.210 106.910 236.030 ;
        RECT 0.100 235.190 107.185 235.210 ;
        RECT 0.610 234.370 107.185 235.190 ;
        RECT 0.100 234.350 107.185 234.370 ;
        RECT 0.100 233.530 106.910 234.350 ;
        RECT 0.100 232.670 107.185 233.530 ;
        RECT 0.100 231.850 106.910 232.670 ;
        RECT 0.100 231.830 107.185 231.850 ;
        RECT 0.610 231.010 107.185 231.830 ;
        RECT 0.100 230.990 107.185 231.010 ;
        RECT 0.100 230.170 106.910 230.990 ;
        RECT 0.100 229.310 107.185 230.170 ;
        RECT 0.100 228.490 106.910 229.310 ;
        RECT 0.100 228.470 107.185 228.490 ;
        RECT 0.610 227.650 107.185 228.470 ;
        RECT 0.100 227.630 107.185 227.650 ;
        RECT 0.100 226.810 106.910 227.630 ;
        RECT 0.100 225.950 107.185 226.810 ;
        RECT 0.100 225.130 106.910 225.950 ;
        RECT 0.100 225.110 107.185 225.130 ;
        RECT 0.610 224.290 107.185 225.110 ;
        RECT 0.100 224.270 107.185 224.290 ;
        RECT 0.100 223.450 106.910 224.270 ;
        RECT 0.100 222.590 107.185 223.450 ;
        RECT 0.100 221.770 106.910 222.590 ;
        RECT 0.100 221.750 107.185 221.770 ;
        RECT 0.610 220.930 107.185 221.750 ;
        RECT 0.100 220.910 107.185 220.930 ;
        RECT 0.100 220.090 106.910 220.910 ;
        RECT 0.100 219.230 107.185 220.090 ;
        RECT 0.100 218.410 106.910 219.230 ;
        RECT 0.100 218.390 107.185 218.410 ;
        RECT 0.610 217.570 107.185 218.390 ;
        RECT 0.100 217.550 107.185 217.570 ;
        RECT 0.100 216.730 106.910 217.550 ;
        RECT 0.100 215.870 107.185 216.730 ;
        RECT 0.100 215.050 106.910 215.870 ;
        RECT 0.100 215.030 107.185 215.050 ;
        RECT 0.610 214.210 107.185 215.030 ;
        RECT 0.100 214.190 107.185 214.210 ;
        RECT 0.100 213.370 106.910 214.190 ;
        RECT 0.100 212.510 107.185 213.370 ;
        RECT 0.100 211.690 106.910 212.510 ;
        RECT 0.100 211.670 107.185 211.690 ;
        RECT 0.610 210.850 107.185 211.670 ;
        RECT 0.100 210.830 107.185 210.850 ;
        RECT 0.100 210.010 106.910 210.830 ;
        RECT 0.100 209.150 107.185 210.010 ;
        RECT 0.100 208.330 106.910 209.150 ;
        RECT 0.100 208.310 107.185 208.330 ;
        RECT 0.610 207.490 107.185 208.310 ;
        RECT 0.100 207.470 107.185 207.490 ;
        RECT 0.100 206.650 106.910 207.470 ;
        RECT 0.100 205.790 107.185 206.650 ;
        RECT 0.100 204.970 106.910 205.790 ;
        RECT 0.100 204.950 107.185 204.970 ;
        RECT 0.610 204.130 107.185 204.950 ;
        RECT 0.100 204.110 107.185 204.130 ;
        RECT 0.100 203.290 106.910 204.110 ;
        RECT 0.100 202.430 107.185 203.290 ;
        RECT 0.100 201.610 106.910 202.430 ;
        RECT 0.100 201.590 107.185 201.610 ;
        RECT 0.610 200.770 107.185 201.590 ;
        RECT 0.100 200.750 107.185 200.770 ;
        RECT 0.100 199.930 106.910 200.750 ;
        RECT 0.100 199.070 107.185 199.930 ;
        RECT 0.100 198.250 106.910 199.070 ;
        RECT 0.100 198.230 107.185 198.250 ;
        RECT 0.610 197.410 107.185 198.230 ;
        RECT 0.100 197.390 107.185 197.410 ;
        RECT 0.100 196.570 106.910 197.390 ;
        RECT 0.100 195.710 107.185 196.570 ;
        RECT 0.100 194.890 106.910 195.710 ;
        RECT 0.100 194.870 107.185 194.890 ;
        RECT 0.610 194.050 107.185 194.870 ;
        RECT 0.100 194.030 107.185 194.050 ;
        RECT 0.100 193.210 106.910 194.030 ;
        RECT 0.100 192.350 107.185 193.210 ;
        RECT 0.100 191.530 106.910 192.350 ;
        RECT 0.100 191.510 107.185 191.530 ;
        RECT 0.610 190.690 107.185 191.510 ;
        RECT 0.100 190.670 107.185 190.690 ;
        RECT 0.100 189.850 106.910 190.670 ;
        RECT 0.100 188.990 107.185 189.850 ;
        RECT 0.100 188.170 106.910 188.990 ;
        RECT 0.100 188.150 107.185 188.170 ;
        RECT 0.610 187.330 107.185 188.150 ;
        RECT 0.100 187.310 107.185 187.330 ;
        RECT 0.100 186.490 106.910 187.310 ;
        RECT 0.100 185.630 107.185 186.490 ;
        RECT 0.100 184.810 106.910 185.630 ;
        RECT 0.100 184.790 107.185 184.810 ;
        RECT 0.610 183.970 107.185 184.790 ;
        RECT 0.100 183.950 107.185 183.970 ;
        RECT 0.100 183.130 106.910 183.950 ;
        RECT 0.100 182.270 107.185 183.130 ;
        RECT 0.100 181.450 106.910 182.270 ;
        RECT 0.100 181.430 107.185 181.450 ;
        RECT 0.610 180.610 107.185 181.430 ;
        RECT 0.100 180.590 107.185 180.610 ;
        RECT 0.100 179.770 106.910 180.590 ;
        RECT 0.100 178.910 107.185 179.770 ;
        RECT 0.100 178.090 106.910 178.910 ;
        RECT 0.100 178.070 107.185 178.090 ;
        RECT 0.610 177.250 107.185 178.070 ;
        RECT 0.100 177.230 107.185 177.250 ;
        RECT 0.100 176.410 106.910 177.230 ;
        RECT 0.100 175.550 107.185 176.410 ;
        RECT 0.100 174.730 106.910 175.550 ;
        RECT 0.100 174.710 107.185 174.730 ;
        RECT 0.610 173.890 107.185 174.710 ;
        RECT 0.100 173.870 107.185 173.890 ;
        RECT 0.100 173.050 106.910 173.870 ;
        RECT 0.100 172.190 107.185 173.050 ;
        RECT 0.100 171.370 106.910 172.190 ;
        RECT 0.100 171.350 107.185 171.370 ;
        RECT 0.610 170.530 107.185 171.350 ;
        RECT 0.100 170.510 107.185 170.530 ;
        RECT 0.100 169.690 106.910 170.510 ;
        RECT 0.100 168.830 107.185 169.690 ;
        RECT 0.100 168.010 106.910 168.830 ;
        RECT 0.100 167.990 107.185 168.010 ;
        RECT 0.610 167.170 107.185 167.990 ;
        RECT 0.100 167.150 107.185 167.170 ;
        RECT 0.100 166.330 106.910 167.150 ;
        RECT 0.100 165.470 107.185 166.330 ;
        RECT 0.100 164.650 106.910 165.470 ;
        RECT 0.100 164.630 107.185 164.650 ;
        RECT 0.610 163.810 107.185 164.630 ;
        RECT 0.100 163.790 107.185 163.810 ;
        RECT 0.100 162.970 106.910 163.790 ;
        RECT 0.100 162.110 107.185 162.970 ;
        RECT 0.100 161.290 106.910 162.110 ;
        RECT 0.100 161.270 107.185 161.290 ;
        RECT 0.610 160.450 107.185 161.270 ;
        RECT 0.100 160.430 107.185 160.450 ;
        RECT 0.100 159.610 106.910 160.430 ;
        RECT 0.100 158.750 107.185 159.610 ;
        RECT 0.100 157.930 106.910 158.750 ;
        RECT 0.100 157.910 107.185 157.930 ;
        RECT 0.610 157.090 107.185 157.910 ;
        RECT 0.100 157.070 107.185 157.090 ;
        RECT 0.100 156.250 106.910 157.070 ;
        RECT 0.100 155.390 107.185 156.250 ;
        RECT 0.100 154.570 106.910 155.390 ;
        RECT 0.100 154.550 107.185 154.570 ;
        RECT 0.610 153.730 107.185 154.550 ;
        RECT 0.100 153.710 107.185 153.730 ;
        RECT 0.100 152.890 106.910 153.710 ;
        RECT 0.100 152.030 107.185 152.890 ;
        RECT 0.100 151.210 106.910 152.030 ;
        RECT 0.100 151.190 107.185 151.210 ;
        RECT 0.610 150.370 107.185 151.190 ;
        RECT 0.100 150.350 107.185 150.370 ;
        RECT 0.100 149.530 106.910 150.350 ;
        RECT 0.100 148.670 107.185 149.530 ;
        RECT 0.100 147.850 106.910 148.670 ;
        RECT 0.100 147.830 107.185 147.850 ;
        RECT 0.610 147.010 107.185 147.830 ;
        RECT 0.100 146.990 107.185 147.010 ;
        RECT 0.100 146.170 106.910 146.990 ;
        RECT 0.100 145.310 107.185 146.170 ;
        RECT 0.100 144.490 106.910 145.310 ;
        RECT 0.100 144.470 107.185 144.490 ;
        RECT 0.610 143.650 107.185 144.470 ;
        RECT 0.100 143.630 107.185 143.650 ;
        RECT 0.100 142.810 106.910 143.630 ;
        RECT 0.100 141.950 107.185 142.810 ;
        RECT 0.100 141.130 106.910 141.950 ;
        RECT 0.100 141.110 107.185 141.130 ;
        RECT 0.610 140.290 107.185 141.110 ;
        RECT 0.100 140.270 107.185 140.290 ;
        RECT 0.100 139.450 106.910 140.270 ;
        RECT 0.100 138.590 107.185 139.450 ;
        RECT 0.100 137.770 106.910 138.590 ;
        RECT 0.100 137.750 107.185 137.770 ;
        RECT 0.610 136.930 107.185 137.750 ;
        RECT 0.100 136.910 107.185 136.930 ;
        RECT 0.100 136.090 106.910 136.910 ;
        RECT 0.100 135.230 107.185 136.090 ;
        RECT 0.100 134.410 106.910 135.230 ;
        RECT 0.100 134.390 107.185 134.410 ;
        RECT 0.610 133.570 107.185 134.390 ;
        RECT 0.100 133.550 107.185 133.570 ;
        RECT 0.100 132.730 106.910 133.550 ;
        RECT 0.100 131.870 107.185 132.730 ;
        RECT 0.100 131.050 106.910 131.870 ;
        RECT 0.100 131.030 107.185 131.050 ;
        RECT 0.610 130.210 107.185 131.030 ;
        RECT 0.100 130.190 107.185 130.210 ;
        RECT 0.100 129.370 106.910 130.190 ;
        RECT 0.100 128.510 107.185 129.370 ;
        RECT 0.100 127.690 106.910 128.510 ;
        RECT 0.100 127.670 107.185 127.690 ;
        RECT 0.610 126.850 107.185 127.670 ;
        RECT 0.100 126.830 107.185 126.850 ;
        RECT 0.100 126.010 106.910 126.830 ;
        RECT 0.100 125.150 107.185 126.010 ;
        RECT 0.100 124.330 106.910 125.150 ;
        RECT 0.100 124.310 107.185 124.330 ;
        RECT 0.610 123.490 107.185 124.310 ;
        RECT 0.100 123.470 107.185 123.490 ;
        RECT 0.100 122.650 106.910 123.470 ;
        RECT 0.100 121.790 107.185 122.650 ;
        RECT 0.100 120.970 106.910 121.790 ;
        RECT 0.100 120.950 107.185 120.970 ;
        RECT 0.610 120.130 107.185 120.950 ;
        RECT 0.100 120.110 107.185 120.130 ;
        RECT 0.100 119.290 106.910 120.110 ;
        RECT 0.100 118.430 107.185 119.290 ;
        RECT 0.100 117.610 106.910 118.430 ;
        RECT 0.100 117.590 107.185 117.610 ;
        RECT 0.610 116.770 107.185 117.590 ;
        RECT 0.100 116.750 107.185 116.770 ;
        RECT 0.100 115.930 106.910 116.750 ;
        RECT 0.100 115.070 107.185 115.930 ;
        RECT 0.100 114.250 106.910 115.070 ;
        RECT 0.100 114.230 107.185 114.250 ;
        RECT 0.610 113.410 107.185 114.230 ;
        RECT 0.100 113.390 107.185 113.410 ;
        RECT 0.100 112.570 106.910 113.390 ;
        RECT 0.100 111.710 107.185 112.570 ;
        RECT 0.100 110.890 106.910 111.710 ;
        RECT 0.100 110.870 107.185 110.890 ;
        RECT 0.610 110.050 107.185 110.870 ;
        RECT 0.100 110.030 107.185 110.050 ;
        RECT 0.100 109.210 106.910 110.030 ;
        RECT 0.100 108.350 107.185 109.210 ;
        RECT 0.100 107.530 106.910 108.350 ;
        RECT 0.100 107.510 107.185 107.530 ;
        RECT 0.610 106.690 107.185 107.510 ;
        RECT 0.100 106.670 107.185 106.690 ;
        RECT 0.100 105.850 106.910 106.670 ;
        RECT 0.100 104.990 107.185 105.850 ;
        RECT 0.100 104.170 106.910 104.990 ;
        RECT 0.100 104.150 107.185 104.170 ;
        RECT 0.610 103.330 107.185 104.150 ;
        RECT 0.100 103.310 107.185 103.330 ;
        RECT 0.100 102.490 106.910 103.310 ;
        RECT 0.100 101.630 107.185 102.490 ;
        RECT 0.100 100.810 106.910 101.630 ;
        RECT 0.100 100.790 107.185 100.810 ;
        RECT 0.610 99.970 107.185 100.790 ;
        RECT 0.100 99.950 107.185 99.970 ;
        RECT 0.100 99.130 106.910 99.950 ;
        RECT 0.100 98.270 107.185 99.130 ;
        RECT 0.100 97.450 106.910 98.270 ;
        RECT 0.100 97.430 107.185 97.450 ;
        RECT 0.610 96.610 107.185 97.430 ;
        RECT 0.100 96.590 107.185 96.610 ;
        RECT 0.100 95.770 106.910 96.590 ;
        RECT 0.100 94.910 107.185 95.770 ;
        RECT 0.100 94.090 106.910 94.910 ;
        RECT 0.100 94.070 107.185 94.090 ;
        RECT 0.610 93.250 107.185 94.070 ;
        RECT 0.100 93.230 107.185 93.250 ;
        RECT 0.100 92.410 106.910 93.230 ;
        RECT 0.100 91.550 107.185 92.410 ;
        RECT 0.100 90.730 106.910 91.550 ;
        RECT 0.100 90.710 107.185 90.730 ;
        RECT 0.610 89.890 107.185 90.710 ;
        RECT 0.100 89.870 107.185 89.890 ;
        RECT 0.100 89.050 106.910 89.870 ;
        RECT 0.100 88.190 107.185 89.050 ;
        RECT 0.100 87.370 106.910 88.190 ;
        RECT 0.100 87.350 107.185 87.370 ;
        RECT 0.610 86.530 107.185 87.350 ;
        RECT 0.100 86.510 107.185 86.530 ;
        RECT 0.100 85.690 106.910 86.510 ;
        RECT 0.100 84.830 107.185 85.690 ;
        RECT 0.100 84.010 106.910 84.830 ;
        RECT 0.100 83.990 107.185 84.010 ;
        RECT 0.610 83.170 107.185 83.990 ;
        RECT 0.100 83.150 107.185 83.170 ;
        RECT 0.100 82.330 106.910 83.150 ;
        RECT 0.100 81.470 107.185 82.330 ;
        RECT 0.100 80.650 106.910 81.470 ;
        RECT 0.100 80.630 107.185 80.650 ;
        RECT 0.610 79.810 107.185 80.630 ;
        RECT 0.100 79.790 107.185 79.810 ;
        RECT 0.100 78.970 106.910 79.790 ;
        RECT 0.100 78.110 107.185 78.970 ;
        RECT 0.100 77.290 106.910 78.110 ;
        RECT 0.100 77.270 107.185 77.290 ;
        RECT 0.610 76.450 107.185 77.270 ;
        RECT 0.100 76.430 107.185 76.450 ;
        RECT 0.100 75.610 106.910 76.430 ;
        RECT 0.100 74.750 107.185 75.610 ;
        RECT 0.100 73.930 106.910 74.750 ;
        RECT 0.100 73.910 107.185 73.930 ;
        RECT 0.610 73.090 107.185 73.910 ;
        RECT 0.100 73.070 107.185 73.090 ;
        RECT 0.100 72.250 106.910 73.070 ;
        RECT 0.100 71.390 107.185 72.250 ;
        RECT 0.100 70.570 106.910 71.390 ;
        RECT 0.100 70.550 107.185 70.570 ;
        RECT 0.610 69.730 107.185 70.550 ;
        RECT 0.100 69.710 107.185 69.730 ;
        RECT 0.100 68.890 106.910 69.710 ;
        RECT 0.100 68.030 107.185 68.890 ;
        RECT 0.100 67.210 106.910 68.030 ;
        RECT 0.100 67.190 107.185 67.210 ;
        RECT 0.610 66.370 107.185 67.190 ;
        RECT 0.100 66.350 107.185 66.370 ;
        RECT 0.100 65.530 106.910 66.350 ;
        RECT 0.100 64.670 107.185 65.530 ;
        RECT 0.100 63.850 106.910 64.670 ;
        RECT 0.100 63.830 107.185 63.850 ;
        RECT 0.610 63.010 107.185 63.830 ;
        RECT 0.100 62.990 107.185 63.010 ;
        RECT 0.100 62.170 106.910 62.990 ;
        RECT 0.100 61.310 107.185 62.170 ;
        RECT 0.100 60.490 106.910 61.310 ;
        RECT 0.100 60.470 107.185 60.490 ;
        RECT 0.610 59.650 107.185 60.470 ;
        RECT 0.100 59.630 107.185 59.650 ;
        RECT 0.100 58.810 106.910 59.630 ;
        RECT 0.100 57.950 107.185 58.810 ;
        RECT 0.100 57.130 106.910 57.950 ;
        RECT 0.100 57.110 107.185 57.130 ;
        RECT 0.610 56.290 107.185 57.110 ;
        RECT 0.100 56.270 107.185 56.290 ;
        RECT 0.100 55.450 106.910 56.270 ;
        RECT 0.100 54.590 107.185 55.450 ;
        RECT 0.100 53.770 106.910 54.590 ;
        RECT 0.100 53.750 107.185 53.770 ;
        RECT 0.610 52.930 107.185 53.750 ;
        RECT 0.100 52.910 107.185 52.930 ;
        RECT 0.100 52.090 106.910 52.910 ;
        RECT 0.100 51.230 107.185 52.090 ;
        RECT 0.100 50.410 106.910 51.230 ;
        RECT 0.100 50.390 107.185 50.410 ;
        RECT 0.610 49.570 107.185 50.390 ;
        RECT 0.100 49.550 107.185 49.570 ;
        RECT 0.100 48.730 106.910 49.550 ;
        RECT 0.100 47.870 107.185 48.730 ;
        RECT 0.100 47.050 106.910 47.870 ;
        RECT 0.100 47.030 107.185 47.050 ;
        RECT 0.610 46.210 107.185 47.030 ;
        RECT 0.100 46.190 107.185 46.210 ;
        RECT 0.100 45.370 106.910 46.190 ;
        RECT 0.100 44.510 107.185 45.370 ;
        RECT 0.100 43.690 106.910 44.510 ;
        RECT 0.100 43.670 107.185 43.690 ;
        RECT 0.610 42.850 107.185 43.670 ;
        RECT 0.100 42.830 107.185 42.850 ;
        RECT 0.100 42.010 106.910 42.830 ;
        RECT 0.100 41.150 107.185 42.010 ;
        RECT 0.100 40.330 106.910 41.150 ;
        RECT 0.100 40.310 107.185 40.330 ;
        RECT 0.610 39.490 107.185 40.310 ;
        RECT 0.100 39.470 107.185 39.490 ;
        RECT 0.100 38.650 106.910 39.470 ;
        RECT 0.100 37.790 107.185 38.650 ;
        RECT 0.100 36.970 106.910 37.790 ;
        RECT 0.100 36.950 107.185 36.970 ;
        RECT 0.610 36.130 107.185 36.950 ;
        RECT 0.100 36.110 107.185 36.130 ;
        RECT 0.100 35.290 106.910 36.110 ;
        RECT 0.100 34.430 107.185 35.290 ;
        RECT 0.100 33.610 106.910 34.430 ;
        RECT 0.100 32.750 107.185 33.610 ;
        RECT 0.100 31.930 106.910 32.750 ;
        RECT 0.100 31.070 107.185 31.930 ;
        RECT 0.100 30.250 106.910 31.070 ;
        RECT 0.100 29.390 107.185 30.250 ;
        RECT 0.100 28.570 106.910 29.390 ;
        RECT 0.100 27.710 107.185 28.570 ;
        RECT 0.100 26.890 106.910 27.710 ;
        RECT 0.100 26.030 107.185 26.890 ;
        RECT 0.100 25.210 106.910 26.030 ;
        RECT 0.100 24.350 107.185 25.210 ;
        RECT 0.100 23.530 106.910 24.350 ;
        RECT 0.100 22.670 107.185 23.530 ;
        RECT 0.100 21.850 106.910 22.670 ;
        RECT 0.100 20.990 107.185 21.850 ;
        RECT 0.100 20.170 106.910 20.990 ;
        RECT 0.100 19.310 107.185 20.170 ;
        RECT 0.100 18.490 106.910 19.310 ;
        RECT 0.100 17.630 107.185 18.490 ;
        RECT 0.100 16.810 106.910 17.630 ;
        RECT 0.100 15.950 107.185 16.810 ;
        RECT 0.100 15.130 106.910 15.950 ;
        RECT 0.100 14.270 107.185 15.130 ;
        RECT 0.100 13.450 106.910 14.270 ;
        RECT 0.100 12.590 107.185 13.450 ;
        RECT 0.100 11.770 106.910 12.590 ;
        RECT 0.100 10.910 107.185 11.770 ;
        RECT 0.100 10.090 106.910 10.910 ;
        RECT 0.100 9.230 107.185 10.090 ;
        RECT 0.100 8.410 106.910 9.230 ;
        RECT 0.100 7.550 107.185 8.410 ;
        RECT 0.100 6.730 106.910 7.550 ;
        RECT 0.100 5.870 107.185 6.730 ;
        RECT 0.100 5.050 106.910 5.870 ;
        RECT 0.100 4.190 107.185 5.050 ;
        RECT 0.100 3.370 106.910 4.190 ;
        RECT 0.100 2.510 107.185 3.370 ;
        RECT 0.100 1.690 106.910 2.510 ;
        RECT 0.100 0.830 107.185 1.690 ;
        RECT 0.100 0.315 106.910 0.830 ;
      LAYER Metal4 ;
        RECT 0.375 0.270 107.140 429.805 ;
      LAYER Metal5 ;
        RECT 0.335 0.320 104.305 429.760 ;
      LAYER TopMetal1 ;
        RECT 5.380 0.020 16.620 430.060 ;
        RECT 22.100 0.020 22.820 430.060 ;
        RECT 28.300 0.020 86.820 430.060 ;
  END
END W_TT_IF2
END LIBRARY

