* NGSPICE file created from E_TT_IF2.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

.subckt E_TT_IF2 CLK_TT_PROJECT ENA_TT_PROJECT RST_N_TT_PROJECT Tile_X0Y0_E1END[0]
+ Tile_X0Y0_E1END[1] Tile_X0Y0_E1END[2] Tile_X0Y0_E1END[3] Tile_X0Y0_E2END[0] Tile_X0Y0_E2END[1]
+ Tile_X0Y0_E2END[2] Tile_X0Y0_E2END[3] Tile_X0Y0_E2END[4] Tile_X0Y0_E2END[5] Tile_X0Y0_E2END[6]
+ Tile_X0Y0_E2END[7] Tile_X0Y0_E2MID[0] Tile_X0Y0_E2MID[1] Tile_X0Y0_E2MID[2] Tile_X0Y0_E2MID[3]
+ Tile_X0Y0_E2MID[4] Tile_X0Y0_E2MID[5] Tile_X0Y0_E2MID[6] Tile_X0Y0_E2MID[7] Tile_X0Y0_E6END[0]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E6END[11] Tile_X0Y0_E6END[1] Tile_X0Y0_E6END[2] Tile_X0Y0_E6END[3]
+ Tile_X0Y0_E6END[4] Tile_X0Y0_E6END[5] Tile_X0Y0_E6END[6] Tile_X0Y0_E6END[7] Tile_X0Y0_E6END[8]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_EE4END[0] Tile_X0Y0_EE4END[10] Tile_X0Y0_EE4END[11]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_EE4END[13] Tile_X0Y0_EE4END[14] Tile_X0Y0_EE4END[15]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_EE4END[2] Tile_X0Y0_EE4END[3] Tile_X0Y0_EE4END[4]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_EE4END[6] Tile_X0Y0_EE4END[7] Tile_X0Y0_EE4END[8]
+ Tile_X0Y0_EE4END[9] Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData[11]
+ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData[15]
+ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData[19]
+ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData[22]
+ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData[26]
+ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData[2]
+ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData[4]
+ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData[8]
+ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[0] Tile_X0Y0_FrameData_O[10] Tile_X0Y0_FrameData_O[11]
+ Tile_X0Y0_FrameData_O[12] Tile_X0Y0_FrameData_O[13] Tile_X0Y0_FrameData_O[14] Tile_X0Y0_FrameData_O[15]
+ Tile_X0Y0_FrameData_O[16] Tile_X0Y0_FrameData_O[17] Tile_X0Y0_FrameData_O[18] Tile_X0Y0_FrameData_O[19]
+ Tile_X0Y0_FrameData_O[1] Tile_X0Y0_FrameData_O[20] Tile_X0Y0_FrameData_O[21] Tile_X0Y0_FrameData_O[22]
+ Tile_X0Y0_FrameData_O[23] Tile_X0Y0_FrameData_O[24] Tile_X0Y0_FrameData_O[25] Tile_X0Y0_FrameData_O[26]
+ Tile_X0Y0_FrameData_O[27] Tile_X0Y0_FrameData_O[28] Tile_X0Y0_FrameData_O[29] Tile_X0Y0_FrameData_O[2]
+ Tile_X0Y0_FrameData_O[30] Tile_X0Y0_FrameData_O[31] Tile_X0Y0_FrameData_O[3] Tile_X0Y0_FrameData_O[4]
+ Tile_X0Y0_FrameData_O[5] Tile_X0Y0_FrameData_O[6] Tile_X0Y0_FrameData_O[7] Tile_X0Y0_FrameData_O[8]
+ Tile_X0Y0_FrameData_O[9] Tile_X0Y0_FrameStrobe_O[0] Tile_X0Y0_FrameStrobe_O[10]
+ Tile_X0Y0_FrameStrobe_O[11] Tile_X0Y0_FrameStrobe_O[12] Tile_X0Y0_FrameStrobe_O[13]
+ Tile_X0Y0_FrameStrobe_O[14] Tile_X0Y0_FrameStrobe_O[15] Tile_X0Y0_FrameStrobe_O[16]
+ Tile_X0Y0_FrameStrobe_O[17] Tile_X0Y0_FrameStrobe_O[18] Tile_X0Y0_FrameStrobe_O[19]
+ Tile_X0Y0_FrameStrobe_O[1] Tile_X0Y0_FrameStrobe_O[2] Tile_X0Y0_FrameStrobe_O[3]
+ Tile_X0Y0_FrameStrobe_O[4] Tile_X0Y0_FrameStrobe_O[5] Tile_X0Y0_FrameStrobe_O[6]
+ Tile_X0Y0_FrameStrobe_O[7] Tile_X0Y0_FrameStrobe_O[8] Tile_X0Y0_FrameStrobe_O[9]
+ Tile_X0Y0_N1BEG[0] Tile_X0Y0_N1BEG[1] Tile_X0Y0_N1BEG[2] Tile_X0Y0_N1BEG[3] Tile_X0Y0_N2BEG[0]
+ Tile_X0Y0_N2BEG[1] Tile_X0Y0_N2BEG[2] Tile_X0Y0_N2BEG[3] Tile_X0Y0_N2BEG[4] Tile_X0Y0_N2BEG[5]
+ Tile_X0Y0_N2BEG[6] Tile_X0Y0_N2BEG[7] Tile_X0Y0_N2BEGb[0] Tile_X0Y0_N2BEGb[1] Tile_X0Y0_N2BEGb[2]
+ Tile_X0Y0_N2BEGb[3] Tile_X0Y0_N2BEGb[4] Tile_X0Y0_N2BEGb[5] Tile_X0Y0_N2BEGb[6]
+ Tile_X0Y0_N2BEGb[7] Tile_X0Y0_N4BEG[0] Tile_X0Y0_N4BEG[10] Tile_X0Y0_N4BEG[11] Tile_X0Y0_N4BEG[12]
+ Tile_X0Y0_N4BEG[13] Tile_X0Y0_N4BEG[14] Tile_X0Y0_N4BEG[15] Tile_X0Y0_N4BEG[1] Tile_X0Y0_N4BEG[2]
+ Tile_X0Y0_N4BEG[3] Tile_X0Y0_N4BEG[4] Tile_X0Y0_N4BEG[5] Tile_X0Y0_N4BEG[6] Tile_X0Y0_N4BEG[7]
+ Tile_X0Y0_N4BEG[8] Tile_X0Y0_N4BEG[9] Tile_X0Y0_S1END[0] Tile_X0Y0_S1END[1] Tile_X0Y0_S1END[2]
+ Tile_X0Y0_S1END[3] Tile_X0Y0_S2END[0] Tile_X0Y0_S2END[1] Tile_X0Y0_S2END[2] Tile_X0Y0_S2END[3]
+ Tile_X0Y0_S2END[4] Tile_X0Y0_S2END[5] Tile_X0Y0_S2END[6] Tile_X0Y0_S2END[7] Tile_X0Y0_S2MID[0]
+ Tile_X0Y0_S2MID[1] Tile_X0Y0_S2MID[2] Tile_X0Y0_S2MID[3] Tile_X0Y0_S2MID[4] Tile_X0Y0_S2MID[5]
+ Tile_X0Y0_S2MID[6] Tile_X0Y0_S2MID[7] Tile_X0Y0_S4END[0] Tile_X0Y0_S4END[10] Tile_X0Y0_S4END[11]
+ Tile_X0Y0_S4END[12] Tile_X0Y0_S4END[13] Tile_X0Y0_S4END[14] Tile_X0Y0_S4END[15]
+ Tile_X0Y0_S4END[1] Tile_X0Y0_S4END[2] Tile_X0Y0_S4END[3] Tile_X0Y0_S4END[4] Tile_X0Y0_S4END[5]
+ Tile_X0Y0_S4END[6] Tile_X0Y0_S4END[7] Tile_X0Y0_S4END[8] Tile_X0Y0_S4END[9] Tile_X0Y0_UserCLKo
+ Tile_X0Y0_W1BEG[0] Tile_X0Y0_W1BEG[1] Tile_X0Y0_W1BEG[2] Tile_X0Y0_W1BEG[3] Tile_X0Y0_W2BEG[0]
+ Tile_X0Y0_W2BEG[1] Tile_X0Y0_W2BEG[2] Tile_X0Y0_W2BEG[3] Tile_X0Y0_W2BEG[4] Tile_X0Y0_W2BEG[5]
+ Tile_X0Y0_W2BEG[6] Tile_X0Y0_W2BEG[7] Tile_X0Y0_W2BEGb[0] Tile_X0Y0_W2BEGb[1] Tile_X0Y0_W2BEGb[2]
+ Tile_X0Y0_W2BEGb[3] Tile_X0Y0_W2BEGb[4] Tile_X0Y0_W2BEGb[5] Tile_X0Y0_W2BEGb[6]
+ Tile_X0Y0_W2BEGb[7] Tile_X0Y0_W6BEG[0] Tile_X0Y0_W6BEG[10] Tile_X0Y0_W6BEG[11] Tile_X0Y0_W6BEG[1]
+ Tile_X0Y0_W6BEG[2] Tile_X0Y0_W6BEG[3] Tile_X0Y0_W6BEG[4] Tile_X0Y0_W6BEG[5] Tile_X0Y0_W6BEG[6]
+ Tile_X0Y0_W6BEG[7] Tile_X0Y0_W6BEG[8] Tile_X0Y0_W6BEG[9] Tile_X0Y0_WW4BEG[0] Tile_X0Y0_WW4BEG[10]
+ Tile_X0Y0_WW4BEG[11] Tile_X0Y0_WW4BEG[12] Tile_X0Y0_WW4BEG[13] Tile_X0Y0_WW4BEG[14]
+ Tile_X0Y0_WW4BEG[15] Tile_X0Y0_WW4BEG[1] Tile_X0Y0_WW4BEG[2] Tile_X0Y0_WW4BEG[3]
+ Tile_X0Y0_WW4BEG[4] Tile_X0Y0_WW4BEG[5] Tile_X0Y0_WW4BEG[6] Tile_X0Y0_WW4BEG[7]
+ Tile_X0Y0_WW4BEG[8] Tile_X0Y0_WW4BEG[9] Tile_X0Y1_E1END[0] Tile_X0Y1_E1END[1] Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E1END[3] Tile_X0Y1_E2END[0] Tile_X0Y1_E2END[1] Tile_X0Y1_E2END[2] Tile_X0Y1_E2END[3]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E2END[5] Tile_X0Y1_E2END[6] Tile_X0Y1_E2END[7] Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2MID[1] Tile_X0Y1_E2MID[2] Tile_X0Y1_E2MID[3] Tile_X0Y1_E2MID[4] Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2MID[6] Tile_X0Y1_E2MID[7] Tile_X0Y1_E6END[0] Tile_X0Y1_E6END[10] Tile_X0Y1_E6END[11]
+ Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[3] Tile_X0Y1_E6END[4] Tile_X0Y1_E6END[5]
+ Tile_X0Y1_E6END[6] Tile_X0Y1_E6END[7] Tile_X0Y1_E6END[8] Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_EE4END[10] Tile_X0Y1_EE4END[11] Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[13]
+ Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[15] Tile_X0Y1_EE4END[1] Tile_X0Y1_EE4END[2]
+ Tile_X0Y1_EE4END[3] Tile_X0Y1_EE4END[4] Tile_X0Y1_EE4END[5] Tile_X0Y1_EE4END[6]
+ Tile_X0Y1_EE4END[7] Tile_X0Y1_EE4END[8] Tile_X0Y1_EE4END[9] Tile_X0Y1_FrameData[0]
+ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData[13]
+ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData[17]
+ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData[20]
+ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData[24]
+ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData[28]
+ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData[31]
+ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData[6]
+ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[0]
+ Tile_X0Y1_FrameData_O[10] Tile_X0Y1_FrameData_O[11] Tile_X0Y1_FrameData_O[12] Tile_X0Y1_FrameData_O[13]
+ Tile_X0Y1_FrameData_O[14] Tile_X0Y1_FrameData_O[15] Tile_X0Y1_FrameData_O[16] Tile_X0Y1_FrameData_O[17]
+ Tile_X0Y1_FrameData_O[18] Tile_X0Y1_FrameData_O[19] Tile_X0Y1_FrameData_O[1] Tile_X0Y1_FrameData_O[20]
+ Tile_X0Y1_FrameData_O[21] Tile_X0Y1_FrameData_O[22] Tile_X0Y1_FrameData_O[23] Tile_X0Y1_FrameData_O[24]
+ Tile_X0Y1_FrameData_O[25] Tile_X0Y1_FrameData_O[26] Tile_X0Y1_FrameData_O[27] Tile_X0Y1_FrameData_O[28]
+ Tile_X0Y1_FrameData_O[29] Tile_X0Y1_FrameData_O[2] Tile_X0Y1_FrameData_O[30] Tile_X0Y1_FrameData_O[31]
+ Tile_X0Y1_FrameData_O[3] Tile_X0Y1_FrameData_O[4] Tile_X0Y1_FrameData_O[5] Tile_X0Y1_FrameData_O[6]
+ Tile_X0Y1_FrameData_O[7] Tile_X0Y1_FrameData_O[8] Tile_X0Y1_FrameData_O[9] Tile_X0Y1_FrameStrobe[0]
+ Tile_X0Y1_FrameStrobe[10] Tile_X0Y1_FrameStrobe[11] Tile_X0Y1_FrameStrobe[12] Tile_X0Y1_FrameStrobe[13]
+ Tile_X0Y1_FrameStrobe[14] Tile_X0Y1_FrameStrobe[15] Tile_X0Y1_FrameStrobe[16] Tile_X0Y1_FrameStrobe[17]
+ Tile_X0Y1_FrameStrobe[18] Tile_X0Y1_FrameStrobe[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_FrameStrobe[2]
+ Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_FrameStrobe[6]
+ Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_FrameStrobe[8] Tile_X0Y1_FrameStrobe[9] Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N1END[1] Tile_X0Y1_N1END[2] Tile_X0Y1_N1END[3] Tile_X0Y1_N2END[0] Tile_X0Y1_N2END[1]
+ Tile_X0Y1_N2END[2] Tile_X0Y1_N2END[3] Tile_X0Y1_N2END[4] Tile_X0Y1_N2END[5] Tile_X0Y1_N2END[6]
+ Tile_X0Y1_N2END[7] Tile_X0Y1_N2MID[0] Tile_X0Y1_N2MID[1] Tile_X0Y1_N2MID[2] Tile_X0Y1_N2MID[3]
+ Tile_X0Y1_N2MID[4] Tile_X0Y1_N2MID[5] Tile_X0Y1_N2MID[6] Tile_X0Y1_N2MID[7] Tile_X0Y1_N4END[0]
+ Tile_X0Y1_N4END[10] Tile_X0Y1_N4END[11] Tile_X0Y1_N4END[12] Tile_X0Y1_N4END[13]
+ Tile_X0Y1_N4END[14] Tile_X0Y1_N4END[15] Tile_X0Y1_N4END[1] Tile_X0Y1_N4END[2] Tile_X0Y1_N4END[3]
+ Tile_X0Y1_N4END[4] Tile_X0Y1_N4END[5] Tile_X0Y1_N4END[6] Tile_X0Y1_N4END[7] Tile_X0Y1_N4END[8]
+ Tile_X0Y1_N4END[9] Tile_X0Y1_S1BEG[0] Tile_X0Y1_S1BEG[1] Tile_X0Y1_S1BEG[2] Tile_X0Y1_S1BEG[3]
+ Tile_X0Y1_S2BEG[0] Tile_X0Y1_S2BEG[1] Tile_X0Y1_S2BEG[2] Tile_X0Y1_S2BEG[3] Tile_X0Y1_S2BEG[4]
+ Tile_X0Y1_S2BEG[5] Tile_X0Y1_S2BEG[6] Tile_X0Y1_S2BEG[7] Tile_X0Y1_S2BEGb[0] Tile_X0Y1_S2BEGb[1]
+ Tile_X0Y1_S2BEGb[2] Tile_X0Y1_S2BEGb[3] Tile_X0Y1_S2BEGb[4] Tile_X0Y1_S2BEGb[5]
+ Tile_X0Y1_S2BEGb[6] Tile_X0Y1_S2BEGb[7] Tile_X0Y1_S4BEG[0] Tile_X0Y1_S4BEG[10] Tile_X0Y1_S4BEG[11]
+ Tile_X0Y1_S4BEG[12] Tile_X0Y1_S4BEG[13] Tile_X0Y1_S4BEG[14] Tile_X0Y1_S4BEG[15]
+ Tile_X0Y1_S4BEG[1] Tile_X0Y1_S4BEG[2] Tile_X0Y1_S4BEG[3] Tile_X0Y1_S4BEG[4] Tile_X0Y1_S4BEG[5]
+ Tile_X0Y1_S4BEG[6] Tile_X0Y1_S4BEG[7] Tile_X0Y1_S4BEG[8] Tile_X0Y1_S4BEG[9] Tile_X0Y1_UserCLK
+ Tile_X0Y1_W1BEG[0] Tile_X0Y1_W1BEG[1] Tile_X0Y1_W1BEG[2] Tile_X0Y1_W1BEG[3] Tile_X0Y1_W2BEG[0]
+ Tile_X0Y1_W2BEG[1] Tile_X0Y1_W2BEG[2] Tile_X0Y1_W2BEG[3] Tile_X0Y1_W2BEG[4] Tile_X0Y1_W2BEG[5]
+ Tile_X0Y1_W2BEG[6] Tile_X0Y1_W2BEG[7] Tile_X0Y1_W2BEGb[0] Tile_X0Y1_W2BEGb[1] Tile_X0Y1_W2BEGb[2]
+ Tile_X0Y1_W2BEGb[3] Tile_X0Y1_W2BEGb[4] Tile_X0Y1_W2BEGb[5] Tile_X0Y1_W2BEGb[6]
+ Tile_X0Y1_W2BEGb[7] Tile_X0Y1_W6BEG[0] Tile_X0Y1_W6BEG[10] Tile_X0Y1_W6BEG[11] Tile_X0Y1_W6BEG[1]
+ Tile_X0Y1_W6BEG[2] Tile_X0Y1_W6BEG[3] Tile_X0Y1_W6BEG[4] Tile_X0Y1_W6BEG[5] Tile_X0Y1_W6BEG[6]
+ Tile_X0Y1_W6BEG[7] Tile_X0Y1_W6BEG[8] Tile_X0Y1_W6BEG[9] Tile_X0Y1_WW4BEG[0] Tile_X0Y1_WW4BEG[10]
+ Tile_X0Y1_WW4BEG[11] Tile_X0Y1_WW4BEG[12] Tile_X0Y1_WW4BEG[13] Tile_X0Y1_WW4BEG[14]
+ Tile_X0Y1_WW4BEG[15] Tile_X0Y1_WW4BEG[1] Tile_X0Y1_WW4BEG[2] Tile_X0Y1_WW4BEG[3]
+ Tile_X0Y1_WW4BEG[4] Tile_X0Y1_WW4BEG[5] Tile_X0Y1_WW4BEG[6] Tile_X0Y1_WW4BEG[7]
+ Tile_X0Y1_WW4BEG[8] Tile_X0Y1_WW4BEG[9] UIO_IN_TT_PROJECT0 UIO_IN_TT_PROJECT1 UIO_IN_TT_PROJECT2
+ UIO_IN_TT_PROJECT3 UIO_IN_TT_PROJECT4 UIO_IN_TT_PROJECT5 UIO_IN_TT_PROJECT6 UIO_IN_TT_PROJECT7
+ UIO_OE_TT_PROJECT0 UIO_OE_TT_PROJECT1 UIO_OE_TT_PROJECT2 UIO_OE_TT_PROJECT3 UIO_OE_TT_PROJECT4
+ UIO_OE_TT_PROJECT5 UIO_OE_TT_PROJECT6 UIO_OE_TT_PROJECT7 UIO_OUT_TT_PROJECT0 UIO_OUT_TT_PROJECT1
+ UIO_OUT_TT_PROJECT2 UIO_OUT_TT_PROJECT3 UIO_OUT_TT_PROJECT4 UIO_OUT_TT_PROJECT5
+ UIO_OUT_TT_PROJECT6 UIO_OUT_TT_PROJECT7 UI_IN_TT_PROJECT0 UI_IN_TT_PROJECT1 UI_IN_TT_PROJECT2
+ UI_IN_TT_PROJECT3 UI_IN_TT_PROJECT4 UI_IN_TT_PROJECT5 UI_IN_TT_PROJECT6 UI_IN_TT_PROJECT7
+ UO_OUT_TT_PROJECT0 UO_OUT_TT_PROJECT1 UO_OUT_TT_PROJECT2 UO_OUT_TT_PROJECT3 UO_OUT_TT_PROJECT4
+ UO_OUT_TT_PROJECT5 UO_OUT_TT_PROJECT6 UO_OUT_TT_PROJECT7 VGND VPWR
XFILLER_36_19 VPWR VGND sg13g2_fill_1
X_0367_ VPWR _0297_ Tile_X0Y1_E6END[3] VGND sg13g2_inv_1
XFILLER_22_188 VPWR VGND sg13g2_decap_8
XFILLER_22_199 VPWR VGND sg13g2_fill_1
XFILLER_13_100 VPWR VGND sg13g2_decap_8
XFILLER_3_23 VPWR VGND sg13g2_fill_2
XFILLER_95_158 VPWR VGND sg13g2_decap_8
XFILLER_95_125 VPWR VGND sg13g2_decap_8
X_1270_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1606_ Tile_X0Y0_S4END[8] Tile_X0Y1_S4BEG[0] VPWR VGND sg13g2_buf_1
X_0985_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1468_ Tile_X0Y1_FrameStrobe[19] Tile_X0Y0_FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_0419_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q Tile_X0Y0_E2MID[6]
+ Tile_X0Y0_E2END[6] Tile_X0Y0_E6END[9] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_86_147 VPWR VGND sg13g2_decap_8
X_1537_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG11 Tile_X0Y0_W6BEG[11]
+ VPWR VGND sg13g2_buf_1
X_1399_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_103_24 VPWR VGND sg13g2_decap_8
XFILLER_77_103 VPWR VGND sg13g2_fill_2
XFILLER_37_40 VPWR VGND sg13g2_fill_1
XFILLER_53_94 VPWR VGND sg13g2_fill_1
XFILLER_5_173 VPWR VGND sg13g2_decap_8
X_0770_ _0162_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q
+ _0163_ VPWR VGND sg13g2_nor2b_1
X_1322_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1253_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1184_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0968_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0899_ VGND VPWR Tile_X0Y1_E2MID[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0275_ _0274_ sg13g2_a21oi_1
XFILLER_74_128 VPWR VGND sg13g2_fill_2
XFILLER_23_31 VPWR VGND sg13g2_fill_1
XFILLER_2_198 VPWR VGND sg13g2_fill_2
XFILLER_2_187 VPWR VGND sg13g2_decap_8
XFILLER_2_121 VPWR VGND sg13g2_fill_1
XFILLER_64_82 VPWR VGND sg13g2_decap_8
XFILLER_0_46 VPWR VGND sg13g2_fill_2
XFILLER_0_79 VPWR VGND sg13g2_fill_2
X_0822_ VGND VPWR Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
+ _0207_ _0208_ _0304_ sg13g2_a21oi_1
X_0684_ _0119_ _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_nand2b_1
X_0753_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q UO_OUT_TT_PROJECT3
+ _0158_ UO_OUT_TT_PROJECT7 _0335_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG15 VPWR VGND sg13g2_mux4_1
X_1305_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_0 VPWR VGND sg13g2_fill_2
X_1236_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1098_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1167_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_85_59 VPWR VGND sg13g2_fill_1
XFILLER_18_64 VPWR VGND sg13g2_fill_2
XFILLER_47_139 VPWR VGND sg13g2_decap_8
XFILLER_55_161 VPWR VGND sg13g2_decap_8
XFILLER_75_70 VPWR VGND sg13g2_decap_4
X_1021_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_46_161 VPWR VGND sg13g2_decap_8
X_0805_ _0153_ _0149_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q
+ _0193_ VPWR VGND sg13g2_mux2_1
X_0598_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q _0065_
+ _0066_ VPWR VGND sg13g2_and2_1
X_0667_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q Tile_X0Y1_E2MID[6]
+ Tile_X0Y1_E2END[6] Tile_X0Y1_E6END[9] _0342_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG1 VPWR VGND sg13g2_mux4_1
X_0736_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0007_ Tile_X0Y0_S4END[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q
+ _0150_ VPWR VGND sg13g2_mux4_1
X_1219_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_161 VPWR VGND sg13g2_fill_2
XFILLER_43_164 VPWR VGND sg13g2_decap_8
XFILLER_45_51 VPWR VGND sg13g2_fill_2
XFILLER_45_95 VPWR VGND sg13g2_fill_1
XANTENNA_5 VPWR VGND Tile_X0Y1_FrameStrobe[13] sg13g2_antennanp
X_0521_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q
+ _0011_ VPWR VGND sg13g2_mux4_1
X_0452_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_E2END[3] Tile_X0Y0_E2MID[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG4
+ VPWR VGND sg13g2_mux4_1
X_1570_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameData_O[16] VPWR VGND sg13g2_buf_1
X_0383_ Tile_X0Y1_N1END[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q _0313_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_96_0 VPWR VGND sg13g2_decap_4
X_1004_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_164 VPWR VGND sg13g2_fill_2
XFILLER_106_68 VPWR VGND sg13g2_decap_8
XFILLER_103_125 VPWR VGND sg13g2_decap_8
XFILLER_66_39 VPWR VGND sg13g2_fill_2
X_0719_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q
+ _0142_ _0141_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb5 _0348_ sg13g2_a221oi_1
XFILLER_17_109 VPWR VGND sg13g2_fill_2
XFILLER_16_120 VPWR VGND sg13g2_decap_4
XFILLER_31_123 VPWR VGND sg13g2_fill_1
XFILLER_31_145 VPWR VGND sg13g2_fill_2
X_1622_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG0 Tile_X0Y1_W1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1484_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb3 Tile_X0Y0_N2BEGb[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_98_134 VPWR VGND sg13g2_decap_8
X_0504_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q UIO_OUT_TT_PROJECT3
+ UIO_OE_TT_PROJECT7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG3 VPWR VGND sg13g2_mux4_1
X_1553_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG15 Tile_X0Y0_WW4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_0435_ _0345_ _0346_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q
+ _0347_ VPWR VGND sg13g2_nand3_1
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_0366_ VPWR _0296_ Tile_X0Y0_S2MID[3] VGND sg13g2_inv_1
XFILLER_22_167 VPWR VGND sg13g2_decap_4
XFILLER_42_85 VPWR VGND sg13g2_decap_8
X_0984_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1536_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG10 Tile_X0Y0_W6BEG[10]
+ VPWR VGND sg13g2_buf_1
XFILLER_8_193 VPWR VGND sg13g2_decap_8
X_1605_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG7 Tile_X0Y1_S2BEGb[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_59_0 VPWR VGND sg13g2_fill_2
X_1467_ Tile_X0Y1_FrameStrobe[18] Tile_X0Y0_FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_0418_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y0_E2MID[7]
+ Tile_X0Y0_E2END[7] Tile_X0Y0_E6END[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG0
+ VPWR VGND sg13g2_mux4_1
X_1398_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_94_192 VPWR VGND sg13g2_decap_8
XFILLER_10_159 VPWR VGND sg13g2_decap_8
XFILLER_83_129 VPWR VGND sg13g2_fill_1
XFILLER_68_115 VPWR VGND sg13g2_fill_2
X_1321_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1252_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1183_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0967_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1519_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb1 Tile_X0Y0_W2BEGb[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_59_126 VPWR VGND sg13g2_fill_1
X_0898_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_N2END[3]
+ _0274_ VPWR VGND sg13g2_nor2b_1
XFILLER_82_195 VPWR VGND sg13g2_decap_4
XFILLER_99_69 VPWR VGND sg13g2_fill_2
XFILLER_65_129 VPWR VGND sg13g2_decap_4
XFILLER_65_107 VPWR VGND sg13g2_fill_1
XFILLER_3_2 VPWR VGND sg13g2_fill_1
XFILLER_2_166 VPWR VGND sg13g2_decap_8
XFILLER_0_36 VPWR VGND sg13g2_decap_4
X_0752_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0007_ Tile_X0Y0_S4END[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q
+ _0158_ VPWR VGND sg13g2_mux4_1
X_0821_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 _0003_
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q _0207_ VPWR
+ VGND sg13g2_mux2_1
X_0683_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q
+ _0118_ _0117_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG1 _0341_ sg13g2_a221oi_1
X_1304_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1235_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1166_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_129 VPWR VGND sg13g2_fill_2
XFILLER_100_26 VPWR VGND sg13g2_decap_8
X_1097_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_184 VPWR VGND sg13g2_fill_1
XFILLER_55_140 VPWR VGND sg13g2_decap_8
XFILLER_70_198 VPWR VGND sg13g2_fill_2
X_1020_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_118 VPWR VGND sg13g2_fill_1
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_61_198 VPWR VGND sg13g2_fill_2
XFILLER_46_184 VPWR VGND sg13g2_fill_1
X_0735_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT6 _0149_ _0342_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG6 VPWR VGND sg13g2_mux4_1
X_0804_ VGND VPWR _0188_ _0190_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG0
+ _0192_ sg13g2_a21oi_1
X_0597_ _0065_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 VPWR VGND sg13g2_nand2b_1
X_0666_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q Tile_X0Y1_E2MID[7]
+ Tile_X0Y1_E2END[7] Tile_X0Y1_E6END[8] _0335_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_41_0 VPWR VGND sg13g2_decap_8
X_1149_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1218_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_176 VPWR VGND sg13g2_decap_8
XFILLER_106_189 VPWR VGND sg13g2_decap_8
XFILLER_106_145 VPWR VGND sg13g2_decap_4
XFILLER_96_26 VPWR VGND sg13g2_decap_8
XFILLER_28_195 VPWR VGND sg13g2_decap_4
XANTENNA_6 VPWR VGND Tile_X0Y1_FrameStrobe[14] sg13g2_antennanp
XFILLER_61_95 VPWR VGND sg13g2_fill_2
X_0451_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q Tile_X0Y0_E2MID[4]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E6END[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG3
+ VPWR VGND sg13g2_mux4_1
X_0520_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q UIO_OUT_TT_PROJECT7
+ UIO_OE_TT_PROJECT3 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG11 VPWR VGND sg13g2_mux4_1
X_0382_ _0312_ _0311_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
X_1003_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_184 VPWR VGND sg13g2_decap_8
XFILLER_89_0 VPWR VGND sg13g2_decap_8
XFILLER_34_198 VPWR VGND sg13g2_fill_2
XFILLER_103_104 VPWR VGND sg13g2_decap_8
X_0718_ UO_OUT_TT_PROJECT5 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q _0142_ VPWR
+ VGND sg13g2_nor3_1
X_0649_ Tile_X0Y0_E6END[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q
+ _0105_ VPWR VGND sg13g2_nor2b_1
XFILLER_25_198 VPWR VGND sg13g2_fill_2
XFILLER_82_7 VPWR VGND sg13g2_decap_8
XFILLER_72_94 VPWR VGND sg13g2_decap_4
XFILLER_72_61 VPWR VGND sg13g2_decap_8
XFILLER_16_198 VPWR VGND sg13g2_fill_2
X_1552_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG14 Tile_X0Y0_WW4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_1621_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG3 Tile_X0Y1_S4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_1483_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb2 Tile_X0Y0_N2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_0503_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_mux4_1
X_0434_ _0346_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y0_S2MID[2] VPWR VGND sg13g2_nand2_1
X_0365_ VPWR _0295_ Tile_X0Y1_E2END[5] VGND sg13g2_inv_1
XFILLER_22_124 VPWR VGND sg13g2_decap_4
XFILLER_89_124 VPWR VGND sg13g2_decap_4
XFILLER_13_168 VPWR VGND sg13g2_decap_4
XFILLER_42_42 VPWR VGND sg13g2_decap_8
X_0983_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_172 VPWR VGND sg13g2_decap_8
X_1535_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG9 Tile_X0Y0_W6BEG[9]
+ VPWR VGND sg13g2_buf_1
X_1604_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG6 Tile_X0Y1_S2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_1466_ Tile_X0Y1_FrameStrobe[17] Tile_X0Y0_FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_0417_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb0
+ Tile_X0Y0_S2MID[0] Tile_X0Y1_N2MID[0] Tile_X0Y0_S2END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_94_171 VPWR VGND sg13g2_decap_8
X_1397_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_12_78 VPWR VGND sg13g2_decap_4
XFILLER_10_127 VPWR VGND sg13g2_decap_8
XFILLER_53_63 VPWR VGND sg13g2_decap_4
X_1320_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1251_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1182_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0966_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_0 VPWR VGND sg13g2_decap_4
X_0897_ VGND VPWR Tile_X0Y1_E2MID[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0273_ _0272_ sg13g2_a21oi_1
X_1449_ Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
X_1518_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb0 Tile_X0Y0_W2BEGb[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_67_171 VPWR VGND sg13g2_decap_4
XFILLER_23_22 VPWR VGND sg13g2_decap_8
XFILLER_23_77 VPWR VGND sg13g2_decap_8
XFILLER_99_37 VPWR VGND sg13g2_fill_1
XFILLER_0_15 VPWR VGND sg13g2_decap_8
XFILLER_58_171 VPWR VGND sg13g2_fill_2
XFILLER_0_48 VPWR VGND sg13g2_fill_1
XFILLER_80_83 VPWR VGND sg13g2_decap_4
X_0751_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT6 _0157_ _0342_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG14 VPWR VGND sg13g2_mux4_1
X_0820_ _0206_ _0205_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_nand2b_1
X_0682_ UO_OUT_TT_PROJECT1 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q _0118_ VPWR
+ VGND sg13g2_nor3_1
X_1303_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_4 VPWR VGND sg13g2_fill_1
X_1096_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1165_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1234_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_193 VPWR VGND sg13g2_decap_8
X_0949_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_66 VPWR VGND sg13g2_fill_1
XFILLER_18_88 VPWR VGND sg13g2_fill_1
XFILLER_34_32 VPWR VGND sg13g2_fill_2
XFILLER_1_0 VPWR VGND sg13g2_fill_2
XFILLER_50_97 VPWR VGND sg13g2_decap_8
XFILLER_59_51 VPWR VGND sg13g2_fill_2
XFILLER_59_84 VPWR VGND sg13g2_fill_1
X_0734_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0311_ Tile_X0Y0_S4END[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q
+ _0149_ VPWR VGND sg13g2_mux4_1
X_0803_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q _0191_
+ _0192_ VPWR VGND sg13g2_nor2_1
X_0665_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_E6END[11] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15
+ _0328_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG3
+ VPWR VGND sg13g2_mux4_1
X_0596_ VPWR _0064_ _0063_ VGND sg13g2_inv_1
XFILLER_34_0 VPWR VGND sg13g2_fill_1
X_1148_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_174 VPWR VGND sg13g2_fill_1
X_1217_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_155 VPWR VGND sg13g2_decap_8
X_1079_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_168 VPWR VGND sg13g2_decap_8
XFILLER_106_124 VPWR VGND sg13g2_decap_8
XFILLER_28_163 VPWR VGND sg13g2_fill_1
XFILLER_28_174 VPWR VGND sg13g2_decap_8
XFILLER_43_199 VPWR VGND sg13g2_fill_1
XFILLER_45_53 VPWR VGND sg13g2_fill_1
XANTENNA_7 VPWR VGND Tile_X0Y1_FrameStrobe[15] sg13g2_antennanp
XFILLER_105_190 VPWR VGND sg13g2_decap_8
X_0450_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb3
+ Tile_X0Y0_S2MID[3] Tile_X0Y1_N2MID[3] Tile_X0Y0_S2END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 VPWR VGND sg13g2_mux4_1
X_0381_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_E6END[9] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13
+ _0310_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q _0311_
+ VPWR VGND sg13g2_mux4_1
X_1002_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_166 VPWR VGND sg13g2_fill_1
X_0648_ VGND VPWR UIO_IN_TT_PROJECT5 _0104_ _0103_ sg13g2_or2_1
X_0717_ _0141_ _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_nand2b_1
X_0579_ _0048_ VPWR _0049_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ _0014_ sg13g2_o21ai_1
XFILLER_15_34 VPWR VGND sg13g2_fill_1
XFILLER_25_177 VPWR VGND sg13g2_decap_8
XFILLER_31_55 VPWR VGND sg13g2_fill_1
XFILLER_102_193 VPWR VGND sg13g2_decap_8
XFILLER_56_41 VPWR VGND sg13g2_decap_8
XFILLER_16_177 VPWR VGND sg13g2_decap_8
XFILLER_31_169 VPWR VGND sg13g2_decap_4
X_1482_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb1 Tile_X0Y0_N2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_1551_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG13 Tile_X0Y0_WW4BEG[13]
+ VPWR VGND sg13g2_buf_1
X_0502_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q UIO_OUT_TT_PROJECT2
+ UIO_OE_TT_PROJECT6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG2 VPWR VGND sg13g2_mux4_1
X_1620_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG2 Tile_X0Y1_S4BEG[14]
+ VPWR VGND sg13g2_buf_1
XFILLER_100_119 VPWR VGND sg13g2_decap_8
XFILLER_98_169 VPWR VGND sg13g2_decap_8
X_0364_ VPWR _0294_ Tile_X0Y0_E6END[11] VGND sg13g2_inv_1
XFILLER_11_2 VPWR VGND sg13g2_fill_1
X_0433_ _0345_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG2 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_101_0 VPWR VGND sg13g2_decap_8
XFILLER_21_191 VPWR VGND sg13g2_decap_8
XFILLER_95_139 VPWR VGND sg13g2_decap_8
XFILLER_67_73 VPWR VGND sg13g2_decap_4
XFILLER_67_40 VPWR VGND sg13g2_decap_8
X_0982_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_12_191 VPWR VGND sg13g2_decap_8
X_1465_ Tile_X0Y1_FrameStrobe[16] Tile_X0Y0_FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
X_1534_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG8 Tile_X0Y0_W6BEG[8]
+ VPWR VGND sg13g2_buf_1
X_1603_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG5 Tile_X0Y1_S2BEGb[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_59_2 VPWR VGND sg13g2_fill_1
X_1396_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_0416_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q Tile_X0Y1_E2MID[7]
+ Tile_X0Y1_E2END[7] Tile_X0Y1_E6END[7] _0335_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb0 VPWR VGND sg13g2_mux4_1
XFILLER_85_183 VPWR VGND sg13g2_decap_8
XFILLER_68_117 VPWR VGND sg13g2_fill_1
XFILLER_5_198 VPWR VGND sg13g2_fill_2
XFILLER_5_187 VPWR VGND sg13g2_decap_8
X_1250_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1181_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0965_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_0 VPWR VGND sg13g2_fill_2
X_0896_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_E2MID[3]
+ _0272_ VPWR VGND sg13g2_nor2b_1
X_1448_ Tile_X0Y0_FrameData[31] Tile_X0Y0_FrameData_O[31] VPWR VGND sg13g2_buf_1
XFILLER_59_117 VPWR VGND sg13g2_decap_4
X_1517_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG7 Tile_X0Y0_W2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1379_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_73_120 VPWR VGND sg13g2_decap_4
X_0750_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0311_ Tile_X0Y0_S4END[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q
+ _0157_ VPWR VGND sg13g2_mux4_1
X_0681_ _0117_ _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_nand2b_1
X_1302_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1233_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1095_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_197 VPWR VGND sg13g2_fill_2
X_1164_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_172 VPWR VGND sg13g2_decap_8
X_0948_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0879_ Tile_X0Y1_E2END[4] Tile_X0Y0_S2MID[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0256_ VPWR VGND sg13g2_mux2_1
XFILLER_70_123 VPWR VGND sg13g2_decap_8
XFILLER_55_175 VPWR VGND sg13g2_decap_4
XFILLER_55_197 VPWR VGND sg13g2_fill_2
XFILLER_109_155 VPWR VGND sg13g2_decap_4
XFILLER_109_100 VPWR VGND sg13g2_decap_4
XFILLER_75_95 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_46_197 VPWR VGND sg13g2_fill_2
X_0802_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_E6END[4] _0158_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
+ _0191_ VPWR VGND sg13g2_mux4_1
X_0733_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q UO_OUT_TT_PROJECT1
+ _0148_ UO_OUT_TT_PROJECT5 _0349_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG5 VPWR VGND sg13g2_mux4_1
X_0664_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14
+ _0321_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG2
+ VPWR VGND sg13g2_mux4_1
X_0595_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q VPWR
+ _0063_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q
+ _0062_ sg13g2_o21ai_1
XFILLER_27_0 VPWR VGND sg13g2_decap_4
XFILLER_37_131 VPWR VGND sg13g2_decap_8
X_1216_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1147_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1078_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_112 VPWR VGND sg13g2_decap_8
XFILLER_52_134 VPWR VGND sg13g2_decap_8
XFILLER_106_103 VPWR VGND sg13g2_decap_8
XFILLER_20_68 VPWR VGND sg13g2_decap_8
XFILLER_61_31 VPWR VGND sg13g2_decap_8
XFILLER_43_178 VPWR VGND sg13g2_decap_8
XANTENNA_8 VPWR VGND Tile_X0Y1_FrameStrobe[16] sg13g2_antennanp
XFILLER_61_97 VPWR VGND sg13g2_fill_1
X_0380_ VPWR VGND _0308_ _0309_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q
+ _0287_ _0310_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a221oi_1
X_1001_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_153 VPWR VGND sg13g2_decap_8
XFILLER_34_134 VPWR VGND sg13g2_fill_1
XFILLER_103_139 VPWR VGND sg13g2_decap_8
X_0647_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q _0100_
+ _0101_ _0104_ VPWR VGND sg13g2_nor3_1
X_0578_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q _0047_
+ _0048_ VPWR VGND sg13g2_and2_1
X_0716_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q
+ _0140_ _0139_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb4 _0355_ sg13g2_a221oi_1
XFILLER_102_172 VPWR VGND sg13g2_decap_8
X_1481_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb0 Tile_X0Y0_N2BEGb[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_98_148 VPWR VGND sg13g2_decap_8
X_1550_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG12 Tile_X0Y0_WW4BEG[12]
+ VPWR VGND sg13g2_buf_1
X_0501_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q UIO_OUT_TT_PROJECT1
+ UIO_OE_TT_PROJECT5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG1 VPWR VGND sg13g2_mux4_1
X_0432_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q _0343_
+ _0344_ VPWR VGND sg13g2_nor2_1
X_0363_ VPWR _0293_ Tile_X0Y0_E6END[10] VGND sg13g2_inv_1
XFILLER_94_0 VPWR VGND sg13g2_decap_8
XFILLER_22_104 VPWR VGND sg13g2_fill_2
XFILLER_89_104 VPWR VGND sg13g2_fill_2
XFILLER_97_192 VPWR VGND sg13g2_decap_8
XFILLER_9_119 VPWR VGND sg13g2_fill_1
XFILLER_13_126 VPWR VGND sg13g2_fill_1
XFILLER_42_99 VPWR VGND sg13g2_decap_8
XFILLER_107_92 VPWR VGND sg13g2_decap_8
XFILLER_95_118 VPWR VGND sg13g2_decap_8
X_0981_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1602_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG4 Tile_X0Y1_S2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_1464_ Tile_X0Y1_FrameStrobe[15] Tile_X0Y0_FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_1533_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG7 Tile_X0Y0_W6BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1395_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0415_ _0330_ _0333_ _0335_ VPWR VGND sg13g2_nor2b_1
XFILLER_37_11 VPWR VGND sg13g2_fill_1
XFILLER_37_33 VPWR VGND sg13g2_decap_8
XFILLER_53_87 VPWR VGND sg13g2_decap_8
XFILLER_5_166 VPWR VGND sg13g2_decap_8
XFILLER_76_151 VPWR VGND sg13g2_fill_1
X_1180_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0964_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0895_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0270_ _0271_ VPWR VGND sg13g2_nor3_1
XFILLER_57_0 VPWR VGND sg13g2_decap_4
X_1516_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG6 Tile_X0Y0_W2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1447_ Tile_X0Y0_FrameData[30] Tile_X0Y0_FrameData_O[30] VPWR VGND sg13g2_buf_1
XFILLER_4_92 VPWR VGND sg13g2_fill_1
X_1378_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_114 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_4
XFILLER_80_30 VPWR VGND sg13g2_decap_8
X_0680_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q
+ _0116_ _0115_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG0 _0334_ sg13g2_a221oi_1
XFILLER_50_7 VPWR VGND sg13g2_fill_1
X_1301_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1232_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_151 VPWR VGND sg13g2_decap_8
X_1094_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1163_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0947_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_109_49 VPWR VGND sg13g2_fill_1
X_0878_ _0305_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 _0255_ VPWR VGND sg13g2_nor3_1
XFILLER_18_57 VPWR VGND sg13g2_decap_8
XFILLER_55_110 VPWR VGND sg13g2_decap_4
XFILLER_55_154 VPWR VGND sg13g2_decap_8
XFILLER_34_89 VPWR VGND sg13g2_fill_2
XFILLER_109_123 VPWR VGND sg13g2_fill_1
XFILLER_1_2 VPWR VGND sg13g2_fill_1
XFILLER_75_52 VPWR VGND sg13g2_fill_1
XFILLER_61_102 VPWR VGND sg13g2_fill_1
XFILLER_46_154 VPWR VGND sg13g2_decap_8
XFILLER_91_62 VPWR VGND sg13g2_decap_8
X_0801_ VGND VPWR Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
+ _0189_ _0190_ _0301_ sg13g2_a21oi_1
X_0594_ _0061_ VPWR _0062_ VGND Tile_X0Y0_E6END[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ sg13g2_o21ai_1
X_0732_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0318_ Tile_X0Y0_S4END[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q
+ _0148_ VPWR VGND sg13g2_mux4_1
X_0663_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13
+ _0314_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1146_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1215_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1077_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_45 VPWR VGND sg13g2_fill_1
XFILLER_28_154 VPWR VGND sg13g2_decap_8
XFILLER_43_113 VPWR VGND sg13g2_fill_2
XFILLER_43_157 VPWR VGND sg13g2_decap_8
XFILLER_45_33 VPWR VGND sg13g2_fill_1
XANTENNA_9 VPWR VGND Tile_X0Y1_FrameStrobe[17] sg13g2_antennanp
XFILLER_86_95 VPWR VGND sg13g2_decap_8
XFILLER_86_84 VPWR VGND sg13g2_fill_1
X_1000_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_4 VPWR VGND sg13g2_fill_1
XFILLER_19_198 VPWR VGND sg13g2_fill_2
XFILLER_34_157 VPWR VGND sg13g2_decap_8
X_0715_ UO_OUT_TT_PROJECT4 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q _0140_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_103_118 VPWR VGND sg13g2_decap_8
X_0646_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q _0102_
+ _0103_ VPWR VGND sg13g2_nor2b_1
X_0577_ _0047_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 VPWR VGND sg13g2_nand2b_1
X_1129_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_31_35 VPWR VGND sg13g2_fill_2
XFILLER_102_151 VPWR VGND sg13g2_decap_8
XFILLER_16_113 VPWR VGND sg13g2_decap_8
XFILLER_16_124 VPWR VGND sg13g2_fill_1
XFILLER_16_146 VPWR VGND sg13g2_decap_8
X_1480_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG7 Tile_X0Y0_N2BEG[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_98_127 VPWR VGND sg13g2_decap_8
X_0362_ VPWR _0292_ Tile_X0Y0_E6END[9] VGND sg13g2_inv_1
X_0500_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q UIO_OUT_TT_PROJECT0
+ UIO_OE_TT_PROJECT4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG0 VPWR VGND sg13g2_mux4_1
X_0431_ Tile_X0Y1_N2MID[2] Tile_X0Y1_N2END[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
+ _0343_ VPWR VGND sg13g2_mux2_1
XFILLER_87_0 VPWR VGND sg13g2_decap_4
XFILLER_97_171 VPWR VGND sg13g2_decap_8
X_0629_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q Tile_X0Y0_EE4END[2]
+ Tile_X0Y0_EE4END[10] _0012_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q _0089_ VPWR
+ VGND sg13g2_mux4_1
XFILLER_42_78 VPWR VGND sg13g2_decap_8
XFILLER_107_71 VPWR VGND sg13g2_decap_8
X_0980_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_83_96 VPWR VGND sg13g2_decap_4
XFILLER_80_7 VPWR VGND sg13g2_fill_2
X_1532_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG6 Tile_X0Y0_W6BEG[6]
+ VPWR VGND sg13g2_buf_1
XFILLER_8_186 VPWR VGND sg13g2_decap_8
X_1601_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG3 Tile_X0Y1_S2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_1463_ Tile_X0Y1_FrameStrobe[14] Tile_X0Y0_FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
X_1394_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0414_ _0334_ _0333_ _0330_ VPWR VGND sg13g2_nand2b_1
XFILLER_94_185 VPWR VGND sg13g2_decap_8
XFILLER_85_130 VPWR VGND sg13g2_decap_8
XFILLER_76_196 VPWR VGND sg13g2_decap_4
X_0963_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_0894_ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2END[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0270_ VPWR VGND sg13g2_mux2_1
XFILLER_64_2 VPWR VGND sg13g2_fill_1
X_1515_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG5 Tile_X0Y0_W2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_1446_ Tile_X0Y0_FrameData[29] Tile_X0Y0_FrameData_O[29] VPWR VGND sg13g2_buf_1
X_1377_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_199 VPWR VGND sg13g2_fill_1
XFILLER_82_188 VPWR VGND sg13g2_decap_8
XFILLER_2_159 VPWR VGND sg13g2_decap_8
XFILLER_58_141 VPWR VGND sg13g2_decap_4
XFILLER_104_94 VPWR VGND sg13g2_decap_8
XFILLER_64_32 VPWR VGND sg13g2_decap_8
XFILLER_0_29 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_4
X_1300_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_181 VPWR VGND sg13g2_decap_8
X_1231_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1162_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_141 VPWR VGND sg13g2_decap_4
XFILLER_49_185 VPWR VGND sg13g2_decap_4
X_1093_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_199 VPWR VGND sg13g2_fill_1
X_0946_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0877_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0251_ _0253_ _0248_ _0254_ _0249_ sg13g2_a221oi_1
X_1429_ Tile_X0Y0_FrameData[12] Tile_X0Y0_FrameData_O[12] VPWR VGND sg13g2_buf_1
XFILLER_55_133 VPWR VGND sg13g2_decap_8
XFILLER_55_199 VPWR VGND sg13g2_fill_1
XFILLER_46_199 VPWR VGND sg13g2_fill_1
X_0731_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT4 _0147_ _0356_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG4 VPWR VGND sg13g2_mux4_1
X_0800_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 _0000_
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q _0189_ VPWR
+ VGND sg13g2_mux2_1
X_0593_ _0061_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_nand2b_1
X_0662_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit4.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_E6END[8] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12
+ _0010_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit5.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1145_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1214_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_155 VPWR VGND sg13g2_fill_1
X_1076_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_169 VPWR VGND sg13g2_decap_8
X_0929_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_149 VPWR VGND sg13g2_fill_1
XFILLER_106_138 VPWR VGND sg13g2_decap_8
XFILLER_20_26 VPWR VGND sg13g2_decap_4
XFILLER_28_188 VPWR VGND sg13g2_decap_8
XFILLER_28_199 VPWR VGND sg13g2_fill_1
XFILLER_101_95 VPWR VGND sg13g2_decap_8
XFILLER_61_88 VPWR VGND sg13g2_decap_8
XFILLER_61_66 VPWR VGND sg13g2_decap_4
XFILLER_51_180 VPWR VGND sg13g2_decap_4
XFILLER_19_177 VPWR VGND sg13g2_decap_8
XFILLER_42_180 VPWR VGND sg13g2_decap_8
X_0645_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_EE4END[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q
+ _0102_ VPWR VGND sg13g2_mux4_1
X_0714_ _0139_ _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_nand2b_1
X_0576_ VPWR _0046_ _0045_ VGND sg13g2_inv_1
XFILLER_32_0 VPWR VGND sg13g2_decap_8
X_1128_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_147 VPWR VGND sg13g2_fill_2
X_1059_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_110_7 VPWR VGND sg13g2_decap_8
XFILLER_102_130 VPWR VGND sg13g2_decap_8
XFILLER_56_11 VPWR VGND sg13g2_fill_2
X_0361_ VPWR _0291_ Tile_X0Y0_E6END[8] VGND sg13g2_inv_1
X_0430_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2END[5] Tile_X0Y0_E6END[10] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_22_106 VPWR VGND sg13g2_fill_1
XFILLER_89_128 VPWR VGND sg13g2_fill_2
XFILLER_89_106 VPWR VGND sg13g2_fill_1
X_0628_ _0087_ VPWR _0088_ VGND Tile_X0Y0_E6END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q
+ sg13g2_o21ai_1
XFILLER_97_150 VPWR VGND sg13g2_decap_8
X_0559_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q VPWR
+ _0031_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q
+ _0030_ sg13g2_o21ai_1
XFILLER_42_35 VPWR VGND sg13g2_decap_8
XFILLER_107_50 VPWR VGND sg13g2_decap_8
XFILLER_83_64 VPWR VGND sg13g2_decap_4
XFILLER_83_42 VPWR VGND sg13g2_fill_1
XFILLER_83_31 VPWR VGND sg13g2_decap_8
X_1462_ Tile_X0Y1_FrameStrobe[13] Tile_X0Y0_FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
X_1531_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG5 Tile_X0Y0_W6BEG[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_8_165 VPWR VGND sg13g2_decap_8
X_1600_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG2 Tile_X0Y1_S2BEGb[2]
+ VPWR VGND sg13g2_buf_1
XFILLER_94_131 VPWR VGND sg13g2_fill_2
XFILLER_86_109 VPWR VGND sg13g2_decap_8
XFILLER_79_194 VPWR VGND sg13g2_decap_4
X_0413_ _0331_ _0332_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q
+ _0333_ VPWR VGND sg13g2_nand3_1
X_1393_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_85_197 VPWR VGND sg13g2_fill_2
XFILLER_37_79 VPWR VGND sg13g2_fill_2
X_0962_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_71_4 VPWR VGND sg13g2_fill_2
X_0893_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q _0268_
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q _0269_ VPWR
+ VGND sg13g2_nand3_1
X_1445_ Tile_X0Y0_FrameData[28] Tile_X0Y0_FrameData_O[28] VPWR VGND sg13g2_buf_1
XFILLER_4_72 VPWR VGND sg13g2_decap_8
XFILLER_4_50 VPWR VGND sg13g2_decap_8
X_1514_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG4 Tile_X0Y0_W2BEG[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_82_123 VPWR VGND sg13g2_fill_2
XFILLER_67_175 VPWR VGND sg13g2_fill_2
X_1376_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_73_167 VPWR VGND sg13g2_fill_1
XFILLER_80_87 VPWR VGND sg13g2_fill_1
XFILLER_1_160 VPWR VGND sg13g2_decap_8
X_1092_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_64_145 VPWR VGND sg13g2_fill_1
X_1230_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1161_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0945_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_62_0 VPWR VGND sg13g2_decap_4
X_0876_ VPWR _0253_ _0252_ VGND sg13g2_inv_1
X_1428_ Tile_X0Y0_FrameData[11] Tile_X0Y0_FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_70_148 VPWR VGND sg13g2_fill_1
X_1359_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_11 VPWR VGND sg13g2_fill_2
XFILLER_59_77 VPWR VGND sg13g2_decap_8
XFILLER_61_137 VPWR VGND sg13g2_decap_4
X_0661_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_E6END[4]
+ _0006_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG0
+ VPWR VGND sg13g2_mux4_1
X_0730_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0325_ Tile_X0Y0_S4END[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q
+ _0147_ VPWR VGND sg13g2_mux4_1
XFILLER_108_191 VPWR VGND sg13g2_fill_1
X_0592_ VGND VPWR _0055_ _0058_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG1
+ _0060_ sg13g2_a21oi_1
X_1213_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1144_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1075_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_1_51 VPWR VGND sg13g2_fill_1
XFILLER_1_95 VPWR VGND sg13g2_fill_2
XFILLER_52_148 VPWR VGND sg13g2_decap_8
XFILLER_60_170 VPWR VGND sg13g2_fill_2
X_0928_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_117 VPWR VGND sg13g2_decap_8
X_0859_ _0238_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_nand2b_1
XFILLER_28_167 VPWR VGND sg13g2_fill_2
XFILLER_43_115 VPWR VGND sg13g2_fill_1
XFILLER_105_183 VPWR VGND sg13g2_decap_8
XFILLER_86_64 VPWR VGND sg13g2_fill_2
XFILLER_19_80 VPWR VGND sg13g2_decap_8
X_0644_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q VPWR
+ _0101_ VGND Tile_X0Y0_EE4END[13] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q
+ sg13g2_o21ai_1
X_0713_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q
+ _0138_ _0137_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb3 _0355_ sg13g2_a221oi_1
X_0575_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q VPWR
+ _0045_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q
+ _0044_ sg13g2_o21ai_1
XFILLER_25_0 VPWR VGND sg13g2_decap_8
X_1127_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1058_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_31_37 VPWR VGND sg13g2_fill_1
XFILLER_102_186 VPWR VGND sg13g2_decap_8
XFILLER_56_34 VPWR VGND sg13g2_decap_8
XFILLER_97_41 VPWR VGND sg13g2_fill_2
X_0360_ VPWR _0290_ Tile_X0Y0_E6END[0] VGND sg13g2_inv_1
XFILLER_30_173 VPWR VGND sg13g2_fill_2
X_0558_ _0029_ VPWR _0030_ VGND Tile_X0Y0_E6END[10] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ sg13g2_o21ai_1
X_0627_ VGND VPWR _0293_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit22.Q
+ _0087_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit24.Q sg13g2_a21oi_1
X_0489_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q UIO_OUT_TT_PROJECT5
+ UIO_OE_TT_PROJECT5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_13_107 VPWR VGND sg13g2_fill_2
XFILLER_21_184 VPWR VGND sg13g2_decap_8
XFILLER_88_140 VPWR VGND sg13g2_fill_1
XFILLER_67_66 VPWR VGND sg13g2_decap_8
XFILLER_67_33 VPWR VGND sg13g2_decap_8
XFILLER_67_11 VPWR VGND sg13g2_fill_1
XFILLER_12_184 VPWR VGND sg13g2_decap_8
X_1461_ Tile_X0Y1_FrameStrobe[12] Tile_X0Y0_FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
X_1530_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG4 Tile_X0Y0_W6BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0412_ _0332_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
+ Tile_X0Y0_S2MID[0] VPWR VGND sg13g2_nand2_1
X_1392_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_0 VPWR VGND sg13g2_decap_8
X_1659_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG5 Tile_X0Y1_WW4BEG[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_85_176 VPWR VGND sg13g2_decap_8
XFILLER_53_24 VPWR VGND sg13g2_fill_1
XFILLER_5_125 VPWR VGND sg13g2_decap_4
XFILLER_91_135 VPWR VGND sg13g2_fill_2
X_0961_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_94_97 VPWR VGND sg13g2_decap_8
XFILLER_91_168 VPWR VGND sg13g2_fill_2
X_0892_ _0268_ Tile_X0Y1_E2END[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_nand2_1
X_1444_ Tile_X0Y0_FrameData[27] Tile_X0Y0_FrameData_O[27] VPWR VGND sg13g2_buf_1
X_1375_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1513_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG3 Tile_X0Y0_W2BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_82_113 VPWR VGND sg13g2_decap_4
XFILLER_67_198 VPWR VGND sg13g2_fill_2
XFILLER_2_139 VPWR VGND sg13g2_fill_2
XFILLER_73_124 VPWR VGND sg13g2_fill_1
XFILLER_58_198 VPWR VGND sg13g2_fill_2
XFILLER_81_190 VPWR VGND sg13g2_decap_8
XFILLER_64_89 VPWR VGND sg13g2_fill_1
XFILLER_80_44 VPWR VGND sg13g2_fill_1
XFILLER_89_97 VPWR VGND sg13g2_decap_8
X_1091_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_165 VPWR VGND sg13g2_decap_8
X_1160_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0944_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0875_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q Tile_X0Y1_N2END[3]
+ Tile_X0Y1_E2END[1] Tile_X0Y1_E2MID[0] Tile_X0Y1_E2END[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0252_ VPWR VGND sg13g2_mux4_1
X_1358_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1427_ Tile_X0Y0_FrameData[10] Tile_X0Y0_FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_70_116 VPWR VGND sg13g2_decap_8
X_1289_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_168 VPWR VGND sg13g2_decap_8
XFILLER_55_179 VPWR VGND sg13g2_fill_2
XFILLER_109_159 VPWR VGND sg13g2_fill_1
XFILLER_109_148 VPWR VGND sg13g2_fill_2
XFILLER_109_104 VPWR VGND sg13g2_fill_1
XFILLER_46_168 VPWR VGND sg13g2_decap_8
X_0660_ VGND VPWR UIO_IN_TT_PROJECT7 _0114_ _0113_ sg13g2_or2_1
X_0591_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q _0059_
+ _0060_ VPWR VGND sg13g2_nor2_1
XFILLER_40_80 VPWR VGND sg13g2_fill_2
X_1212_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_4 VPWR VGND sg13g2_fill_1
X_1143_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1074_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_105 VPWR VGND sg13g2_decap_8
XFILLER_52_127 VPWR VGND sg13g2_decap_8
X_0927_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0858_ _0237_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q VPWR VGND
+ sg13g2_nand2b_1
X_0789_ VGND VPWR _0174_ _0177_ Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_10.A _0179_ sg13g2_a21oi_1
XFILLER_6_19 VPWR VGND sg13g2_fill_1
XFILLER_105_162 VPWR VGND sg13g2_decap_8
XFILLER_86_21 VPWR VGND sg13g2_fill_2
XFILLER_10_72 VPWR VGND sg13g2_fill_2
X_0643_ Tile_X0Y0_E6END[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q
+ _0100_ VPWR VGND sg13g2_nor2b_1
X_0574_ _0043_ VPWR _0044_ VGND Tile_X0Y0_E6END[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ sg13g2_o21ai_1
X_0712_ UO_OUT_TT_PROJECT3 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q _0138_ VPWR
+ VGND sg13g2_nor3_1
X_1126_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_0 VPWR VGND sg13g2_fill_2
X_1057_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_25_149 VPWR VGND sg13g2_fill_1
XFILLER_33_193 VPWR VGND sg13g2_decap_8
XFILLER_102_165 VPWR VGND sg13g2_decap_8
XFILLER_24_193 VPWR VGND sg13g2_decap_8
XFILLER_97_97 VPWR VGND sg13g2_fill_2
XFILLER_15_193 VPWR VGND sg13g2_decap_8
XFILLER_97_185 VPWR VGND sg13g2_decap_8
X_0557_ _0029_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_nand2b_1
X_0626_ VGND VPWR Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q
+ _0084_ UIO_IN_TT_PROJECT1 _0086_ sg13g2_a21oi_1
X_1109_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0488_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q UIO_OUT_TT_PROJECT4
+ UIO_OE_TT_PROJECT4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG4 VPWR VGND sg13g2_mux4_1
XFILLER_107_85 VPWR VGND sg13g2_decap_8
XFILLER_88_130 VPWR VGND sg13g2_decap_4
X_1460_ Tile_X0Y1_FrameStrobe[11] Tile_X0Y0_FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
X_1391_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0411_ _0331_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_94_199 VPWR VGND sg13g2_fill_1
XFILLER_85_0 VPWR VGND sg13g2_fill_2
X_1658_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG4 Tile_X0Y1_WW4BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0609_ _0075_ VPWR _0076_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ _0011_ sg13g2_o21ai_1
X_1589_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG3 Tile_X0Y1_S1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_85_199 VPWR VGND sg13g2_fill_1
XFILLER_5_148 VPWR VGND sg13g2_fill_1
XFILLER_76_133 VPWR VGND sg13g2_fill_1
X_0960_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1512_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG2 Tile_X0Y0_W2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0891_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q Tile_X0Y1_E2END[1]
+ _0267_ VPWR VGND sg13g2_nor2b_1
XFILLER_57_4 VPWR VGND sg13g2_fill_2
X_1443_ Tile_X0Y0_FrameData[26] Tile_X0Y0_FrameData_O[26] VPWR VGND sg13g2_buf_1
XFILLER_4_181 VPWR VGND sg13g2_decap_8
X_1374_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_107 VPWR VGND sg13g2_decap_8
XFILLER_58_111 VPWR VGND sg13g2_fill_2
XFILLER_64_46 VPWR VGND sg13g2_fill_2
XFILLER_1_195 VPWR VGND sg13g2_decap_4
X_1090_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_80 VPWR VGND sg13g2_fill_1
X_0943_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0874_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ _0250_ _0251_ VPWR VGND sg13g2_nor3_1
XFILLER_48_0 VPWR VGND sg13g2_decap_8
X_1288_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_28 VPWR VGND sg13g2_fill_1
X_1357_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_55_103 VPWR VGND sg13g2_decap_8
XFILLER_55_114 VPWR VGND sg13g2_fill_2
XFILLER_55_147 VPWR VGND sg13g2_decap_8
X_1426_ Tile_X0Y0_FrameData[9] Tile_X0Y0_FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_109_116 VPWR VGND sg13g2_decap_8
Xclkbuf_1_1__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_1__leaf_Tile_X0Y1_UserCLK
+ VPWR VGND sg13g2_buf_8
XFILLER_75_45 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_108_171 VPWR VGND sg13g2_fill_1
X_0590_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_EE4END[13] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ _0059_ VPWR VGND sg13g2_mux4_1
XFILLER_41_7 VPWR VGND sg13g2_decap_4
X_1142_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1211_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1073_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_172 VPWR VGND sg13g2_fill_1
X_0857_ _0233_ VPWR UI_IN_TT_PROJECT5 VGND _0234_ _0236_ sg13g2_o21ai_1
X_0926_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0788_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q _0178_
+ _0179_ VPWR VGND sg13g2_nor2_1
X_1409_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_147 VPWR VGND sg13g2_decap_8
XFILLER_105_141 VPWR VGND sg13g2_decap_8
XFILLER_86_66 VPWR VGND sg13g2_fill_1
XFILLER_42_150 VPWR VGND sg13g2_decap_4
XFILLER_89_7 VPWR VGND sg13g2_decap_4
X_0711_ _0137_ _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_42_194 VPWR VGND sg13g2_decap_4
X_0642_ VGND VPWR UIO_IN_TT_PROJECT4 _0099_ _0098_ sg13g2_or2_1
X_0573_ _0043_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_nand2b_1
X_1125_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1056_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0909_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q _0282_
+ _0284_ _0285_ VPWR VGND sg13g2_nor3_1
XFILLER_102_144 VPWR VGND sg13g2_decap_8
XFILLER_72_68 VPWR VGND sg13g2_fill_1
XFILLER_16_106 VPWR VGND sg13g2_decap_8
XFILLER_97_76 VPWR VGND sg13g2_fill_1
XFILLER_97_43 VPWR VGND sg13g2_fill_1
XFILLER_87_4 VPWR VGND sg13g2_fill_1
X_0625_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q _0085_
+ _0086_ VPWR VGND sg13g2_nor2_1
XFILLER_30_175 VPWR VGND sg13g2_fill_1
XFILLER_97_164 VPWR VGND sg13g2_decap_8
X_0556_ _0026_ _0028_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG1
+ VPWR VGND sg13g2_nor2_1
X_0487_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit30.Q UIO_OUT_TT_PROJECT3
+ UIO_OE_TT_PROJECT3 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG3 VPWR VGND sg13g2_mux4_1
X_1108_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1039_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_42_49 VPWR VGND sg13g2_fill_2
XFILLER_107_64 VPWR VGND sg13g2_decap_8
XFILLER_12_120 VPWR VGND sg13g2_decap_4
XFILLER_8_179 VPWR VGND sg13g2_decap_8
XFILLER_79_175 VPWR VGND sg13g2_fill_2
X_1390_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0410_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit9.Q _0329_
+ _0330_ VPWR VGND sg13g2_nor2_1
XFILLER_94_178 VPWR VGND sg13g2_decap_8
XFILLER_78_0 VPWR VGND sg13g2_fill_2
X_0608_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q _0074_
+ _0075_ VPWR VGND sg13g2_and2_1
X_1657_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG3 Tile_X0Y1_WW4BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_7_190 VPWR VGND sg13g2_decap_8
X_1588_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG2 Tile_X0Y1_S1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0539_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q UIO_OUT_TT_PROJECT2
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 _0013_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG10
+ VPWR VGND sg13g2_mux4_1
XFILLER_43_70 VPWR VGND sg13g2_decap_4
X_0890_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0266_ VPWR VGND sg13g2_nor2b_1
X_1442_ Tile_X0Y0_FrameData[25] Tile_X0Y0_FrameData_O[25] VPWR VGND sg13g2_buf_1
X_1511_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG1 Tile_X0Y0_W2BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_4_160 VPWR VGND sg13g2_decap_8
XFILLER_4_42 VPWR VGND sg13g2_fill_2
XFILLER_67_145 VPWR VGND sg13g2_decap_4
XFILLER_4_86 VPWR VGND sg13g2_fill_1
X_1373_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_29 VPWR VGND sg13g2_fill_2
XFILLER_104_87 VPWR VGND sg13g2_decap_8
XFILLER_58_134 VPWR VGND sg13g2_decap_8
XFILLER_58_145 VPWR VGND sg13g2_fill_1
XFILLER_58_167 VPWR VGND sg13g2_decap_4
XFILLER_89_11 VPWR VGND sg13g2_fill_1
XFILLER_8_0 VPWR VGND sg13g2_fill_2
XFILLER_1_174 VPWR VGND sg13g2_decap_8
XFILLER_49_145 VPWR VGND sg13g2_fill_2
X_0942_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0873_ Tile_X0Y1_N2MID[6] Tile_X0Y1_N2END[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0250_ VPWR VGND sg13g2_mux2_1
X_1425_ Tile_X0Y0_FrameData[8] Tile_X0Y0_FrameData_O[8] VPWR VGND sg13g2_buf_1
X_1287_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1356_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_46_104 VPWR VGND sg13g2_fill_1
XFILLER_59_47 VPWR VGND sg13g2_decap_4
XFILLER_91_56 VPWR VGND sg13g2_fill_2
XFILLER_108_150 VPWR VGND sg13g2_decap_8
X_1141_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1072_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1210_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0925_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0856_ _0235_ VPWR _0236_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
+ _0153_ sg13g2_o21ai_1
X_0787_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E6END[10] Tile_X0Y1_EE4END[2] _0156_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ _0178_ VPWR VGND sg13g2_mux4_1
XFILLER_28_104 VPWR VGND sg13g2_decap_4
X_1408_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1339_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_88 VPWR VGND sg13g2_decap_8
XFILLER_61_59 VPWR VGND sg13g2_decap_8
XFILLER_51_173 VPWR VGND sg13g2_decap_8
XFILLER_51_184 VPWR VGND sg13g2_fill_1
XFILLER_105_120 VPWR VGND sg13g2_decap_8
XFILLER_105_197 VPWR VGND sg13g2_fill_2
XFILLER_19_94 VPWR VGND sg13g2_decap_4
XFILLER_34_107 VPWR VGND sg13g2_fill_2
XFILLER_42_173 VPWR VGND sg13g2_decap_8
X_0641_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q _0095_
+ _0096_ _0099_ VPWR VGND sg13g2_nor3_1
X_0710_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q
+ _0136_ _0135_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb2 _0348_ sg13g2_a221oi_1
X_0572_ _0040_ _0042_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG3
+ VPWR VGND sg13g2_nor2_1
X_1124_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_18_192 VPWR VGND sg13g2_decap_8
X_1055_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0839_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q _0219_
+ _0220_ _0222_ VPWR VGND sg13g2_nor3_1
X_0908_ Tile_X0Y0_S2MID[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ _0284_ VPWR VGND sg13g2_nor2b_1
XFILLER_102_123 VPWR VGND sg13g2_decap_8
XFILLER_56_48 VPWR VGND sg13g2_decap_4
XFILLER_24_162 VPWR VGND sg13g2_decap_8
XFILLER_108_0 VPWR VGND sg13g2_decap_8
X_0624_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q Tile_X0Y0_EE4END[1]
+ Tile_X0Y0_EE4END[9] _0013_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q _0085_ VPWR
+ VGND sg13g2_mux4_1
XFILLER_30_198 VPWR VGND sg13g2_fill_2
XFILLER_97_143 VPWR VGND sg13g2_decap_8
X_0555_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q _0027_
+ _0028_ VPWR VGND sg13g2_nor2_1
X_0486_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit28.Q UIO_OUT_TT_PROJECT2
+ UIO_OE_TT_PROJECT2 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit29.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG2 VPWR VGND sg13g2_mux4_1
X_1107_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1038_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_198 VPWR VGND sg13g2_fill_2
XFILLER_107_43 VPWR VGND sg13g2_decap_8
XFILLER_101_7 VPWR VGND sg13g2_decap_8
XFILLER_67_47 VPWR VGND sg13g2_fill_2
XFILLER_83_68 VPWR VGND sg13g2_fill_1
XFILLER_12_198 VPWR VGND sg13g2_fill_2
XFILLER_8_158 VPWR VGND sg13g2_decap_8
XFILLER_79_198 VPWR VGND sg13g2_fill_2
XFILLER_85_2 VPWR VGND sg13g2_fill_1
X_0607_ _0074_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 VPWR VGND sg13g2_nand2b_1
X_0538_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q UIO_OUT_TT_PROJECT1
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 _0012_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG9
+ VPWR VGND sg13g2_mux4_1
X_1656_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG2 Tile_X0Y1_WW4BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1587_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG1 Tile_X0Y1_S1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_0469_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit22.Q Tile_X0Y1_E2MID[0]
+ Tile_X0Y1_E2END[0] Tile_X0Y1_E6END[0] _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit23.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb7 VPWR VGND sg13g2_mux4_1
XFILLER_76_102 VPWR VGND sg13g2_fill_1
XFILLER_84_190 VPWR VGND sg13g2_decap_8
X_1441_ Tile_X0Y0_FrameData[24] Tile_X0Y0_FrameData_O[24] VPWR VGND sg13g2_buf_1
X_1510_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG0 Tile_X0Y0_W2BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_4_98 VPWR VGND sg13g2_fill_1
X_1372_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_90_0 VPWR VGND sg13g2_decap_4
X_1639_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb5 Tile_X0Y1_W2BEGb[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_66 VPWR VGND sg13g2_decap_4
XFILLER_13_30 VPWR VGND sg13g2_fill_2
XFILLER_13_74 VPWR VGND sg13g2_decap_4
XFILLER_1_131 VPWR VGND sg13g2_fill_1
XFILLER_49_179 VPWR VGND sg13g2_fill_2
XFILLER_72_193 VPWR VGND sg13g2_decap_8
X_0941_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_0872_ VGND VPWR Tile_X0Y1_E2MID[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
+ _0249_ _0247_ sg13g2_a21oi_1
X_1355_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1424_ Tile_X0Y0_FrameData[7] Tile_X0Y0_FrameData_O[7] VPWR VGND sg13g2_buf_1
X_1286_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_195 VPWR VGND sg13g2_fill_1
X_1140_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1071_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_52_119 VPWR VGND sg13g2_decap_4
X_0924_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_163 VPWR VGND sg13g2_decap_8
XFILLER_45_193 VPWR VGND sg13g2_decap_8
X_0855_ _0235_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_nand2b_1
X_0786_ _0176_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q
+ _0177_ VPWR VGND sg13g2_nor2b_1
XFILLER_53_0 VPWR VGND sg13g2_decap_8
X_1338_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1407_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1269_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_152 VPWR VGND sg13g2_decap_8
XFILLER_105_176 VPWR VGND sg13g2_decap_8
X_0571_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q _0041_
+ _0042_ VPWR VGND sg13g2_nor2_1
X_0640_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q _0097_
+ _0098_ VPWR VGND sg13g2_nor2b_1
X_1123_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1054_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0907_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q VPWR
+ _0283_ VGND _0295_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q
+ sg13g2_o21ai_1
XFILLER_102_102 VPWR VGND sg13g2_decap_8
X_0769_ VGND VPWR Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ _0334_ _0162_ _0161_ sg13g2_a21oi_1
X_0838_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y1_EE4END[2]
+ Tile_X0Y1_EE4END[10] Tile_X0Y1_E6END[2] Tile_X0Y1_E6END[10] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q
+ _0221_ VPWR VGND sg13g2_mux4_1
XFILLER_102_179 VPWR VGND sg13g2_decap_8
XFILLER_97_34 VPWR VGND sg13g2_decap_8
XFILLER_97_122 VPWR VGND sg13g2_decap_8
X_0623_ _0083_ VPWR _0084_ VGND Tile_X0Y0_E6END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q
+ sg13g2_o21ai_1
X_0554_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_EE4END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ _0027_ VPWR VGND sg13g2_mux4_1
XFILLER_97_199 VPWR VGND sg13g2_fill_1
X_1106_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0485_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit26.Q UIO_OUT_TT_PROJECT1
+ UIO_OE_TT_PROJECT1 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit27.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG1 VPWR VGND sg13g2_mux4_1
X_1037_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_21_122 VPWR VGND sg13g2_decap_8
XFILLER_107_99 VPWR VGND sg13g2_decap_8
XFILLER_88_111 VPWR VGND sg13g2_fill_2
XFILLER_32_84 VPWR VGND sg13g2_decap_4
X_0606_ VPWR _0073_ _0072_ VGND sg13g2_inv_1
X_0537_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q UIO_OUT_TT_PROJECT0
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 _0011_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG8
+ VPWR VGND sg13g2_mux4_1
X_1655_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG1 Tile_X0Y1_WW4BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1586_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S1BEG0 Tile_X0Y1_S1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0399_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3 _0323_ VPWR VGND sg13g2_nor3_1
X_0468_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q Tile_X0Y1_N2MID[7]
+ Tile_X0Y1_N2END[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG7
+ Tile_X0Y0_S2MID[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q
+ _0003_ VPWR VGND sg13g2_mux4_1
XFILLER_78_36 VPWR VGND sg13g2_decap_8
XFILLER_5_129 VPWR VGND sg13g2_fill_2
XFILLER_91_128 VPWR VGND sg13g2_decap_8
X_1440_ Tile_X0Y0_FrameData[23] Tile_X0Y0_FrameData_O[23] VPWR VGND sg13g2_buf_1
XFILLER_4_195 VPWR VGND sg13g2_decap_4
XFILLER_4_44 VPWR VGND sg13g2_fill_1
XFILLER_4_22 VPWR VGND sg13g2_fill_2
X_1371_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_117 VPWR VGND sg13g2_fill_1
XFILLER_82_106 VPWR VGND sg13g2_decap_8
XFILLER_75_180 VPWR VGND sg13g2_decap_8
XFILLER_83_0 VPWR VGND sg13g2_decap_8
X_1638_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb4 Tile_X0Y1_W2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_1569_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameData_O[15] VPWR VGND sg13g2_buf_1
XFILLER_81_183 VPWR VGND sg13g2_decap_8
XFILLER_80_37 VPWR VGND sg13g2_decap_8
XFILLER_8_2 VPWR VGND sg13g2_fill_1
XFILLER_49_103 VPWR VGND sg13g2_decap_4
XFILLER_49_158 VPWR VGND sg13g2_decap_8
X_0940_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0871_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q _0306_
+ _0248_ VPWR VGND sg13g2_nor2_1
X_1285_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1354_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1423_ Tile_X0Y0_FrameData[6] Tile_X0Y0_FrameData_O[6] VPWR VGND sg13g2_buf_1
XFILLER_91_69 VPWR VGND sg13g2_decap_4
XFILLER_108_130 VPWR VGND sg13g2_decap_4
XFILLER_45_183 VPWR VGND sg13g2_fill_2
X_1070_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0923_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0854_ _0234_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q VPWR VGND
+ sg13g2_nand2b_1
X_0785_ VGND VPWR Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ _0348_ _0176_ _0175_ sg13g2_a21oi_1
X_1337_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1268_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_128 VPWR VGND sg13g2_fill_2
X_1406_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1199_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_131 VPWR VGND sg13g2_decap_8
XFILLER_51_197 VPWR VGND sg13g2_fill_2
XFILLER_105_199 VPWR VGND sg13g2_fill_1
XFILLER_105_155 VPWR VGND sg13g2_decap_8
XFILLER_27_194 VPWR VGND sg13g2_decap_4
XFILLER_35_73 VPWR VGND sg13g2_fill_2
X_0570_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_EE4END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ _0041_ VPWR VGND sg13g2_mux4_1
XFILLER_51_94 VPWR VGND sg13g2_fill_2
X_1122_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1053_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0837_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q _0156_
+ _0220_ VPWR VGND sg13g2_nor2_1
X_0906_ Tile_X0Y1_E2END[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q _0282_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_102_158 VPWR VGND sg13g2_decap_8
X_0699_ _0129_ _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
X_0768_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q VPWR
+ _0161_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 sg13g2_o21ai_1
XFILLER_110_191 VPWR VGND sg13g2_decap_8
XFILLER_24_186 VPWR VGND sg13g2_decap_8
XFILLER_15_175 VPWR VGND sg13g2_fill_1
XFILLER_62_93 VPWR VGND sg13g2_fill_1
XFILLER_7_77 VPWR VGND sg13g2_fill_1
XFILLER_7_22 VPWR VGND sg13g2_fill_2
X_0622_ VGND VPWR _0292_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q
+ _0083_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q sg13g2_a21oi_1
X_0553_ VGND VPWR Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q
+ _0025_ _0026_ _0024_ sg13g2_a21oi_1
X_0484_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit24.Q UIO_OUT_TT_PROJECT0
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit25.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG0 VPWR VGND sg13g2_mux4_1
XFILLER_97_178 VPWR VGND sg13g2_decap_8
X_1105_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1036_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_78 VPWR VGND sg13g2_decap_8
XFILLER_88_167 VPWR VGND sg13g2_fill_2
XFILLER_16_86 VPWR VGND sg13g2_fill_2
XFILLER_12_145 VPWR VGND sg13g2_fill_1
XFILLER_8_105 VPWR VGND sg13g2_fill_2
XFILLER_94_104 VPWR VGND sg13g2_decap_4
XFILLER_73_92 VPWR VGND sg13g2_fill_2
X_1654_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG0 Tile_X0Y1_WW4BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0605_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q VPWR
+ _0072_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q
+ _0071_ sg13g2_o21ai_1
XFILLER_85_137 VPWR VGND sg13g2_fill_1
X_0467_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E2MID[0] Tile_X0Y0_E2END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG7
+ VPWR VGND sg13g2_mux4_1
X_0536_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit6.Q UIO_OUT_TT_PROJECT7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit7.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG7 VPWR VGND sg13g2_mux4_1
X_1585_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameData_O[31] VPWR VGND sg13g2_buf_1
X_0398_ _0322_ Tile_X0Y0_S1END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_93_192 VPWR VGND sg13g2_decap_8
X_1019_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_4_174 VPWR VGND sg13g2_decap_8
X_1370_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1637_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb3 Tile_X0Y1_W2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_1499_ Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_10.A Tile_X0Y0_N4BEG[10] VPWR VGND sg13g2_buf_1
X_0519_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 VPWR VGND sg13g2_mux4_1
X_1568_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameData_O[14] VPWR VGND sg13g2_buf_1
XFILLER_58_104 VPWR VGND sg13g2_decap_8
XFILLER_64_39 VPWR VGND sg13g2_decap_8
XFILLER_1_188 VPWR VGND sg13g2_decap_8
XFILLER_1_199 VPWR VGND sg13g2_fill_1
XFILLER_38_95 VPWR VGND sg13g2_fill_1
X_0870_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q Tile_X0Y1_E2MID[3]
+ _0247_ VPWR VGND sg13g2_nor2b_1
X_1422_ Tile_X0Y0_FrameData[5] Tile_X0Y0_FrameData_O[5] VPWR VGND sg13g2_buf_1
X_1284_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1353_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_181 VPWR VGND sg13g2_decap_4
XFILLER_109_109 VPWR VGND sg13g2_decap_8
X_0999_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_97 VPWR VGND sg13g2_decap_8
XFILLER_108_164 VPWR VGND sg13g2_decap_4
XFILLER_6_0 VPWR VGND sg13g2_fill_2
XFILLER_40_30 VPWR VGND sg13g2_fill_2
XFILLER_60_110 VPWR VGND sg13g2_fill_1
XFILLER_45_151 VPWR VGND sg13g2_decap_8
XFILLER_45_162 VPWR VGND sg13g2_decap_8
X_0922_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_81_92 VPWR VGND sg13g2_fill_2
XFILLER_60_198 VPWR VGND sg13g2_fill_2
X_0853_ _0233_ _0232_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit25.Q
+ VPWR VGND sg13g2_nand2b_1
X_1405_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_39_0 VPWR VGND sg13g2_decap_4
X_0784_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q VPWR
+ _0175_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 sg13g2_o21ai_1
X_1336_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1267_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1198_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_14 VPWR VGND sg13g2_fill_2
XFILLER_105_134 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_fill_2
XFILLER_42_154 VPWR VGND sg13g2_fill_2
XFILLER_42_187 VPWR VGND sg13g2_decap_8
XFILLER_42_198 VPWR VGND sg13g2_fill_2
XFILLER_51_62 VPWR VGND sg13g2_decap_4
XFILLER_32_7 VPWR VGND sg13g2_fill_2
X_1121_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1052_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_91 VPWR VGND sg13g2_fill_2
XFILLER_18_162 VPWR VGND sg13g2_fill_2
XFILLER_33_110 VPWR VGND sg13g2_fill_2
X_0767_ _0160_ _0159_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q
+ VPWR VGND sg13g2_nand2b_1
X_0836_ _0148_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q
+ _0219_ VPWR VGND sg13g2_nor2b_1
X_0905_ _0278_ _0280_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit4.Q
+ _0281_ VPWR VGND sg13g2_nand3_1
XFILLER_102_137 VPWR VGND sg13g2_decap_8
X_0698_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q
+ _0128_ _0127_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG6 _0341_ sg13g2_a221oi_1
X_1319_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_121 VPWR VGND sg13g2_decap_4
XFILLER_97_69 VPWR VGND sg13g2_decap_8
XFILLER_21_43 VPWR VGND sg13g2_decap_8
X_0621_ VGND VPWR Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q
+ _0080_ UIO_IN_TT_PROJECT0 _0082_ sg13g2_a21oi_1
XFILLER_97_157 VPWR VGND sg13g2_decap_8
XFILLER_97_102 VPWR VGND sg13g2_fill_2
XFILLER_87_91 VPWR VGND sg13g2_fill_2
X_0552_ _0013_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ _0025_ VPWR VGND sg13g2_mux2_1
X_0483_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3
+ UIO_OUT_TT_PROJECT1 Tile_X0Y0_S1END[3] UIO_OUT_TT_PROJECT4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG3 VPWR VGND sg13g2_mux4_1
X_1104_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1035_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_57 VPWR VGND sg13g2_decap_8
XFILLER_107_24 VPWR VGND sg13g2_fill_2
X_0819_ _0151_ _0147_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q
+ _0205_ VPWR VGND sg13g2_mux2_1
XFILLER_83_38 VPWR VGND sg13g2_decap_4
XFILLER_79_157 VPWR VGND sg13g2_fill_1
XFILLER_57_72 VPWR VGND sg13g2_decap_8
X_0604_ _0070_ VPWR _0071_ VGND Tile_X0Y0_E6END[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ sg13g2_o21ai_1
XFILLER_7_183 VPWR VGND sg13g2_decap_8
X_1653_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG11 Tile_X0Y1_W6BEG[11]
+ VPWR VGND sg13g2_buf_1
X_1584_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameData_O[30] VPWR VGND sg13g2_buf_1
X_0397_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E6END[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14
+ _0317_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux4_1
X_0466_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q Tile_X0Y0_E2MID[1]
+ Tile_X0Y0_E2END[1] Tile_X0Y0_E6END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG6
+ VPWR VGND sg13g2_mux4_1
XFILLER_78_190 VPWR VGND sg13g2_decap_8
X_0535_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit4.Q UIO_OUT_TT_PROJECT6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit5.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG6 VPWR VGND sg13g2_mux4_1
X_1018_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_4_120 VPWR VGND sg13g2_fill_2
XFILLER_4_24 VPWR VGND sg13g2_fill_1
XFILLER_68_93 VPWR VGND sg13g2_fill_1
XFILLER_67_149 VPWR VGND sg13g2_fill_1
XFILLER_4_79 VPWR VGND sg13g2_decap_8
XFILLER_4_57 VPWR VGND sg13g2_fill_2
XFILLER_69_0 VPWR VGND sg13g2_fill_2
X_0518_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q UIO_OUT_TT_PROJECT6
+ UIO_OE_TT_PROJECT2 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG10 VPWR VGND sg13g2_mux4_1
X_1636_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb2 Tile_X0Y1_W2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_1567_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameData_O[13] VPWR VGND sg13g2_buf_1
X_1498_ Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_9.A Tile_X0Y0_N4BEG[9] VPWR VGND sg13g2_buf_1
X_0449_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y1_E2MID[4]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E6END[4] _0356_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb3 VPWR VGND sg13g2_mux4_1
XFILLER_1_167 VPWR VGND sg13g2_decap_8
XFILLER_38_52 VPWR VGND sg13g2_decap_8
XFILLER_72_185 VPWR VGND sg13g2_decap_4
XFILLER_72_141 VPWR VGND sg13g2_fill_2
XFILLER_57_171 VPWR VGND sg13g2_decap_4
XFILLER_110_90 VPWR VGND sg13g2_decap_8
X_1421_ Tile_X0Y0_FrameData[4] Tile_X0Y0_FrameData_O[4] VPWR VGND sg13g2_buf_1
X_1283_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1352_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_160 VPWR VGND sg13g2_decap_8
X_0998_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1619_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG1 Tile_X0Y1_S4BEG[13]
+ VPWR VGND sg13g2_buf_1
XFILLER_54_152 VPWR VGND sg13g2_decap_8
XFILLER_54_163 VPWR VGND sg13g2_fill_1
XFILLER_108_143 VPWR VGND sg13g2_decap_8
XFILLER_37_108 VPWR VGND sg13g2_fill_2
XFILLER_49_73 VPWR VGND sg13g2_fill_2
X_0921_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0852_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit24.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_EE4END[13] Tile_X0Y1_EE4END[5] Tile_X0Y1_E6END[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit23.Q
+ _0232_ VPWR VGND sg13g2_mux4_1
X_0783_ _0174_ _0173_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_nand2b_1
X_1335_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1404_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1197_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1266_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_130 VPWR VGND sg13g2_decap_8
XFILLER_101_37 VPWR VGND sg13g2_fill_2
XFILLER_51_166 VPWR VGND sg13g2_decap_8
XFILLER_51_199 VPWR VGND sg13g2_fill_1
XFILLER_105_113 VPWR VGND sg13g2_decap_8
XFILLER_19_87 VPWR VGND sg13g2_decap_8
XFILLER_35_75 VPWR VGND sg13g2_fill_1
XFILLER_35_97 VPWR VGND sg13g2_decap_4
XFILLER_25_7 VPWR VGND sg13g2_decap_4
X_1120_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_76_60 VPWR VGND sg13g2_decap_4
XFILLER_18_185 VPWR VGND sg13g2_decap_8
X_1051_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0904_ VGND VPWR _0296_ _0266_ _0280_ _0279_ sg13g2_a21oi_1
X_0697_ UO_OUT_TT_PROJECT6 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit29.Q _0128_ VPWR
+ VGND sg13g2_nor3_1
X_0766_ _0154_ _0150_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ _0159_ VPWR VGND sg13g2_mux2_1
X_0835_ _0216_ VPWR UI_IN_TT_PROJECT1 VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q
+ _0218_ sg13g2_o21ai_1
XFILLER_51_0 VPWR VGND sg13g2_decap_8
XFILLER_110_160 VPWR VGND sg13g2_decap_8
XFILLER_102_116 VPWR VGND sg13g2_decap_8
X_1318_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1249_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_155 VPWR VGND sg13g2_decap_8
XFILLER_101_193 VPWR VGND sg13g2_decap_8
XFILLER_30_103 VPWR VGND sg13g2_decap_4
X_0620_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q _0081_
+ _0082_ VPWR VGND sg13g2_nor2_1
X_0551_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q VPWR
+ _0024_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q
+ _0023_ sg13g2_o21ai_1
XFILLER_7_24 VPWR VGND sg13g2_fill_1
XFILLER_97_136 VPWR VGND sg13g2_decap_8
X_0482_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2
+ UIO_OUT_TT_PROJECT0 Tile_X0Y0_S1END[2] UIO_OUT_TT_PROJECT5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG2 VPWR VGND sg13g2_mux4_1
X_1103_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1034_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_0 VPWR VGND sg13g2_fill_2
X_0749_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q UO_OUT_TT_PROJECT1
+ _0156_ UO_OUT_TT_PROJECT5 _0349_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG13 VPWR VGND sg13g2_mux4_1
X_0818_ VGND VPWR _0200_ _0202_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG2
+ _0204_ sg13g2_a21oi_1
XFILLER_96_180 VPWR VGND sg13g2_decap_8
XFILLER_16_55 VPWR VGND sg13g2_fill_2
XFILLER_16_88 VPWR VGND sg13g2_fill_1
XFILLER_79_125 VPWR VGND sg13g2_decap_4
XFILLER_92_7 VPWR VGND sg13g2_decap_4
XFILLER_73_94 VPWR VGND sg13g2_fill_1
XFILLER_98_80 VPWR VGND sg13g2_fill_2
X_0603_ _0070_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_nand2b_1
X_0534_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit3.Q UIO_OUT_TT_PROJECT5
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG5 VPWR VGND sg13g2_mux4_1
X_1652_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG10 Tile_X0Y1_W6BEG[10]
+ VPWR VGND sg13g2_buf_1
X_1583_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameData_O[29] VPWR VGND sg13g2_buf_1
X_0465_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit21.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb6
+ Tile_X0Y0_S2MID[6] Tile_X0Y1_N2MID[6] Tile_X0Y0_S2END[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit20.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 VPWR VGND sg13g2_mux4_1
X_0396_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_mux4_1
XFILLER_14_0 VPWR VGND sg13g2_fill_2
X_1017_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_84_183 VPWR VGND sg13g2_decap_8
XFILLER_75_150 VPWR VGND sg13g2_fill_2
XFILLER_90_197 VPWR VGND sg13g2_fill_2
XFILLER_90_175 VPWR VGND sg13g2_fill_2
XFILLER_90_4 VPWR VGND sg13g2_fill_2
XFILLER_75_194 VPWR VGND sg13g2_decap_4
X_1497_ Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_8.A Tile_X0Y0_N4BEG[8] VPWR VGND sg13g2_buf_1
X_0517_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG5 VPWR VGND sg13g2_mux4_1
X_1635_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb1 Tile_X0Y1_W2BEGb[1]
+ VPWR VGND sg13g2_buf_1
X_1566_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameData_O[12] VPWR VGND sg13g2_buf_1
X_0379_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1 _0309_ VPWR VGND sg13g2_nor3_1
X_0448_ _0351_ _0354_ _0356_ VPWR VGND sg13g2_nor2b_1
XFILLER_81_197 VPWR VGND sg13g2_fill_2
XFILLER_1_124 VPWR VGND sg13g2_fill_1
XFILLER_54_41 VPWR VGND sg13g2_fill_1
X_1351_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1420_ Tile_X0Y0_FrameData[3] Tile_X0Y0_FrameData_O[3] VPWR VGND sg13g2_buf_1
X_1282_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_81_0 VPWR VGND sg13g2_decap_4
X_0997_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1618_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG0 Tile_X0Y1_S4BEG[12]
+ VPWR VGND sg13g2_buf_1
X_1549_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG11 Tile_X0Y0_WW4BEG[11]
+ VPWR VGND sg13g2_buf_1
XFILLER_54_131 VPWR VGND sg13g2_decap_8
XFILLER_54_175 VPWR VGND sg13g2_fill_2
XFILLER_40_32 VPWR VGND sg13g2_fill_1
XFILLER_40_54 VPWR VGND sg13g2_fill_1
XFILLER_108_199 VPWR VGND sg13g2_fill_1
XFILLER_40_76 VPWR VGND sg13g2_decap_4
XFILLER_45_120 VPWR VGND sg13g2_fill_2
XFILLER_49_96 VPWR VGND sg13g2_decap_8
X_0920_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_145 VPWR VGND sg13g2_fill_1
X_0851_ _0228_ VPWR UI_IN_TT_PROJECT4 VGND _0229_ _0231_ sg13g2_o21ai_1
X_0782_ _0152_ _0148_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ _0173_ VPWR VGND sg13g2_mux2_1
X_1334_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1265_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1403_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1196_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_175 VPWR VGND sg13g2_fill_2
XFILLER_51_145 VPWR VGND sg13g2_decap_8
XFILLER_105_169 VPWR VGND sg13g2_decap_8
XFILLER_86_17 VPWR VGND sg13g2_decap_4
XFILLER_10_68 VPWR VGND sg13g2_decap_4
XFILLER_42_123 VPWR VGND sg13g2_fill_2
XFILLER_104_191 VPWR VGND sg13g2_decap_8
XFILLER_32_9 VPWR VGND sg13g2_fill_1
X_1050_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_93 VPWR VGND sg13g2_fill_1
X_0834_ VPWR _0218_ _0217_ VGND sg13g2_inv_1
X_0903_ Tile_X0Y1_E2END[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q _0279_ VPWR
+ VGND sg13g2_nor3_1
X_0696_ _0127_ _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_0765_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q UO_OUT_TT_PROJECT3
+ _0154_ _0158_ _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit6.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG11 VPWR VGND sg13g2_mux4_1
XFILLER_44_0 VPWR VGND sg13g2_decap_8
XFILLER_110_183 VPWR VGND sg13g2_fill_1
X_1317_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1248_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1179_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_172 VPWR VGND sg13g2_decap_8
XFILLER_62_63 VPWR VGND sg13g2_decap_4
XFILLER_30_126 VPWR VGND sg13g2_fill_1
XFILLER_30_148 VPWR VGND sg13g2_fill_1
XFILLER_97_104 VPWR VGND sg13g2_fill_1
X_0550_ _0022_ VPWR _0023_ VGND Tile_X0Y0_E6END[9] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ sg13g2_o21ai_1
XFILLER_87_93 VPWR VGND sg13g2_fill_1
X_1102_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0481_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1
+ UIO_OUT_TT_PROJECT3 Tile_X0Y0_S1END[1] UIO_OUT_TT_PROJECT6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG1 VPWR VGND sg13g2_mux4_1
X_1033_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0817_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q _0203_
+ _0204_ VPWR VGND sg13g2_nor2_1
X_0748_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0318_ Tile_X0Y0_S4END[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit13.Q
+ _0156_ VPWR VGND sg13g2_mux4_1
X_0679_ UO_OUT_TT_PROJECT0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit17.Q _0116_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_20_181 VPWR VGND sg13g2_decap_8
XFILLER_32_77 VPWR VGND sg13g2_decap_8
XFILLER_32_88 VPWR VGND sg13g2_fill_1
XFILLER_57_85 VPWR VGND sg13g2_fill_2
XFILLER_73_40 VPWR VGND sg13g2_decap_8
X_1651_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG9 Tile_X0Y1_W6BEG[9]
+ VPWR VGND sg13g2_buf_1
X_0602_ VGND VPWR _0064_ _0067_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG2
+ _0069_ sg13g2_a21oi_1
X_0533_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q UIO_OUT_TT_PROJECT4
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG4 VPWR VGND sg13g2_mux4_1
X_0464_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit20.Q Tile_X0Y1_E2MID[1]
+ Tile_X0Y1_E2END[1] Tile_X0Y1_E6END[1] _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit21.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb6 VPWR VGND sg13g2_mux4_1
X_1582_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameData_O[28] VPWR VGND sg13g2_buf_1
X_0395_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 Tile_X0Y1_E6END[6]
+ _0321_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2
+ VPWR VGND sg13g2_mux4_1
X_1016_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_94_28 VPWR VGND sg13g2_decap_8
XFILLER_27_22 VPWR VGND sg13g2_fill_2
XFILLER_68_51 VPWR VGND sg13g2_decap_8
XFILLER_4_199 VPWR VGND sg13g2_fill_1
XFILLER_4_188 VPWR VGND sg13g2_decap_8
XFILLER_4_15 VPWR VGND sg13g2_fill_2
XFILLER_75_173 VPWR VGND sg13g2_decap_8
XFILLER_69_2 VPWR VGND sg13g2_fill_1
X_1634_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb0 Tile_X0Y1_W2BEGb[0]
+ VPWR VGND sg13g2_buf_1
X_0516_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q UIO_OUT_TT_PROJECT5
+ UIO_OE_TT_PROJECT1 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG9 VPWR VGND sg13g2_mux4_1
X_1496_ Tile_X0Y1_N4END[15] Tile_X0Y0_N4BEG[7] VPWR VGND sg13g2_buf_1
X_0447_ _0355_ _0354_ _0351_ VPWR VGND sg13g2_nand2b_1
X_1565_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_81_176 VPWR VGND sg13g2_decap_8
XFILLER_81_132 VPWR VGND sg13g2_decap_8
X_0378_ _0308_ Tile_X0Y0_S1END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_66_173 VPWR VGND sg13g2_fill_1
XFILLER_72_143 VPWR VGND sg13g2_fill_1
X_1281_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1350_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_7 VPWR VGND sg13g2_decap_4
XFILLER_0_191 VPWR VGND sg13g2_decap_8
XFILLER_74_0 VPWR VGND sg13g2_decap_4
X_0996_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1617_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG3 Tile_X0Y1_S4BEG[11]
+ VPWR VGND sg13g2_buf_1
X_1479_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG6 Tile_X0Y0_N2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1548_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG10 Tile_X0Y0_WW4BEG[10]
+ VPWR VGND sg13g2_buf_1
XFILLER_54_198 VPWR VGND sg13g2_fill_2
XFILLER_108_134 VPWR VGND sg13g2_fill_1
XFILLER_108_123 VPWR VGND sg13g2_decap_8
XFILLER_49_64 VPWR VGND sg13g2_fill_1
XFILLER_105_92 VPWR VGND sg13g2_decap_8
XFILLER_45_132 VPWR VGND sg13g2_fill_2
XFILLER_45_176 VPWR VGND sg13g2_decap_8
X_0850_ _0230_ VPWR _0231_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
+ _0154_ sg13g2_o21ai_1
X_0781_ VGND VPWR _0167_ _0170_ Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_9.A _0172_ sg13g2_a21oi_1
X_1402_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1333_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1264_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_39 VPWR VGND sg13g2_fill_1
X_1195_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_113 VPWR VGND sg13g2_decap_4
XFILLER_51_124 VPWR VGND sg13g2_decap_8
X_0979_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_105_148 VPWR VGND sg13g2_decap_8
XFILLER_27_187 VPWR VGND sg13g2_decap_8
XFILLER_27_198 VPWR VGND sg13g2_fill_2
XFILLER_35_66 VPWR VGND sg13g2_decap_8
XFILLER_42_113 VPWR VGND sg13g2_fill_2
XFILLER_4_0 VPWR VGND sg13g2_fill_2
XFILLER_51_87 VPWR VGND sg13g2_decap_8
XFILLER_104_170 VPWR VGND sg13g2_decap_8
X_0833_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q Tile_X0Y1_EE4END[1]
+ Tile_X0Y1_EE4END[9] Tile_X0Y1_E6END[1] Tile_X0Y1_E6END[9] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q
+ _0217_ VPWR VGND sg13g2_mux4_1
X_0902_ _0278_ _0265_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0
+ VPWR VGND sg13g2_nand2b_1
X_0764_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit5.Q UO_OUT_TT_PROJECT2
+ _0153_ _0157_ _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit4.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG10 VPWR VGND sg13g2_mux4_1
X_0695_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q
+ _0126_ _0125_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG5 _0348_ sg13g2_a221oi_1
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_2_70 VPWR VGND sg13g2_fill_2
X_1316_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1247_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1178_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_101_151 VPWR VGND sg13g2_decap_8
XFILLER_15_124 VPWR VGND sg13g2_decap_4
X_0480_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0
+ UIO_OUT_TT_PROJECT2 Tile_X0Y0_S1END[0] UIO_OUT_TT_PROJECT7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
X_1101_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1032_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_190 VPWR VGND sg13g2_decap_8
X_0747_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT4 _0155_ _0356_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG12 VPWR VGND sg13g2_mux4_1
X_0816_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_EE4END[14] Tile_X0Y1_E6END[6] _0156_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
+ _0203_ VPWR VGND sg13g2_mux4_1
XFILLER_88_138 VPWR VGND sg13g2_fill_2
X_0678_ _0115_ _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_16_57 VPWR VGND sg13g2_fill_1
XFILLER_16_79 VPWR VGND sg13g2_decap_8
XFILLER_94_108 VPWR VGND sg13g2_fill_2
XFILLER_73_85 VPWR VGND sg13g2_decap_8
X_0601_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit11.Q _0068_
+ _0069_ VPWR VGND sg13g2_nor2_1
XFILLER_11_171 VPWR VGND sg13g2_fill_1
XFILLER_7_197 VPWR VGND sg13g2_fill_2
X_1650_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG8 Tile_X0Y1_W6BEG[8]
+ VPWR VGND sg13g2_buf_1
X_1581_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameData_O[27] VPWR VGND sg13g2_buf_1
X_0532_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q Tile_X0Y1_N4END[7]
+ Tile_X0Y0_S4END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG3 VPWR VGND sg13g2_mux4_1
X_0394_ VPWR VGND _0319_ _0320_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q
+ _0298_ _0321_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
+ sg13g2_a221oi_1
X_0463_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q Tile_X0Y1_N2MID[6]
+ Tile_X0Y1_N2END[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG6
+ Tile_X0Y0_S2MID[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q
+ _0002_ VPWR VGND sg13g2_mux4_1
X_1015_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_45 VPWR VGND sg13g2_fill_2
XFILLER_43_22 VPWR VGND sg13g2_fill_2
XFILLER_108_81 VPWR VGND sg13g2_decap_8
XFILLER_4_167 VPWR VGND sg13g2_decap_8
XFILLER_90_111 VPWR VGND sg13g2_fill_1
XFILLER_75_152 VPWR VGND sg13g2_fill_1
XFILLER_90_199 VPWR VGND sg13g2_fill_1
X_1633_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG7 Tile_X0Y1_W2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1564_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameData_O[10] VPWR VGND sg13g2_buf_1
XFILLER_104_17 VPWR VGND sg13g2_decap_8
X_0515_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_66_152 VPWR VGND sg13g2_decap_4
X_1495_ Tile_X0Y1_N4END[14] Tile_X0Y0_N4BEG[6] VPWR VGND sg13g2_buf_1
X_0446_ _0352_ _0353_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q
+ _0354_ VPWR VGND sg13g2_nand3_1
X_0377_ VPWR _0307_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit7.Q
+ VGND sg13g2_inv_1
XFILLER_81_199 VPWR VGND sg13g2_fill_1
XFILLER_89_29 VPWR VGND sg13g2_fill_1
XFILLER_54_32 VPWR VGND sg13g2_decap_4
XFILLER_57_130 VPWR VGND sg13g2_fill_2
XFILLER_70_42 VPWR VGND sg13g2_decap_8
X_1280_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_170 VPWR VGND sg13g2_decap_8
XFILLER_63_199 VPWR VGND sg13g2_fill_1
XFILLER_48_174 VPWR VGND sg13g2_decap_8
X_0995_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_0 VPWR VGND sg13g2_fill_2
X_1547_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG9 Tile_X0Y0_WW4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_1616_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG2 Tile_X0Y1_S4BEG[10]
+ VPWR VGND sg13g2_buf_1
X_1478_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG5 Tile_X0Y0_N2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0429_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y0_E2MID[6]
+ Tile_X0Y0_E2END[6] Tile_X0Y0_E6END[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit19.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_54_177 VPWR VGND sg13g2_fill_1
XFILLER_108_157 VPWR VGND sg13g2_decap_8
XFILLER_108_102 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_4
XFILLER_105_71 VPWR VGND sg13g2_decap_8
XFILLER_65_64 VPWR VGND sg13g2_fill_2
X_0780_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q _0171_
+ _0172_ VPWR VGND sg13g2_nor2_1
XFILLER_107_190 VPWR VGND sg13g2_decap_8
X_1401_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1332_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1194_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1263_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_199 VPWR VGND sg13g2_fill_1
X_0978_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_105_127 VPWR VGND sg13g2_decap_8
XFILLER_19_35 VPWR VGND sg13g2_decap_8
XFILLER_51_66 VPWR VGND sg13g2_fill_1
XFILLER_18_155 VPWR VGND sg13g2_decap_8
XFILLER_18_199 VPWR VGND sg13g2_fill_1
X_0763_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit3.Q UO_OUT_TT_PROJECT1
+ _0152_ _0156_ _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit2.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG9 VPWR VGND sg13g2_mux4_1
X_0832_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q _0215_
+ _0216_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q
+ sg13g2_nand3b_1
X_0901_ _0276_ VPWR _0277_ VGND _0267_ _0269_ sg13g2_o21ai_1
X_1315_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0694_ UO_OUT_TT_PROJECT5 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q _0126_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_110_174 VPWR VGND sg13g2_fill_2
XFILLER_24_125 VPWR VGND sg13g2_fill_2
X_1246_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1177_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_10 VPWR VGND Tile_X0Y1_FrameStrobe[18] sg13g2_antennanp
XFILLER_32_191 VPWR VGND sg13g2_decap_8
XFILLER_21_25 VPWR VGND sg13g2_fill_1
XFILLER_101_130 VPWR VGND sg13g2_decap_8
XFILLER_15_147 VPWR VGND sg13g2_decap_8
XFILLER_23_191 VPWR VGND sg13g2_decap_8
X_1100_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1031_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_17 VPWR VGND sg13g2_decap_8
X_0815_ VGND VPWR Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
+ _0201_ _0202_ _0303_ sg13g2_a21oi_1
X_0746_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0325_ Tile_X0Y0_S4END[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q
+ _0155_ VPWR VGND sg13g2_mux4_1
XFILLER_96_194 VPWR VGND sg13g2_decap_4
X_0677_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit15.Q Tile_X0Y1_N1END[3]
+ UO_OUT_TT_PROJECT1 _0325_ UO_OUT_TT_PROJECT4 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit14.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG3 VPWR VGND sg13g2_mux4_1
X_1229_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_87_172 VPWR VGND sg13g2_fill_2
XFILLER_57_65 VPWR VGND sg13g2_decap_8
XFILLER_57_87 VPWR VGND sg13g2_fill_1
XFILLER_11_150 VPWR VGND sg13g2_fill_2
X_0600_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit10.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_EE4END[14] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ _0068_ VPWR VGND sg13g2_mux4_1
X_0531_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q Tile_X0Y1_N4END[6]
+ Tile_X0Y0_S4END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG2 VPWR VGND sg13g2_mux4_1
XFILLER_7_165 VPWR VGND sg13g2_fill_1
X_1580_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameData_O[26] VPWR VGND sg13g2_buf_1
X_0462_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit0.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E2MID[1] Tile_X0Y0_E2END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit1.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG6
+ VPWR VGND sg13g2_mux4_1
X_0393_ Tile_X0Y1_N1END[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit29.Q _0320_ VPWR
+ VGND sg13g2_nor3_1
X_1014_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_81 VPWR VGND sg13g2_fill_2
X_0729_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q UO_OUT_TT_PROJECT3
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 UO_OUT_TT_PROJECT7
+ _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_84_197 VPWR VGND sg13g2_fill_2
XFILLER_68_86 VPWR VGND sg13g2_decap_8
XFILLER_84_85 VPWR VGND sg13g2_fill_2
X_0514_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit8.Q UIO_OUT_TT_PROJECT4
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG8 VPWR VGND sg13g2_mux4_1
X_1632_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG6 Tile_X0Y1_W2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1494_ Tile_X0Y1_N4END[13] Tile_X0Y0_N4BEG[5] VPWR VGND sg13g2_buf_1
X_1563_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_66_120 VPWR VGND sg13g2_decap_4
XFILLER_12_0 VPWR VGND sg13g2_fill_2
X_0376_ VPWR _0306_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ VGND sg13g2_inv_1
X_0445_ _0353_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
+ Tile_X0Y0_S2MID[3] VPWR VGND sg13g2_nand2_1
XFILLER_81_156 VPWR VGND sg13g2_fill_2
XFILLER_13_26 VPWR VGND sg13g2_decap_4
XFILLER_72_178 VPWR VGND sg13g2_decap_8
XFILLER_72_123 VPWR VGND sg13g2_fill_1
XFILLER_38_78 VPWR VGND sg13g2_fill_2
XFILLER_57_175 VPWR VGND sg13g2_fill_1
XFILLER_57_197 VPWR VGND sg13g2_fill_2
XFILLER_110_83 VPWR VGND sg13g2_decap_8
XFILLER_95_51 VPWR VGND sg13g2_fill_2
XFILLER_48_153 VPWR VGND sg13g2_decap_8
XFILLER_63_167 VPWR VGND sg13g2_decap_8
XFILLER_63_145 VPWR VGND sg13g2_decap_4
XFILLER_48_197 VPWR VGND sg13g2_fill_2
X_0994_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1477_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG4 Tile_X0Y0_N2BEG[4]
+ VPWR VGND sg13g2_buf_1
X_1546_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG8 Tile_X0Y0_WW4BEG[8]
+ VPWR VGND sg13g2_buf_1
X_1615_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG1 Tile_X0Y1_S4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_0359_ VPWR _0289_ Tile_X0Y0_E6END[3] VGND sg13g2_inv_1
X_0428_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb1
+ Tile_X0Y0_S2MID[1] Tile_X0Y1_N2MID[1] Tile_X0Y0_S2END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_54_145 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_decap_4
XFILLER_24_69 VPWR VGND sg13g2_decap_8
XFILLER_60_115 VPWR VGND sg13g2_fill_2
X_1331_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1400_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1262_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_112 VPWR VGND sg13g2_fill_1
X_1193_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_159 VPWR VGND sg13g2_decap_8
XFILLER_105_106 VPWR VGND sg13g2_decap_8
X_0977_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1529_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG3 Tile_X0Y0_W6BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_27_123 VPWR VGND sg13g2_decap_4
XFILLER_50_170 VPWR VGND sg13g2_decap_8
XFILLER_104_150 VPWR VGND sg13g2_fill_2
XFILLER_4_2 VPWR VGND sg13g2_fill_1
XFILLER_41_192 VPWR VGND sg13g2_decap_8
X_0900_ VPWR VGND _0265_ _0271_ _0275_ _0266_ _0276_ _0273_ sg13g2_a221oi_1
X_0693_ _0125_ _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_nand2b_1
X_0762_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q UO_OUT_TT_PROJECT0
+ _0151_ _0155_ _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG8 VPWR VGND sg13g2_mux4_1
X_0831_ _0157_ _0149_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q
+ _0215_ VPWR VGND sg13g2_mux2_1
XFILLER_110_153 VPWR VGND sg13g2_decap_8
XFILLER_102_109 VPWR VGND sg13g2_decap_8
X_1314_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_24_148 VPWR VGND sg13g2_decap_8
X_1245_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1176_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_11 VPWR VGND Tile_X0Y1_FrameStrobe[8] sg13g2_antennanp
XFILLER_32_170 VPWR VGND sg13g2_decap_8
XFILLER_101_186 VPWR VGND sg13g2_decap_8
XFILLER_102_95 VPWR VGND sg13g2_decap_8
XFILLER_97_129 VPWR VGND sg13g2_decap_8
XFILLER_11_92 VPWR VGND sg13g2_fill_2
X_1030_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0814_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 _0002_
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q _0201_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_88_107 VPWR VGND sg13g2_decap_4
X_0676_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit13.Q Tile_X0Y1_N1END[2]
+ UO_OUT_TT_PROJECT0 _0318_ UO_OUT_TT_PROJECT5 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit12.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG2 VPWR VGND sg13g2_mux4_1
X_0745_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit7.Q UO_OUT_TT_PROJECT3
+ _0154_ UO_OUT_TT_PROJECT7 _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit6.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG11 VPWR VGND sg13g2_mux4_1
XFILLER_42_0 VPWR VGND sg13g2_decap_8
XFILLER_96_173 VPWR VGND sg13g2_decap_8
X_1228_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1159_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_195 VPWR VGND sg13g2_decap_4
XFILLER_79_129 VPWR VGND sg13g2_fill_2
X_0530_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q Tile_X0Y1_N4END[5]
+ Tile_X0Y0_S4END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG1 VPWR VGND sg13g2_mux4_1
XFILLER_7_199 VPWR VGND sg13g2_fill_1
X_0461_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit26.Q Tile_X0Y0_E2MID[2]
+ Tile_X0Y0_E2END[2] Tile_X0Y0_E6END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit27.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG5
+ VPWR VGND sg13g2_mux4_1
X_0392_ _0319_ _0318_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_93_187 VPWR VGND sg13g2_fill_2
X_1013_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0659_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q _0110_
+ _0111_ _0114_ VPWR VGND sg13g2_nor3_1
X_0728_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT6 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13
+ _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_84_176 VPWR VGND sg13g2_decap_8
XFILLER_108_61 VPWR VGND sg13g2_fill_2
XFILLER_75_143 VPWR VGND sg13g2_decap_8
XFILLER_90_157 VPWR VGND sg13g2_fill_1
XFILLER_75_198 VPWR VGND sg13g2_fill_2
XFILLER_75_187 VPWR VGND sg13g2_decap_8
XFILLER_83_7 VPWR VGND sg13g2_fill_2
X_1631_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG5 Tile_X0Y1_W2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0513_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7 VPWR VGND sg13g2_mux4_1
X_1493_ Tile_X0Y1_N4END[12] Tile_X0Y0_N4BEG[4] VPWR VGND sg13g2_buf_1
X_1562_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameData_O[8] VPWR VGND sg13g2_buf_1
X_0444_ _0352_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG3 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
+ VPWR VGND sg13g2_nand2b_1
X_0375_ VPWR _0305_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ VGND sg13g2_inv_1
XFILLER_1_117 VPWR VGND sg13g2_fill_2
XFILLER_57_132 VPWR VGND sg13g2_fill_1
XFILLER_110_62 VPWR VGND sg13g2_decap_8
XFILLER_28_90 VPWR VGND sg13g2_decap_8
XFILLER_81_4 VPWR VGND sg13g2_fill_1
X_0993_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_67_2 VPWR VGND sg13g2_fill_1
X_1614_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG0 Tile_X0Y1_S4BEG[8]
+ VPWR VGND sg13g2_buf_1
X_1476_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG3 Tile_X0Y0_N2BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1545_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG7 Tile_X0Y0_WW4BEG[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_5_72 VPWR VGND sg13g2_fill_2
X_0427_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y1_E2MID[6]
+ Tile_X0Y1_E2END[6] Tile_X0Y1_E6END[6] _0342_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit11.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb1 VPWR VGND sg13g2_mux4_1
X_0358_ VPWR _0288_ Tile_X0Y0_E6END[2] VGND sg13g2_inv_1
XFILLER_39_176 VPWR VGND sg13g2_fill_2
XFILLER_39_198 VPWR VGND sg13g2_fill_2
XFILLER_54_124 VPWR VGND sg13g2_decap_8
XFILLER_54_168 VPWR VGND sg13g2_decap_8
XFILLER_1_19 VPWR VGND sg13g2_fill_1
XFILLER_60_138 VPWR VGND sg13g2_decap_8
X_1330_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1261_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1192_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_0976_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_72_0 VPWR VGND sg13g2_fill_2
XFILLER_51_138 VPWR VGND sg13g2_decap_8
X_1459_ Tile_X0Y1_FrameStrobe[10] Tile_X0Y0_FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
X_1528_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG2 Tile_X0Y0_W6BEG[2]
+ VPWR VGND sg13g2_buf_1
XFILLER_50_193 VPWR VGND sg13g2_decap_8
XFILLER_104_184 VPWR VGND sg13g2_decap_8
XFILLER_76_98 VPWR VGND sg13g2_decap_4
X_0830_ _0213_ _0214_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit10.Q
+ UI_IN_TT_PROJECT0 VPWR VGND sg13g2_mux2_1
XFILLER_41_171 VPWR VGND sg13g2_decap_8
X_0692_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q
+ _0124_ _0123_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG4 _0355_ sg13g2_a221oi_1
X_0761_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q UO_OUT_TT_PROJECT7
+ _0150_ _0154_ _0356_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG7 VPWR VGND sg13g2_mux4_1
XFILLER_110_198 VPWR VGND sg13g2_fill_2
XFILLER_110_187 VPWR VGND sg13g2_fill_1
XFILLER_110_132 VPWR VGND sg13g2_decap_8
X_1313_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_1244_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1175_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_12 VPWR VGND Tile_X0Y1_FrameStrobe[9] sg13g2_antennanp
X_0959_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_182 VPWR VGND sg13g2_decap_8
XFILLER_101_165 VPWR VGND sg13g2_decap_8
XFILLER_62_89 VPWR VGND sg13g2_decap_4
XFILLER_62_67 VPWR VGND sg13g2_fill_1
XFILLER_2_0 VPWR VGND sg13g2_fill_2
XFILLER_87_75 VPWR VGND sg13g2_fill_2
X_0813_ _0200_ _0199_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_nand2b_1
X_0675_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q Tile_X0Y1_N1END[1]
+ UO_OUT_TT_PROJECT3 _0311_ UO_OUT_TT_PROJECT6 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG1 VPWR VGND sg13g2_mux4_1
X_0744_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0007_ Tile_X0Y0_S4END[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q
+ _0154_ VPWR VGND sg13g2_mux4_1
XFILLER_96_152 VPWR VGND sg13g2_decap_8
X_1158_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1227_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_1089_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_87_174 VPWR VGND sg13g2_fill_1
XFILLER_11_196 VPWR VGND sg13g2_decap_4
XFILLER_7_145 VPWR VGND sg13g2_fill_2
X_0460_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit19.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb5
+ Tile_X0Y0_S2MID[5] Tile_X0Y1_N2MID[5] Tile_X0Y0_S2END[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit18.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 VPWR VGND sg13g2_mux4_1
X_0391_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_E6END[10] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14
+ _0317_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q _0318_
+ VPWR VGND sg13g2_mux4_1
X_1012_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_93_199 VPWR VGND sg13g2_fill_1
X_0727_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit19.Q UO_OUT_TT_PROJECT1
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 UO_OUT_TT_PROJECT5
+ _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit18.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG1
+ VPWR VGND sg13g2_mux4_1
X_0658_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q _0112_
+ _0113_ VPWR VGND sg13g2_nor2b_1
X_0589_ _0057_ VPWR _0058_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ _0013_ sg13g2_o21ai_1
XFILLER_84_199 VPWR VGND sg13g2_fill_1
XFILLER_108_95 VPWR VGND sg13g2_decap_8
XFILLER_68_44 VPWR VGND sg13g2_decap_8
XFILLER_17_81 VPWR VGND sg13g2_fill_2
X_1630_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG4 Tile_X0Y1_W2BEG[4]
+ VPWR VGND sg13g2_buf_1
X_0512_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit6.Q UIO_OUT_TT_PROJECT7
+ UIO_OE_TT_PROJECT3 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit7.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG7 VPWR VGND sg13g2_mux4_1
X_1492_ Tile_X0Y1_N4END[11] Tile_X0Y0_N4BEG[3] VPWR VGND sg13g2_buf_1
X_0374_ VPWR _0304_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q
+ VGND sg13g2_inv_1
X_0443_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit15.Q _0350_
+ _0351_ VPWR VGND sg13g2_nor2_1
X_1561_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameData_O[7] VPWR VGND sg13g2_buf_1
XFILLER_81_158 VPWR VGND sg13g2_fill_1
XFILLER_66_199 VPWR VGND sg13g2_fill_1
XFILLER_1_129 VPWR VGND sg13g2_fill_2
XFILLER_110_41 VPWR VGND sg13g2_decap_8
XFILLER_57_199 VPWR VGND sg13g2_fill_1
XFILLER_70_56 VPWR VGND sg13g2_fill_1
XFILLER_0_140 VPWR VGND sg13g2_fill_2
XFILLER_0_151 VPWR VGND sg13g2_fill_1
XFILLER_0_184 VPWR VGND sg13g2_decap_8
XFILLER_48_199 VPWR VGND sg13g2_fill_1
X_0992_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1613_ Tile_X0Y0_S4END[15] Tile_X0Y1_S4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_74_4 VPWR VGND sg13g2_fill_2
X_1544_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG6 Tile_X0Y0_WW4BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1475_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG2 Tile_X0Y0_N2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0357_ VPWR _0287_ Tile_X0Y0_E6END[1] VGND sg13g2_inv_1
X_0426_ _0337_ _0340_ _0342_ VPWR VGND sg13g2_nor2b_1
XFILLER_39_111 VPWR VGND sg13g2_fill_1
XFILLER_39_155 VPWR VGND sg13g2_decap_4
XFILLER_108_116 VPWR VGND sg13g2_decap_8
XFILLER_105_85 VPWR VGND sg13g2_decap_8
XFILLER_45_169 VPWR VGND sg13g2_decap_8
XFILLER_81_22 VPWR VGND sg13g2_decap_8
XFILLER_53_180 VPWR VGND sg13g2_decap_4
XFILLER_107_182 VPWR VGND sg13g2_fill_1
X_1260_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1191_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_117 VPWR VGND sg13g2_fill_2
X_0975_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_0 VPWR VGND sg13g2_fill_2
X_1527_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG1 Tile_X0Y0_W6BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1458_ Tile_X0Y1_FrameStrobe[9] Tile_X0Y0_FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
X_1389_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0409_ Tile_X0Y1_N2MID[0] Tile_X0Y1_N2END[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit8.Q
+ _0329_ VPWR VGND sg13g2_mux2_1
XFILLER_35_48 VPWR VGND sg13g2_fill_1
XFILLER_42_106 VPWR VGND sg13g2_decap_8
XFILLER_104_163 VPWR VGND sg13g2_decap_8
XFILLER_26_191 VPWR VGND sg13g2_decap_8
XFILLER_33_106 VPWR VGND sg13g2_decap_4
X_0760_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q UO_OUT_TT_PROJECT6
+ _0149_ _0153_ _0349_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG6 VPWR VGND sg13g2_mux4_1
X_0691_ UO_OUT_TT_PROJECT4 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q _0124_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_41_80 VPWR VGND sg13g2_fill_2
XFILLER_110_111 VPWR VGND sg13g2_decap_8
X_1312_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_1243_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1174_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_13 VPWR VGND Tile_X0Y1_N2MID[5] sg13g2_antennanp
X_0958_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0889_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit6.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit5.Q
+ _0265_ VPWR VGND sg13g2_nor2b_1
XFILLER_101_144 VPWR VGND sg13g2_decap_8
XFILLER_99_161 VPWR VGND sg13g2_decap_8
XFILLER_15_128 VPWR VGND sg13g2_fill_2
XFILLER_11_94 VPWR VGND sg13g2_fill_1
XFILLER_11_50 VPWR VGND sg13g2_fill_2
X_0743_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit4.Q UO_OUT_TT_PROJECT2
+ UO_OUT_TT_PROJECT6 _0153_ _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit5.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG10 VPWR VGND sg13g2_mux4_1
X_0812_ _0152_ _0148_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q
+ _0199_ VPWR VGND sg13g2_mux2_1
XFILLER_96_131 VPWR VGND sg13g2_decap_8
X_0674_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q Tile_X0Y1_N1END[0]
+ UO_OUT_TT_PROJECT2 _0007_ UO_OUT_TT_PROJECT7 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG0 VPWR VGND sg13g2_mux4_1
X_1157_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1226_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1088_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_87_197 VPWR VGND sg13g2_fill_2
XFILLER_57_79 VPWR VGND sg13g2_fill_2
X_0390_ VPWR VGND _0315_ _0316_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q
+ _0288_ _0317_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q
+ sg13g2_a221oi_1
XFILLER_78_197 VPWR VGND sg13g2_fill_2
X_1011_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0726_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit16.Q UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT4 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15
+ _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit17.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG0
+ VPWR VGND sg13g2_mux4_1
X_0657_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_EE4END[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit7.Q
+ _0112_ VPWR VGND sg13g2_mux4_1
X_0588_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q _0056_
+ _0057_ VPWR VGND sg13g2_and2_1
XFILLER_69_197 VPWR VGND sg13g2_fill_2
X_1209_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_48 VPWR VGND sg13g2_fill_2
XFILLER_108_74 VPWR VGND sg13g2_decap_8
XFILLER_4_116 VPWR VGND sg13g2_decap_4
XFILLER_83_9 VPWR VGND sg13g2_fill_1
X_0511_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 VPWR VGND sg13g2_mux4_1
X_1560_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameData_O[6] VPWR VGND sg13g2_buf_1
XFILLER_66_145 VPWR VGND sg13g2_decap_8
XFILLER_3_193 VPWR VGND sg13g2_decap_8
X_1491_ Tile_X0Y1_N4END[10] Tile_X0Y0_N4BEG[2] VPWR VGND sg13g2_buf_1
X_0373_ VPWR _0303_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q
+ VGND sg13g2_inv_1
X_0442_ Tile_X0Y1_N2MID[3] Tile_X0Y1_N2END[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit14.Q
+ _0350_ VPWR VGND sg13g2_mux2_1
X_0709_ UO_OUT_TT_PROJECT2 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit5.Q _0136_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_1_119 VPWR VGND sg13g2_fill_1
XFILLER_38_59 VPWR VGND sg13g2_fill_2
XFILLER_54_36 VPWR VGND sg13g2_fill_2
XFILLER_110_97 VPWR VGND sg13g2_decap_8
XFILLER_0_163 VPWR VGND sg13g2_decap_8
XFILLER_48_167 VPWR VGND sg13g2_decap_8
X_0991_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1474_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG1 Tile_X0Y0_N2BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1612_ Tile_X0Y0_S4END[14] Tile_X0Y1_S4BEG[6] VPWR VGND sg13g2_buf_1
X_1543_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG5 Tile_X0Y0_WW4BEG[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_5_74 VPWR VGND sg13g2_fill_1
XFILLER_10_0 VPWR VGND sg13g2_fill_2
X_0425_ _0341_ _0340_ _0337_ VPWR VGND sg13g2_nand2b_1
XFILLER_54_159 VPWR VGND sg13g2_decap_4
XFILLER_49_25 VPWR VGND sg13g2_fill_1
XFILLER_105_64 VPWR VGND sg13g2_decap_8
XFILLER_65_57 VPWR VGND sg13g2_decap_8
XFILLER_14_94 VPWR VGND sg13g2_fill_2
X_1190_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_44_170 VPWR VGND sg13g2_decap_8
X_0974_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1457_ Tile_X0Y1_FrameStrobe[8] Tile_X0Y0_FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_1526_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG0 Tile_X0Y0_W6BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_58_0 VPWR VGND sg13g2_fill_2
X_0408_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q Tile_X0Y0_E2MID[7]
+ Tile_X0Y0_E2END[7] Tile_X0Y0_E6END[8] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0
+ VPWR VGND sg13g2_mux4_1
XFILLER_27_104 VPWR VGND sg13g2_fill_2
X_1388_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_27_148 VPWR VGND sg13g2_fill_1
XFILLER_35_170 VPWR VGND sg13g2_decap_4
XFILLER_50_184 VPWR VGND sg13g2_decap_4
XFILLER_92_33 VPWR VGND sg13g2_decap_4
XFILLER_92_11 VPWR VGND sg13g2_fill_1
XFILLER_18_148 VPWR VGND sg13g2_decap_8
XFILLER_33_129 VPWR VGND sg13g2_decap_4
X_0690_ _0123_ _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
X_1311_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_110_167 VPWR VGND sg13g2_decap_8
X_1242_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1173_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_14 VPWR VGND Tile_X0Y1_N2MID[5] sg13g2_antennanp
XFILLER_17_170 VPWR VGND sg13g2_fill_2
XFILLER_32_184 VPWR VGND sg13g2_decap_8
X_0957_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0888_ VPWR ENA_TT_PROJECT _0264_ VGND sg13g2_inv_1
XFILLER_101_123 VPWR VGND sg13g2_decap_8
XFILLER_99_140 VPWR VGND sg13g2_decap_8
X_1509_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG3 Tile_X0Y0_W1BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_102_21 VPWR VGND sg13g2_fill_1
XFILLER_23_184 VPWR VGND sg13g2_decap_8
XFILLER_87_22 VPWR VGND sg13g2_fill_2
XFILLER_2_2 VPWR VGND sg13g2_fill_1
XFILLER_14_151 VPWR VGND sg13g2_fill_1
XFILLER_36_70 VPWR VGND sg13g2_fill_1
X_0742_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0311_ Tile_X0Y0_S4END[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q
+ _0153_ VPWR VGND sg13g2_mux4_1
X_0673_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit27.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_E2END[0] Tile_X0Y1_E2MID[0] _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit26.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG7 VPWR VGND sg13g2_mux4_1
X_0811_ VGND VPWR _0194_ _0196_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG1
+ _0198_ sg13g2_a21oi_1
XFILLER_96_187 VPWR VGND sg13g2_decap_8
XFILLER_96_198 VPWR VGND sg13g2_fill_2
X_1156_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1225_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1087_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_7_147 VPWR VGND sg13g2_fill_1
XFILLER_98_76 VPWR VGND sg13g2_decap_4
XFILLER_93_113 VPWR VGND sg13g2_fill_1
XFILLER_93_102 VPWR VGND sg13g2_decap_8
XFILLER_78_110 VPWR VGND sg13g2_fill_1
X_1010_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0656_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q VPWR
+ _0111_ VGND Tile_X0Y0_EE4END[15] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q
+ sg13g2_o21ai_1
X_0725_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q
+ _0146_ _0145_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb7 _0334_ sg13g2_a221oi_1
X_0587_ _0056_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 VPWR VGND sg13g2_nand2b_1
XFILLER_69_176 VPWR VGND sg13g2_decap_4
X_1208_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1139_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_75_102 VPWR VGND sg13g2_fill_2
XFILLER_68_79 VPWR VGND sg13g2_decap_8
XFILLER_17_83 VPWR VGND sg13g2_fill_1
X_0510_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit4.Q UIO_OUT_TT_PROJECT6
+ UIO_OE_TT_PROJECT2 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit5.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_3_172 VPWR VGND sg13g2_decap_8
X_1490_ Tile_X0Y1_N4END[9] Tile_X0Y0_N4BEG[1] VPWR VGND sg13g2_buf_1
X_0441_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit26.Q Tile_X0Y0_E2MID[4]
+ Tile_X0Y0_E2END[4] Tile_X0Y0_E6END[11] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit27.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG3
+ VPWR VGND sg13g2_mux4_1
X_0372_ VPWR _0302_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q
+ VGND sg13g2_inv_1
XFILLER_88_0 VPWR VGND sg13g2_decap_8
X_0639_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_EE4END[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit30.Q
+ _0097_ VPWR VGND sg13g2_mux4_1
X_0708_ _0135_ _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_110_76 VPWR VGND sg13g2_decap_8
XFILLER_80_182 VPWR VGND sg13g2_decap_8
XFILLER_54_59 VPWR VGND sg13g2_decap_8
XFILLER_0_142 VPWR VGND sg13g2_fill_1
XFILLER_48_102 VPWR VGND sg13g2_fill_1
XFILLER_48_146 VPWR VGND sg13g2_decap_8
XFILLER_63_149 VPWR VGND sg13g2_fill_1
XFILLER_28_60 VPWR VGND sg13g2_decap_8
X_1611_ Tile_X0Y0_S4END[13] Tile_X0Y1_S4BEG[5] VPWR VGND sg13g2_buf_1
X_0990_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1473_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG0 Tile_X0Y0_N2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1542_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG4 Tile_X0Y0_WW4BEG[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_5_97 VPWR VGND sg13g2_fill_1
X_0424_ _0338_ _0339_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q
+ _0340_ VPWR VGND sg13g2_nand3_1
XFILLER_54_138 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_24_29 VPWR VGND sg13g2_fill_2
XFILLER_105_21 VPWR VGND sg13g2_decap_4
XFILLER_107_173 VPWR VGND sg13g2_fill_2
XFILLER_107_162 VPWR VGND sg13g2_decap_8
X_0973_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1456_ Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
X_0407_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E6END[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15
+ _0324_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG3
+ VPWR VGND sg13g2_mux4_1
X_1525_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb7 Tile_X0Y0_W2BEGb[7]
+ VPWR VGND sg13g2_buf_1
X_1387_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_42_119 VPWR VGND sg13g2_decap_4
XFILLER_50_163 VPWR VGND sg13g2_decap_8
XFILLER_104_143 VPWR VGND sg13g2_decap_8
XFILLER_104_198 VPWR VGND sg13g2_fill_2
XFILLER_76_24 VPWR VGND sg13g2_fill_2
XFILLER_41_185 VPWR VGND sg13g2_decap_8
XFILLER_110_146 VPWR VGND sg13g2_decap_8
X_1310_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1241_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_44_7 VPWR VGND sg13g2_fill_2
XFILLER_110_179 VPWR VGND sg13g2_fill_1
X_1172_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_0956_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_32_141 VPWR VGND sg13g2_fill_2
XANTENNA_15 VPWR VGND Tile_X0Y1_N2MID[5] sg13g2_antennanp
X_0887_ _0263_ VPWR _0264_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q
+ _0254_ sg13g2_o21ai_1
XFILLER_101_179 VPWR VGND sg13g2_decap_8
XFILLER_101_102 VPWR VGND sg13g2_decap_8
XFILLER_99_196 VPWR VGND sg13g2_decap_4
X_1439_ Tile_X0Y0_FrameData[22] Tile_X0Y0_FrameData_O[22] VPWR VGND sg13g2_buf_1
X_1508_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG2 Tile_X0Y0_W1BEG[2]
+ VPWR VGND sg13g2_buf_1
XFILLER_11_52 VPWR VGND sg13g2_fill_1
X_0810_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit1.Q _0197_
+ _0198_ VPWR VGND sg13g2_nor2_1
X_0741_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit3.Q UO_OUT_TT_PROJECT1
+ _0152_ UO_OUT_TT_PROJECT5 _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit2.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG9 VPWR VGND sg13g2_mux4_1
X_0672_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit25.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_E2END[1] Tile_X0Y1_E2MID[1] _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit24.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG6 VPWR VGND sg13g2_mux4_1
XFILLER_96_166 VPWR VGND sg13g2_decap_8
X_1224_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1155_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1086_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_0939_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_111 VPWR VGND sg13g2_decap_4
XFILLER_20_188 VPWR VGND sg13g2_decap_8
XFILLER_20_199 VPWR VGND sg13g2_fill_1
XFILLER_87_111 VPWR VGND sg13g2_fill_1
XFILLER_87_199 VPWR VGND sg13g2_fill_1
XFILLER_78_199 VPWR VGND sg13g2_fill_1
XFILLER_0_0 VPWR VGND sg13g2_fill_2
X_0655_ Tile_X0Y0_E6END[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q
+ _0110_ VPWR VGND sg13g2_nor2b_1
X_0586_ VPWR _0055_ _0054_ VGND sg13g2_inv_1
X_0724_ UO_OUT_TT_PROJECT7 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit15.Q _0146_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_33_0 VPWR VGND sg13g2_fill_2
XFILLER_69_199 VPWR VGND sg13g2_fill_1
X_1207_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_1138_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1069_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_54 VPWR VGND sg13g2_decap_8
XFILLER_84_79 VPWR VGND sg13g2_fill_1
XFILLER_83_180 VPWR VGND sg13g2_decap_8
XFILLER_17_62 VPWR VGND sg13g2_fill_2
XFILLER_33_50 VPWR VGND sg13g2_fill_1
X_0440_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit20.Q Tile_X0Y0_E2MID[5]
+ Tile_X0Y0_E2END[5] Tile_X0Y0_E6END[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit21.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG2
+ VPWR VGND sg13g2_mux4_1
X_0371_ VPWR _0301_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit30.Q
+ VGND sg13g2_inv_1
XFILLER_81_139 VPWR VGND sg13g2_fill_2
X_0707_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q
+ _0134_ _0133_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb1 _0341_ sg13g2_a221oi_1
X_0569_ VGND VPWR Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q
+ _0039_ _0040_ _0038_ sg13g2_a21oi_1
X_0638_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit29.Q VPWR
+ _0096_ VGND Tile_X0Y0_EE4END[12] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q
+ sg13g2_o21ai_1
XFILLER_38_17 VPWR VGND sg13g2_fill_1
XFILLER_110_55 VPWR VGND sg13g2_decap_8
XFILLER_63_106 VPWR VGND sg13g2_fill_1
XFILLER_0_198 VPWR VGND sg13g2_fill_2
XFILLER_28_83 VPWR VGND sg13g2_decap_8
X_1610_ Tile_X0Y0_S4END[12] Tile_X0Y1_S4BEG[4] VPWR VGND sg13g2_buf_1
X_1472_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG3 Tile_X0Y0_N1BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1541_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG3 Tile_X0Y0_WW4BEG[3]
+ VPWR VGND sg13g2_buf_1
X_0423_ _0339_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
+ Tile_X0Y0_S2MID[1] VPWR VGND sg13g2_nand2_1
XFILLER_10_2 VPWR VGND sg13g2_fill_1
XFILLER_54_117 VPWR VGND sg13g2_decap_8
XFILLER_105_99 VPWR VGND sg13g2_decap_8
XFILLER_14_96 VPWR VGND sg13g2_fill_1
XFILLER_107_141 VPWR VGND sg13g2_decap_8
XFILLER_100_0 VPWR VGND sg13g2_decap_8
XFILLER_55_70 VPWR VGND sg13g2_fill_2
X_0972_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1524_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb6 Tile_X0Y0_W2BEGb[6]
+ VPWR VGND sg13g2_buf_1
XFILLER_58_2 VPWR VGND sg13g2_fill_1
X_1455_ Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
X_0406_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_mux4_1
X_1386_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_50_142 VPWR VGND sg13g2_decap_8
XFILLER_104_177 VPWR VGND sg13g2_decap_8
XFILLER_104_122 VPWR VGND sg13g2_decap_8
XFILLER_18_106 VPWR VGND sg13g2_decap_4
XFILLER_41_164 VPWR VGND sg13g2_decap_8
XFILLER_110_125 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_fill_1
X_1240_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1171_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_32_120 VPWR VGND sg13g2_decap_4
XANTENNA_16 VPWR VGND Tile_X0Y1_N2MID[5] sg13g2_antennanp
X_0955_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0886_ _0262_ VPWR _0263_ VGND _0255_ _0257_ sg13g2_o21ai_1
XFILLER_99_175 VPWR VGND sg13g2_decap_8
X_1507_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG1 Tile_X0Y0_W1BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_101_158 VPWR VGND sg13g2_decap_8
X_1438_ Tile_X0Y0_FrameData[21] Tile_X0Y0_FrameData_O[21] VPWR VGND sg13g2_buf_1
X_1369_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_102_56 VPWR VGND sg13g2_fill_1
XFILLER_14_197 VPWR VGND sg13g2_fill_2
X_0740_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0318_ Tile_X0Y0_S4END[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q
+ _0152_ VPWR VGND sg13g2_mux4_1
X_0671_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_E2END[2] Tile_X0Y1_E2MID[2] _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG5 VPWR VGND sg13g2_mux4_1
XFILLER_96_145 VPWR VGND sg13g2_decap_8
X_1154_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1223_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1085_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_0938_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_134 VPWR VGND sg13g2_decap_4
X_0869_ _0243_ VPWR UI_IN_TT_PROJECT7 VGND _0244_ _0246_ sg13g2_o21ai_1
XFILLER_11_189 VPWR VGND sg13g2_decap_8
XFILLER_7_138 VPWR VGND sg13g2_decap_8
XFILLER_7_116 VPWR VGND sg13g2_fill_1
XFILLER_93_148 VPWR VGND sg13g2_fill_1
XFILLER_47_82 VPWR VGND sg13g2_decap_8
XFILLER_47_93 VPWR VGND sg13g2_fill_1
X_0723_ _0145_ _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit14.Q
+ VPWR VGND sg13g2_nand2b_1
X_0654_ VGND VPWR UIO_IN_TT_PROJECT6 _0109_ _0108_ sg13g2_or2_1
X_0585_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit8.Q VPWR
+ _0054_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit7.Q
+ _0053_ sg13g2_o21ai_1
XFILLER_6_193 VPWR VGND sg13g2_decap_8
XFILLER_26_0 VPWR VGND sg13g2_fill_2
XFILLER_92_170 VPWR VGND sg13g2_fill_1
X_1137_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_1206_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_29 VPWR VGND sg13g2_fill_2
X_1068_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_88 VPWR VGND sg13g2_decap_8
XFILLER_75_104 VPWR VGND sg13g2_fill_1
XFILLER_90_129 VPWR VGND sg13g2_fill_1
XFILLER_3_141 VPWR VGND sg13g2_decap_8
X_0370_ VPWR _0300_ Tile_X0Y1_E6END[0] VGND sg13g2_inv_1
X_0706_ UO_OUT_TT_PROJECT1 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit3.Q _0134_ VPWR
+ VGND sg13g2_nor3_1
X_0568_ _0011_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ _0039_ VPWR VGND sg13g2_mux2_1
X_0637_ Tile_X0Y0_E6END[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit28.Q
+ _0095_ VPWR VGND sg13g2_nor2b_1
X_0499_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q UIO_OUT_TT_PROJECT7
+ UIO_OE_TT_PROJECT7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb7 VPWR VGND sg13g2_mux4_1
XFILLER_110_34 VPWR VGND sg13g2_decap_8
XFILLER_70_49 VPWR VGND sg13g2_decap_8
XFILLER_79_14 VPWR VGND sg13g2_fill_2
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_0_177 VPWR VGND sg13g2_decap_8
X_1540_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG2 Tile_X0Y0_WW4BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1471_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG2 Tile_X0Y0_N1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0422_ _0338_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG1 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_47_181 VPWR VGND sg13g2_decap_4
XFILLER_108_109 VPWR VGND sg13g2_decap_8
X_1669_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG15 Tile_X0Y1_WW4BEG[15]
+ VPWR VGND sg13g2_buf_1
XFILLER_105_78 VPWR VGND sg13g2_decap_8
XFILLER_53_173 VPWR VGND sg13g2_decap_8
XFILLER_107_120 VPWR VGND sg13g2_decap_8
XFILLER_107_197 VPWR VGND sg13g2_fill_2
XFILLER_107_186 VPWR VGND sg13g2_fill_1
XFILLER_39_50 VPWR VGND sg13g2_decap_8
X_0971_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_44_184 VPWR VGND sg13g2_decap_4
X_1454_ Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
X_1523_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb5 Tile_X0Y0_W2BEGb[5]
+ VPWR VGND sg13g2_buf_1
X_1385_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0405_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit7.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 Tile_X0Y1_E6END[7]
+ _0328_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit6.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3
+ VPWR VGND sg13g2_mux4_1
XFILLER_35_140 VPWR VGND sg13g2_decap_8
XFILLER_104_156 VPWR VGND sg13g2_decap_8
XFILLER_104_101 VPWR VGND sg13g2_decap_8
XFILLER_92_69 VPWR VGND sg13g2_fill_1
XFILLER_25_30 VPWR VGND sg13g2_fill_2
XFILLER_26_184 VPWR VGND sg13g2_decap_8
XFILLER_110_104 VPWR VGND sg13g2_decap_8
XFILLER_2_23 VPWR VGND sg13g2_fill_1
X_1170_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XANTENNA_17 VPWR VGND Tile_X0Y1_FrameStrobe[19] sg13g2_antennanp
X_0954_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_32_198 VPWR VGND sg13g2_fill_2
X_0885_ _0261_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q
+ _0262_ VPWR VGND sg13g2_nor2b_1
XFILLER_101_137 VPWR VGND sg13g2_decap_8
XFILLER_99_154 VPWR VGND sg13g2_decap_8
X_1437_ Tile_X0Y0_FrameData[20] Tile_X0Y0_FrameData_O[20] VPWR VGND sg13g2_buf_1
XFILLER_56_0 VPWR VGND sg13g2_decap_8
X_1506_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W1BEG0 Tile_X0Y0_W1BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1299_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1368_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_198 VPWR VGND sg13g2_fill_2
XFILLER_11_43 VPWR VGND sg13g2_decap_8
XFILLER_14_121 VPWR VGND sg13g2_fill_2
X_0670_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_E2END[3] Tile_X0Y1_E2MID[3] _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG4 VPWR VGND sg13g2_mux4_1
XFILLER_52_83 VPWR VGND sg13g2_fill_1
XFILLER_96_124 VPWR VGND sg13g2_decap_8
X_1153_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1084_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1222_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0937_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0799_ _0188_ _0187_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit29.Q
+ VPWR VGND sg13g2_nand2b_1
X_0868_ _0245_ VPWR _0246_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0151_ sg13g2_o21ai_1
XFILLER_11_146 VPWR VGND sg13g2_decap_4
XFILLER_98_24 VPWR VGND sg13g2_decap_8
XFILLER_0_2 VPWR VGND sg13g2_fill_1
XFILLER_22_97 VPWR VGND sg13g2_decap_8
X_0653_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q _0105_
+ _0106_ _0109_ VPWR VGND sg13g2_nor3_1
X_0722_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q
+ _0144_ _0143_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb6 _0341_ sg13g2_a221oi_1
X_0584_ _0052_ VPWR _0053_ VGND Tile_X0Y0_E6END[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ sg13g2_o21ai_1
XFILLER_33_2 VPWR VGND sg13g2_fill_1
X_1136_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_77_190 VPWR VGND sg13g2_decap_8
X_1205_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_19_0 VPWR VGND sg13g2_fill_2
X_1067_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_67 VPWR VGND sg13g2_decap_8
XFILLER_3_186 VPWR VGND sg13g2_decap_8
X_0636_ VGND VPWR Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q
+ _0092_ UIO_IN_TT_PROJECT3 _0094_ sg13g2_a21oi_1
X_0705_ _0133_ _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
X_0567_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit10.Q VPWR
+ _0038_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit9.Q
+ _0037_ sg13g2_o21ai_1
XFILLER_72_119 VPWR VGND sg13g2_decap_4
X_0498_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit20.Q UIO_OUT_TT_PROJECT6
+ UIO_OE_TT_PROJECT6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit21.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb6 VPWR VGND sg13g2_mux4_1
X_1119_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_196 VPWR VGND sg13g2_decap_4
XFILLER_70_17 VPWR VGND sg13g2_decap_4
XFILLER_79_37 VPWR VGND sg13g2_fill_2
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_0_156 VPWR VGND sg13g2_decap_8
XFILLER_56_193 VPWR VGND sg13g2_decap_8
XFILLER_44_95 VPWR VGND sg13g2_fill_1
X_1470_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG1 Tile_X0Y0_N1BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_5_45 VPWR VGND sg13g2_fill_2
X_0421_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit11.Q _0336_
+ _0337_ VPWR VGND sg13g2_nor2_1
XFILLER_39_127 VPWR VGND sg13g2_fill_2
XFILLER_47_160 VPWR VGND sg13g2_decap_8
XFILLER_47_193 VPWR VGND sg13g2_decap_8
X_0619_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q Tile_X0Y0_EE4END[0]
+ Tile_X0Y0_EE4END[8] _0014_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q _0081_ VPWR
+ VGND sg13g2_mux4_1
X_1668_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG14 Tile_X0Y1_WW4BEG[14]
+ VPWR VGND sg13g2_buf_1
X_1599_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG1 Tile_X0Y1_S2BEGb[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_53_152 VPWR VGND sg13g2_decap_8
XFILLER_53_196 VPWR VGND sg13g2_decap_4
XFILLER_29_160 VPWR VGND sg13g2_fill_2
XFILLER_44_163 VPWR VGND sg13g2_decap_8
XFILLER_44_196 VPWR VGND sg13g2_decap_4
X_0970_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1453_ Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
X_0404_ VPWR VGND _0326_ _0327_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q
+ _0297_ _0328_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a221oi_1
X_1522_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb4 Tile_X0Y0_W2BEGb[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_96_90 VPWR VGND sg13g2_fill_2
X_1384_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_174 VPWR VGND sg13g2_fill_2
XFILLER_50_177 VPWR VGND sg13g2_decap_8
XFILLER_50_188 VPWR VGND sg13g2_fill_1
XFILLER_92_37 VPWR VGND sg13g2_fill_2
XFILLER_41_133 VPWR VGND sg13g2_decap_4
XFILLER_41_199 VPWR VGND sg13g2_fill_1
XFILLER_66_93 VPWR VGND sg13g2_fill_2
XFILLER_17_196 VPWR VGND sg13g2_decap_4
XFILLER_32_177 VPWR VGND sg13g2_decap_8
X_0953_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0884_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q _0259_
+ _0260_ _0261_ VPWR VGND sg13g2_nor3_1
X_1505_ clknet_1_1__leaf_Tile_X0Y1_UserCLK Tile_X0Y0_UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_101_116 VPWR VGND sg13g2_decap_8
XFILLER_99_133 VPWR VGND sg13g2_decap_8
X_1436_ Tile_X0Y0_FrameData[19] Tile_X0Y0_FrameData_O[19] VPWR VGND sg13g2_buf_1
X_1367_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_0 VPWR VGND sg13g2_decap_4
X_1298_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_122 VPWR VGND sg13g2_decap_8
XFILLER_100_182 VPWR VGND sg13g2_decap_8
XFILLER_14_144 VPWR VGND sg13g2_decap_8
XFILLER_14_199 VPWR VGND sg13g2_fill_1
XFILLER_42_7 VPWR VGND sg13g2_decap_8
X_1221_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1152_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_1083_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_0936_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_192 VPWR VGND sg13g2_decap_8
X_0798_ _0154_ _0150_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit28.Q
+ _0187_ VPWR VGND sg13g2_mux2_1
X_0867_ _0245_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_nand2b_1
X_1419_ Tile_X0Y0_FrameData[2] Tile_X0Y0_FrameData_O[2] VPWR VGND sg13g2_buf_1
XFILLER_11_169 VPWR VGND sg13g2_fill_2
XFILLER_98_69 VPWR VGND sg13g2_decap_8
XFILLER_78_103 VPWR VGND sg13g2_decap_8
X_0652_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q _0107_
+ _0108_ VPWR VGND sg13g2_nor2b_1
X_0583_ _0052_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit9.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_nand2b_1
X_0721_ UO_OUT_TT_PROJECT6 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q _0144_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_69_169 VPWR VGND sg13g2_decap_8
X_1204_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1135_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1066_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_0919_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_108_24 VPWR VGND sg13g2_fill_1
XFILLER_83_194 VPWR VGND sg13g2_decap_4
XFILLER_33_20 VPWR VGND sg13g2_decap_4
XFILLER_3_165 VPWR VGND sg13g2_decap_8
XFILLER_74_82 VPWR VGND sg13g2_decap_4
X_0566_ _0036_ VPWR _0037_ VGND Tile_X0Y0_E6END[11] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ sg13g2_o21ai_1
X_0635_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit26.Q _0093_
+ _0094_ VPWR VGND sg13g2_nor2_1
X_0704_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q
+ _0132_ _0131_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb0 _0334_ sg13g2_a221oi_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
XFILLER_65_150 VPWR VGND sg13g2_fill_2
X_0497_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit18.Q UIO_OUT_TT_PROJECT5
+ UIO_OE_TT_PROJECT5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit19.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb5 VPWR VGND sg13g2_mux4_1
XFILLER_110_69 VPWR VGND sg13g2_decap_8
XFILLER_110_14 VPWR VGND sg13g2_decap_4
X_1118_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_175 VPWR VGND sg13g2_decap_8
XFILLER_80_131 VPWR VGND sg13g2_decap_4
X_1049_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_48_128 VPWR VGND sg13g2_fill_1
XFILLER_71_164 VPWR VGND sg13g2_fill_2
XFILLER_28_97 VPWR VGND sg13g2_decap_8
XFILLER_56_150 VPWR VGND sg13g2_fill_2
X_0420_ Tile_X0Y1_N2MID[1] Tile_X0Y1_N2END[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit10.Q
+ _0336_ VPWR VGND sg13g2_mux2_1
XFILLER_62_153 VPWR VGND sg13g2_fill_2
XFILLER_79_0 VPWR VGND sg13g2_decap_8
XFILLER_105_25 VPWR VGND sg13g2_fill_1
X_0618_ _0079_ VPWR _0080_ VGND Tile_X0Y0_E6END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q
+ sg13g2_o21ai_1
X_0549_ _0022_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_nand2b_1
X_1598_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG0 Tile_X0Y1_S2BEGb[0]
+ VPWR VGND sg13g2_buf_1
X_1667_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG13 Tile_X0Y1_WW4BEG[13]
+ VPWR VGND sg13g2_buf_1
XFILLER_53_131 VPWR VGND sg13g2_decap_8
XFILLER_107_199 VPWR VGND sg13g2_fill_1
XFILLER_107_155 VPWR VGND sg13g2_decap_8
XFILLER_71_61 VPWR VGND sg13g2_decap_8
X_1452_ Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
X_1521_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb3 Tile_X0Y0_W2BEGb[3]
+ VPWR VGND sg13g2_buf_1
X_1383_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_0403_ Tile_X0Y1_N1END[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit31.Q _0327_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_50_156 VPWR VGND sg13g2_decap_8
XFILLER_104_136 VPWR VGND sg13g2_decap_8
XFILLER_76_17 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_fill_1
XFILLER_41_178 VPWR VGND sg13g2_decap_8
XFILLER_110_139 VPWR VGND sg13g2_decap_8
XFILLER_103_180 VPWR VGND sg13g2_decap_8
X_0952_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1504_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG3 Tile_X0Y0_N4BEG[15]
+ VPWR VGND sg13g2_buf_1
X_0883_ Tile_X0Y1_E2END[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q _0260_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_99_189 VPWR VGND sg13g2_decap_8
X_1435_ Tile_X0Y0_FrameData[18] Tile_X0Y0_FrameData_O[18] VPWR VGND sg13g2_buf_1
X_1366_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1297_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_156 VPWR VGND sg13g2_decap_8
XFILLER_100_161 VPWR VGND sg13g2_fill_2
XFILLER_14_101 VPWR VGND sg13g2_fill_2
X_1151_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_159 VPWR VGND sg13g2_decap_8
X_1220_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1082_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_0935_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_104 VPWR VGND sg13g2_decap_8
XFILLER_20_115 VPWR VGND sg13g2_fill_2
X_0866_ _0244_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q VPWR VGND
+ sg13g2_nand2b_1
XFILLER_61_0 VPWR VGND sg13g2_decap_4
X_0797_ VGND VPWR _0181_ _0184_ Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_11.A _0186_ sg13g2_a21oi_1
X_1349_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1418_ Tile_X0Y0_FrameData[1] Tile_X0Y0_FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_22_44 VPWR VGND sg13g2_fill_2
XFILLER_8_46 VPWR VGND sg13g2_fill_1
X_0720_ _0143_ _0002_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_nand2b_1
X_0651_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_EE4END[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG14 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit4.Q
+ _0107_ VPWR VGND sg13g2_mux4_1
X_0582_ VGND VPWR _0046_ _0049_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG0
+ _0051_ sg13g2_a21oi_1
XFILLER_92_140 VPWR VGND sg13g2_fill_1
X_1134_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_69_137 VPWR VGND sg13g2_decap_8
X_1203_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1065_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0918_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0849_ _0230_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_nand2b_1
XFILLER_108_47 VPWR VGND sg13g2_decap_8
XFILLER_84_17 VPWR VGND sg13g2_decap_8
XFILLER_17_55 VPWR VGND sg13g2_decap_8
XFILLER_109_0 VPWR VGND sg13g2_decap_4
XFILLER_58_40 VPWR VGND sg13g2_decap_4
XFILLER_74_151 VPWR VGND sg13g2_fill_1
X_0703_ UO_OUT_TT_PROJECT0 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit1.Q _0132_ VPWR
+ VGND sg13g2_nor3_1
X_0565_ _0036_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit11.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_nand2b_1
X_0634_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q Tile_X0Y0_EE4END[3]
+ Tile_X0Y0_EE4END[11] _0011_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q _0093_ VPWR
+ VGND sg13g2_mux4_1
XFILLER_24_0 VPWR VGND sg13g2_fill_1
X_0496_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit16.Q UIO_OUT_TT_PROJECT4
+ UIO_OE_TT_PROJECT4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit17.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb4 VPWR VGND sg13g2_mux4_1
X_1117_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_110_48 VPWR VGND sg13g2_decap_8
X_1048_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_79_39 VPWR VGND sg13g2_fill_1
XFILLER_0_147 VPWR VGND sg13g2_decap_4
XFILLER_56_140 VPWR VGND sg13g2_fill_2
XFILLER_28_76 VPWR VGND sg13g2_decap_8
XFILLER_56_184 VPWR VGND sg13g2_fill_1
Xclkbuf_1_0__f_Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK clknet_1_0__leaf_Tile_X0Y1_UserCLK
+ VPWR VGND sg13g2_buf_8
XFILLER_62_198 VPWR VGND sg13g2_fill_2
X_1666_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG12 Tile_X0Y1_WW4BEG[12]
+ VPWR VGND sg13g2_buf_1
X_0617_ VGND VPWR _0291_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit16.Q
+ _0079_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q sg13g2_a21oi_1
X_0548_ _0019_ _0021_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG0
+ VPWR VGND sg13g2_nor2_1
X_1597_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG7 Tile_X0Y1_S2BEG[7]
+ VPWR VGND sg13g2_buf_1
X_0479_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 Tile_X0Y1_E6END[4]
+ _0010_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0
+ VPWR VGND sg13g2_mux4_1
XFILLER_81_29 VPWR VGND sg13g2_fill_2
XFILLER_107_178 VPWR VGND sg13g2_fill_1
XFILLER_107_134 VPWR VGND sg13g2_decap_8
XFILLER_29_184 VPWR VGND sg13g2_fill_2
XFILLER_55_96 VPWR VGND sg13g2_decap_8
X_1520_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb2 Tile_X0Y0_W2BEGb[2]
+ VPWR VGND sg13g2_buf_1
X_1451_ Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
X_1382_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_0402_ _0326_ _0325_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_35_198 VPWR VGND sg13g2_fill_2
XFILLER_104_115 VPWR VGND sg13g2_decap_8
X_1649_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG7 Tile_X0Y1_W6BEG[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_25_11 VPWR VGND sg13g2_fill_2
XFILLER_26_132 VPWR VGND sg13g2_decap_4
XFILLER_26_154 VPWR VGND sg13g2_fill_1
XFILLER_26_198 VPWR VGND sg13g2_fill_2
XFILLER_110_118 VPWR VGND sg13g2_decap_8
XFILLER_32_113 VPWR VGND sg13g2_decap_8
X_0951_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_0882_ _0259_ _0258_ _0305_ _0306_ Tile_X0Y1_E2END[5] VPWR VGND sg13g2_a22oi_1
X_1503_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG2 Tile_X0Y0_N4BEG[14]
+ VPWR VGND sg13g2_buf_1
XFILLER_99_168 VPWR VGND sg13g2_decap_8
X_1434_ Tile_X0Y0_FrameData[17] Tile_X0Y0_FrameData_O[17] VPWR VGND sg13g2_buf_1
X_1296_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1365_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_98_190 VPWR VGND sg13g2_decap_8
XFILLER_100_140 VPWR VGND sg13g2_decap_8
X_1150_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_96_138 VPWR VGND sg13g2_decap_8
XFILLER_77_83 VPWR VGND sg13g2_fill_2
X_1081_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_0934_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0865_ _0243_ _0242_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit31.Q
+ VPWR VGND sg13g2_nand2b_1
X_0796_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q _0185_
+ _0186_ VPWR VGND sg13g2_nor2_1
X_1417_ Tile_X0Y0_FrameData[0] Tile_X0Y0_FrameData_O[0] VPWR VGND sg13g2_buf_1
XFILLER_54_0 VPWR VGND sg13g2_decap_8
XFILLER_95_193 VPWR VGND sg13g2_decap_8
X_1279_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1348_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_0650_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit3.Q VPWR
+ _0106_ VGND Tile_X0Y0_EE4END[14] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit2.Q
+ sg13g2_o21ai_1
X_0581_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit5.Q _0050_
+ _0051_ VPWR VGND sg13g2_nor2_1
XFILLER_6_186 VPWR VGND sg13g2_decap_8
X_1133_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1202_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1064_ Tile_X0Y0_FrameData[7] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
X_0917_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_0779_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_E6END[9] Tile_X0Y1_EE4END[1] _0157_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ _0171_ VPWR VGND sg13g2_mux4_1
X_0848_ _0229_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q VPWR VGND
+ sg13g2_nand2b_1
XFILLER_59_182 VPWR VGND sg13g2_fill_1
XFILLER_99_92 VPWR VGND sg13g2_fill_2
X_0633_ _0091_ VPWR _0092_ VGND Tile_X0Y0_E6END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q
+ sg13g2_o21ai_1
X_0702_ _0131_ _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit0.Q
+ VPWR VGND sg13g2_nand2b_1
X_0564_ _0033_ _0035_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG2
+ VPWR VGND sg13g2_nor2_1
X_0495_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit14.Q UIO_OUT_TT_PROJECT3
+ UIO_OE_TT_PROJECT3 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit15.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb3 VPWR VGND sg13g2_mux4_1
X_1116_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1047_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_17_0 VPWR VGND sg13g2_fill_1
XFILLER_110_27 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_71_166 VPWR VGND sg13g2_fill_1
XFILLER_60_31 VPWR VGND sg13g2_fill_2
XFILLER_109_91 VPWR VGND sg13g2_fill_1
XFILLER_62_155 VPWR VGND sg13g2_fill_1
XFILLER_62_111 VPWR VGND sg13g2_decap_8
XFILLER_47_174 VPWR VGND sg13g2_decap_8
X_1596_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG6 Tile_X0Y1_S2BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1665_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG11 Tile_X0Y1_WW4BEG[11]
+ VPWR VGND sg13g2_buf_1
X_0616_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0325_ Tile_X0Y0_S4END[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit7.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 VPWR VGND sg13g2_mux4_1
X_0547_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q _0020_
+ _0021_ VPWR VGND sg13g2_nor2_1
X_0478_ VPWR VGND _0008_ _0009_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q
+ _0300_ _0010_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_a221oi_1
XFILLER_53_166 VPWR VGND sg13g2_decap_8
XFILLER_107_113 VPWR VGND sg13g2_decap_8
XFILLER_29_130 VPWR VGND sg13g2_fill_2
XFILLER_44_177 VPWR VGND sg13g2_decap_8
XFILLER_44_188 VPWR VGND sg13g2_fill_1
X_1450_ Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
X_0401_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit18.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_E6END[11] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15
+ _0324_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit19.Q _0325_
+ VPWR VGND sg13g2_mux4_1
X_1381_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_35_122 VPWR VGND sg13g2_fill_1
XFILLER_50_136 VPWR VGND sg13g2_fill_2
X_1648_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG6 Tile_X0Y1_W6BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1579_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameData_O[25] VPWR VGND sg13g2_buf_1
XFILLER_26_111 VPWR VGND sg13g2_decap_4
XFILLER_41_11 VPWR VGND sg13g2_fill_2
XFILLER_103_160 VPWR VGND sg13g2_fill_2
XFILLER_66_63 VPWR VGND sg13g2_fill_2
XFILLER_66_41 VPWR VGND sg13g2_fill_1
XFILLER_2_49 VPWR VGND sg13g2_decap_4
XFILLER_2_16 VPWR VGND sg13g2_decap_8
X_0950_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_0881_ _0258_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit2.Q
+ Tile_X0Y0_S2MID[2] VPWR VGND sg13g2_nand2b_1
X_1502_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG1 Tile_X0Y0_N4BEG[13]
+ VPWR VGND sg13g2_buf_1
XFILLER_99_147 VPWR VGND sg13g2_decap_8
X_1433_ Tile_X0Y0_FrameData[16] Tile_X0Y0_FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_102_17 VPWR VGND sg13g2_decap_4
X_1295_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
X_1364_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_100_196 VPWR VGND sg13g2_decap_4
XFILLER_100_163 VPWR VGND sg13g2_fill_1
XFILLER_14_103 VPWR VGND sg13g2_fill_1
XFILLER_36_88 VPWR VGND sg13g2_fill_2
XFILLER_96_117 VPWR VGND sg13g2_decap_8
XFILLER_89_191 VPWR VGND sg13g2_decap_8
X_1080_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_0933_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0864_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit30.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_EE4END[15] Tile_X0Y1_EE4END[7] Tile_X0Y1_E6END[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit29.Q
+ _0242_ VPWR VGND sg13g2_mux4_1
X_0795_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_E6END[11] Tile_X0Y1_EE4END[3] _0155_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ _0185_ VPWR VGND sg13g2_mux4_1
X_1347_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1416_ clknet_1_0__leaf_Tile_X0Y1_UserCLK CLK_TT_PROJECT VPWR VGND sg13g2_buf_1
XFILLER_95_172 VPWR VGND sg13g2_decap_8
X_1278_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_98_17 VPWR VGND sg13g2_decap_8
XFILLER_93_109 VPWR VGND sg13g2_decap_4
XFILLER_47_43 VPWR VGND sg13g2_decap_4
XFILLER_63_75 VPWR VGND sg13g2_fill_2
XFILLER_6_143 VPWR VGND sg13g2_fill_1
X_0580_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_EE4END[12] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit6.Q
+ _0050_ VPWR VGND sg13g2_mux4_1
X_1201_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1132_ Tile_X0Y0_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1063_ Tile_X0Y0_FrameData[8] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_0916_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_0778_ _0169_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit29.Q
+ _0170_ VPWR VGND sg13g2_nor2b_1
X_0847_ _0228_ _0227_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit22.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_3_179 VPWR VGND sg13g2_decap_8
XFILLER_88_7 VPWR VGND sg13g2_decap_4
X_0563_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit7.Q _0034_
+ _0035_ VPWR VGND sg13g2_nor2_1
X_0632_ VGND VPWR _0294_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit25.Q
+ _0091_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit27.Q sg13g2_a21oi_1
X_0701_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q
+ _0130_ _0129_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG7 _0334_ sg13g2_a221oi_1
X_0494_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit12.Q UIO_OUT_TT_PROJECT2
+ UIO_OE_TT_PROJECT2 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit13.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb2 VPWR VGND sg13g2_mux4_1
X_1115_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_189 VPWR VGND sg13g2_decap_8
XFILLER_80_112 VPWR VGND sg13g2_fill_2
X_1046_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_80 VPWR VGND sg13g2_fill_2
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_28_67 VPWR VGND sg13g2_decap_4
XFILLER_56_131 VPWR VGND sg13g2_fill_1
XFILLER_69_41 VPWR VGND sg13g2_decap_8
XFILLER_39_109 VPWR VGND sg13g2_fill_2
XFILLER_47_153 VPWR VGND sg13g2_decap_8
X_0546_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_EE4END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG8 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ _0020_ VPWR VGND sg13g2_mux4_1
X_1664_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG10 Tile_X0Y1_WW4BEG[10]
+ VPWR VGND sg13g2_buf_1
X_1595_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG5 Tile_X0Y1_S2BEG[5]
+ VPWR VGND sg13g2_buf_1
X_0615_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q Tile_X0Y1_N1END[2]
+ Tile_X0Y1_N4END[2] _0318_ Tile_X0Y0_S4END[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14 VPWR VGND sg13g2_mux4_1
XFILLER_38_164 VPWR VGND sg13g2_decap_4
X_0477_ Tile_X0Y1_N1END[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit25.Q _0009_ VPWR
+ VGND sg13g2_nor3_1
X_1029_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_14_69 VPWR VGND sg13g2_decap_4
XFILLER_53_145 VPWR VGND sg13g2_decap_8
XFILLER_107_169 VPWR VGND sg13g2_decap_4
XFILLER_29_186 VPWR VGND sg13g2_fill_1
XFILLER_29_197 VPWR VGND sg13g2_fill_2
XFILLER_44_156 VPWR VGND sg13g2_decap_8
XFILLER_71_42 VPWR VGND sg13g2_fill_2
XFILLER_71_31 VPWR VGND sg13g2_decap_8
X_0400_ VPWR VGND _0322_ _0323_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q
+ _0289_ _0324_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a221oi_1
X_1380_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_50_104 VPWR VGND sg13g2_fill_2
XFILLER_77_0 VPWR VGND sg13g2_decap_8
X_0529_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit24.Q Tile_X0Y1_N4END[4]
+ Tile_X0Y0_S4END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG15 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit25.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG0 VPWR VGND sg13g2_mux4_1
X_1647_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG5 Tile_X0Y1_W6BEG[5]
+ VPWR VGND sg13g2_buf_1
X_1578_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameData_O[24] VPWR VGND sg13g2_buf_1
XFILLER_41_126 VPWR VGND sg13g2_decap_4
XFILLER_106_82 VPWR VGND sg13g2_decap_8
XFILLER_103_194 VPWR VGND sg13g2_decap_4
XFILLER_66_86 VPWR VGND sg13g2_decap_8
XFILLER_17_189 VPWR VGND sg13g2_decap_8
XFILLER_32_159 VPWR VGND sg13g2_fill_1
X_0880_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit0.Q VPWR
+ _0257_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit1.Q
+ _0256_ sg13g2_o21ai_1
X_1501_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N4BEG0 Tile_X0Y0_N4BEG[12]
+ VPWR VGND sg13g2_buf_1
XFILLER_101_109 VPWR VGND sg13g2_decap_8
XFILLER_99_126 VPWR VGND sg13g2_decap_8
X_1432_ Tile_X0Y0_FrameData[15] Tile_X0Y0_FrameData_O[15] VPWR VGND sg13g2_buf_1
X_1363_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
X_1294_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_31_192 VPWR VGND sg13g2_decap_8
XFILLER_11_26 VPWR VGND sg13g2_decap_4
XFILLER_11_15 VPWR VGND sg13g2_fill_1
XFILLER_100_175 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_fill_1
XFILLER_77_85 VPWR VGND sg13g2_fill_1
X_0932_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_141 VPWR VGND sg13g2_fill_2
XFILLER_9_185 VPWR VGND sg13g2_decap_8
X_0863_ _0241_ VPWR UI_IN_TT_PROJECT6 VGND _0237_ _0239_ sg13g2_o21ai_1
X_0794_ _0183_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit3.Q
+ _0184_ VPWR VGND sg13g2_nor2b_1
X_1415_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1346_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1277_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_86_173 VPWR VGND sg13g2_decap_4
XFILLER_86_140 VPWR VGND sg13g2_decap_8
XFILLER_63_21 VPWR VGND sg13g2_fill_2
X_1200_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[1] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_92_198 VPWR VGND sg13g2_fill_2
X_1131_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1062_ Tile_X0Y0_FrameData[9] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_0915_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
X_0777_ VGND VPWR Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ _0341_ _0169_ _0168_ sg13g2_a21oi_1
X_0846_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit21.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_EE4END[12] Tile_X0Y1_EE4END[4] Tile_X0Y1_E6END[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit20.Q
+ _0227_ VPWR VGND sg13g2_mux4_1
X_1329_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_83_198 VPWR VGND sg13g2_fill_2
XFILLER_83_187 VPWR VGND sg13g2_decap_8
XFILLER_33_46 VPWR VGND sg13g2_decap_4
XFILLER_59_195 VPWR VGND sg13g2_decap_4
X_0700_ UO_OUT_TT_PROJECT7 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit30.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit31.Q _0130_ VPWR
+ VGND sg13g2_nor3_1
XFILLER_99_94 VPWR VGND sg13g2_fill_1
X_0562_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q Tile_X0Y0_E1END[2]
+ Tile_X0Y0_EE4END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG6
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ _0034_ VPWR VGND sg13g2_mux4_1
X_0631_ VGND VPWR Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q
+ _0088_ UIO_IN_TT_PROJECT2 _0090_ sg13g2_a21oi_1
X_1114_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_180 VPWR VGND sg13g2_decap_8
X_0493_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q UIO_OUT_TT_PROJECT1
+ UIO_OE_TT_PROJECT1 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb1 VPWR VGND sg13g2_mux4_1
XFILLER_110_18 VPWR VGND sg13g2_fill_1
XFILLER_80_168 VPWR VGND sg13g2_decap_8
XFILLER_80_135 VPWR VGND sg13g2_fill_2
X_1045_ Tile_X0Y0_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_198 VPWR VGND sg13g2_fill_2
XFILLER_0_61 VPWR VGND sg13g2_fill_2
XFILLER_0_72 VPWR VGND sg13g2_decap_8
X_0829_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q _0211_
+ _0212_ _0214_ VPWR VGND sg13g2_nor3_1
XFILLER_60_33 VPWR VGND sg13g2_fill_1
XFILLER_62_146 VPWR VGND sg13g2_decap_8
X_1663_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG9 Tile_X0Y1_WW4BEG[9]
+ VPWR VGND sg13g2_buf_1
X_0545_ VGND VPWR Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q
+ _0018_ _0019_ _0017_ sg13g2_a21oi_1
X_0614_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y1_N1END[1]
+ Tile_X0Y1_N4END[1] _0311_ Tile_X0Y0_S4END[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_mux4_1
X_1594_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG4 Tile_X0Y1_S2BEG[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_22_0 VPWR VGND sg13g2_fill_1
X_0476_ _0008_ _0007_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_53_124 VPWR VGND sg13g2_decap_8
X_1028_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_148 VPWR VGND sg13g2_decap_8
XFILLER_100_7 VPWR VGND sg13g2_fill_2
XFILLER_29_132 VPWR VGND sg13g2_fill_1
XFILLER_55_66 VPWR VGND sg13g2_decap_4
XFILLER_50_149 VPWR VGND sg13g2_decap_8
X_1646_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG4 Tile_X0Y1_W6BEG[4]
+ VPWR VGND sg13g2_buf_1
XFILLER_104_129 VPWR VGND sg13g2_decap_8
X_0528_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit22.Q UIO_OUT_TT_PROJECT3
+ UIO_OE_TT_PROJECT7 _0014_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit23.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG15
+ VPWR VGND sg13g2_mux4_1
X_0459_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit18.Q Tile_X0Y1_E2MID[2]
+ Tile_X0Y1_E2END[2] Tile_X0Y1_E6END[2] _0001_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit19.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb5 VPWR VGND sg13g2_mux4_1
X_1577_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameData_O[23] VPWR VGND sg13g2_buf_1
XFILLER_41_68 VPWR VGND sg13g2_fill_2
XFILLER_103_173 VPWR VGND sg13g2_decap_8
XFILLER_66_21 VPWR VGND sg13g2_fill_1
X_1500_ Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_11.A Tile_X0Y0_N4BEG[11] VPWR VGND sg13g2_buf_1
X_1431_ Tile_X0Y0_FrameData[14] Tile_X0Y0_FrameData_O[14] VPWR VGND sg13g2_buf_1
X_1293_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1362_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
X_1629_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG3 Tile_X0Y1_W2BEG[3]
+ VPWR VGND sg13g2_buf_1
XFILLER_100_154 VPWR VGND sg13g2_decap_8
XFILLER_36_68 VPWR VGND sg13g2_fill_2
XFILLER_52_45 VPWR VGND sg13g2_decap_4
XFILLER_93_41 VPWR VGND sg13g2_fill_2
X_0931_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_193 VPWR VGND sg13g2_decap_8
X_0862_ _0241_ _0240_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_61_4 VPWR VGND sg13g2_fill_2
X_0793_ VGND VPWR Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ _0355_ _0183_ _0182_ sg13g2_a21oi_1
XFILLER_3_50 VPWR VGND sg13g2_decap_4
X_1276_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1414_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1345_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_86_196 VPWR VGND sg13g2_decap_4
XFILLER_47_89 VPWR VGND sg13g2_decap_4
XFILLER_63_99 VPWR VGND sg13g2_decap_8
XFILLER_63_77 VPWR VGND sg13g2_fill_1
XFILLER_10_152 VPWR VGND sg13g2_decap_8
XFILLER_6_101 VPWR VGND sg13g2_decap_4
XFILLER_10_196 VPWR VGND sg13g2_decap_4
X_1130_ Tile_X0Y0_FrameData[5] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
X_1061_ Tile_X0Y0_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_0914_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0845_ _0225_ _0226_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit19.Q
+ UI_IN_TT_PROJECT3 VPWR VGND sg13g2_mux2_1
XFILLER_108_29 VPWR VGND sg13g2_fill_1
X_0776_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q VPWR
+ _0168_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 sg13g2_o21ai_1
XFILLER_83_166 VPWR VGND sg13g2_fill_1
XFILLER_68_163 VPWR VGND sg13g2_decap_4
X_1328_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1259_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_17_48 VPWR VGND sg13g2_decap_8
XFILLER_109_4 VPWR VGND sg13g2_fill_1
XFILLER_58_11 VPWR VGND sg13g2_fill_1
XFILLER_58_33 VPWR VGND sg13g2_decap_8
XFILLER_58_44 VPWR VGND sg13g2_fill_1
XFILLER_58_66 VPWR VGND sg13g2_decap_4
XFILLER_74_199 VPWR VGND sg13g2_fill_1
X_0561_ VGND VPWR Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit6.Q
+ _0032_ _0033_ _0031_ sg13g2_a21oi_1
X_0630_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit23.Q _0089_
+ _0090_ VPWR VGND sg13g2_nor2_1
X_0492_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit8.Q UIO_OUT_TT_PROJECT0
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit9.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEGb0 VPWR VGND sg13g2_mux4_1
X_1113_ Tile_X0Y0_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
X_1044_ Tile_X0Y0_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_65_100 VPWR VGND sg13g2_decap_8
XFILLER_0_40 VPWR VGND sg13g2_fill_1
XFILLER_9_82 VPWR VGND sg13g2_fill_1
X_0759_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit27.Q UO_OUT_TT_PROJECT5
+ _0148_ _0152_ _0342_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit26.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG5 VPWR VGND sg13g2_mux4_1
X_0828_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q Tile_X0Y1_EE4END[0]
+ Tile_X0Y1_EE4END[8] Tile_X0Y1_E6END[0] Tile_X0Y1_E6END[8] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit9.Q
+ _0213_ VPWR VGND sg13g2_mux4_1
XFILLER_44_35 VPWR VGND sg13g2_decap_4
XFILLER_56_177 VPWR VGND sg13g2_decap_8
XFILLER_109_83 VPWR VGND sg13g2_decap_4
XFILLER_85_31 VPWR VGND sg13g2_fill_1
XFILLER_62_125 VPWR VGND sg13g2_decap_4
X_1662_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG8 Tile_X0Y1_WW4BEG[8]
+ VPWR VGND sg13g2_buf_1
X_0613_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit0.Q Tile_X0Y1_N1END[0]
+ Tile_X0Y1_N4END[0] _0007_ Tile_X0Y0_S4END[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit1.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_mux4_1
X_0544_ _0014_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ _0018_ VPWR VGND sg13g2_mux2_1
X_0475_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit13.Q Tile_X0Y0_E1END[0]
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 Tile_X0Y0_E6END[8]
+ _0006_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit12.Q _0007_
+ VPWR VGND sg13g2_mux4_1
X_1593_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG3 Tile_X0Y1_S2BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1027_ Tile_X0Y0_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_107_127 VPWR VGND sg13g2_decap_8
XFILLER_39_57 VPWR VGND sg13g2_decap_4
XFILLER_29_199 VPWR VGND sg13g2_fill_1
XFILLER_55_89 VPWR VGND sg13g2_decap_8
XFILLER_106_182 VPWR VGND sg13g2_decap_8
XFILLER_29_90 VPWR VGND sg13g2_fill_2
XFILLER_35_147 VPWR VGND sg13g2_fill_2
XFILLER_50_106 VPWR VGND sg13g2_fill_1
XFILLER_104_108 VPWR VGND sg13g2_decap_8
X_1645_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG3 Tile_X0Y1_W6BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1576_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameData_O[22] VPWR VGND sg13g2_buf_1
X_0389_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit29.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2 _0316_ VPWR VGND sg13g2_nor3_1
X_0527_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit8.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0
+ Tile_X0Y1_N4END[4] Tile_X0Y0_S1END[0] Tile_X0Y0_S4END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit9.Q
+ _0014_ VPWR VGND sg13g2_mux4_1
X_0458_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit18.Q Tile_X0Y1_N2MID[5]
+ Tile_X0Y1_N2END[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG5
+ Tile_X0Y0_S2MID[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit19.Q
+ _0001_ VPWR VGND sg13g2_mux4_1
XFILLER_26_136 VPWR VGND sg13g2_fill_1
XFILLER_82_87 VPWR VGND sg13g2_fill_2
XFILLER_82_43 VPWR VGND sg13g2_decap_4
XFILLER_25_191 VPWR VGND sg13g2_decap_8
XFILLER_32_106 VPWR VGND sg13g2_decap_8
X_1430_ Tile_X0Y0_FrameData[13] Tile_X0Y0_FrameData_O[13] VPWR VGND sg13g2_buf_1
XFILLER_56_7 VPWR VGND sg13g2_decap_4
X_1292_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1361_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_16_191 VPWR VGND sg13g2_decap_8
XFILLER_82_0 VPWR VGND sg13g2_decap_8
XFILLER_98_183 VPWR VGND sg13g2_decap_8
X_1628_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG2 Tile_X0Y1_W2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1559_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameData_O[5] VPWR VGND sg13g2_buf_1
XFILLER_100_133 VPWR VGND sg13g2_decap_8
XFILLER_52_24 VPWR VGND sg13g2_decap_4
X_0930_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_161 VPWR VGND sg13g2_decap_8
X_0861_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit27.Q Tile_X0Y1_E1END[2]
+ Tile_X0Y1_EE4END[14] Tile_X0Y1_EE4END[6] Tile_X0Y1_E6END[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
+ _0240_ VPWR VGND sg13g2_mux4_1
X_0792_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q VPWR
+ _0182_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15 sg13g2_o21ai_1
X_1413_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_186 VPWR VGND sg13g2_decap_8
XFILLER_95_153 VPWR VGND sg13g2_fill_1
X_1275_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1344_ Tile_X0Y1_FrameData[7] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_103_74 VPWR VGND sg13g2_decap_4
XFILLER_10_120 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_fill_1
XFILLER_77_197 VPWR VGND sg13g2_fill_2
X_1060_ Tile_X0Y0_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_0913_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0775_ _0167_ _0166_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_0844_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q _0223_
+ _0224_ _0226_ VPWR VGND sg13g2_nor3_1
XFILLER_45_0 VPWR VGND sg13g2_fill_2
XFILLER_68_197 VPWR VGND sg13g2_fill_2
XFILLER_68_186 VPWR VGND sg13g2_fill_2
X_1189_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
X_1258_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_1327_ Tile_X0Y1_FrameData[24] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_74_156 VPWR VGND sg13g2_fill_1
XFILLER_99_30 VPWR VGND sg13g2_decap_8
XFILLER_23_70 VPWR VGND sg13g2_decap_8
X_0560_ _0012_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit8.Q
+ _0032_ VPWR VGND sg13g2_mux2_1
X_0491_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit6.Q UIO_OUT_TT_PROJECT7
+ UIO_OE_TT_PROJECT7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG0
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit7.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG7 VPWR VGND sg13g2_mux4_1
X_1112_ Tile_X0Y0_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1043_ Tile_X0Y0_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_63 VPWR VGND sg13g2_fill_1
X_0758_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit25.Q UO_OUT_TT_PROJECT4
+ _0147_ _0151_ _0335_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit24.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG4 VPWR VGND sg13g2_mux4_1
X_0827_ _0150_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q
+ _0212_ VPWR VGND sg13g2_nor2b_1
X_0689_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q
+ _0122_ _0121_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG3 _0355_ sg13g2_a221oi_1
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_71_104 VPWR VGND sg13g2_fill_1
XFILLER_60_68 VPWR VGND sg13g2_decap_4
XFILLER_60_24 VPWR VGND sg13g2_decap_8
XFILLER_47_167 VPWR VGND sg13g2_decap_8
XFILLER_70_170 VPWR VGND sg13g2_fill_2
XFILLER_34_91 VPWR VGND sg13g2_fill_1
X_0612_ VGND VPWR _0073_ _0076_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S4BEG3
+ _0078_ sg13g2_a21oi_1
X_1661_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG7 Tile_X0Y1_WW4BEG[7]
+ VPWR VGND sg13g2_buf_1
X_1592_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG2 Tile_X0Y1_S2BEG[2]
+ VPWR VGND sg13g2_buf_1
X_0543_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit1.Q VPWR
+ _0017_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit0.Q
+ _0016_ sg13g2_o21ai_1
X_0474_ VPWR VGND _0004_ _0005_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q
+ _0290_ _0006_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q
+ sg13g2_a221oi_1
X_1026_ Tile_X0Y0_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_53_159 VPWR VGND sg13g2_decap_8
XFILLER_107_106 VPWR VGND sg13g2_decap_8
XFILLER_106_161 VPWR VGND sg13g2_decap_8
XFILLER_20_82 VPWR VGND sg13g2_fill_1
XFILLER_50_129 VPWR VGND sg13g2_decap_8
XFILLER_43_192 VPWR VGND sg13g2_decap_8
X_0526_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit20.Q UIO_OUT_TT_PROJECT2
+ UIO_OE_TT_PROJECT6 _0013_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit21.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG14
+ VPWR VGND sg13g2_mux4_1
X_1644_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG2 Tile_X0Y1_W6BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1575_ Tile_X0Y1_FrameData[21] Tile_X0Y1_FrameData_O[21] VPWR VGND sg13g2_buf_1
X_0388_ _0315_ Tile_X0Y0_S1END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit28.Q
+ VPWR VGND sg13g2_nand2b_1
X_0457_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit30.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_E2MID[2] Tile_X0Y0_E2END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG5
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit31.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG5
+ VPWR VGND sg13g2_mux4_1
XFILLER_26_104 VPWR VGND sg13g2_decap_8
X_1009_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_96 VPWR VGND sg13g2_decap_8
XFILLER_103_153 VPWR VGND sg13g2_decap_8
X_1360_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[6] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
X_1291_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_16_170 VPWR VGND sg13g2_decap_8
XFILLER_23_129 VPWR VGND sg13g2_fill_2
XFILLER_75_0 VPWR VGND sg13g2_decap_8
XFILLER_31_173 VPWR VGND sg13g2_fill_2
XFILLER_100_112 VPWR VGND sg13g2_decap_8
XFILLER_98_162 VPWR VGND sg13g2_decap_8
X_0509_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit26.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit27.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG9 VPWR VGND sg13g2_mux4_1
X_1627_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG1 Tile_X0Y1_W2BEG[1]
+ VPWR VGND sg13g2_buf_1
X_1489_ Tile_X0Y1_N4END[8] Tile_X0Y0_N4BEG[0] VPWR VGND sg13g2_buf_1
X_1558_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_100_189 VPWR VGND sg13g2_decap_8
XFILLER_22_195 VPWR VGND sg13g2_decap_4
XFILLER_77_11 VPWR VGND sg13g2_fill_2
XFILLER_93_43 VPWR VGND sg13g2_fill_1
XFILLER_9_100 VPWR VGND sg13g2_fill_2
XFILLER_9_199 VPWR VGND sg13g2_fill_1
X_0860_ _0238_ VPWR _0239_ VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit26.Q
+ _0152_ sg13g2_o21ai_1
X_0791_ _0181_ _0180_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit2.Q
+ VPWR VGND sg13g2_nand2b_1
XFILLER_95_132 VPWR VGND sg13g2_decap_8
X_1343_ Tile_X0Y1_FrameData[8] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit8.Q
+ VPWR VGND sg13g2_dlhq_1
X_1412_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_165 VPWR VGND sg13g2_decap_8
X_1274_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_0989_ Tile_X0Y0_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_47_47 VPWR VGND sg13g2_fill_1
XFILLER_103_97 VPWR VGND sg13g2_decap_8
XFILLER_63_57 VPWR VGND sg13g2_fill_1
XFILLER_5_0 VPWR VGND sg13g2_fill_2
XFILLER_92_168 VPWR VGND sg13g2_fill_2
X_0912_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_5_180 VPWR VGND sg13g2_decap_8
X_0774_ _0153_ _0149_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit27.Q
+ _0166_ VPWR VGND sg13g2_mux2_1
X_0843_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q Tile_X0Y1_EE4END[3]
+ Tile_X0Y1_EE4END[11] Tile_X0Y1_E6END[3] Tile_X0Y1_E6END[11] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q
+ _0225_ VPWR VGND sg13g2_mux4_1
X_1326_ Tile_X0Y1_FrameData[25] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
X_1188_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit3.Q
+ VPWR VGND sg13g2_dlhq_1
X_1257_ Tile_X0Y1_FrameData[30] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_121 VPWR VGND sg13g2_fill_1
XFILLER_59_110 VPWR VGND sg13g2_decap_8
XFILLER_90_66 VPWR VGND sg13g2_decap_8
XFILLER_2_194 VPWR VGND sg13g2_decap_4
X_0490_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit4.Q UIO_OUT_TT_PROJECT6
+ UIO_OE_TT_PROJECT6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG1
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG6 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit5.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W2BEG6 VPWR VGND sg13g2_mux4_1
X_1111_ Tile_X0Y0_FrameData[24] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit24.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_105 VPWR VGND sg13g2_decap_8
X_1042_ Tile_X0Y0_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
X_0688_ UO_OUT_TT_PROJECT3 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit23.Q _0122_ VPWR
+ VGND sg13g2_nor3_1
X_0826_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit8.Q _0158_
+ _0211_ VPWR VGND sg13g2_nor2_1
X_0757_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit22.Q Tile_X0Y1_N4END[3]
+ Tile_X0Y0_S4END[7] _0150_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG12
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit23.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG3
+ VPWR VGND sg13g2_mux4_1
X_1309_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_146 VPWR VGND sg13g2_decap_4
XFILLER_109_74 VPWR VGND sg13g2_fill_1
XFILLER_47_146 VPWR VGND sg13g2_decap_8
XFILLER_79_7 VPWR VGND sg13g2_decap_8
X_0611_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit14.Q _0077_
+ _0078_ VPWR VGND sg13g2_nor2_1
X_0542_ _0015_ VPWR _0016_ VGND Tile_X0Y0_E6END[8] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ sg13g2_o21ai_1
X_1660_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG6 Tile_X0Y1_WW4BEG[6]
+ VPWR VGND sg13g2_buf_1
X_1591_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG1 Tile_X0Y1_S2BEG[1]
+ VPWR VGND sg13g2_buf_1
X_0473_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit25.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END0 _0005_ VPWR VGND sg13g2_nor3_1
XFILLER_38_124 VPWR VGND sg13g2_fill_1
XFILLER_38_157 VPWR VGND sg13g2_decap_8
XFILLER_38_168 VPWR VGND sg13g2_fill_1
X_1025_ Tile_X0Y0_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_53_116 VPWR VGND sg13g2_decap_4
XFILLER_53_138 VPWR VGND sg13g2_decap_8
X_0809_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_EE4END[13] Tile_X0Y1_E6END[5] _0157_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
+ _0197_ VPWR VGND sg13g2_mux4_1
XFILLER_30_17 VPWR VGND sg13g2_fill_2
XFILLER_71_68 VPWR VGND sg13g2_fill_2
XFILLER_105_0 VPWR VGND sg13g2_decap_4
XFILLER_35_149 VPWR VGND sg13g2_fill_1
XFILLER_43_171 VPWR VGND sg13g2_decap_8
X_1643_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG1 Tile_X0Y1_W6BEG[1]
+ VPWR VGND sg13g2_buf_1
XANTENNA_1 VPWR VGND Tile_X0Y0_S2END[4] sg13g2_antennanp
X_0456_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit24.Q Tile_X0Y0_E2MID[3]
+ Tile_X0Y0_E2END[3] Tile_X0Y0_E6END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit25.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG4
+ VPWR VGND sg13g2_mux4_1
X_0525_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit10.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit11.Q
+ _0013_ VPWR VGND sg13g2_mux4_1
X_1574_ Tile_X0Y1_FrameData[20] Tile_X0Y1_FrameData_O[20] VPWR VGND sg13g2_buf_1
X_0387_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit10.Q Tile_X0Y0_E1END[1]
+ Tile_X0Y0_E6END[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13
+ _0310_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit11.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1008_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_106_75 VPWR VGND sg13g2_decap_8
XFILLER_103_198 VPWR VGND sg13g2_fill_2
XFILLER_103_187 VPWR VGND sg13g2_decap_8
XFILLER_103_132 VPWR VGND sg13g2_decap_8
XFILLER_17_105 VPWR VGND sg13g2_decap_4
XFILLER_99_119 VPWR VGND sg13g2_decap_8
X_1290_ Tile_X0Y1_FrameData[29] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit29.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_90 VPWR VGND sg13g2_fill_1
XFILLER_31_141 VPWR VGND sg13g2_decap_4
XFILLER_68_0 VPWR VGND sg13g2_fill_2
X_1626_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG0 Tile_X0Y1_W2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1488_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb7 Tile_X0Y0_N2BEGb[7]
+ VPWR VGND sg13g2_buf_1
XFILLER_100_168 VPWR VGND sg13g2_decap_8
XFILLER_98_141 VPWR VGND sg13g2_decap_8
X_0439_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit13.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb2
+ Tile_X0Y0_S2MID[2] Tile_X0Y1_N2MID[2] Tile_X0Y0_S2END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit12.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 VPWR VGND sg13g2_mux4_1
X_0508_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit2.Q UIO_OUT_TT_PROJECT5
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit3.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG5 VPWR VGND sg13g2_mux4_1
X_1557_ Tile_X0Y1_FrameData[3] Tile_X0Y1_FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_77_34 VPWR VGND sg13g2_decap_8
XFILLER_93_66 VPWR VGND sg13g2_fill_2
XFILLER_42_92 VPWR VGND sg13g2_decap_8
X_0790_ _0151_ _0147_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit1.Q
+ _0180_ VPWR VGND sg13g2_mux2_1
X_1342_ Tile_X0Y1_FrameData[9] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit9.Q
+ VPWR VGND sg13g2_dlhq_1
X_1273_ Tile_X0Y1_FrameData[14] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit14.Q
+ VPWR VGND sg13g2_dlhq_1
X_1411_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_0988_ Tile_X0Y0_FrameData[19] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit19.Q
+ VPWR VGND sg13g2_dlhq_1
X_1609_ Tile_X0Y0_S4END[11] Tile_X0Y1_S4BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_86_177 VPWR VGND sg13g2_fill_2
XFILLER_86_166 VPWR VGND sg13g2_decap_8
XFILLER_86_133 VPWR VGND sg13g2_fill_2
XFILLER_10_166 VPWR VGND sg13g2_fill_2
XFILLER_88_66 VPWR VGND sg13g2_fill_2
XFILLER_77_199 VPWR VGND sg13g2_fill_1
X_0842_ _0147_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q
+ _0224_ VPWR VGND sg13g2_nor2b_1
X_0911_ RST_N_TT_PROJECT _0281_ _0286_ _0277_ _0307_ VPWR VGND sg13g2_a22oi_1
X_0773_ VGND VPWR _0160_ _0163_ Tile_X0Y0_E_TT_IF2_top.N4BEG_outbuf_8.A _0165_ sg13g2_a21oi_1
XFILLER_68_199 VPWR VGND sg13g2_fill_1
XFILLER_68_188 VPWR VGND sg13g2_fill_1
X_1325_ Tile_X0Y1_FrameData[26] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit26.Q
+ VPWR VGND sg13g2_dlhq_1
X_1256_ Tile_X0Y1_FrameData[31] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
X_1187_ Tile_X0Y1_FrameData[4] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_59_199 VPWR VGND sg13g2_fill_1
X_1110_ Tile_X0Y0_FrameData[25] Tile_X0Y1_FrameStrobe[6] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit25.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_2_173 VPWR VGND sg13g2_decap_8
X_1041_ Tile_X0Y0_FrameData[30] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit30.Q
+ VPWR VGND sg13g2_dlhq_1
X_0825_ VGND VPWR _0206_ _0208_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S4BEG3
+ _0210_ sg13g2_a21oi_1
X_0687_ _0121_ _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit22.Q
+ VPWR VGND sg13g2_nand2b_1
X_0756_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit20.Q Tile_X0Y1_N4END[2]
+ Tile_X0Y0_S4END[6] _0149_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit21.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_50_0 VPWR VGND sg13g2_decap_8
X_1308_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
X_1239_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_56_136 VPWR VGND sg13g2_decap_4
XFILLER_100_55 VPWR VGND sg13g2_fill_2
XFILLER_70_172 VPWR VGND sg13g2_fill_1
XFILLER_18_50 VPWR VGND sg13g2_decap_8
X_0610_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit13.Q Tile_X0Y0_E1END[3]
+ Tile_X0Y0_EE4END[15] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit15.Q
+ _0077_ VPWR VGND sg13g2_mux4_1
X_0541_ _0015_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame6_bit2.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG12 VPWR VGND sg13g2_nand2b_1
X_0472_ _0004_ Tile_X0Y0_S1END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
X_1590_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG0 Tile_X0Y1_S2BEG[0]
+ VPWR VGND sg13g2_buf_1
X_1024_ Tile_X0Y0_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0808_ VGND VPWR Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
+ _0195_ _0196_ _0302_ sg13g2_a21oi_1
X_0739_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit0.Q UO_OUT_TT_PROJECT0
+ UO_OUT_TT_PROJECT4 _0151_ _0003_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG8 VPWR VGND sg13g2_mux4_1
XFILLER_55_59 VPWR VGND sg13g2_decap_8
XFILLER_52_183 VPWR VGND sg13g2_fill_1
XFILLER_106_196 VPWR VGND sg13g2_decap_4
XFILLER_96_33 VPWR VGND sg13g2_fill_2
XFILLER_96_66 VPWR VGND sg13g2_fill_2
XANTENNA_2 VPWR VGND Tile_X0Y1_FrameStrobe[10] sg13g2_antennanp
XFILLER_6_75 VPWR VGND sg13g2_fill_1
X_1642_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG0 Tile_X0Y1_W6BEG[0]
+ VPWR VGND sg13g2_buf_1
X_0524_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit18.Q UIO_OUT_TT_PROJECT1
+ UIO_OE_TT_PROJECT5 _0012_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG2
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit19.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG13
+ VPWR VGND sg13g2_mux4_1
X_1573_ Tile_X0Y1_FrameData[19] Tile_X0Y1_FrameData_O[19] VPWR VGND sg13g2_buf_1
X_0455_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit17.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb4
+ Tile_X0Y0_S2MID[4] Tile_X0Y1_N2MID[4] Tile_X0Y0_S2END[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit16.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG4 VPWR VGND sg13g2_mux4_1
X_0386_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit2.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1
+ Tile_X0Y1_N4END[5] Tile_X0Y0_S1END[1] Tile_X0Y0_S4END[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit3.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG13 VPWR VGND sg13g2_mux4_1
X_1007_ Tile_X0Y0_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_0 VPWR VGND sg13g2_fill_1
XFILLER_19_191 VPWR VGND sg13g2_decap_8
XFILLER_103_111 VPWR VGND sg13g2_decap_8
XFILLER_103_166 VPWR VGND sg13g2_decap_8
XFILLER_17_128 VPWR VGND sg13g2_decap_4
XFILLER_40_175 VPWR VGND sg13g2_fill_2
XFILLER_98_120 VPWR VGND sg13g2_decap_8
X_1625_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG3 Tile_X0Y1_W1BEG[3]
+ VPWR VGND sg13g2_buf_1
X_1556_ Tile_X0Y1_FrameData[2] Tile_X0Y1_FrameData_O[2] VPWR VGND sg13g2_buf_1
X_1487_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb6 Tile_X0Y0_N2BEGb[6]
+ VPWR VGND sg13g2_buf_1
XFILLER_100_147 VPWR VGND sg13g2_decap_8
XFILLER_98_197 VPWR VGND sg13g2_fill_2
X_0507_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit28.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit29.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG10 VPWR VGND sg13g2_mux4_1
X_0369_ VPWR _0299_ Tile_X0Y1_E6END[1] VGND sg13g2_inv_1
XFILLER_36_17 VPWR VGND sg13g2_fill_2
X_0438_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit12.Q Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2END[5] Tile_X0Y1_E6END[5] _0349_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit13.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb2 VPWR VGND sg13g2_mux4_1
XFILLER_93_34 VPWR VGND sg13g2_decap_8
XFILLER_26_83 VPWR VGND sg13g2_decap_4
X_1410_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_3_76 VPWR VGND sg13g2_fill_1
X_1341_ Tile_X0Y1_FrameData[10] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit10.Q
+ VPWR VGND sg13g2_dlhq_1
X_1272_ Tile_X0Y1_FrameData[15] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit15.Q
+ VPWR VGND sg13g2_dlhq_1
X_0987_ Tile_X0Y0_FrameData[20] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit20.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_80_0 VPWR VGND sg13g2_decap_8
X_1608_ Tile_X0Y0_S4END[10] Tile_X0Y1_S4BEG[2] VPWR VGND sg13g2_buf_1
X_1539_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG1 Tile_X0Y0_WW4BEG[1]
+ VPWR VGND sg13g2_buf_1
XFILLER_10_134 VPWR VGND sg13g2_fill_1
XFILLER_10_189 VPWR VGND sg13g2_decap_8
X_0772_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit26.Q _0164_
+ _0165_ VPWR VGND sg13g2_nor2_1
X_0841_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q _0155_
+ _0223_ VPWR VGND sg13g2_nor2_1
X_0910_ VGND VPWR _0283_ _0285_ _0286_ _0307_ sg13g2_a21oi_1
XFILLER_68_167 VPWR VGND sg13g2_fill_2
XFILLER_68_156 VPWR VGND sg13g2_decap_8
X_1324_ Tile_X0Y1_FrameData[27] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit27.Q
+ VPWR VGND sg13g2_dlhq_1
X_1255_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit0.Q
+ VPWR VGND sg13g2_dlhq_1
X_1186_ Tile_X0Y1_FrameData[5] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit5.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_181 VPWR VGND sg13g2_decap_8
XFILLER_2_141 VPWR VGND sg13g2_fill_1
X_1040_ Tile_X0Y0_FrameData[31] Tile_X0Y1_FrameStrobe[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame4_bit31.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_22 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
X_0755_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit18.Q Tile_X0Y1_N4END[1]
+ Tile_X0Y0_S4END[5] _0148_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG14
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit19.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG1
+ VPWR VGND sg13g2_mux4_1
X_0824_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit7.Q _0209_
+ _0210_ VPWR VGND sg13g2_nor2_1
X_0686_ VPWR VGND Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q
+ _0120_ _0119_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEG2 _0348_ sg13g2_a221oi_1
XFILLER_43_0 VPWR VGND sg13g2_decap_4
X_1307_ Tile_X0Y1_FrameData[12] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit12.Q
+ VPWR VGND sg13g2_dlhq_1
X_1238_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
X_1169_ Tile_X0Y1_FrameData[22] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit22.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_85_24 VPWR VGND sg13g2_decap_8
XFILLER_62_118 VPWR VGND sg13g2_decap_8
XFILLER_109_150 VPWR VGND sg13g2_fill_1
X_0471_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit30.Q Tile_X0Y0_E2MID[0]
+ Tile_X0Y0_E2END[0] Tile_X0Y0_E6END[0] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame7_bit31.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEG7
+ VPWR VGND sg13g2_mux4_1
X_0540_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit15.Q UIO_OUT_TT_PROJECT3
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG4 _0014_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit14.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.W6BEG11
+ VPWR VGND sg13g2_mux4_1
X_1023_ Tile_X0Y0_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
X_0807_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 _0001_
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit31.Q _0195_ VPWR
+ VGND sg13g2_mux2_1
X_0738_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit22.Q Tile_X0Y1_N1END[3]
+ Tile_X0Y1_N4END[3] _0325_ Tile_X0Y0_S4END[7] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame1_bit23.Q
+ _0151_ VPWR VGND sg13g2_mux4_1
X_0669_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit18.Q Tile_X0Y1_E2MID[4]
+ Tile_X0Y1_E2END[4] Tile_X0Y1_E6END[11] _0356_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit19.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG3 VPWR VGND sg13g2_mux4_1
XFILLER_52_162 VPWR VGND sg13g2_decap_8
XFILLER_106_175 VPWR VGND sg13g2_decap_8
XFILLER_106_131 VPWR VGND sg13g2_decap_8
XFILLER_29_83 VPWR VGND sg13g2_decap_8
XFILLER_28_181 VPWR VGND sg13g2_decap_8
XFILLER_35_118 VPWR VGND sg13g2_decap_4
XFILLER_61_70 VPWR VGND sg13g2_fill_1
XFILLER_45_93 VPWR VGND sg13g2_fill_2
XANTENNA_3 VPWR VGND Tile_X0Y1_FrameStrobe[11] sg13g2_antennanp
X_1641_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb7 Tile_X0Y1_W2BEGb[7]
+ VPWR VGND sg13g2_buf_1
X_1572_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameData_O[18] VPWR VGND sg13g2_buf_1
X_0523_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit12.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END2
+ Tile_X0Y1_N4END[6] Tile_X0Y0_S1END[2] Tile_X0Y0_S4END[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit13.Q
+ _0012_ VPWR VGND sg13g2_mux4_1
X_0385_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit3.Q Tile_X0Y1_E1END[1]
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG13 Tile_X0Y1_E6END[5]
+ _0314_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit2.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END1
+ VPWR VGND sg13g2_mux4_1
X_0454_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit16.Q Tile_X0Y1_E2MID[3]
+ Tile_X0Y1_E2END[3] Tile_X0Y1_E6END[3] _0000_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit17.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb4 VPWR VGND sg13g2_mux4_1
X_1006_ Tile_X0Y0_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_82_14 VPWR VGND sg13g2_fill_1
XFILLER_82_47 VPWR VGND sg13g2_fill_2
XFILLER_82_36 VPWR VGND sg13g2_decap_8
XFILLER_15_30 VPWR VGND sg13g2_decap_4
XFILLER_25_140 VPWR VGND sg13g2_decap_8
XFILLER_25_184 VPWR VGND sg13g2_decap_8
XFILLER_110_0 VPWR VGND sg13g2_decap_8
XFILLER_40_198 VPWR VGND sg13g2_fill_2
XFILLER_16_184 VPWR VGND sg13g2_decap_8
XFILLER_31_121 VPWR VGND sg13g2_fill_2
X_0506_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit0.Q UIO_OUT_TT_PROJECT4
+ UIO_OE_TT_PROJECT0 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3 Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit1.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG4 VPWR VGND sg13g2_mux4_1
X_1624_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG2 Tile_X0Y1_W1BEG[2]
+ VPWR VGND sg13g2_buf_1
X_1555_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameData_O[1] VPWR VGND sg13g2_buf_1
X_1486_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb5 Tile_X0Y0_N2BEGb[5]
+ VPWR VGND sg13g2_buf_1
XFILLER_100_126 VPWR VGND sg13g2_decap_8
XFILLER_98_176 VPWR VGND sg13g2_decap_8
X_0368_ VPWR _0298_ Tile_X0Y1_E6END[2] VGND sg13g2_inv_1
X_0437_ _0344_ _0347_ _0349_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_17 VPWR VGND sg13g2_decap_8
XFILLER_89_198 VPWR VGND sg13g2_fill_2
X_1340_ Tile_X0Y1_FrameData[11] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit11.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_95_179 VPWR VGND sg13g2_decap_8
XFILLER_95_146 VPWR VGND sg13g2_decap_8
X_1271_ Tile_X0Y1_FrameData[16] Tile_X0Y1_FrameStrobe[3] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q
+ VPWR VGND sg13g2_dlhq_1
Xclkbuf_0_Tile_X0Y1_UserCLK Tile_X0Y1_UserCLK clknet_0_Tile_X0Y1_UserCLK VPWR VGND
+ sg13g2_buf_8
X_0986_ Tile_X0Y0_FrameData[21] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit21.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_73_0 VPWR VGND sg13g2_fill_2
X_1607_ Tile_X0Y0_S4END[9] Tile_X0Y1_S4BEG[1] VPWR VGND sg13g2_buf_1
X_1469_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1BEG0 Tile_X0Y0_N1BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_86_102 VPWR VGND sg13g2_decap_8
X_1538_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG0 Tile_X0Y0_WW4BEG[0]
+ VPWR VGND sg13g2_buf_1
XFILLER_103_78 VPWR VGND sg13g2_fill_2
XFILLER_88_68 VPWR VGND sg13g2_fill_1
XFILLER_12_53 VPWR VGND sg13g2_decap_8
XFILLER_6_139 VPWR VGND sg13g2_decap_4
XFILLER_92_116 VPWR VGND sg13g2_decap_8
XFILLER_85_190 VPWR VGND sg13g2_decap_8
X_0771_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit25.Q Tile_X0Y1_E1END[0]
+ Tile_X0Y1_E6END[8] Tile_X0Y1_EE4END[0] _0158_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame7_bit24.Q
+ _0164_ VPWR VGND sg13g2_mux4_1
X_0840_ _0221_ _0222_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit16.Q
+ UI_IN_TT_PROJECT2 VPWR VGND sg13g2_mux2_1
XFILLER_5_194 VPWR VGND sg13g2_decap_4
X_1323_ Tile_X0Y1_FrameData[28] Tile_X0Y1_FrameStrobe[5] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit28.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_83_127 VPWR VGND sg13g2_fill_2
X_1254_ Tile_X0Y1_FrameData[1] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit1.Q
+ VPWR VGND sg13g2_dlhq_1
X_1185_ Tile_X0Y1_FrameData[6] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
X_0969_ Tile_X0Y0_FrameData[6] Tile_X0Y1_FrameStrobe[1] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit6.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_99_23 VPWR VGND sg13g2_decap_8
XFILLER_3_0 VPWR VGND sg13g2_fill_2
XFILLER_73_193 VPWR VGND sg13g2_decap_8
X_0685_ UO_OUT_TT_PROJECT2 Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit20.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit21.Q _0120_ VPWR
+ VGND sg13g2_nor3_1
X_0754_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit16.Q Tile_X0Y1_N4END[0]
+ Tile_X0Y0_S4END[4] _0147_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.J_NS4_BEG15
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame3_bit17.Q Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W6BEG0
+ VPWR VGND sg13g2_mux4_1
X_0823_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit5.Q Tile_X0Y1_E1END[3]
+ Tile_X0Y1_EE4END[15] Tile_X0Y1_E6END[7] _0155_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit6.Q
+ _0209_ VPWR VGND sg13g2_mux4_1
X_1306_ Tile_X0Y1_FrameData[13] Tile_X0Y1_FrameStrobe[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit13.Q
+ VPWR VGND sg13g2_dlhq_1
X_1099_ Tile_X0Y0_FrameData[4] Tile_X0Y1_FrameStrobe[5] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit4.Q
+ VPWR VGND sg13g2_dlhq_1
X_1237_ Tile_X0Y1_FrameData[18] Tile_X0Y1_FrameStrobe[2] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame2_bit18.Q
+ VPWR VGND sg13g2_dlhq_1
X_1168_ Tile_X0Y1_FrameData[23] Tile_X0Y1_FrameStrobe[0] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit23.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_60_17 VPWR VGND sg13g2_decap_8
XFILLER_70_130 VPWR VGND sg13g2_fill_1
X_0470_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit23.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb7
+ Tile_X0Y0_S2MID[7] Tile_X0Y1_N2MID[7] Tile_X0Y0_S2END[7] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame0_bit22.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG7 VPWR VGND sg13g2_mux4_1
XFILLER_59_70 VPWR VGND sg13g2_decap_8
X_1022_ Tile_X0Y0_FrameData[17] Tile_X0Y1_FrameStrobe[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_61_141 VPWR VGND sg13g2_fill_2
XFILLER_46_182 VPWR VGND sg13g2_fill_2
X_0737_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit31.Q UO_OUT_TT_PROJECT3
+ _0150_ UO_OUT_TT_PROJECT7 _0335_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame4_bit30.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.WW4BEG7 VPWR VGND sg13g2_mux4_1
X_0806_ _0194_ _0193_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame5_bit0.Q
+ VPWR VGND sg13g2_nand2b_1
X_0668_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit16.Q Tile_X0Y1_E2MID[5]
+ Tile_X0Y1_E2END[5] Tile_X0Y1_E6END[10] _0349_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame6_bit17.Q
+ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.S2BEG2 VPWR VGND sg13g2_mux4_1
X_0599_ _0066_ VPWR _0067_ VGND Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame5_bit12.Q
+ _0012_ sg13g2_o21ai_1
XFILLER_55_17 VPWR VGND sg13g2_decap_4
XFILLER_71_38 VPWR VGND sg13g2_decap_4
XFILLER_52_141 VPWR VGND sg13g2_decap_8
XFILLER_106_110 VPWR VGND sg13g2_decap_8
XFILLER_106_154 VPWR VGND sg13g2_decap_8
XFILLER_96_57 VPWR VGND sg13g2_fill_1
XFILLER_96_35 VPWR VGND sg13g2_fill_1
XFILLER_20_75 VPWR VGND sg13g2_decap_8
XFILLER_43_185 VPWR VGND sg13g2_decap_8
XANTENNA_4 VPWR VGND Tile_X0Y1_FrameStrobe[12] sg13g2_antennanp
X_0522_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit16.Q UIO_OUT_TT_PROJECT0
+ UIO_OE_TT_PROJECT4 _0011_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS2_BEG3
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame3_bit17.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.WW4BEG12
+ VPWR VGND sg13g2_mux4_1
X_1640_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W2BEGb6 Tile_X0Y1_W2BEGb[6]
+ VPWR VGND sg13g2_buf_1
X_1571_ Tile_X0Y1_FrameData[17] Tile_X0Y1_FrameData_O[17] VPWR VGND sg13g2_buf_1
X_0384_ VPWR VGND _0312_ _0313_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit27.Q
+ _0299_ _0314_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a221oi_1
X_0453_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit16.Q Tile_X0Y1_N2MID[4]
+ Tile_X0Y1_N2END[4] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.S2BEG4
+ Tile_X0Y0_S2MID[4] Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_ConfigMem.Inst_frame0_bit17.Q
+ _0000_ VPWR VGND sg13g2_mux4_1
X_1005_ Tile_X0Y0_FrameData[2] Tile_X0Y1_FrameStrobe[2] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame2_bit2.Q
+ VPWR VGND sg13g2_dlhq_1
XFILLER_34_130 VPWR VGND sg13g2_decap_4
XFILLER_103_146 VPWR VGND sg13g2_decap_8
XFILLER_106_89 VPWR VGND sg13g2_decap_8
XFILLER_103_0 VPWR VGND sg13g2_decap_8
XFILLER_31_199 VPWR VGND sg13g2_fill_1
X_1485_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N2BEGb4 Tile_X0Y0_N2BEGb[4]
+ VPWR VGND sg13g2_buf_1
X_0505_ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit30.Q Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.N1END3
+ Tile_X0Y1_N4END[7] Tile_X0Y0_S1END[3] Tile_X0Y0_S4END[3] Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_ConfigMem.Inst_frame1_bit31.Q
+ Tile_X0Y0_E_TT_IF2_top.Inst_E_TT_IF2_top_switch_matrix.J_NS4_BEG11 VPWR VGND sg13g2_mux4_1
XFILLER_98_199 VPWR VGND sg13g2_fill_1
XFILLER_98_155 VPWR VGND sg13g2_decap_8
X_1623_ Tile_X0Y1_E_TT_IF2_bot.Inst_E_TT_IF2_bot_switch_matrix.W1BEG1 Tile_X0Y1_W1BEG[1]
+ VPWR VGND sg13g2_buf_1
X_0436_ _0348_ _0347_ _0344_ VPWR VGND sg13g2_nand2b_1
X_1554_ Tile_X0Y1_FrameData[0] Tile_X0Y1_FrameData_O[0] VPWR VGND sg13g2_buf_1
.ends

