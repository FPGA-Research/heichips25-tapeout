* NGSPICE file created from heichips25_example_small.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xor2_1 abstract view
.subckt sg13g2_xor2_1 B A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_xnor2_1 abstract view
.subckt sg13g2_xnor2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tielo abstract view
.subckt sg13g2_tielo VDD VSS L_LO
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_a21oi_2 abstract view
.subckt sg13g2_a21oi_2 VSS VDD B1 Y A2 A1
.ends

.subckt heichips25_example_small VGND VPWR clk ena rst_n ui_in[0] ui_in[1] ui_in[2]
+ ui_in[3] ui_in[4] ui_in[5] ui_in[6] ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3]
+ uio_in[4] uio_in[5] uio_in[6] uio_in[7] uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3]
+ uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7] uio_out[0] uio_out[1] uio_out[2] uio_out[3]
+ uio_out[4] uio_out[5] uio_out[6] uio_out[7] uo_out[0] uo_out[1] uo_out[2] uo_out[3]
+ uo_out[4] uo_out[5] uo_out[6] uo_out[7]
XFILLER_27_406 VPWR VGND sg13g2_decap_8
XFILLER_39_266 VPWR VGND sg13g2_decap_8
XFILLER_35_450 VPWR VGND sg13g2_decap_8
XFILLER_23_634 VPWR VGND sg13g2_decap_8
XFILLER_22_144 VPWR VGND sg13g2_decap_8
XFILLER_7_7 VPWR VGND sg13g2_decap_8
XFILLER_19_907 VPWR VGND sg13g2_decap_8
XFILLER_18_417 VPWR VGND sg13g2_decap_8
XFILLER_45_214 VPWR VGND sg13g2_decap_8
XFILLER_14_634 VPWR VGND sg13g2_decap_8
XFILLER_26_494 VPWR VGND sg13g2_decap_8
XFILLER_13_144 VPWR VGND sg13g2_decap_8
XFILLER_41_464 VPWR VGND sg13g2_decap_8
XFILLER_9_137 VPWR VGND sg13g2_decap_8
XFILLER_10_851 VPWR VGND sg13g2_decap_8
XFILLER_6_844 VPWR VGND sg13g2_decap_8
XFILLER_5_354 VPWR VGND sg13g2_decap_8
XFILLER_1_560 VPWR VGND sg13g2_decap_8
XFILLER_3_67 VPWR VGND sg13g2_decap_8
XFILLER_49_553 VPWR VGND sg13g2_decap_8
XFILLER_36_214 VPWR VGND sg13g2_decap_8
XFILLER_17_483 VPWR VGND sg13g2_decap_8
XFILLER_45_781 VPWR VGND sg13g2_decap_8
XFILLER_32_431 VPWR VGND sg13g2_decap_8
XFILLER_44_291 VPWR VGND sg13g2_decap_8
XFILLER_20_648 VPWR VGND sg13g2_decap_8
XFILLER_27_203 VPWR VGND sg13g2_decap_8
XFILLER_28_748 VPWR VGND sg13g2_decap_8
XFILLER_43_718 VPWR VGND sg13g2_decap_8
XFILLER_36_781 VPWR VGND sg13g2_decap_8
XFILLER_23_431 VPWR VGND sg13g2_decap_8
XFILLER_42_239 VPWR VGND sg13g2_decap_8
XFILLER_11_648 VPWR VGND sg13g2_decap_8
XFILLER_10_158 VPWR VGND sg13g2_decap_8
XFILLER_12_32 VPWR VGND sg13g2_decap_8
XFILLER_5_4 VPWR VGND sg13g2_decap_8
XFILLER_3_858 VPWR VGND sg13g2_decap_8
XFILLER_2_368 VPWR VGND sg13g2_decap_8
XFILLER_19_704 VPWR VGND sg13g2_decap_8
XFILLER_18_214 VPWR VGND sg13g2_decap_8
XFILLER_46_567 VPWR VGND sg13g2_decap_8
XFILLER_37_84 VPWR VGND sg13g2_decap_8
XFILLER_15_921 VPWR VGND sg13g2_decap_4
XFILLER_27_770 VPWR VGND sg13g2_decap_8
XFILLER_14_431 VPWR VGND sg13g2_decap_8
XFILLER_26_291 VPWR VGND sg13g2_decap_8
XFILLER_41_261 VPWR VGND sg13g2_decap_8
XFILLER_6_641 VPWR VGND sg13g2_decap_8
XFILLER_5_151 VPWR VGND sg13g2_decap_8
XFILLER_38_4 VPWR VGND sg13g2_decap_8
XFILLER_49_350 VPWR VGND sg13g2_decap_8
XFILLER_37_567 VPWR VGND sg13g2_decap_8
XFILLER_18_781 VPWR VGND sg13g2_decap_8
XFILLER_17_280 VPWR VGND sg13g2_decap_8
XFILLER_33_751 VPWR VGND sg13g2_decap_8
XFILLER_20_445 VPWR VGND sg13g2_decap_8
XFILLER_28_545 VPWR VGND sg13g2_decap_8
XFILLER_16_718 VPWR VGND sg13g2_decap_8
XFILLER_43_515 VPWR VGND sg13g2_decap_8
XFILLER_15_228 VPWR VGND sg13g2_decap_8
XFILLER_24_740 VPWR VGND sg13g2_decap_8
XFILLER_11_445 VPWR VGND sg13g2_decap_8
XFILLER_23_53 VPWR VGND sg13g2_decap_8
XFILLER_7_427 VPWR VGND sg13g2_decap_8
XFILLER_3_655 VPWR VGND sg13g2_decap_8
XFILLER_2_165 VPWR VGND sg13g2_decap_8
XFILLER_19_501 VPWR VGND sg13g2_decap_8
XFILLER_47_854 VPWR VGND sg13g2_decap_8
XFILLER_0_35 VPWR VGND sg13g2_decap_8
XFILLER_46_364 VPWR VGND sg13g2_decap_8
XFILLER_19_578 VPWR VGND sg13g2_decap_8
XFILLER_34_559 VPWR VGND sg13g2_decap_8
XFILLER_9_11 VPWR VGND sg13g2_decap_8
XFILLER_15_795 VPWR VGND sg13g2_decap_8
XFILLER_9_88 VPWR VGND sg13g2_decap_8
XFILLER_30_765 VPWR VGND sg13g2_decap_8
XFILLER_38_810 VPWR VGND sg13g2_decap_8
X_49_ _17_ _13_ _15_ VPWR VGND sg13g2_nand2_1
XFILLER_37_364 VPWR VGND sg13g2_decap_8
XFILLER_38_887 VPWR VGND sg13g2_decap_8
XFILLER_25_559 VPWR VGND sg13g2_decap_8
XFILLER_21_732 VPWR VGND sg13g2_decap_8
XFILLER_40_529 VPWR VGND sg13g2_decap_8
XFILLER_20_242 VPWR VGND sg13g2_decap_8
XFILLER_0_658 VPWR VGND sg13g2_decap_8
XFILLER_29_810 VPWR VGND sg13g2_decap_8
XFILLER_18_53 VPWR VGND sg13g2_decap_8
XFILLER_28_342 VPWR VGND sg13g2_decap_8
XFILLER_16_515 VPWR VGND sg13g2_decap_8
XFILLER_29_887 VPWR VGND sg13g2_decap_8
XFILLER_44_802 VPWR VGND sg13g2_decap_8
XFILLER_43_312 VPWR VGND sg13g2_decap_8
XFILLER_31_507 VPWR VGND sg13g2_decap_8
XFILLER_44_879 VPWR VGND sg13g2_decap_8
XFILLER_34_63 VPWR VGND sg13g2_decap_8
XFILLER_43_389 VPWR VGND sg13g2_decap_8
XFILLER_12_732 VPWR VGND sg13g2_decap_8
XFILLER_11_242 VPWR VGND sg13g2_decap_8
XFILLER_8_725 VPWR VGND sg13g2_decap_8
XFILLER_7_224 VPWR VGND sg13g2_decap_8
XFILLER_3_452 VPWR VGND sg13g2_decap_8
XFILLER_38_117 VPWR VGND sg13g2_decap_8
XFILLER_47_651 VPWR VGND sg13g2_decap_8
XFILLER_19_375 VPWR VGND sg13g2_decap_8
XFILLER_46_161 VPWR VGND sg13g2_decap_8
XFILLER_35_835 VPWR VGND sg13g2_decap_8
XFILLER_34_356 VPWR VGND sg13g2_decap_8
XFILLER_22_529 VPWR VGND sg13g2_decap_8
XFILLER_15_592 VPWR VGND sg13g2_decap_8
XFILLER_30_562 VPWR VGND sg13g2_decap_8
XFILLER_7_791 VPWR VGND sg13g2_decap_8
XFILLER_26_802 VPWR VGND sg13g2_decap_8
XFILLER_44_109 VPWR VGND sg13g2_decap_8
XFILLER_37_161 VPWR VGND sg13g2_decap_8
XFILLER_38_684 VPWR VGND sg13g2_decap_8
XFILLER_25_356 VPWR VGND sg13g2_decap_8
XFILLER_26_879 VPWR VGND sg13g2_decap_8
XFILLER_13_529 VPWR VGND sg13g2_decap_8
XFILLER_40_326 VPWR VGND sg13g2_decap_8
XFILLER_41_849 VPWR VGND sg13g2_decap_8
XFILLER_5_739 VPWR VGND sg13g2_decap_8
XFILLER_4_249 VPWR VGND sg13g2_decap_8
XFILLER_20_32 VPWR VGND sg13g2_decap_8
XFILLER_0_455 VPWR VGND sg13g2_decap_8
XFILLER_48_448 VPWR VGND sg13g2_decap_8
XFILLER_29_74 VPWR VGND sg13g2_decap_8
XFILLER_16_312 VPWR VGND sg13g2_decap_8
XFILLER_29_684 VPWR VGND sg13g2_decap_8
XFILLER_17_868 VPWR VGND sg13g2_decap_8
XFILLER_32_816 VPWR VGND sg13g2_decap_8
XFILLER_44_676 VPWR VGND sg13g2_decap_8
XFILLER_16_389 VPWR VGND sg13g2_decap_8
XFILLER_31_304 VPWR VGND sg13g2_decap_8
XFILLER_43_186 VPWR VGND sg13g2_decap_8
XFILLER_45_95 VPWR VGND sg13g2_decap_8
XFILLER_8_522 VPWR VGND sg13g2_decap_8
XFILLER_40_893 VPWR VGND sg13g2_decap_8
XFILLER_8_599 VPWR VGND sg13g2_decap_8
XFILLER_6_67 VPWR VGND sg13g2_decap_8
XFILLER_20_4 VPWR VGND sg13g2_decap_8
XFILLER_39_448 VPWR VGND sg13g2_decap_8
XFILLER_26_109 VPWR VGND sg13g2_decap_8
XFILLER_19_172 VPWR VGND sg13g2_decap_8
XFILLER_35_632 VPWR VGND sg13g2_decap_8
XFILLER_23_816 VPWR VGND sg13g2_decap_8
XFILLER_34_153 VPWR VGND sg13g2_decap_8
XFILLER_22_326 VPWR VGND sg13g2_decap_8
XFILLER_31_871 VPWR VGND sg13g2_decap_8
XFILLER_38_481 VPWR VGND sg13g2_decap_8
XFILLER_14_816 VPWR VGND sg13g2_decap_8
XFILLER_15_32 VPWR VGND sg13g2_decap_8
XFILLER_25_153 VPWR VGND sg13g2_decap_8
XFILLER_26_676 VPWR VGND sg13g2_decap_8
XFILLER_13_326 VPWR VGND sg13g2_decap_8
XFILLER_40_123 VPWR VGND sg13g2_decap_8
XFILLER_41_646 VPWR VGND sg13g2_decap_8
XFILLER_9_319 VPWR VGND sg13g2_decap_8
XFILLER_22_893 VPWR VGND sg13g2_decap_8
XFILLER_5_536 VPWR VGND sg13g2_decap_8
Xoutput20 net20 uo_out[3] VPWR VGND sg13g2_buf_1
XFILLER_1_742 VPWR VGND sg13g2_decap_8
XFILLER_0_252 VPWR VGND sg13g2_decap_8
XFILLER_49_735 VPWR VGND sg13g2_decap_8
XFILLER_48_245 VPWR VGND sg13g2_decap_8
XFILLER_29_481 VPWR VGND sg13g2_decap_8
XFILLER_17_665 VPWR VGND sg13g2_decap_8
XFILLER_32_613 VPWR VGND sg13g2_decap_8
XFILLER_44_473 VPWR VGND sg13g2_decap_8
XFILLER_16_186 VPWR VGND sg13g2_decap_8
XFILLER_13_893 VPWR VGND sg13g2_decap_8
XFILLER_31_178 VPWR VGND sg13g2_decap_8
XFILLER_40_690 VPWR VGND sg13g2_decap_8
XFILLER_9_886 VPWR VGND sg13g2_decap_8
XFILLER_8_396 VPWR VGND sg13g2_decap_8
XFILLER_39_245 VPWR VGND sg13g2_decap_8
XFILLER_23_613 VPWR VGND sg13g2_decap_8
XFILLER_22_123 VPWR VGND sg13g2_decap_8
XFILLER_46_749 VPWR VGND sg13g2_decap_8
XFILLER_14_613 VPWR VGND sg13g2_decap_8
XFILLER_26_75 VPWR VGND sg13g2_decap_4
XFILLER_26_473 VPWR VGND sg13g2_decap_8
XFILLER_42_911 VPWR VGND sg13g2_decap_8
XFILLER_13_123 VPWR VGND sg13g2_decap_8
XFILLER_9_116 VPWR VGND sg13g2_decap_8
XFILLER_41_443 VPWR VGND sg13g2_decap_8
XFILLER_10_830 VPWR VGND sg13g2_decap_8
XFILLER_22_690 VPWR VGND sg13g2_decap_8
XFILLER_42_85 VPWR VGND sg13g2_decap_8
XFILLER_6_823 VPWR VGND sg13g2_decap_8
XFILLER_5_333 VPWR VGND sg13g2_decap_8
XFILLER_3_46 VPWR VGND sg13g2_decap_8
XFILLER_49_532 VPWR VGND sg13g2_decap_8
XFILLER_37_749 VPWR VGND sg13g2_decap_8
XFILLER_17_462 VPWR VGND sg13g2_decap_8
XFILLER_45_760 VPWR VGND sg13g2_decap_8
XFILLER_32_410 VPWR VGND sg13g2_decap_8
XFILLER_44_270 VPWR VGND sg13g2_decap_8
XFILLER_20_627 VPWR VGND sg13g2_decap_8
XFILLER_32_487 VPWR VGND sg13g2_decap_8
XFILLER_13_690 VPWR VGND sg13g2_decap_8
XFILLER_9_683 VPWR VGND sg13g2_decap_8
XFILLER_8_193 VPWR VGND sg13g2_decap_8
XFILLER_28_727 VPWR VGND sg13g2_decap_8
XFILLER_27_259 VPWR VGND sg13g2_decap_8
XFILLER_24_922 VPWR VGND sg13g2_fill_2
XFILLER_36_760 VPWR VGND sg13g2_decap_8
XFILLER_42_218 VPWR VGND sg13g2_decap_8
XFILLER_23_410 VPWR VGND sg13g2_decap_8
XFILLER_11_627 VPWR VGND sg13g2_decap_8
XFILLER_23_487 VPWR VGND sg13g2_decap_8
XFILLER_10_137 VPWR VGND sg13g2_decap_8
XFILLER_7_609 VPWR VGND sg13g2_decap_8
XFILLER_12_11 VPWR VGND sg13g2_decap_8
XFILLER_12_88 VPWR VGND sg13g2_decap_8
XFILLER_3_837 VPWR VGND sg13g2_decap_8
XFILLER_2_347 VPWR VGND sg13g2_decap_8
XFILLER_46_546 VPWR VGND sg13g2_decap_8
XFILLER_37_63 VPWR VGND sg13g2_decap_8
XFILLER_15_900 VPWR VGND sg13g2_decap_8
XFILLER_14_410 VPWR VGND sg13g2_decap_8
XFILLER_26_270 VPWR VGND sg13g2_decap_8
XFILLER_41_240 VPWR VGND sg13g2_decap_8
XFILLER_14_487 VPWR VGND sg13g2_decap_8
XFILLER_42_785 VPWR VGND sg13g2_decap_8
XFILLER_6_620 VPWR VGND sg13g2_decap_8
XFILLER_5_130 VPWR VGND sg13g2_decap_8
XFILLER_6_697 VPWR VGND sg13g2_decap_8
X_65_ net9 net1 net17 VPWR VGND sg13g2_xor2_1
XFILLER_37_546 VPWR VGND sg13g2_decap_8
XFILLER_18_760 VPWR VGND sg13g2_decap_8
XFILLER_24_229 VPWR VGND sg13g2_decap_8
XFILLER_33_730 VPWR VGND sg13g2_decap_8
XFILLER_21_914 VPWR VGND sg13g2_decap_8
XFILLER_20_424 VPWR VGND sg13g2_decap_8
XFILLER_32_284 VPWR VGND sg13g2_decap_8
XFILLER_9_480 VPWR VGND sg13g2_decap_8
XFILLER_28_524 VPWR VGND sg13g2_decap_8
XFILLER_15_207 VPWR VGND sg13g2_decap_8
XFILLER_12_914 VPWR VGND sg13g2_decap_8
XFILLER_11_424 VPWR VGND sg13g2_decap_8
XFILLER_24_796 VPWR VGND sg13g2_decap_8
XFILLER_8_907 VPWR VGND sg13g2_decap_8
XFILLER_7_406 VPWR VGND sg13g2_decap_8
XFILLER_23_32 VPWR VGND sg13g2_decap_8
XFILLER_23_284 VPWR VGND sg13g2_decap_8
XFILLER_3_634 VPWR VGND sg13g2_decap_8
XFILLER_2_144 VPWR VGND sg13g2_decap_8
XFILLER_47_833 VPWR VGND sg13g2_decap_8
XFILLER_48_84 VPWR VGND sg13g2_decap_8
XFILLER_46_343 VPWR VGND sg13g2_decap_8
XFILLER_0_14 VPWR VGND sg13g2_decap_8
XFILLER_19_557 VPWR VGND sg13g2_decap_8
XFILLER_34_538 VPWR VGND sg13g2_decap_8
XFILLER_15_774 VPWR VGND sg13g2_decap_8
XFILLER_42_582 VPWR VGND sg13g2_decap_8
XFILLER_9_67 VPWR VGND sg13g2_decap_8
XFILLER_14_284 VPWR VGND sg13g2_decap_8
XFILLER_30_744 VPWR VGND sg13g2_decap_8
XFILLER_6_494 VPWR VGND sg13g2_decap_8
XFILLER_38_866 VPWR VGND sg13g2_decap_8
X_48_ VPWR _16_ _15_ VGND sg13g2_inv_1
XFILLER_37_343 VPWR VGND sg13g2_decap_8
XFILLER_25_538 VPWR VGND sg13g2_decap_8
XFILLER_40_508 VPWR VGND sg13g2_decap_8
XFILLER_21_711 VPWR VGND sg13g2_decap_8
XFILLER_20_221 VPWR VGND sg13g2_decap_8
XFILLER_21_788 VPWR VGND sg13g2_decap_8
XFILLER_20_298 VPWR VGND sg13g2_decap_8
XFILLER_0_637 VPWR VGND sg13g2_decap_8
XFILLER_18_32 VPWR VGND sg13g2_decap_8
XFILLER_28_321 VPWR VGND sg13g2_decap_8
XFILLER_29_866 VPWR VGND sg13g2_decap_8
XFILLER_28_398 VPWR VGND sg13g2_decap_8
XFILLER_44_858 VPWR VGND sg13g2_decap_8
XFILLER_43_368 VPWR VGND sg13g2_decap_8
XFILLER_12_711 VPWR VGND sg13g2_decap_8
XFILLER_11_221 VPWR VGND sg13g2_decap_8
XFILLER_8_704 VPWR VGND sg13g2_decap_8
XFILLER_24_593 VPWR VGND sg13g2_decap_8
XFILLER_7_203 VPWR VGND sg13g2_decap_8
XFILLER_12_788 VPWR VGND sg13g2_decap_8
XFILLER_11_298 VPWR VGND sg13g2_decap_8
XFILLER_4_921 VPWR VGND sg13g2_decap_4
XFILLER_3_431 VPWR VGND sg13g2_decap_8
XFILLER_47_630 VPWR VGND sg13g2_decap_8
XFILLER_46_140 VPWR VGND sg13g2_decap_8
XFILLER_19_354 VPWR VGND sg13g2_decap_8
XFILLER_35_814 VPWR VGND sg13g2_decap_8
XFILLER_22_508 VPWR VGND sg13g2_decap_8
XFILLER_34_335 VPWR VGND sg13g2_decap_8
XFILLER_15_571 VPWR VGND sg13g2_decap_8
XFILLER_30_541 VPWR VGND sg13g2_decap_8
XFILLER_7_770 VPWR VGND sg13g2_decap_8
XFILLER_6_291 VPWR VGND sg13g2_decap_8
XFILLER_29_118 VPWR VGND sg13g2_fill_1
XFILLER_37_140 VPWR VGND sg13g2_decap_8
XFILLER_38_663 VPWR VGND sg13g2_decap_8
XFILLER_25_335 VPWR VGND sg13g2_decap_8
XFILLER_26_858 VPWR VGND sg13g2_decap_8
XFILLER_13_508 VPWR VGND sg13g2_decap_8
XFILLER_40_305 VPWR VGND sg13g2_decap_8
XFILLER_41_828 VPWR VGND sg13g2_decap_8
XFILLER_21_585 VPWR VGND sg13g2_decap_8
XFILLER_5_718 VPWR VGND sg13g2_decap_8
XFILLER_4_228 VPWR VGND sg13g2_decap_8
XFILLER_20_11 VPWR VGND sg13g2_decap_8
XFILLER_1_924 VPWR VGND sg13g2_fill_1
XFILLER_20_88 VPWR VGND sg13g2_decap_8
XFILLER_49_917 VPWR VGND sg13g2_decap_8
XFILLER_0_434 VPWR VGND sg13g2_decap_8
XFILLER_48_427 VPWR VGND sg13g2_decap_8
XFILLER_29_53 VPWR VGND sg13g2_decap_8
XFILLER_29_663 VPWR VGND sg13g2_decap_8
XFILLER_17_847 VPWR VGND sg13g2_decap_8
XFILLER_28_195 VPWR VGND sg13g2_decap_8
XFILLER_44_655 VPWR VGND sg13g2_decap_8
XFILLER_45_74 VPWR VGND sg13g2_decap_8
XFILLER_16_368 VPWR VGND sg13g2_decap_8
XFILLER_43_165 VPWR VGND sg13g2_decap_8
XFILLER_24_390 VPWR VGND sg13g2_decap_8
XFILLER_8_501 VPWR VGND sg13g2_decap_8
XFILLER_40_872 VPWR VGND sg13g2_decap_8
XFILLER_12_585 VPWR VGND sg13g2_decap_8
XFILLER_8_578 VPWR VGND sg13g2_decap_8
XFILLER_6_46 VPWR VGND sg13g2_decap_8
XFILLER_4_795 VPWR VGND sg13g2_decap_8
XFILLER_13_4 VPWR VGND sg13g2_decap_8
XFILLER_39_427 VPWR VGND sg13g2_decap_8
XFILLER_19_151 VPWR VGND sg13g2_decap_8
XFILLER_35_611 VPWR VGND sg13g2_decap_8
XFILLER_34_132 VPWR VGND sg13g2_decap_8
XFILLER_22_305 VPWR VGND sg13g2_decap_8
XFILLER_35_688 VPWR VGND sg13g2_decap_8
XFILLER_31_850 VPWR VGND sg13g2_decap_8
XFILLER_38_460 VPWR VGND sg13g2_decap_8
XFILLER_25_132 VPWR VGND sg13g2_decap_8
XFILLER_26_655 VPWR VGND sg13g2_decap_8
XFILLER_13_305 VPWR VGND sg13g2_decap_8
XFILLER_15_11 VPWR VGND sg13g2_decap_8
XFILLER_41_625 VPWR VGND sg13g2_decap_8
XFILLER_40_102 VPWR VGND sg13g2_decap_8
XFILLER_15_88 VPWR VGND sg13g2_decap_8
XFILLER_22_872 VPWR VGND sg13g2_decap_8
XFILLER_21_382 VPWR VGND sg13g2_decap_8
XFILLER_40_179 VPWR VGND sg13g2_decap_8
XFILLER_31_32 VPWR VGND sg13g2_decap_4
XFILLER_5_515 VPWR VGND sg13g2_decap_8
Xoutput21 net21 uo_out[4] VPWR VGND sg13g2_buf_1
XFILLER_1_721 VPWR VGND sg13g2_decap_8
XFILLER_49_714 VPWR VGND sg13g2_decap_8
XFILLER_0_231 VPWR VGND sg13g2_decap_8
XFILLER_48_224 VPWR VGND sg13g2_decap_8
XFILLER_1_798 VPWR VGND sg13g2_decap_8
XFILLER_29_460 VPWR VGND sg13g2_decap_8
XFILLER_17_644 VPWR VGND sg13g2_decap_8
XFILLER_16_165 VPWR VGND sg13g2_decap_8
XFILLER_44_452 VPWR VGND sg13g2_decap_8
XFILLER_13_872 VPWR VGND sg13g2_decap_8
XFILLER_20_809 VPWR VGND sg13g2_decap_8
XFILLER_31_157 VPWR VGND sg13g2_decap_8
XFILLER_32_669 VPWR VGND sg13g2_decap_8
XFILLER_12_382 VPWR VGND sg13g2_decap_8
XFILLER_9_865 VPWR VGND sg13g2_decap_8
XFILLER_8_375 VPWR VGND sg13g2_decap_8
XFILLER_4_592 VPWR VGND sg13g2_decap_8
XFILLER_39_224 VPWR VGND sg13g2_decap_8
XFILLER_28_909 VPWR VGND sg13g2_decap_8
XFILLER_48_791 VPWR VGND sg13g2_decap_8
XFILLER_22_102 VPWR VGND sg13g2_decap_8
XFILLER_35_485 VPWR VGND sg13g2_decap_8
XFILLER_11_809 VPWR VGND sg13g2_decap_8
XFILLER_23_669 VPWR VGND sg13g2_decap_8
XFILLER_10_319 VPWR VGND sg13g2_decap_8
XFILLER_22_179 VPWR VGND sg13g2_decap_8
XFILLER_2_529 VPWR VGND sg13g2_decap_8
XFILLER_46_728 VPWR VGND sg13g2_decap_8
XFILLER_39_791 VPWR VGND sg13g2_decap_8
XFILLER_45_249 VPWR VGND sg13g2_decap_8
XFILLER_26_54 VPWR VGND sg13g2_decap_8
XFILLER_26_452 VPWR VGND sg13g2_decap_8
XFILLER_13_102 VPWR VGND sg13g2_decap_8
XFILLER_41_422 VPWR VGND sg13g2_decap_8
XFILLER_14_669 VPWR VGND sg13g2_decap_8
XFILLER_13_179 VPWR VGND sg13g2_decap_8
XFILLER_41_499 VPWR VGND sg13g2_decap_8
XFILLER_6_802 VPWR VGND sg13g2_decap_8
XFILLER_42_64 VPWR VGND sg13g2_decap_8
XFILLER_10_886 VPWR VGND sg13g2_decap_8
XFILLER_5_312 VPWR VGND sg13g2_decap_8
XFILLER_6_879 VPWR VGND sg13g2_decap_8
XFILLER_5_389 VPWR VGND sg13g2_decap_8
XFILLER_3_25 VPWR VGND sg13g2_decap_8
XFILLER_49_511 VPWR VGND sg13g2_decap_8
XFILLER_1_595 VPWR VGND sg13g2_decap_8
XFILLER_49_588 VPWR VGND sg13g2_decap_8
XFILLER_37_728 VPWR VGND sg13g2_decap_8
XFILLER_36_249 VPWR VGND sg13g2_decap_8
XFILLER_17_441 VPWR VGND sg13g2_decap_8
XFILLER_33_912 VPWR VGND sg13g2_decap_8
XFILLER_33_923 VPWR VGND sg13g2_fill_2
XFILLER_20_606 VPWR VGND sg13g2_decap_8
XFILLER_32_466 VPWR VGND sg13g2_decap_8
XFILLER_9_662 VPWR VGND sg13g2_decap_8
XFILLER_8_172 VPWR VGND sg13g2_decap_8
XFILLER_28_706 VPWR VGND sg13g2_decap_8
XFILLER_27_238 VPWR VGND sg13g2_decap_8
XFILLER_24_901 VPWR VGND sg13g2_decap_8
XFILLER_35_282 VPWR VGND sg13g2_decap_8
XFILLER_11_606 VPWR VGND sg13g2_decap_8
XFILLER_23_466 VPWR VGND sg13g2_decap_8
XFILLER_10_116 VPWR VGND sg13g2_decap_8
XFILLER_6_109 VPWR VGND sg13g2_decap_8
XFILLER_12_67 VPWR VGND sg13g2_decap_8
XFILLER_3_816 VPWR VGND sg13g2_decap_8
XFILLER_2_326 VPWR VGND sg13g2_decap_8
XFILLER_46_525 VPWR VGND sg13g2_decap_8
XFILLER_19_739 VPWR VGND sg13g2_decap_8
XFILLER_37_42 VPWR VGND sg13g2_decap_8
XFILLER_18_249 VPWR VGND sg13g2_decap_8
XFILLER_33_219 VPWR VGND sg13g2_decap_8
XFILLER_42_764 VPWR VGND sg13g2_decap_8
XFILLER_14_466 VPWR VGND sg13g2_decap_8
XFILLER_41_296 VPWR VGND sg13g2_decap_8
XFILLER_10_683 VPWR VGND sg13g2_decap_8
XFILLER_6_676 VPWR VGND sg13g2_decap_8
XFILLER_5_186 VPWR VGND sg13g2_decap_8
XFILLER_2_893 VPWR VGND sg13g2_decap_8
XFILLER_1_392 VPWR VGND sg13g2_decap_8
XFILLER_37_525 VPWR VGND sg13g2_decap_8
X_64_ net24 _27_ _28_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_385 VPWR VGND sg13g2_decap_8
XFILLER_24_208 VPWR VGND sg13g2_decap_8
XFILLER_20_403 VPWR VGND sg13g2_decap_8
XFILLER_32_263 VPWR VGND sg13g2_decap_8
XFILLER_33_786 VPWR VGND sg13g2_decap_8
XFILLER_0_819 VPWR VGND sg13g2_decap_8
XFILLER_28_503 VPWR VGND sg13g2_decap_8
XFILLER_11_403 VPWR VGND sg13g2_decap_8
XFILLER_23_11 VPWR VGND sg13g2_decap_8
XFILLER_23_263 VPWR VGND sg13g2_decap_8
XFILLER_24_775 VPWR VGND sg13g2_decap_8
XFILLER_23_88 VPWR VGND sg13g2_decap_8
XFILLER_3_613 VPWR VGND sg13g2_decap_8
XFILLER_2_123 VPWR VGND sg13g2_decap_8
XFILLER_47_812 VPWR VGND sg13g2_decap_8
XFILLER_48_63 VPWR VGND sg13g2_decap_8
XFILLER_46_322 VPWR VGND sg13g2_decap_8
XFILLER_19_536 VPWR VGND sg13g2_decap_8
XFILLER_47_889 VPWR VGND sg13g2_decap_8
XFILLER_34_517 VPWR VGND sg13g2_decap_8
XFILLER_46_399 VPWR VGND sg13g2_decap_8
XFILLER_15_753 VPWR VGND sg13g2_decap_8
XFILLER_14_263 VPWR VGND sg13g2_decap_8
XFILLER_30_723 VPWR VGND sg13g2_decap_8
XFILLER_42_561 VPWR VGND sg13g2_decap_8
XFILLER_9_46 VPWR VGND sg13g2_decap_8
XFILLER_10_480 VPWR VGND sg13g2_decap_8
XFILLER_6_473 VPWR VGND sg13g2_decap_8
XFILLER_43_4 VPWR VGND sg13g2_decap_8
XFILLER_2_690 VPWR VGND sg13g2_decap_8
XFILLER_49_182 VPWR VGND sg13g2_decap_8
XFILLER_37_322 VPWR VGND sg13g2_decap_8
XFILLER_38_845 VPWR VGND sg13g2_decap_8
X_47_ net13 net5 _15_ VPWR VGND sg13g2_xor2_1
XFILLER_25_517 VPWR VGND sg13g2_decap_8
XFILLER_37_399 VPWR VGND sg13g2_decap_8
XFILLER_20_200 VPWR VGND sg13g2_decap_8
XFILLER_33_583 VPWR VGND sg13g2_decap_8
XFILLER_21_767 VPWR VGND sg13g2_decap_8
XFILLER_20_277 VPWR VGND sg13g2_decap_8
XFILLER_0_616 VPWR VGND sg13g2_decap_8
XFILLER_48_609 VPWR VGND sg13g2_decap_8
XFILLER_47_119 VPWR VGND sg13g2_decap_8
XFILLER_18_11 VPWR VGND sg13g2_decap_8
XFILLER_28_300 VPWR VGND sg13g2_decap_8
XFILLER_29_845 VPWR VGND sg13g2_decap_8
XFILLER_18_88 VPWR VGND sg13g2_decap_8
XFILLER_28_377 VPWR VGND sg13g2_decap_8
XFILLER_44_837 VPWR VGND sg13g2_decap_8
XFILLER_43_347 VPWR VGND sg13g2_decap_8
XFILLER_24_572 VPWR VGND sg13g2_decap_8
XFILLER_11_200 VPWR VGND sg13g2_decap_8
XFILLER_34_98 VPWR VGND sg13g2_decap_8
XFILLER_12_767 VPWR VGND sg13g2_decap_8
XFILLER_11_277 VPWR VGND sg13g2_decap_8
XFILLER_7_259 VPWR VGND sg13g2_decap_8
XFILLER_4_900 VPWR VGND sg13g2_decap_8
XFILLER_3_410 VPWR VGND sg13g2_decap_8
XFILLER_3_487 VPWR VGND sg13g2_decap_8
XFILLER_1_0 VPWR VGND sg13g2_decap_8
XFILLER_39_609 VPWR VGND sg13g2_decap_8
XFILLER_19_333 VPWR VGND sg13g2_decap_8
XFILLER_47_686 VPWR VGND sg13g2_decap_8
XFILLER_34_314 VPWR VGND sg13g2_decap_8
XFILLER_46_196 VPWR VGND sg13g2_decap_8
XFILLER_15_550 VPWR VGND sg13g2_decap_8
XFILLER_30_520 VPWR VGND sg13g2_decap_8
XFILLER_30_597 VPWR VGND sg13g2_decap_8
XFILLER_6_270 VPWR VGND sg13g2_decap_8
XFILLER_38_642 VPWR VGND sg13g2_decap_8
XFILLER_1_91 VPWR VGND sg13g2_decap_8
XFILLER_25_314 VPWR VGND sg13g2_decap_8
XFILLER_26_837 VPWR VGND sg13g2_decap_8
XFILLER_37_196 VPWR VGND sg13g2_decap_8
XFILLER_41_807 VPWR VGND sg13g2_decap_8
XFILLER_34_881 VPWR VGND sg13g2_decap_8
XFILLER_33_380 VPWR VGND sg13g2_decap_8
XFILLER_21_564 VPWR VGND sg13g2_decap_8
XFILLER_4_207 VPWR VGND sg13g2_decap_8
XFILLER_1_903 VPWR VGND sg13g2_decap_8
XFILLER_20_67 VPWR VGND sg13g2_decap_8
XFILLER_0_413 VPWR VGND sg13g2_decap_8
XFILLER_48_406 VPWR VGND sg13g2_decap_8
XFILLER_29_32 VPWR VGND sg13g2_decap_8
XFILLER_29_642 VPWR VGND sg13g2_decap_8
XFILLER_17_826 VPWR VGND sg13g2_decap_8
XFILLER_28_174 VPWR VGND sg13g2_decap_8
XFILLER_16_347 VPWR VGND sg13g2_decap_8
XFILLER_44_634 VPWR VGND sg13g2_decap_8
XFILLER_45_53 VPWR VGND sg13g2_decap_8
XFILLER_43_144 VPWR VGND sg13g2_decap_8
XFILLER_25_881 VPWR VGND sg13g2_decap_8
XFILLER_31_339 VPWR VGND sg13g2_decap_8
XFILLER_12_564 VPWR VGND sg13g2_decap_8
XFILLER_40_851 VPWR VGND sg13g2_decap_8
XFILLER_8_557 VPWR VGND sg13g2_decap_8
XFILLER_6_25 VPWR VGND sg13g2_decap_8
XFILLER_4_774 VPWR VGND sg13g2_decap_8
XFILLER_3_284 VPWR VGND sg13g2_decap_8
XFILLER_39_406 VPWR VGND sg13g2_decap_8
XFILLER_19_130 VPWR VGND sg13g2_decap_8
XFILLER_47_483 VPWR VGND sg13g2_decap_8
XFILLER_35_667 VPWR VGND sg13g2_decap_8
XFILLER_34_188 VPWR VGND sg13g2_decap_8
XFILLER_30_394 VPWR VGND sg13g2_decap_8
XFILLER_25_111 VPWR VGND sg13g2_decap_8
XFILLER_26_634 VPWR VGND sg13g2_decap_8
XFILLER_41_604 VPWR VGND sg13g2_decap_8
XFILLER_25_188 VPWR VGND sg13g2_decap_8
XFILLER_15_67 VPWR VGND sg13g2_decap_8
XFILLER_22_851 VPWR VGND sg13g2_decap_8
XFILLER_40_158 VPWR VGND sg13g2_decap_8
XFILLER_21_361 VPWR VGND sg13g2_decap_8
XFILLER_31_11 VPWR VGND sg13g2_decap_8
XFILLER_31_88 VPWR VGND sg13g2_decap_8
Xoutput22 net22 uo_out[5] VPWR VGND sg13g2_buf_1
XFILLER_1_700 VPWR VGND sg13g2_decap_8
XFILLER_0_210 VPWR VGND sg13g2_decap_8
XFILLER_1_777 VPWR VGND sg13g2_decap_8
XFILLER_48_203 VPWR VGND sg13g2_decap_8
XFILLER_0_287 VPWR VGND sg13g2_decap_8
XFILLER_45_921 VPWR VGND sg13g2_decap_4
XFILLER_17_623 VPWR VGND sg13g2_decap_8
XFILLER_44_431 VPWR VGND sg13g2_decap_8
XFILLER_16_144 VPWR VGND sg13g2_decap_8
XFILLER_32_648 VPWR VGND sg13g2_decap_8
XFILLER_13_851 VPWR VGND sg13g2_decap_8
XFILLER_31_136 VPWR VGND sg13g2_decap_8
XFILLER_9_844 VPWR VGND sg13g2_decap_8
XFILLER_12_361 VPWR VGND sg13g2_decap_8
XFILLER_8_354 VPWR VGND sg13g2_decap_8
XFILLER_4_571 VPWR VGND sg13g2_decap_8
XFILLER_39_203 VPWR VGND sg13g2_decap_8
XFILLER_48_770 VPWR VGND sg13g2_decap_8
XFILLER_36_921 VPWR VGND sg13g2_decap_4
XFILLER_47_280 VPWR VGND sg13g2_decap_8
XFILLER_35_464 VPWR VGND sg13g2_decap_8
XFILLER_23_648 VPWR VGND sg13g2_decap_8
XFILLER_22_158 VPWR VGND sg13g2_decap_8
XFILLER_30_191 VPWR VGND sg13g2_decap_8
XFILLER_2_508 VPWR VGND sg13g2_decap_8
XFILLER_46_707 VPWR VGND sg13g2_decap_8
XFILLER_27_910 VPWR VGND sg13g2_decap_8
XFILLER_39_770 VPWR VGND sg13g2_decap_8
XFILLER_26_11 VPWR VGND sg13g2_decap_8
XFILLER_26_431 VPWR VGND sg13g2_decap_8
XFILLER_45_228 VPWR VGND sg13g2_decap_8
XFILLER_14_648 VPWR VGND sg13g2_decap_8
XFILLER_26_88 VPWR VGND sg13g2_decap_8
XFILLER_41_401 VPWR VGND sg13g2_decap_8
XFILLER_13_158 VPWR VGND sg13g2_decap_8
XFILLER_41_478 VPWR VGND sg13g2_decap_8
XFILLER_42_32 VPWR VGND sg13g2_fill_2
XFILLER_42_43 VPWR VGND sg13g2_decap_8
XFILLER_10_865 VPWR VGND sg13g2_decap_8
XFILLER_6_858 VPWR VGND sg13g2_decap_8
XFILLER_5_368 VPWR VGND sg13g2_decap_8
XFILLER_1_574 VPWR VGND sg13g2_decap_8
XFILLER_49_567 VPWR VGND sg13g2_decap_8
XFILLER_37_707 VPWR VGND sg13g2_decap_8
XFILLER_18_921 VPWR VGND sg13g2_decap_4
XFILLER_17_420 VPWR VGND sg13g2_decap_8
XFILLER_36_228 VPWR VGND sg13g2_decap_8
XFILLER_17_497 VPWR VGND sg13g2_decap_8
XFILLER_45_795 VPWR VGND sg13g2_decap_8
XFILLER_32_445 VPWR VGND sg13g2_decap_8
XFILLER_9_641 VPWR VGND sg13g2_decap_8
XFILLER_8_151 VPWR VGND sg13g2_decap_8
XFILLER_27_217 VPWR VGND sg13g2_decap_8
XFILLER_24_924 VPWR VGND sg13g2_fill_1
XFILLER_35_261 VPWR VGND sg13g2_decap_8
XFILLER_36_795 VPWR VGND sg13g2_decap_8
XFILLER_23_445 VPWR VGND sg13g2_decap_8
XFILLER_12_46 VPWR VGND sg13g2_decap_8
XFILLER_2_305 VPWR VGND sg13g2_decap_8
XFILLER_46_504 VPWR VGND sg13g2_decap_8
XFILLER_19_718 VPWR VGND sg13g2_decap_8
XFILLER_37_21 VPWR VGND sg13g2_decap_8
XFILLER_18_228 VPWR VGND sg13g2_decap_8
XFILLER_37_98 VPWR VGND sg13g2_decap_8
XFILLER_27_784 VPWR VGND sg13g2_decap_8
XFILLER_14_445 VPWR VGND sg13g2_decap_8
XFILLER_30_905 VPWR VGND sg13g2_decap_8
XFILLER_42_743 VPWR VGND sg13g2_decap_8
XFILLER_41_275 VPWR VGND sg13g2_decap_8
XFILLER_10_662 VPWR VGND sg13g2_decap_8
XFILLER_6_655 VPWR VGND sg13g2_decap_8
XFILLER_5_165 VPWR VGND sg13g2_decap_8
XFILLER_2_872 VPWR VGND sg13g2_decap_8
XFILLER_1_371 VPWR VGND sg13g2_decap_8
XFILLER_49_364 VPWR VGND sg13g2_decap_8
XFILLER_37_504 VPWR VGND sg13g2_decap_8
X_63_ _28_ net8 net16 VPWR VGND sg13g2_xnor2_1
XFILLER_18_795 VPWR VGND sg13g2_decap_8
XFILLER_17_294 VPWR VGND sg13g2_decap_8
XFILLER_33_765 VPWR VGND sg13g2_decap_8
XFILLER_45_592 VPWR VGND sg13g2_decap_8
XFILLER_32_242 VPWR VGND sg13g2_decap_8
XFILLER_20_459 VPWR VGND sg13g2_decap_8
XFILLER_28_559 VPWR VGND sg13g2_decap_8
XFILLER_43_529 VPWR VGND sg13g2_decap_8
XFILLER_24_754 VPWR VGND sg13g2_decap_8
XFILLER_36_592 VPWR VGND sg13g2_decap_8
XFILLER_23_242 VPWR VGND sg13g2_decap_8
XFILLER_11_459 VPWR VGND sg13g2_decap_8
XFILLER_23_67 VPWR VGND sg13g2_decap_8
XFILLER_2_102 VPWR VGND sg13g2_decap_8
XFILLER_3_669 VPWR VGND sg13g2_decap_8
XFILLER_3_4 VPWR VGND sg13g2_decap_8
XFILLER_2_179 VPWR VGND sg13g2_decap_8
XFILLER_48_42 VPWR VGND sg13g2_decap_8
XFILLER_19_515 VPWR VGND sg13g2_decap_8
XFILLER_46_301 VPWR VGND sg13g2_decap_8
XFILLER_47_868 VPWR VGND sg13g2_decap_8
XFILLER_0_49 VPWR VGND sg13g2_decap_8
XFILLER_46_378 VPWR VGND sg13g2_decap_8
XFILLER_27_581 VPWR VGND sg13g2_decap_8
XFILLER_15_732 VPWR VGND sg13g2_decap_8
XFILLER_42_540 VPWR VGND sg13g2_decap_8
XFILLER_9_25 VPWR VGND sg13g2_decap_8
XFILLER_14_242 VPWR VGND sg13g2_decap_8
XFILLER_30_702 VPWR VGND sg13g2_decap_8
XFILLER_30_779 VPWR VGND sg13g2_decap_8
XFILLER_6_452 VPWR VGND sg13g2_decap_8
XFILLER_36_4 VPWR VGND sg13g2_decap_8
XFILLER_49_161 VPWR VGND sg13g2_decap_8
XFILLER_37_301 VPWR VGND sg13g2_decap_8
XFILLER_38_824 VPWR VGND sg13g2_decap_8
X_46_ _14_ net5 net13 VPWR VGND sg13g2_nand2_1
XFILLER_37_378 VPWR VGND sg13g2_decap_8
XFILLER_18_592 VPWR VGND sg13g2_decap_8
XFILLER_33_562 VPWR VGND sg13g2_decap_8
XFILLER_21_746 VPWR VGND sg13g2_decap_8
XFILLER_20_256 VPWR VGND sg13g2_decap_8
XFILLER_29_824 VPWR VGND sg13g2_decap_8
XFILLER_18_67 VPWR VGND sg13g2_decap_8
XFILLER_28_356 VPWR VGND sg13g2_decap_8
XFILLER_44_816 VPWR VGND sg13g2_decap_8
XFILLER_16_529 VPWR VGND sg13g2_decap_8
XFILLER_43_326 VPWR VGND sg13g2_decap_8
XFILLER_34_11 VPWR VGND sg13g2_decap_8
XFILLER_24_551 VPWR VGND sg13g2_decap_8
XFILLER_12_746 VPWR VGND sg13g2_decap_8
XFILLER_34_77 VPWR VGND sg13g2_decap_8
XFILLER_11_256 VPWR VGND sg13g2_decap_8
XFILLER_8_739 VPWR VGND sg13g2_decap_8
XFILLER_7_238 VPWR VGND sg13g2_decap_8
XFILLER_3_466 VPWR VGND sg13g2_decap_8
XFILLER_19_312 VPWR VGND sg13g2_decap_8
XFILLER_47_665 VPWR VGND sg13g2_decap_8
XFILLER_46_175 VPWR VGND sg13g2_decap_8
XFILLER_19_389 VPWR VGND sg13g2_decap_8
XFILLER_35_849 VPWR VGND sg13g2_decap_8
XFILLER_43_893 VPWR VGND sg13g2_decap_8
XFILLER_30_576 VPWR VGND sg13g2_decap_8
XFILLER_27_0 VPWR VGND sg13g2_decap_8
XFILLER_29_109 VPWR VGND sg13g2_decap_8
XFILLER_38_621 VPWR VGND sg13g2_decap_8
XFILLER_1_70 VPWR VGND sg13g2_decap_8
X_29_ net1 net9 _00_ VPWR VGND sg13g2_and2_1
XFILLER_26_816 VPWR VGND sg13g2_decap_8
XFILLER_37_175 VPWR VGND sg13g2_decap_8
XFILLER_38_698 VPWR VGND sg13g2_decap_8
XFILLER_34_860 VPWR VGND sg13g2_decap_8
XFILLER_21_543 VPWR VGND sg13g2_decap_8
XFILLER_20_46 VPWR VGND sg13g2_decap_8
XFILLER_29_11 VPWR VGND sg13g2_decap_8
XFILLER_0_469 VPWR VGND sg13g2_decap_8
XFILLER_29_621 VPWR VGND sg13g2_decap_8
XFILLER_17_805 VPWR VGND sg13g2_decap_8
XFILLER_29_88 VPWR VGND sg13g2_decap_8
XFILLER_28_153 VPWR VGND sg13g2_decap_8
XFILLER_29_698 VPWR VGND sg13g2_decap_8
XFILLER_44_613 VPWR VGND sg13g2_decap_8
XFILLER_16_326 VPWR VGND sg13g2_decap_8
XFILLER_43_123 VPWR VGND sg13g2_decap_8
XFILLER_45_32 VPWR VGND sg13g2_decap_8
XFILLER_25_860 VPWR VGND sg13g2_decap_8
XFILLER_31_318 VPWR VGND sg13g2_decap_8
XFILLER_40_830 VPWR VGND sg13g2_decap_8
XFILLER_12_543 VPWR VGND sg13g2_decap_8
XFILLER_8_536 VPWR VGND sg13g2_decap_8
XFILLER_4_753 VPWR VGND sg13g2_decap_8
XFILLER_3_263 VPWR VGND sg13g2_decap_8
XFILLER_47_462 VPWR VGND sg13g2_decap_8
XFILLER_19_186 VPWR VGND sg13g2_decap_8
XFILLER_35_646 VPWR VGND sg13g2_decap_8
XFILLER_34_167 VPWR VGND sg13g2_decap_8
XFILLER_16_893 VPWR VGND sg13g2_decap_8
XFILLER_43_690 VPWR VGND sg13g2_decap_8
XFILLER_30_373 VPWR VGND sg13g2_decap_8
XFILLER_31_885 VPWR VGND sg13g2_decap_8
XFILLER_26_613 VPWR VGND sg13g2_decap_8
XFILLER_38_495 VPWR VGND sg13g2_decap_8
XFILLER_25_167 VPWR VGND sg13g2_decap_8
XFILLER_15_46 VPWR VGND sg13g2_decap_8
XFILLER_22_830 VPWR VGND sg13g2_decap_8
XFILLER_40_137 VPWR VGND sg13g2_decap_8
XFILLER_21_340 VPWR VGND sg13g2_decap_8
XFILLER_31_45 VPWR VGND sg13g2_fill_2
XFILLER_31_56 VPWR VGND sg13g2_fill_2
XFILLER_31_67 VPWR VGND sg13g2_decap_8
Xoutput23 net23 uo_out[6] VPWR VGND sg13g2_buf_1
XFILLER_1_756 VPWR VGND sg13g2_decap_8
XFILLER_49_749 VPWR VGND sg13g2_decap_8
XFILLER_0_266 VPWR VGND sg13g2_decap_8
XFILLER_48_259 VPWR VGND sg13g2_decap_8
XFILLER_45_900 VPWR VGND sg13g2_decap_8
XFILLER_17_602 VPWR VGND sg13g2_decap_8
XFILLER_16_123 VPWR VGND sg13g2_decap_8
XFILLER_29_495 VPWR VGND sg13g2_decap_8
XFILLER_44_410 VPWR VGND sg13g2_decap_8
XFILLER_17_679 VPWR VGND sg13g2_decap_8
XFILLER_31_104 VPWR VGND sg13g2_fill_2
XFILLER_32_627 VPWR VGND sg13g2_decap_8
XFILLER_44_487 VPWR VGND sg13g2_decap_8
XFILLER_13_830 VPWR VGND sg13g2_decap_8
XFILLER_9_823 VPWR VGND sg13g2_decap_8
XFILLER_12_340 VPWR VGND sg13g2_decap_8
XFILLER_8_333 VPWR VGND sg13g2_decap_8
XFILLER_4_550 VPWR VGND sg13g2_decap_8
XFILLER_39_259 VPWR VGND sg13g2_decap_8
XFILLER_36_900 VPWR VGND sg13g2_decap_8
XFILLER_35_443 VPWR VGND sg13g2_decap_8
XFILLER_23_627 VPWR VGND sg13g2_decap_8
XFILLER_16_690 VPWR VGND sg13g2_decap_8
XFILLER_22_137 VPWR VGND sg13g2_decap_8
XFILLER_30_170 VPWR VGND sg13g2_decap_8
XFILLER_31_682 VPWR VGND sg13g2_decap_8
XFILLER_7_91 VPWR VGND sg13g2_decap_8
XFILLER_45_207 VPWR VGND sg13g2_decap_8
XFILLER_26_410 VPWR VGND sg13g2_decap_8
XFILLER_38_292 VPWR VGND sg13g2_decap_8
XFILLER_14_627 VPWR VGND sg13g2_decap_8
XFILLER_26_487 VPWR VGND sg13g2_decap_8
XFILLER_13_137 VPWR VGND sg13g2_decap_8
XFILLER_41_457 VPWR VGND sg13g2_decap_8
XFILLER_42_11 VPWR VGND sg13g2_decap_8
XFILLER_10_844 VPWR VGND sg13g2_decap_8
XFILLER_6_837 VPWR VGND sg13g2_decap_8
XFILLER_42_99 VPWR VGND sg13g2_decap_8
XFILLER_5_347 VPWR VGND sg13g2_decap_8
XFILLER_1_553 VPWR VGND sg13g2_decap_8
XFILLER_49_546 VPWR VGND sg13g2_decap_8
XFILLER_18_900 VPWR VGND sg13g2_decap_8
XFILLER_36_207 VPWR VGND sg13g2_decap_8
XFILLER_29_292 VPWR VGND sg13g2_decap_8
XFILLER_17_476 VPWR VGND sg13g2_decap_8
XFILLER_32_424 VPWR VGND sg13g2_decap_8
XFILLER_45_774 VPWR VGND sg13g2_decap_8
XFILLER_44_284 VPWR VGND sg13g2_decap_8
XFILLER_9_620 VPWR VGND sg13g2_decap_8
XFILLER_8_130 VPWR VGND sg13g2_decap_8
XFILLER_9_697 VPWR VGND sg13g2_decap_8
XFILLER_35_240 VPWR VGND sg13g2_decap_8
XFILLER_36_774 VPWR VGND sg13g2_decap_8
XFILLER_23_424 VPWR VGND sg13g2_decap_8
XFILLER_12_25 VPWR VGND sg13g2_decap_8
XFILLER_18_207 VPWR VGND sg13g2_decap_8
XFILLER_27_763 VPWR VGND sg13g2_decap_8
XFILLER_37_77 VPWR VGND sg13g2_decap_8
XFILLER_15_914 VPWR VGND sg13g2_decap_8
XFILLER_42_722 VPWR VGND sg13g2_decap_8
XFILLER_14_424 VPWR VGND sg13g2_decap_8
XFILLER_26_284 VPWR VGND sg13g2_decap_8
XFILLER_41_254 VPWR VGND sg13g2_decap_8
XFILLER_42_799 VPWR VGND sg13g2_decap_8
XFILLER_10_641 VPWR VGND sg13g2_decap_8
XFILLER_6_634 VPWR VGND sg13g2_decap_8
XFILLER_5_144 VPWR VGND sg13g2_decap_8
XFILLER_2_851 VPWR VGND sg13g2_decap_8
XFILLER_1_350 VPWR VGND sg13g2_decap_8
XFILLER_49_343 VPWR VGND sg13g2_decap_8
X_62_ _24_ VPWR _27_ VGND _23_ _25_ sg13g2_o21ai_1
XFILLER_17_273 VPWR VGND sg13g2_decap_8
XFILLER_18_774 VPWR VGND sg13g2_decap_8
XFILLER_45_571 VPWR VGND sg13g2_decap_8
XFILLER_32_221 VPWR VGND sg13g2_decap_8
XFILLER_33_744 VPWR VGND sg13g2_decap_8
XFILLER_20_438 VPWR VGND sg13g2_decap_8
XFILLER_32_298 VPWR VGND sg13g2_decap_8
XFILLER_9_494 VPWR VGND sg13g2_decap_8
XFILLER_4_81 VPWR VGND sg13g2_decap_8
XFILLER_28_538 VPWR VGND sg13g2_decap_8
XFILLER_43_508 VPWR VGND sg13g2_decap_8
XFILLER_36_571 VPWR VGND sg13g2_decap_8
XFILLER_23_221 VPWR VGND sg13g2_decap_8
XFILLER_24_733 VPWR VGND sg13g2_decap_8
XFILLER_11_438 VPWR VGND sg13g2_decap_8
XFILLER_23_46 VPWR VGND sg13g2_decap_8
XFILLER_23_298 VPWR VGND sg13g2_decap_8
XFILLER_3_648 VPWR VGND sg13g2_decap_8
XFILLER_2_158 VPWR VGND sg13g2_decap_8
XFILLER_48_21 VPWR VGND sg13g2_decap_8
XFILLER_47_847 VPWR VGND sg13g2_decap_8
XFILLER_48_98 VPWR VGND sg13g2_decap_8
XFILLER_46_357 VPWR VGND sg13g2_decap_8
XFILLER_0_28 VPWR VGND sg13g2_decap_8
XFILLER_15_711 VPWR VGND sg13g2_decap_8
XFILLER_27_560 VPWR VGND sg13g2_decap_8
XFILLER_14_221 VPWR VGND sg13g2_decap_8
XFILLER_15_788 VPWR VGND sg13g2_decap_8
XFILLER_14_298 VPWR VGND sg13g2_decap_8
XFILLER_42_596 VPWR VGND sg13g2_decap_8
XFILLER_7_910 VPWR VGND sg13g2_decap_8
XFILLER_30_758 VPWR VGND sg13g2_decap_8
XFILLER_6_431 VPWR VGND sg13g2_decap_8
XFILLER_49_140 VPWR VGND sg13g2_decap_8
XFILLER_29_4 VPWR VGND sg13g2_decap_8
XFILLER_38_803 VPWR VGND sg13g2_decap_8
X_45_ _12_ VPWR _13_ VGND _03_ _11_ sg13g2_o21ai_1
XFILLER_37_357 VPWR VGND sg13g2_decap_8
XFILLER_18_571 VPWR VGND sg13g2_decap_8
XFILLER_33_541 VPWR VGND sg13g2_decap_8
XFILLER_21_725 VPWR VGND sg13g2_decap_8
XFILLER_20_235 VPWR VGND sg13g2_decap_8
XFILLER_9_291 VPWR VGND sg13g2_decap_8
XFILLER_29_803 VPWR VGND sg13g2_decap_8
XFILLER_18_46 VPWR VGND sg13g2_decap_8
XFILLER_28_335 VPWR VGND sg13g2_decap_8
XFILLER_16_508 VPWR VGND sg13g2_decap_8
XFILLER_43_305 VPWR VGND sg13g2_decap_8
XFILLER_24_530 VPWR VGND sg13g2_decap_8
XFILLER_12_725 VPWR VGND sg13g2_decap_8
XFILLER_34_56 VPWR VGND sg13g2_decap_8
XFILLER_11_235 VPWR VGND sg13g2_decap_8
XFILLER_8_718 VPWR VGND sg13g2_decap_8
XFILLER_7_217 VPWR VGND sg13g2_decap_8
XFILLER_3_445 VPWR VGND sg13g2_decap_8
XFILLER_47_644 VPWR VGND sg13g2_decap_8
XFILLER_46_154 VPWR VGND sg13g2_decap_8
XFILLER_19_368 VPWR VGND sg13g2_decap_8
XFILLER_35_828 VPWR VGND sg13g2_decap_8
XFILLER_34_349 VPWR VGND sg13g2_decap_8
XFILLER_43_872 VPWR VGND sg13g2_decap_8
XFILLER_15_585 VPWR VGND sg13g2_decap_8
XFILLER_30_555 VPWR VGND sg13g2_decap_8
XFILLER_42_393 VPWR VGND sg13g2_decap_8
XFILLER_7_784 VPWR VGND sg13g2_decap_8
XFILLER_38_600 VPWR VGND sg13g2_decap_8
XFILLER_37_154 VPWR VGND sg13g2_decap_8
XFILLER_38_677 VPWR VGND sg13g2_decap_8
XFILLER_25_349 VPWR VGND sg13g2_decap_8
XFILLER_21_522 VPWR VGND sg13g2_decap_8
XFILLER_40_319 VPWR VGND sg13g2_decap_8
XFILLER_21_599 VPWR VGND sg13g2_decap_8
XFILLER_20_25 VPWR VGND sg13g2_decap_8
XFILLER_0_448 VPWR VGND sg13g2_decap_8
XFILLER_29_67 VPWR VGND sg13g2_decap_8
XFILLER_29_600 VPWR VGND sg13g2_decap_8
XFILLER_28_132 VPWR VGND sg13g2_decap_8
XFILLER_16_305 VPWR VGND sg13g2_decap_8
XFILLER_29_677 VPWR VGND sg13g2_decap_8
XFILLER_45_11 VPWR VGND sg13g2_decap_8
XFILLER_43_102 VPWR VGND sg13g2_decap_8
XFILLER_32_809 VPWR VGND sg13g2_decap_8
XFILLER_44_669 VPWR VGND sg13g2_decap_8
XFILLER_45_88 VPWR VGND sg13g2_decap_8
XFILLER_43_179 VPWR VGND sg13g2_decap_8
XFILLER_12_522 VPWR VGND sg13g2_decap_8
XFILLER_8_515 VPWR VGND sg13g2_decap_8
XFILLER_40_886 VPWR VGND sg13g2_decap_8
XFILLER_12_599 VPWR VGND sg13g2_decap_8
XFILLER_4_732 VPWR VGND sg13g2_decap_8
XFILLER_3_242 VPWR VGND sg13g2_decap_8
XFILLER_47_441 VPWR VGND sg13g2_decap_8
XFILLER_19_165 VPWR VGND sg13g2_decap_8
XFILLER_35_625 VPWR VGND sg13g2_decap_8
XFILLER_23_809 VPWR VGND sg13g2_decap_8
XFILLER_34_146 VPWR VGND sg13g2_decap_8
XFILLER_16_872 VPWR VGND sg13g2_decap_8
XFILLER_22_319 VPWR VGND sg13g2_decap_8
XFILLER_15_382 VPWR VGND sg13g2_decap_8
XFILLER_31_864 VPWR VGND sg13g2_decap_8
XFILLER_42_190 VPWR VGND sg13g2_decap_8
XFILLER_30_352 VPWR VGND sg13g2_decap_8
XFILLER_7_581 VPWR VGND sg13g2_decap_8
XFILLER_38_474 VPWR VGND sg13g2_decap_8
XFILLER_14_809 VPWR VGND sg13g2_decap_8
XFILLER_25_146 VPWR VGND sg13g2_decap_8
XFILLER_26_669 VPWR VGND sg13g2_decap_8
XFILLER_13_319 VPWR VGND sg13g2_decap_8
XFILLER_15_25 VPWR VGND sg13g2_decap_8
XFILLER_40_116 VPWR VGND sg13g2_decap_8
XFILLER_41_639 VPWR VGND sg13g2_decap_8
XFILLER_22_886 VPWR VGND sg13g2_decap_8
XFILLER_21_396 VPWR VGND sg13g2_decap_8
XFILLER_5_529 VPWR VGND sg13g2_decap_8
Xoutput24 net24 uo_out[7] VPWR VGND sg13g2_buf_1
XFILLER_1_735 VPWR VGND sg13g2_decap_8
XFILLER_0_245 VPWR VGND sg13g2_decap_8
XFILLER_49_728 VPWR VGND sg13g2_decap_8
XFILLER_48_238 VPWR VGND sg13g2_decap_8
XFILLER_16_102 VPWR VGND sg13g2_decap_8
XFILLER_29_474 VPWR VGND sg13g2_decap_8
XFILLER_17_658 VPWR VGND sg13g2_decap_8
XFILLER_32_606 VPWR VGND sg13g2_decap_8
XFILLER_44_466 VPWR VGND sg13g2_decap_8
XFILLER_16_179 VPWR VGND sg13g2_decap_8
XFILLER_9_802 VPWR VGND sg13g2_decap_8
XFILLER_8_312 VPWR VGND sg13g2_decap_8
XFILLER_13_886 VPWR VGND sg13g2_decap_8
XFILLER_12_396 VPWR VGND sg13g2_decap_8
XFILLER_40_683 VPWR VGND sg13g2_decap_8
XFILLER_9_879 VPWR VGND sg13g2_decap_8
XFILLER_8_389 VPWR VGND sg13g2_decap_8
XFILLER_39_238 VPWR VGND sg13g2_decap_8
XFILLER_11_4 VPWR VGND sg13g2_decap_8
XFILLER_35_422 VPWR VGND sg13g2_decap_8
XFILLER_23_606 VPWR VGND sg13g2_decap_8
XFILLER_22_116 VPWR VGND sg13g2_decap_8
XFILLER_35_499 VPWR VGND sg13g2_decap_8
XFILLER_31_661 VPWR VGND sg13g2_decap_8
XFILLER_7_70 VPWR VGND sg13g2_decap_8
XFILLER_38_271 VPWR VGND sg13g2_decap_8
XFILLER_42_904 VPWR VGND sg13g2_decap_8
XFILLER_14_606 VPWR VGND sg13g2_decap_8
XFILLER_26_68 VPWR VGND sg13g2_decap_8
XFILLER_26_79 VPWR VGND sg13g2_fill_1
XFILLER_26_466 VPWR VGND sg13g2_decap_8
XFILLER_13_116 VPWR VGND sg13g2_decap_8
XFILLER_41_436 VPWR VGND sg13g2_decap_8
XFILLER_9_109 VPWR VGND sg13g2_decap_8
XFILLER_42_34 VPWR VGND sg13g2_fill_1
XFILLER_10_823 VPWR VGND sg13g2_decap_8
XFILLER_22_683 VPWR VGND sg13g2_decap_8
XFILLER_42_78 VPWR VGND sg13g2_decap_8
XFILLER_6_816 VPWR VGND sg13g2_decap_8
XFILLER_21_193 VPWR VGND sg13g2_decap_8
XFILLER_5_326 VPWR VGND sg13g2_decap_8
XFILLER_1_532 VPWR VGND sg13g2_decap_8
XFILLER_3_39 VPWR VGND sg13g2_decap_8
XFILLER_49_525 VPWR VGND sg13g2_decap_8
XFILLER_29_271 VPWR VGND sg13g2_decap_8
XFILLER_17_455 VPWR VGND sg13g2_decap_8
XFILLER_45_753 VPWR VGND sg13g2_decap_8
XFILLER_32_403 VPWR VGND sg13g2_decap_8
XFILLER_44_263 VPWR VGND sg13g2_decap_8
XFILLER_13_683 VPWR VGND sg13g2_decap_8
XFILLER_40_480 VPWR VGND sg13g2_decap_8
XFILLER_9_676 VPWR VGND sg13g2_decap_8
XFILLER_12_193 VPWR VGND sg13g2_decap_8
XFILLER_8_186 VPWR VGND sg13g2_decap_8
XFILLER_5_893 VPWR VGND sg13g2_decap_8
XFILLER_36_753 VPWR VGND sg13g2_decap_8
XFILLER_23_403 VPWR VGND sg13g2_decap_8
XFILLER_24_915 VPWR VGND sg13g2_decap_8
XFILLER_35_296 VPWR VGND sg13g2_decap_8
XFILLER_46_539 VPWR VGND sg13g2_decap_8
XFILLER_37_56 VPWR VGND sg13g2_decap_8
XFILLER_27_742 VPWR VGND sg13g2_decap_8
XFILLER_14_403 VPWR VGND sg13g2_decap_8
XFILLER_26_263 VPWR VGND sg13g2_decap_8
XFILLER_42_701 VPWR VGND sg13g2_decap_8
XFILLER_41_233 VPWR VGND sg13g2_decap_8
XFILLER_42_778 VPWR VGND sg13g2_decap_8
XFILLER_10_620 VPWR VGND sg13g2_decap_8
XFILLER_22_480 VPWR VGND sg13g2_decap_8
XFILLER_6_613 VPWR VGND sg13g2_decap_8
XFILLER_10_697 VPWR VGND sg13g2_decap_8
XFILLER_5_123 VPWR VGND sg13g2_decap_8
XFILLER_2_830 VPWR VGND sg13g2_decap_8
XFILLER_49_322 VPWR VGND sg13g2_decap_8
X_61_ net23 _23_ _26_ VPWR VGND sg13g2_xnor2_1
XFILLER_49_399 VPWR VGND sg13g2_decap_8
XFILLER_37_539 VPWR VGND sg13g2_decap_8
XFILLER_18_753 VPWR VGND sg13g2_decap_8
XFILLER_17_252 VPWR VGND sg13g2_decap_8
XFILLER_45_550 VPWR VGND sg13g2_decap_8
XFILLER_32_200 VPWR VGND sg13g2_decap_8
XFILLER_33_723 VPWR VGND sg13g2_decap_8
XFILLER_21_907 VPWR VGND sg13g2_decap_8
XFILLER_20_417 VPWR VGND sg13g2_decap_8
XFILLER_32_277 VPWR VGND sg13g2_decap_8
XFILLER_13_480 VPWR VGND sg13g2_decap_8
XFILLER_9_473 VPWR VGND sg13g2_decap_8
XFILLER_5_690 VPWR VGND sg13g2_decap_8
XFILLER_4_60 VPWR VGND sg13g2_decap_8
XFILLER_28_517 VPWR VGND sg13g2_decap_8
XFILLER_24_712 VPWR VGND sg13g2_decap_8
XFILLER_36_550 VPWR VGND sg13g2_decap_8
XFILLER_23_200 VPWR VGND sg13g2_decap_8
XFILLER_12_907 VPWR VGND sg13g2_decap_8
XFILLER_24_789 VPWR VGND sg13g2_decap_8
XFILLER_11_417 VPWR VGND sg13g2_decap_8
XFILLER_23_25 VPWR VGND sg13g2_decap_8
XFILLER_23_277 VPWR VGND sg13g2_decap_8
XFILLER_3_627 VPWR VGND sg13g2_decap_8
XFILLER_2_137 VPWR VGND sg13g2_decap_8
XFILLER_47_826 VPWR VGND sg13g2_decap_8
XFILLER_48_77 VPWR VGND sg13g2_decap_8
XFILLER_46_336 VPWR VGND sg13g2_decap_8
XFILLER_14_200 VPWR VGND sg13g2_decap_8
XFILLER_15_767 VPWR VGND sg13g2_decap_8
XFILLER_14_277 VPWR VGND sg13g2_decap_8
XFILLER_30_737 VPWR VGND sg13g2_decap_8
XFILLER_42_575 VPWR VGND sg13g2_decap_8
XFILLER_6_410 VPWR VGND sg13g2_decap_8
XFILLER_10_494 VPWR VGND sg13g2_decap_8
XFILLER_6_487 VPWR VGND sg13g2_decap_8
XFILLER_49_196 VPWR VGND sg13g2_decap_8
X_44_ VGND VPWR _04_ _07_ _12_ _08_ sg13g2_a21oi_1
XFILLER_37_336 VPWR VGND sg13g2_decap_8
XFILLER_38_859 VPWR VGND sg13g2_decap_8
XFILLER_18_550 VPWR VGND sg13g2_decap_8
XFILLER_33_520 VPWR VGND sg13g2_decap_8
XFILLER_21_704 VPWR VGND sg13g2_decap_8
XFILLER_20_214 VPWR VGND sg13g2_decap_8
XFILLER_33_597 VPWR VGND sg13g2_decap_8
XFILLER_9_270 VPWR VGND sg13g2_decap_8
XFILLER_18_25 VPWR VGND sg13g2_decap_8
XFILLER_28_314 VPWR VGND sg13g2_decap_8
XFILLER_29_859 VPWR VGND sg13g2_decap_8
XFILLER_12_704 VPWR VGND sg13g2_decap_8
XFILLER_11_214 VPWR VGND sg13g2_decap_8
XFILLER_24_586 VPWR VGND sg13g2_decap_8
XFILLER_20_781 VPWR VGND sg13g2_decap_8
XFILLER_4_914 VPWR VGND sg13g2_decap_8
XFILLER_3_424 VPWR VGND sg13g2_decap_8
XFILLER_47_623 VPWR VGND sg13g2_decap_8
XFILLER_46_133 VPWR VGND sg13g2_decap_8
XFILLER_19_347 VPWR VGND sg13g2_decap_8
XFILLER_35_807 VPWR VGND sg13g2_decap_8
XFILLER_28_881 VPWR VGND sg13g2_decap_8
XFILLER_34_328 VPWR VGND sg13g2_decap_8
XFILLER_43_851 VPWR VGND sg13g2_decap_8
XFILLER_15_564 VPWR VGND sg13g2_decap_8
XFILLER_42_372 VPWR VGND sg13g2_decap_8
XFILLER_30_534 VPWR VGND sg13g2_decap_8
XFILLER_11_781 VPWR VGND sg13g2_decap_8
XFILLER_10_291 VPWR VGND sg13g2_decap_8
XFILLER_7_763 VPWR VGND sg13g2_decap_8
XFILLER_6_284 VPWR VGND sg13g2_decap_8
XFILLER_41_4 VPWR VGND sg13g2_decap_8
XFILLER_37_133 VPWR VGND sg13g2_decap_8
XFILLER_38_656 VPWR VGND sg13g2_decap_8
XFILLER_25_328 VPWR VGND sg13g2_decap_8
XFILLER_21_501 VPWR VGND sg13g2_decap_8
XFILLER_34_895 VPWR VGND sg13g2_decap_8
XFILLER_33_394 VPWR VGND sg13g2_decap_8
XFILLER_21_578 VPWR VGND sg13g2_decap_8
XFILLER_1_917 VPWR VGND sg13g2_decap_8
XFILLER_0_427 VPWR VGND sg13g2_decap_8
XFILLER_29_46 VPWR VGND sg13g2_decap_8
XFILLER_29_656 VPWR VGND sg13g2_decap_8
XFILLER_28_188 VPWR VGND sg13g2_decap_8
XFILLER_44_648 VPWR VGND sg13g2_decap_8
XFILLER_43_158 VPWR VGND sg13g2_decap_8
XFILLER_45_67 VPWR VGND sg13g2_decap_8
XFILLER_12_501 VPWR VGND sg13g2_decap_8
XFILLER_25_895 VPWR VGND sg13g2_decap_8
XFILLER_24_383 VPWR VGND sg13g2_decap_8
XFILLER_12_578 VPWR VGND sg13g2_decap_8
XFILLER_40_865 VPWR VGND sg13g2_decap_8
XFILLER_6_39 VPWR VGND sg13g2_decap_8
XFILLER_4_711 VPWR VGND sg13g2_decap_8
XFILLER_3_221 VPWR VGND sg13g2_decap_8
XFILLER_10_81 VPWR VGND sg13g2_decap_8
XFILLER_4_788 VPWR VGND sg13g2_decap_8
XFILLER_3_298 VPWR VGND sg13g2_decap_8
XFILLER_48_910 VPWR VGND sg13g2_decap_8
XFILLER_47_420 VPWR VGND sg13g2_decap_8
XFILLER_19_144 VPWR VGND sg13g2_decap_8
XFILLER_35_604 VPWR VGND sg13g2_decap_8
XFILLER_47_497 VPWR VGND sg13g2_decap_8
XFILLER_16_851 VPWR VGND sg13g2_decap_8
XFILLER_34_125 VPWR VGND sg13g2_decap_8
XFILLER_15_361 VPWR VGND sg13g2_decap_8
XFILLER_30_331 VPWR VGND sg13g2_decap_8
XFILLER_31_843 VPWR VGND sg13g2_decap_8
XFILLER_7_560 VPWR VGND sg13g2_decap_8
XFILLER_39_910 VPWR VGND sg13g2_decap_8
XFILLER_38_453 VPWR VGND sg13g2_decap_8
XFILLER_26_648 VPWR VGND sg13g2_decap_8
XFILLER_25_125 VPWR VGND sg13g2_decap_8
XFILLER_41_618 VPWR VGND sg13g2_decap_8
XFILLER_34_692 VPWR VGND sg13g2_decap_8
XFILLER_22_865 VPWR VGND sg13g2_decap_8
XFILLER_33_191 VPWR VGND sg13g2_decap_8
XFILLER_21_375 VPWR VGND sg13g2_decap_8
XFILLER_31_25 VPWR VGND sg13g2_decap_8
XFILLER_5_508 VPWR VGND sg13g2_decap_8
XFILLER_31_47 VPWR VGND sg13g2_fill_1
XFILLER_31_58 VPWR VGND sg13g2_fill_1
XFILLER_1_714 VPWR VGND sg13g2_decap_8
XFILLER_49_707 VPWR VGND sg13g2_decap_8
XFILLER_0_224 VPWR VGND sg13g2_decap_8
XFILLER_48_217 VPWR VGND sg13g2_decap_8
XFILLER_29_453 VPWR VGND sg13g2_decap_8
XFILLER_17_637 VPWR VGND sg13g2_decap_8
XFILLER_44_445 VPWR VGND sg13g2_decap_8
XFILLER_16_158 VPWR VGND sg13g2_decap_8
XFILLER_24_180 VPWR VGND sg13g2_decap_8
XFILLER_25_692 VPWR VGND sg13g2_decap_8
XFILLER_13_865 VPWR VGND sg13g2_decap_8
XFILLER_40_662 VPWR VGND sg13g2_decap_8
XFILLER_9_858 VPWR VGND sg13g2_decap_8
XFILLER_12_375 VPWR VGND sg13g2_decap_8
XFILLER_8_368 VPWR VGND sg13g2_decap_8
XFILLER_4_585 VPWR VGND sg13g2_decap_8
XFILLER_0_791 VPWR VGND sg13g2_decap_8
XFILLER_39_217 VPWR VGND sg13g2_decap_8
XFILLER_48_784 VPWR VGND sg13g2_decap_8
XFILLER_35_401 VPWR VGND sg13g2_decap_8
XFILLER_47_294 VPWR VGND sg13g2_decap_8
XFILLER_35_478 VPWR VGND sg13g2_decap_8
XFILLER_31_640 VPWR VGND sg13g2_decap_8
XFILLER_27_924 VPWR VGND sg13g2_fill_1
XFILLER_38_250 VPWR VGND sg13g2_decap_8
XFILLER_39_784 VPWR VGND sg13g2_decap_8
XFILLER_26_25 VPWR VGND sg13g2_fill_2
XFILLER_26_47 VPWR VGND sg13g2_decap_8
XFILLER_26_445 VPWR VGND sg13g2_decap_8
XFILLER_41_415 VPWR VGND sg13g2_decap_8
XFILLER_10_802 VPWR VGND sg13g2_decap_8
XFILLER_22_662 VPWR VGND sg13g2_decap_8
XFILLER_21_172 VPWR VGND sg13g2_decap_8
XFILLER_42_57 VPWR VGND sg13g2_decap_8
XFILLER_10_879 VPWR VGND sg13g2_decap_8
XFILLER_5_305 VPWR VGND sg13g2_decap_8
XFILLER_1_511 VPWR VGND sg13g2_decap_8
XFILLER_3_18 VPWR VGND sg13g2_decap_8
XFILLER_49_504 VPWR VGND sg13g2_decap_8
XFILLER_1_588 VPWR VGND sg13g2_decap_8
XFILLER_29_250 VPWR VGND sg13g2_decap_8
XFILLER_17_434 VPWR VGND sg13g2_decap_8
XFILLER_33_905 VPWR VGND sg13g2_decap_8
XFILLER_45_732 VPWR VGND sg13g2_decap_8
XFILLER_44_242 VPWR VGND sg13g2_decap_8
XFILLER_13_662 VPWR VGND sg13g2_decap_8
XFILLER_32_459 VPWR VGND sg13g2_decap_8
XFILLER_12_172 VPWR VGND sg13g2_decap_8
XFILLER_9_655 VPWR VGND sg13g2_decap_8
XFILLER_8_165 VPWR VGND sg13g2_decap_8
XFILLER_5_872 VPWR VGND sg13g2_decap_8
XFILLER_4_382 VPWR VGND sg13g2_decap_8
XFILLER_48_581 VPWR VGND sg13g2_decap_8
XFILLER_36_732 VPWR VGND sg13g2_decap_8
XFILLER_35_275 VPWR VGND sg13g2_decap_8
XFILLER_23_459 VPWR VGND sg13g2_decap_8
XFILLER_10_109 VPWR VGND sg13g2_decap_8
XFILLER_3_809 VPWR VGND sg13g2_decap_8
XFILLER_2_319 VPWR VGND sg13g2_decap_8
XFILLER_46_518 VPWR VGND sg13g2_decap_8
XFILLER_27_721 VPWR VGND sg13g2_decap_8
XFILLER_37_35 VPWR VGND sg13g2_decap_8
XFILLER_39_581 VPWR VGND sg13g2_decap_8
XFILLER_26_242 VPWR VGND sg13g2_decap_8
XFILLER_27_798 VPWR VGND sg13g2_decap_8
XFILLER_41_212 VPWR VGND sg13g2_decap_8
XFILLER_14_459 VPWR VGND sg13g2_decap_8
XFILLER_30_919 VPWR VGND sg13g2_decap_4
XFILLER_42_757 VPWR VGND sg13g2_decap_8
XFILLER_41_289 VPWR VGND sg13g2_decap_8
XFILLER_10_676 VPWR VGND sg13g2_decap_8
XFILLER_5_102 VPWR VGND sg13g2_decap_8
XFILLER_6_669 VPWR VGND sg13g2_decap_8
XFILLER_5_179 VPWR VGND sg13g2_decap_8
XFILLER_49_301 VPWR VGND sg13g2_decap_8
XFILLER_2_886 VPWR VGND sg13g2_decap_8
XFILLER_1_385 VPWR VGND sg13g2_decap_8
X_60_ net15 net7 _26_ VPWR VGND sg13g2_xor2_1
XFILLER_49_378 VPWR VGND sg13g2_decap_8
XFILLER_37_518 VPWR VGND sg13g2_decap_8
XFILLER_18_732 VPWR VGND sg13g2_decap_8
XFILLER_17_231 VPWR VGND sg13g2_decap_8
XFILLER_33_702 VPWR VGND sg13g2_decap_8
XFILLER_32_256 VPWR VGND sg13g2_decap_8
XFILLER_33_779 VPWR VGND sg13g2_decap_8
XFILLER_9_452 VPWR VGND sg13g2_decap_8
XFILLER_23_256 VPWR VGND sg13g2_decap_8
XFILLER_24_768 VPWR VGND sg13g2_decap_8
XFILLER_3_606 VPWR VGND sg13g2_decap_8
XFILLER_2_116 VPWR VGND sg13g2_decap_8
XFILLER_47_805 VPWR VGND sg13g2_decap_8
XFILLER_48_56 VPWR VGND sg13g2_decap_8
XFILLER_46_315 VPWR VGND sg13g2_decap_8
XFILLER_19_529 VPWR VGND sg13g2_decap_8
XFILLER_15_746 VPWR VGND sg13g2_decap_8
XFILLER_27_595 VPWR VGND sg13g2_decap_8
XFILLER_14_256 VPWR VGND sg13g2_decap_8
XFILLER_42_554 VPWR VGND sg13g2_decap_8
XFILLER_9_39 VPWR VGND sg13g2_decap_8
XFILLER_30_716 VPWR VGND sg13g2_decap_8
XFILLER_10_473 VPWR VGND sg13g2_decap_8
XFILLER_13_81 VPWR VGND sg13g2_decap_8
XFILLER_6_466 VPWR VGND sg13g2_decap_8
XFILLER_2_683 VPWR VGND sg13g2_decap_8
XFILLER_1_182 VPWR VGND sg13g2_decap_8
XFILLER_49_175 VPWR VGND sg13g2_decap_8
X_43_ _11_ _09_ _05_ VPWR VGND sg13g2_nand2b_1
XFILLER_37_315 VPWR VGND sg13g2_decap_8
XFILLER_38_838 VPWR VGND sg13g2_decap_8
XFILLER_46_882 VPWR VGND sg13g2_decap_8
XFILLER_33_576 VPWR VGND sg13g2_decap_8
XFILLER_0_609 VPWR VGND sg13g2_decap_8
XFILLER_29_838 VPWR VGND sg13g2_decap_8
XFILLER_37_882 VPWR VGND sg13g2_decap_8
XFILLER_34_25 VPWR VGND sg13g2_decap_4
XFILLER_24_565 VPWR VGND sg13g2_decap_8
XFILLER_20_760 VPWR VGND sg13g2_decap_8
XFILLER_3_403 VPWR VGND sg13g2_decap_8
XFILLER_47_602 VPWR VGND sg13g2_decap_8
XFILLER_46_112 VPWR VGND sg13g2_decap_8
XFILLER_19_326 VPWR VGND sg13g2_decap_8
XFILLER_47_679 VPWR VGND sg13g2_decap_8
XFILLER_28_860 VPWR VGND sg13g2_decap_8
XFILLER_34_307 VPWR VGND sg13g2_decap_8
XFILLER_46_189 VPWR VGND sg13g2_decap_8
XFILLER_43_830 VPWR VGND sg13g2_decap_8
XFILLER_15_543 VPWR VGND sg13g2_decap_8
XFILLER_27_392 VPWR VGND sg13g2_decap_8
XFILLER_30_513 VPWR VGND sg13g2_decap_8
XFILLER_42_351 VPWR VGND sg13g2_decap_8
XFILLER_11_760 VPWR VGND sg13g2_decap_8
XFILLER_10_270 VPWR VGND sg13g2_decap_8
XFILLER_7_742 VPWR VGND sg13g2_decap_8
XFILLER_6_263 VPWR VGND sg13g2_decap_8
XFILLER_34_4 VPWR VGND sg13g2_decap_8
XFILLER_2_480 VPWR VGND sg13g2_decap_8
XFILLER_37_112 VPWR VGND sg13g2_decap_8
XFILLER_38_635 VPWR VGND sg13g2_decap_8
XFILLER_25_307 VPWR VGND sg13g2_decap_8
XFILLER_1_84 VPWR VGND sg13g2_decap_8
XFILLER_19_893 VPWR VGND sg13g2_decap_8
XFILLER_37_189 VPWR VGND sg13g2_decap_8
XFILLER_33_373 VPWR VGND sg13g2_decap_8
XFILLER_34_874 VPWR VGND sg13g2_decap_8
XFILLER_21_557 VPWR VGND sg13g2_decap_8
XFILLER_0_406 VPWR VGND sg13g2_decap_8
XFILLER_29_25 VPWR VGND sg13g2_decap_8
XFILLER_29_635 VPWR VGND sg13g2_decap_8
XFILLER_17_819 VPWR VGND sg13g2_decap_8
XFILLER_28_167 VPWR VGND sg13g2_decap_8
XFILLER_44_627 VPWR VGND sg13g2_decap_8
XFILLER_45_46 VPWR VGND sg13g2_decap_8
XFILLER_43_137 VPWR VGND sg13g2_decap_8
XFILLER_24_362 VPWR VGND sg13g2_decap_8
XFILLER_25_874 VPWR VGND sg13g2_decap_8
XFILLER_40_844 VPWR VGND sg13g2_decap_8
XFILLER_12_557 VPWR VGND sg13g2_decap_8
XFILLER_6_18 VPWR VGND sg13g2_decap_8
XFILLER_3_200 VPWR VGND sg13g2_decap_8
XFILLER_4_767 VPWR VGND sg13g2_decap_8
XFILLER_10_60 VPWR VGND sg13g2_decap_8
XFILLER_3_277 VPWR VGND sg13g2_decap_8
XFILLER_19_123 VPWR VGND sg13g2_decap_8
XFILLER_47_476 VPWR VGND sg13g2_decap_8
XFILLER_16_830 VPWR VGND sg13g2_decap_8
XFILLER_15_340 VPWR VGND sg13g2_decap_8
XFILLER_30_310 VPWR VGND sg13g2_decap_8
XFILLER_31_822 VPWR VGND sg13g2_decap_8
XFILLER_30_387 VPWR VGND sg13g2_decap_8
XFILLER_31_899 VPWR VGND sg13g2_decap_8
XFILLER_38_432 VPWR VGND sg13g2_decap_8
XFILLER_25_104 VPWR VGND sg13g2_decap_8
XFILLER_26_627 VPWR VGND sg13g2_decap_8
XFILLER_19_690 VPWR VGND sg13g2_decap_8
XFILLER_34_671 VPWR VGND sg13g2_decap_8
XFILLER_22_844 VPWR VGND sg13g2_decap_8
XFILLER_33_170 VPWR VGND sg13g2_decap_8
XFILLER_21_354 VPWR VGND sg13g2_decap_8
XFILLER_0_203 VPWR VGND sg13g2_decap_8
XFILLER_29_432 VPWR VGND sg13g2_decap_8
XFILLER_45_914 VPWR VGND sg13g2_decap_8
XFILLER_17_616 VPWR VGND sg13g2_decap_8
XFILLER_16_137 VPWR VGND sg13g2_decap_8
XFILLER_44_424 VPWR VGND sg13g2_decap_8
XFILLER_25_671 VPWR VGND sg13g2_decap_8
XFILLER_13_844 VPWR VGND sg13g2_decap_8
XFILLER_31_129 VPWR VGND sg13g2_decap_8
XFILLER_12_354 VPWR VGND sg13g2_decap_8
XFILLER_40_641 VPWR VGND sg13g2_decap_8
XFILLER_9_837 VPWR VGND sg13g2_decap_8
XFILLER_8_347 VPWR VGND sg13g2_decap_8
XFILLER_21_81 VPWR VGND sg13g2_decap_8
XFILLER_4_564 VPWR VGND sg13g2_decap_8
XFILLER_0_770 VPWR VGND sg13g2_decap_8
XFILLER_48_763 VPWR VGND sg13g2_decap_8
XFILLER_47_273 VPWR VGND sg13g2_decap_8
XFILLER_36_914 VPWR VGND sg13g2_decap_8
XFILLER_35_457 VPWR VGND sg13g2_decap_8
XFILLER_31_696 VPWR VGND sg13g2_decap_8
XFILLER_30_184 VPWR VGND sg13g2_decap_8
XFILLER_27_903 VPWR VGND sg13g2_decap_8
XFILLER_39_763 VPWR VGND sg13g2_decap_8
XFILLER_26_424 VPWR VGND sg13g2_decap_8
XFILLER_22_641 VPWR VGND sg13g2_decap_8
XFILLER_42_25 VPWR VGND sg13g2_decap_8
XFILLER_21_151 VPWR VGND sg13g2_decap_8
XFILLER_10_858 VPWR VGND sg13g2_decap_8
XFILLER_1_567 VPWR VGND sg13g2_decap_8
XFILLER_17_413 VPWR VGND sg13g2_decap_8
XFILLER_18_914 VPWR VGND sg13g2_decap_8
XFILLER_45_711 VPWR VGND sg13g2_decap_8
XFILLER_44_221 VPWR VGND sg13g2_decap_8
XFILLER_45_788 VPWR VGND sg13g2_decap_8
XFILLER_32_438 VPWR VGND sg13g2_decap_8
XFILLER_44_298 VPWR VGND sg13g2_decap_8
XFILLER_13_641 VPWR VGND sg13g2_decap_8
XFILLER_16_81 VPWR VGND sg13g2_decap_8
XFILLER_9_634 VPWR VGND sg13g2_decap_8
XFILLER_12_151 VPWR VGND sg13g2_decap_8
XFILLER_8_144 VPWR VGND sg13g2_decap_8
XFILLER_5_851 VPWR VGND sg13g2_decap_8
XFILLER_4_361 VPWR VGND sg13g2_decap_8
XFILLER_48_560 VPWR VGND sg13g2_decap_8
XFILLER_36_711 VPWR VGND sg13g2_decap_8
XFILLER_35_254 VPWR VGND sg13g2_decap_8
XFILLER_36_788 VPWR VGND sg13g2_decap_8
XFILLER_23_438 VPWR VGND sg13g2_decap_8
XFILLER_31_493 VPWR VGND sg13g2_decap_8
XFILLER_12_39 VPWR VGND sg13g2_decap_8
XFILLER_37_14 VPWR VGND sg13g2_decap_8
XFILLER_27_700 VPWR VGND sg13g2_decap_8
XFILLER_39_560 VPWR VGND sg13g2_decap_8
XFILLER_26_221 VPWR VGND sg13g2_decap_8
XFILLER_27_777 VPWR VGND sg13g2_decap_8
XFILLER_14_438 VPWR VGND sg13g2_decap_8
XFILLER_26_298 VPWR VGND sg13g2_decap_8
XFILLER_42_736 VPWR VGND sg13g2_decap_8
XFILLER_41_268 VPWR VGND sg13g2_decap_8
XFILLER_10_655 VPWR VGND sg13g2_decap_8
XFILLER_6_648 VPWR VGND sg13g2_decap_8
XFILLER_5_158 VPWR VGND sg13g2_decap_8
XFILLER_2_865 VPWR VGND sg13g2_decap_8
XFILLER_1_364 VPWR VGND sg13g2_decap_8
XFILLER_49_357 VPWR VGND sg13g2_decap_8
XFILLER_18_711 VPWR VGND sg13g2_decap_8
XFILLER_17_210 VPWR VGND sg13g2_decap_8
XFILLER_18_788 VPWR VGND sg13g2_decap_8
XFILLER_17_287 VPWR VGND sg13g2_decap_8
XFILLER_27_91 VPWR VGND sg13g2_decap_8
XFILLER_45_585 VPWR VGND sg13g2_decap_8
XFILLER_32_235 VPWR VGND sg13g2_decap_8
XFILLER_33_758 VPWR VGND sg13g2_decap_8
XFILLER_9_431 VPWR VGND sg13g2_decap_8
XFILLER_4_95 VPWR VGND sg13g2_decap_8
XFILLER_36_585 VPWR VGND sg13g2_decap_8
XFILLER_23_235 VPWR VGND sg13g2_decap_8
XFILLER_24_747 VPWR VGND sg13g2_decap_8
XFILLER_31_290 VPWR VGND sg13g2_decap_8
XFILLER_48_35 VPWR VGND sg13g2_decap_8
XFILLER_19_508 VPWR VGND sg13g2_decap_8
XFILLER_15_725 VPWR VGND sg13g2_decap_8
XFILLER_27_574 VPWR VGND sg13g2_decap_8
XFILLER_9_18 VPWR VGND sg13g2_decap_8
XFILLER_14_235 VPWR VGND sg13g2_decap_8
XFILLER_42_533 VPWR VGND sg13g2_decap_8
XFILLER_10_452 VPWR VGND sg13g2_decap_8
XFILLER_7_924 VPWR VGND sg13g2_fill_1
XFILLER_13_60 VPWR VGND sg13g2_decap_8
XFILLER_6_445 VPWR VGND sg13g2_decap_8
XFILLER_1_161 VPWR VGND sg13g2_decap_8
XFILLER_2_662 VPWR VGND sg13g2_decap_8
XFILLER_49_154 VPWR VGND sg13g2_decap_8
X_42_ net20 _09_ _10_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_817 VPWR VGND sg13g2_decap_8
XFILLER_46_861 VPWR VGND sg13g2_decap_8
XFILLER_18_585 VPWR VGND sg13g2_decap_8
XFILLER_33_555 VPWR VGND sg13g2_decap_8
XFILLER_45_382 VPWR VGND sg13g2_decap_8
XFILLER_21_739 VPWR VGND sg13g2_decap_8
XFILLER_20_249 VPWR VGND sg13g2_decap_8
XFILLER_29_817 VPWR VGND sg13g2_decap_8
XFILLER_28_349 VPWR VGND sg13g2_decap_8
XFILLER_37_861 VPWR VGND sg13g2_decap_8
XFILLER_44_809 VPWR VGND sg13g2_decap_8
XFILLER_43_319 VPWR VGND sg13g2_decap_8
XFILLER_24_544 VPWR VGND sg13g2_decap_8
XFILLER_36_382 VPWR VGND sg13g2_decap_8
XFILLER_12_739 VPWR VGND sg13g2_decap_8
XFILLER_11_249 VPWR VGND sg13g2_decap_8
XFILLER_3_459 VPWR VGND sg13g2_decap_8
XFILLER_19_305 VPWR VGND sg13g2_decap_8
XFILLER_47_658 VPWR VGND sg13g2_decap_8
XFILLER_46_168 VPWR VGND sg13g2_decap_8
XFILLER_27_371 VPWR VGND sg13g2_decap_8
XFILLER_15_522 VPWR VGND sg13g2_decap_8
XFILLER_42_330 VPWR VGND sg13g2_decap_8
XFILLER_43_886 VPWR VGND sg13g2_decap_8
XFILLER_15_599 VPWR VGND sg13g2_decap_8
XFILLER_30_569 VPWR VGND sg13g2_decap_8
XFILLER_7_721 VPWR VGND sg13g2_decap_8
XFILLER_6_242 VPWR VGND sg13g2_decap_8
XFILLER_7_798 VPWR VGND sg13g2_decap_8
XFILLER_38_614 VPWR VGND sg13g2_decap_8
XFILLER_1_63 VPWR VGND sg13g2_decap_8
XFILLER_26_809 VPWR VGND sg13g2_decap_8
XFILLER_19_872 VPWR VGND sg13g2_decap_8
XFILLER_37_168 VPWR VGND sg13g2_decap_8
XFILLER_18_382 VPWR VGND sg13g2_decap_8
XFILLER_34_853 VPWR VGND sg13g2_decap_8
XFILLER_33_352 VPWR VGND sg13g2_decap_8
XFILLER_21_536 VPWR VGND sg13g2_decap_8
XFILLER_20_39 VPWR VGND sg13g2_decap_8
XFILLER_28_102 VPWR VGND sg13g2_decap_4
XFILLER_29_614 VPWR VGND sg13g2_decap_8
XFILLER_28_146 VPWR VGND sg13g2_decap_8
XFILLER_44_606 VPWR VGND sg13g2_decap_8
XFILLER_16_319 VPWR VGND sg13g2_decap_8
XFILLER_43_116 VPWR VGND sg13g2_decap_8
XFILLER_45_25 VPWR VGND sg13g2_decap_8
XFILLER_25_853 VPWR VGND sg13g2_decap_8
XFILLER_24_341 VPWR VGND sg13g2_decap_8
XFILLER_12_536 VPWR VGND sg13g2_decap_8
XFILLER_40_823 VPWR VGND sg13g2_decap_8
XFILLER_8_529 VPWR VGND sg13g2_decap_8
XFILLER_4_746 VPWR VGND sg13g2_decap_8
XFILLER_3_256 VPWR VGND sg13g2_decap_8
XFILLER_19_102 VPWR VGND sg13g2_decap_8
XFILLER_47_455 VPWR VGND sg13g2_decap_8
XFILLER_19_81 VPWR VGND sg13g2_decap_8
XFILLER_19_179 VPWR VGND sg13g2_decap_8
XFILLER_35_639 VPWR VGND sg13g2_decap_8
XFILLER_16_886 VPWR VGND sg13g2_decap_8
XFILLER_31_801 VPWR VGND sg13g2_decap_8
XFILLER_15_396 VPWR VGND sg13g2_decap_8
XFILLER_43_683 VPWR VGND sg13g2_decap_8
XFILLER_31_878 VPWR VGND sg13g2_decap_8
XFILLER_30_366 VPWR VGND sg13g2_decap_8
XFILLER_7_595 VPWR VGND sg13g2_decap_8
XFILLER_38_411 VPWR VGND sg13g2_decap_8
XFILLER_26_606 VPWR VGND sg13g2_decap_8
XFILLER_38_488 VPWR VGND sg13g2_decap_8
XFILLER_15_39 VPWR VGND sg13g2_decap_8
XFILLER_34_650 VPWR VGND sg13g2_decap_8
XFILLER_22_823 VPWR VGND sg13g2_decap_8
XFILLER_21_333 VPWR VGND sg13g2_decap_8
XFILLER_1_749 VPWR VGND sg13g2_decap_8
XFILLER_0_259 VPWR VGND sg13g2_decap_8
XFILLER_29_411 VPWR VGND sg13g2_decap_8
XFILLER_29_488 VPWR VGND sg13g2_decap_8
XFILLER_44_403 VPWR VGND sg13g2_decap_8
XFILLER_16_116 VPWR VGND sg13g2_decap_8
XFILLER_25_650 VPWR VGND sg13g2_decap_8
XFILLER_13_823 VPWR VGND sg13g2_decap_8
XFILLER_40_620 VPWR VGND sg13g2_decap_8
XFILLER_9_816 VPWR VGND sg13g2_decap_8
XFILLER_12_333 VPWR VGND sg13g2_decap_8
XFILLER_8_326 VPWR VGND sg13g2_decap_8
XFILLER_40_697 VPWR VGND sg13g2_decap_8
XFILLER_4_543 VPWR VGND sg13g2_decap_8
XFILLER_21_60 VPWR VGND sg13g2_decap_8
XFILLER_48_742 VPWR VGND sg13g2_decap_8
XFILLER_47_252 VPWR VGND sg13g2_decap_8
XFILLER_35_436 VPWR VGND sg13g2_decap_8
XFILLER_16_683 VPWR VGND sg13g2_decap_8
XFILLER_43_480 VPWR VGND sg13g2_decap_8
XFILLER_15_193 VPWR VGND sg13g2_decap_8
XFILLER_30_163 VPWR VGND sg13g2_decap_8
XFILLER_31_675 VPWR VGND sg13g2_decap_8
XFILLER_8_893 VPWR VGND sg13g2_decap_8
XFILLER_7_392 VPWR VGND sg13g2_decap_8
XFILLER_7_84 VPWR VGND sg13g2_decap_8
XFILLER_39_742 VPWR VGND sg13g2_decap_8
XFILLER_26_403 VPWR VGND sg13g2_decap_8
XFILLER_38_285 VPWR VGND sg13g2_decap_8
XFILLER_42_918 VPWR VGND sg13g2_decap_8
XFILLER_22_620 VPWR VGND sg13g2_decap_8
XFILLER_21_130 VPWR VGND sg13g2_decap_8
XFILLER_10_837 VPWR VGND sg13g2_decap_8
XFILLER_22_697 VPWR VGND sg13g2_decap_8
XFILLER_1_546 VPWR VGND sg13g2_decap_8
XFILLER_49_539 VPWR VGND sg13g2_decap_8
XFILLER_29_285 VPWR VGND sg13g2_decap_8
XFILLER_44_200 VPWR VGND sg13g2_decap_8
XFILLER_17_469 VPWR VGND sg13g2_decap_8
XFILLER_45_767 VPWR VGND sg13g2_decap_8
XFILLER_16_60 VPWR VGND sg13g2_decap_8
XFILLER_32_417 VPWR VGND sg13g2_decap_8
XFILLER_44_277 VPWR VGND sg13g2_decap_8
XFILLER_13_620 VPWR VGND sg13g2_decap_8
XFILLER_9_613 VPWR VGND sg13g2_decap_8
XFILLER_12_130 VPWR VGND sg13g2_decap_8
XFILLER_8_123 VPWR VGND sg13g2_decap_8
XFILLER_13_697 VPWR VGND sg13g2_decap_8
XFILLER_40_494 VPWR VGND sg13g2_decap_8
XFILLER_32_81 VPWR VGND sg13g2_decap_8
XFILLER_5_830 VPWR VGND sg13g2_decap_8
XFILLER_4_340 VPWR VGND sg13g2_decap_8
XFILLER_35_233 VPWR VGND sg13g2_decap_8
XFILLER_36_767 VPWR VGND sg13g2_decap_8
XFILLER_23_417 VPWR VGND sg13g2_decap_8
XFILLER_16_480 VPWR VGND sg13g2_decap_8
XFILLER_12_18 VPWR VGND sg13g2_decap_8
XFILLER_31_472 VPWR VGND sg13g2_decap_8
XFILLER_8_690 VPWR VGND sg13g2_decap_8
XFILLER_26_200 VPWR VGND sg13g2_decap_8
XFILLER_15_907 VPWR VGND sg13g2_decap_8
XFILLER_27_756 VPWR VGND sg13g2_decap_8
XFILLER_14_417 VPWR VGND sg13g2_decap_8
XFILLER_26_277 VPWR VGND sg13g2_decap_8
XFILLER_42_715 VPWR VGND sg13g2_decap_8
XFILLER_41_247 VPWR VGND sg13g2_decap_8
XFILLER_10_634 VPWR VGND sg13g2_decap_8
XFILLER_22_494 VPWR VGND sg13g2_decap_8
XFILLER_6_627 VPWR VGND sg13g2_decap_8
XFILLER_5_137 VPWR VGND sg13g2_decap_8
XFILLER_2_844 VPWR VGND sg13g2_decap_8
XFILLER_1_343 VPWR VGND sg13g2_decap_8
XFILLER_49_336 VPWR VGND sg13g2_decap_8
XFILLER_18_767 VPWR VGND sg13g2_decap_8
XFILLER_27_70 VPWR VGND sg13g2_decap_8
XFILLER_45_564 VPWR VGND sg13g2_decap_8
XFILLER_17_266 VPWR VGND sg13g2_decap_8
XFILLER_32_214 VPWR VGND sg13g2_decap_8
XFILLER_33_737 VPWR VGND sg13g2_decap_8
XFILLER_9_410 VPWR VGND sg13g2_decap_8
XFILLER_13_494 VPWR VGND sg13g2_decap_8
XFILLER_40_291 VPWR VGND sg13g2_decap_8
XFILLER_9_487 VPWR VGND sg13g2_decap_8
XFILLER_4_74 VPWR VGND sg13g2_decap_8
XFILLER_23_214 VPWR VGND sg13g2_decap_8
XFILLER_24_726 VPWR VGND sg13g2_decap_8
XFILLER_36_564 VPWR VGND sg13g2_decap_8
XFILLER_20_921 VPWR VGND sg13g2_decap_4
XFILLER_23_39 VPWR VGND sg13g2_decap_8
XFILLER_32_781 VPWR VGND sg13g2_decap_8
XFILLER_48_14 VPWR VGND sg13g2_decap_8
XFILLER_27_553 VPWR VGND sg13g2_decap_8
XFILLER_15_704 VPWR VGND sg13g2_decap_8
XFILLER_42_512 VPWR VGND sg13g2_decap_8
XFILLER_14_214 VPWR VGND sg13g2_decap_8
XFILLER_42_589 VPWR VGND sg13g2_decap_8
XFILLER_11_921 VPWR VGND sg13g2_decap_4
XFILLER_23_781 VPWR VGND sg13g2_decap_8
XFILLER_10_431 VPWR VGND sg13g2_decap_8
XFILLER_7_903 VPWR VGND sg13g2_decap_8
XFILLER_22_291 VPWR VGND sg13g2_decap_8
XFILLER_6_424 VPWR VGND sg13g2_decap_8
XFILLER_2_641 VPWR VGND sg13g2_decap_8
XFILLER_1_140 VPWR VGND sg13g2_decap_8
XFILLER_49_133 VPWR VGND sg13g2_decap_8
X_41_ _04_ _06_ _10_ VPWR VGND sg13g2_nor2_1
XFILLER_46_840 VPWR VGND sg13g2_decap_8
XFILLER_18_564 VPWR VGND sg13g2_decap_8
XFILLER_45_361 VPWR VGND sg13g2_decap_8
XFILLER_33_534 VPWR VGND sg13g2_decap_8
XFILLER_21_718 VPWR VGND sg13g2_decap_8
XFILLER_14_781 VPWR VGND sg13g2_decap_8
XFILLER_20_228 VPWR VGND sg13g2_decap_8
XFILLER_13_291 VPWR VGND sg13g2_decap_8
XFILLER_9_284 VPWR VGND sg13g2_decap_8
XFILLER_48_0 VPWR VGND sg13g2_decap_8
XFILLER_18_39 VPWR VGND sg13g2_decap_8
XFILLER_28_328 VPWR VGND sg13g2_decap_8
XFILLER_37_840 VPWR VGND sg13g2_decap_8
XFILLER_36_361 VPWR VGND sg13g2_decap_8
XFILLER_24_523 VPWR VGND sg13g2_decap_8
XFILLER_12_718 VPWR VGND sg13g2_decap_8
XFILLER_34_49 VPWR VGND sg13g2_decap_8
XFILLER_11_228 VPWR VGND sg13g2_decap_8
XFILLER_20_795 VPWR VGND sg13g2_decap_8
XFILLER_3_438 VPWR VGND sg13g2_decap_8
XFILLER_47_637 VPWR VGND sg13g2_decap_8
XFILLER_46_147 VPWR VGND sg13g2_decap_8
XFILLER_15_501 VPWR VGND sg13g2_decap_8
XFILLER_27_350 VPWR VGND sg13g2_decap_8
XFILLER_28_895 VPWR VGND sg13g2_decap_8
XFILLER_15_578 VPWR VGND sg13g2_decap_8
XFILLER_43_865 VPWR VGND sg13g2_decap_8
XFILLER_24_60 VPWR VGND sg13g2_decap_8
XFILLER_42_386 VPWR VGND sg13g2_decap_8
XFILLER_7_700 VPWR VGND sg13g2_decap_8
XFILLER_24_82 VPWR VGND sg13g2_decap_8
XFILLER_30_548 VPWR VGND sg13g2_decap_8
XFILLER_7_777 VPWR VGND sg13g2_decap_8
XFILLER_6_221 VPWR VGND sg13g2_decap_8
XFILLER_11_795 VPWR VGND sg13g2_decap_8
XFILLER_40_81 VPWR VGND sg13g2_decap_8
XFILLER_6_298 VPWR VGND sg13g2_decap_8
XFILLER_1_42 VPWR VGND sg13g2_decap_8
XFILLER_19_851 VPWR VGND sg13g2_decap_8
XFILLER_37_147 VPWR VGND sg13g2_decap_8
XFILLER_18_361 VPWR VGND sg13g2_decap_8
XFILLER_34_832 VPWR VGND sg13g2_decap_8
XFILLER_33_331 VPWR VGND sg13g2_decap_8
XFILLER_21_515 VPWR VGND sg13g2_decap_8
XFILLER_20_18 VPWR VGND sg13g2_decap_8
XFILLER_28_125 VPWR VGND sg13g2_decap_8
XFILLER_24_320 VPWR VGND sg13g2_decap_8
XFILLER_25_832 VPWR VGND sg13g2_decap_8
XFILLER_40_802 VPWR VGND sg13g2_decap_8
XFILLER_12_515 VPWR VGND sg13g2_decap_8
XFILLER_24_397 VPWR VGND sg13g2_decap_8
XFILLER_8_508 VPWR VGND sg13g2_decap_8
XFILLER_40_879 VPWR VGND sg13g2_decap_8
XFILLER_20_592 VPWR VGND sg13g2_decap_8
XFILLER_4_725 VPWR VGND sg13g2_decap_8
XFILLER_3_235 VPWR VGND sg13g2_decap_8
XFILLER_10_95 VPWR VGND sg13g2_decap_8
XFILLER_48_924 VPWR VGND sg13g2_fill_1
XFILLER_47_434 VPWR VGND sg13g2_decap_8
XFILLER_19_60 VPWR VGND sg13g2_decap_8
XFILLER_19_158 VPWR VGND sg13g2_decap_8
XFILLER_35_618 VPWR VGND sg13g2_decap_8
XFILLER_28_692 VPWR VGND sg13g2_decap_8
XFILLER_34_139 VPWR VGND sg13g2_decap_8
XFILLER_16_865 VPWR VGND sg13g2_decap_8
XFILLER_43_662 VPWR VGND sg13g2_decap_8
XFILLER_15_375 VPWR VGND sg13g2_decap_8
XFILLER_35_81 VPWR VGND sg13g2_decap_8
XFILLER_30_345 VPWR VGND sg13g2_decap_8
XFILLER_31_857 VPWR VGND sg13g2_decap_8
XFILLER_42_183 VPWR VGND sg13g2_decap_8
XFILLER_11_592 VPWR VGND sg13g2_decap_8
XFILLER_7_574 VPWR VGND sg13g2_decap_8
XFILLER_39_924 VPWR VGND sg13g2_fill_1
XFILLER_38_467 VPWR VGND sg13g2_decap_8
XFILLER_25_139 VPWR VGND sg13g2_decap_8
XFILLER_15_18 VPWR VGND sg13g2_decap_8
XFILLER_22_802 VPWR VGND sg13g2_decap_8
XFILLER_21_312 VPWR VGND sg13g2_decap_8
XFILLER_40_109 VPWR VGND sg13g2_decap_8
XFILLER_22_879 VPWR VGND sg13g2_decap_8
XFILLER_21_389 VPWR VGND sg13g2_decap_8
Xoutput17 net17 uo_out[0] VPWR VGND sg13g2_buf_1
XFILLER_1_728 VPWR VGND sg13g2_decap_8
XFILLER_0_238 VPWR VGND sg13g2_decap_8
XFILLER_29_467 VPWR VGND sg13g2_decap_8
XFILLER_13_802 VPWR VGND sg13g2_decap_8
XFILLER_44_459 VPWR VGND sg13g2_decap_8
XFILLER_12_312 VPWR VGND sg13g2_decap_8
XFILLER_24_194 VPWR VGND sg13g2_decap_8
XFILLER_8_305 VPWR VGND sg13g2_decap_8
XFILLER_13_879 VPWR VGND sg13g2_decap_8
XFILLER_40_676 VPWR VGND sg13g2_decap_8
XFILLER_12_389 VPWR VGND sg13g2_decap_8
XFILLER_4_522 VPWR VGND sg13g2_decap_8
XFILLER_4_599 VPWR VGND sg13g2_decap_8
XFILLER_48_721 VPWR VGND sg13g2_decap_8
XFILLER_47_231 VPWR VGND sg13g2_decap_8
XFILLER_48_798 VPWR VGND sg13g2_decap_8
XFILLER_35_415 VPWR VGND sg13g2_decap_8
XFILLER_46_91 VPWR VGND sg13g2_decap_8
XFILLER_16_662 VPWR VGND sg13g2_decap_8
XFILLER_22_109 VPWR VGND sg13g2_decap_8
XFILLER_15_172 VPWR VGND sg13g2_decap_8
XFILLER_31_654 VPWR VGND sg13g2_decap_8
XFILLER_30_142 VPWR VGND sg13g2_decap_8
XFILLER_8_872 VPWR VGND sg13g2_decap_8
XFILLER_7_63 VPWR VGND sg13g2_decap_8
XFILLER_7_371 VPWR VGND sg13g2_decap_8
XFILLER_39_721 VPWR VGND sg13g2_decap_8
XFILLER_38_264 VPWR VGND sg13g2_decap_8
XFILLER_39_798 VPWR VGND sg13g2_decap_8
XFILLER_26_459 VPWR VGND sg13g2_decap_8
XFILLER_13_109 VPWR VGND sg13g2_decap_8
XFILLER_41_429 VPWR VGND sg13g2_decap_8
XFILLER_10_816 VPWR VGND sg13g2_decap_8
XFILLER_22_676 VPWR VGND sg13g2_decap_8
XFILLER_6_809 VPWR VGND sg13g2_decap_8
XFILLER_21_186 VPWR VGND sg13g2_decap_8
XFILLER_5_319 VPWR VGND sg13g2_decap_8
XFILLER_1_525 VPWR VGND sg13g2_decap_8
XFILLER_49_518 VPWR VGND sg13g2_decap_8
XFILLER_29_264 VPWR VGND sg13g2_decap_8
XFILLER_45_746 VPWR VGND sg13g2_decap_8
XFILLER_17_448 VPWR VGND sg13g2_decap_8
XFILLER_33_919 VPWR VGND sg13g2_decap_4
XFILLER_44_256 VPWR VGND sg13g2_decap_8
XFILLER_8_102 VPWR VGND sg13g2_decap_8
XFILLER_13_676 VPWR VGND sg13g2_decap_8
XFILLER_9_669 VPWR VGND sg13g2_decap_8
XFILLER_12_186 VPWR VGND sg13g2_decap_8
XFILLER_40_473 VPWR VGND sg13g2_decap_8
XFILLER_8_179 VPWR VGND sg13g2_decap_8
XFILLER_32_60 VPWR VGND sg13g2_decap_8
XFILLER_5_886 VPWR VGND sg13g2_decap_8
XFILLER_4_396 VPWR VGND sg13g2_decap_8
XFILLER_48_595 VPWR VGND sg13g2_decap_8
XFILLER_35_212 VPWR VGND sg13g2_decap_8
XFILLER_36_746 VPWR VGND sg13g2_decap_8
XFILLER_24_908 VPWR VGND sg13g2_decap_8
XFILLER_35_289 VPWR VGND sg13g2_decap_8
XFILLER_31_451 VPWR VGND sg13g2_decap_8
XFILLER_37_49 VPWR VGND sg13g2_decap_8
XFILLER_27_735 VPWR VGND sg13g2_decap_8
XFILLER_39_595 VPWR VGND sg13g2_decap_8
XFILLER_26_256 VPWR VGND sg13g2_decap_8
XFILLER_41_226 VPWR VGND sg13g2_decap_8
XFILLER_10_613 VPWR VGND sg13g2_decap_8
XFILLER_22_473 VPWR VGND sg13g2_decap_8
XFILLER_6_606 VPWR VGND sg13g2_decap_8
XFILLER_5_116 VPWR VGND sg13g2_decap_8
XFILLER_2_823 VPWR VGND sg13g2_decap_8
XFILLER_1_322 VPWR VGND sg13g2_decap_8
XFILLER_49_315 VPWR VGND sg13g2_decap_8
XFILLER_1_399 VPWR VGND sg13g2_decap_8
XFILLER_17_245 VPWR VGND sg13g2_decap_8
XFILLER_18_746 VPWR VGND sg13g2_decap_8
XFILLER_45_543 VPWR VGND sg13g2_decap_8
XFILLER_33_716 VPWR VGND sg13g2_decap_8
XFILLER_13_473 VPWR VGND sg13g2_decap_8
XFILLER_40_270 VPWR VGND sg13g2_decap_8
XFILLER_41_793 VPWR VGND sg13g2_decap_8
XFILLER_43_81 VPWR VGND sg13g2_decap_8
XFILLER_9_466 VPWR VGND sg13g2_decap_8
XFILLER_5_683 VPWR VGND sg13g2_decap_8
XFILLER_4_193 VPWR VGND sg13g2_decap_8
XFILLER_4_53 VPWR VGND sg13g2_decap_8
XFILLER_49_882 VPWR VGND sg13g2_decap_8
XFILLER_48_392 VPWR VGND sg13g2_decap_8
XFILLER_36_543 VPWR VGND sg13g2_decap_8
XFILLER_24_705 VPWR VGND sg13g2_decap_8
XFILLER_20_900 VPWR VGND sg13g2_decap_8
XFILLER_23_18 VPWR VGND sg13g2_decap_8
XFILLER_32_760 VPWR VGND sg13g2_decap_8
XFILLER_47_819 VPWR VGND sg13g2_decap_8
XFILLER_46_329 VPWR VGND sg13g2_decap_8
XFILLER_27_532 VPWR VGND sg13g2_decap_8
XFILLER_39_392 VPWR VGND sg13g2_decap_8
XFILLER_11_900 VPWR VGND sg13g2_decap_8
XFILLER_23_760 VPWR VGND sg13g2_decap_8
XFILLER_42_568 VPWR VGND sg13g2_decap_8
XFILLER_10_410 VPWR VGND sg13g2_decap_8
XFILLER_22_270 VPWR VGND sg13g2_decap_8
XFILLER_10_487 VPWR VGND sg13g2_decap_8
XFILLER_6_403 VPWR VGND sg13g2_decap_8
XFILLER_13_95 VPWR VGND sg13g2_decap_8
XFILLER_2_620 VPWR VGND sg13g2_decap_8
XFILLER_49_112 VPWR VGND sg13g2_decap_8
XFILLER_2_697 VPWR VGND sg13g2_decap_8
XFILLER_1_196 VPWR VGND sg13g2_decap_8
X_40_ net12 net4 _09_ VPWR VGND sg13g2_xor2_1
XFILLER_49_189 VPWR VGND sg13g2_decap_8
XFILLER_37_329 VPWR VGND sg13g2_decap_8
XFILLER_18_543 VPWR VGND sg13g2_decap_8
XFILLER_46_896 VPWR VGND sg13g2_decap_8
XFILLER_33_513 VPWR VGND sg13g2_decap_8
XFILLER_45_340 VPWR VGND sg13g2_decap_8
XFILLER_14_760 VPWR VGND sg13g2_decap_8
XFILLER_13_270 VPWR VGND sg13g2_decap_8
XFILLER_20_207 VPWR VGND sg13g2_decap_8
XFILLER_41_590 VPWR VGND sg13g2_decap_8
XFILLER_9_263 VPWR VGND sg13g2_decap_8
XFILLER_5_480 VPWR VGND sg13g2_decap_8
XFILLER_18_18 VPWR VGND sg13g2_decap_8
XFILLER_28_307 VPWR VGND sg13g2_decap_8
XFILLER_24_502 VPWR VGND sg13g2_decap_8
XFILLER_36_340 VPWR VGND sg13g2_decap_8
XFILLER_37_896 VPWR VGND sg13g2_decap_8
XFILLER_24_579 VPWR VGND sg13g2_decap_8
XFILLER_11_207 VPWR VGND sg13g2_decap_8
XFILLER_20_774 VPWR VGND sg13g2_decap_8
XFILLER_4_907 VPWR VGND sg13g2_decap_8
XFILLER_3_417 VPWR VGND sg13g2_decap_8
XFILLER_1_7 VPWR VGND sg13g2_decap_8
XFILLER_47_616 VPWR VGND sg13g2_decap_8
XFILLER_46_126 VPWR VGND sg13g2_decap_8
XFILLER_28_874 VPWR VGND sg13g2_decap_8
XFILLER_43_844 VPWR VGND sg13g2_decap_8
XFILLER_15_557 VPWR VGND sg13g2_decap_8
XFILLER_30_527 VPWR VGND sg13g2_decap_8
XFILLER_42_365 VPWR VGND sg13g2_decap_8
XFILLER_6_200 VPWR VGND sg13g2_decap_8
XFILLER_11_774 VPWR VGND sg13g2_decap_8
XFILLER_10_284 VPWR VGND sg13g2_decap_8
XFILLER_7_756 VPWR VGND sg13g2_decap_8
XFILLER_6_277 VPWR VGND sg13g2_decap_8
XFILLER_40_60 VPWR VGND sg13g2_decap_8
XFILLER_49_91 VPWR VGND sg13g2_decap_8
XFILLER_2_494 VPWR VGND sg13g2_decap_8
XFILLER_1_21 VPWR VGND sg13g2_decap_8
XFILLER_19_830 VPWR VGND sg13g2_decap_8
XFILLER_37_126 VPWR VGND sg13g2_decap_8
XFILLER_38_649 VPWR VGND sg13g2_decap_8
XFILLER_1_98 VPWR VGND sg13g2_decap_8
XFILLER_18_340 VPWR VGND sg13g2_decap_8
XFILLER_34_811 VPWR VGND sg13g2_decap_8
XFILLER_46_693 VPWR VGND sg13g2_decap_8
XFILLER_33_310 VPWR VGND sg13g2_decap_8
XFILLER_33_387 VPWR VGND sg13g2_decap_8
XFILLER_34_888 VPWR VGND sg13g2_decap_8
XFILLER_29_39 VPWR VGND sg13g2_decap_8
XFILLER_29_649 VPWR VGND sg13g2_decap_8
XFILLER_25_811 VPWR VGND sg13g2_decap_8
XFILLER_37_693 VPWR VGND sg13g2_decap_8
XFILLER_24_376 VPWR VGND sg13g2_decap_8
XFILLER_25_888 VPWR VGND sg13g2_decap_8
XFILLER_40_858 VPWR VGND sg13g2_decap_8
XFILLER_20_571 VPWR VGND sg13g2_decap_8
XFILLER_4_704 VPWR VGND sg13g2_decap_8
XFILLER_3_214 VPWR VGND sg13g2_decap_8
XFILLER_10_74 VPWR VGND sg13g2_decap_8
XFILLER_0_910 VPWR VGND sg13g2_decap_8
XFILLER_48_903 VPWR VGND sg13g2_decap_8
XFILLER_47_413 VPWR VGND sg13g2_decap_8
XFILLER_19_137 VPWR VGND sg13g2_decap_8
XFILLER_16_844 VPWR VGND sg13g2_decap_8
XFILLER_28_671 VPWR VGND sg13g2_decap_8
XFILLER_34_118 VPWR VGND sg13g2_decap_8
XFILLER_15_354 VPWR VGND sg13g2_decap_8
XFILLER_35_60 VPWR VGND sg13g2_decap_8
XFILLER_43_641 VPWR VGND sg13g2_decap_8
XFILLER_31_836 VPWR VGND sg13g2_decap_8
XFILLER_42_162 VPWR VGND sg13g2_decap_8
XFILLER_30_324 VPWR VGND sg13g2_decap_8
XFILLER_11_571 VPWR VGND sg13g2_decap_8
XFILLER_7_553 VPWR VGND sg13g2_decap_8
XFILLER_3_781 VPWR VGND sg13g2_decap_8
XFILLER_2_291 VPWR VGND sg13g2_decap_8
XFILLER_32_4 VPWR VGND sg13g2_decap_8
XFILLER_39_903 VPWR VGND sg13g2_decap_8
XFILLER_38_446 VPWR VGND sg13g2_decap_8
XFILLER_25_118 VPWR VGND sg13g2_decap_8
XFILLER_46_490 VPWR VGND sg13g2_decap_8
XFILLER_34_685 VPWR VGND sg13g2_decap_8
XFILLER_22_858 VPWR VGND sg13g2_decap_8
XFILLER_33_184 VPWR VGND sg13g2_decap_8
XFILLER_21_368 VPWR VGND sg13g2_decap_8
XFILLER_30_891 VPWR VGND sg13g2_decap_8
XFILLER_31_18 VPWR VGND sg13g2_decap_8
Xoutput18 net18 uo_out[1] VPWR VGND sg13g2_buf_1
XFILLER_1_707 VPWR VGND sg13g2_decap_8
XFILLER_0_217 VPWR VGND sg13g2_decap_8
XFILLER_29_446 VPWR VGND sg13g2_decap_8
XFILLER_44_438 VPWR VGND sg13g2_decap_8
XFILLER_37_490 VPWR VGND sg13g2_decap_8
XFILLER_25_685 VPWR VGND sg13g2_decap_8
XFILLER_13_858 VPWR VGND sg13g2_decap_8
XFILLER_24_173 VPWR VGND sg13g2_decap_8
XFILLER_12_368 VPWR VGND sg13g2_decap_8
XFILLER_40_655 VPWR VGND sg13g2_decap_8
XFILLER_4_501 VPWR VGND sg13g2_decap_8
XFILLER_21_95 VPWR VGND sg13g2_decap_8
XFILLER_4_578 VPWR VGND sg13g2_decap_8
XFILLER_48_700 VPWR VGND sg13g2_decap_8
XFILLER_47_210 VPWR VGND sg13g2_decap_8
XFILLER_0_784 VPWR VGND sg13g2_decap_8
XFILLER_48_777 VPWR VGND sg13g2_decap_8
XFILLER_47_287 VPWR VGND sg13g2_decap_8
XFILLER_46_70 VPWR VGND sg13g2_decap_8
XFILLER_16_641 VPWR VGND sg13g2_decap_8
XFILLER_15_151 VPWR VGND sg13g2_decap_8
XFILLER_30_121 VPWR VGND sg13g2_decap_8
XFILLER_31_633 VPWR VGND sg13g2_decap_8
XFILLER_8_851 VPWR VGND sg13g2_decap_8
XFILLER_7_350 VPWR VGND sg13g2_decap_8
XFILLER_7_42 VPWR VGND sg13g2_decap_8
XFILLER_30_198 VPWR VGND sg13g2_decap_8
XFILLER_39_700 VPWR VGND sg13g2_decap_8
XFILLER_27_917 VPWR VGND sg13g2_decap_8
XFILLER_38_243 VPWR VGND sg13g2_decap_8
XFILLER_39_777 VPWR VGND sg13g2_decap_8
XFILLER_26_18 VPWR VGND sg13g2_decap_8
XFILLER_26_438 VPWR VGND sg13g2_decap_8
XFILLER_41_408 VPWR VGND sg13g2_decap_8
XFILLER_34_482 VPWR VGND sg13g2_decap_8
XFILLER_22_655 VPWR VGND sg13g2_decap_8
XFILLER_21_165 VPWR VGND sg13g2_decap_8
XFILLER_1_504 VPWR VGND sg13g2_decap_8
XFILLER_29_243 VPWR VGND sg13g2_decap_8
XFILLER_17_427 VPWR VGND sg13g2_decap_8
XFILLER_45_725 VPWR VGND sg13g2_decap_8
XFILLER_44_235 VPWR VGND sg13g2_decap_8
XFILLER_16_95 VPWR VGND sg13g2_decap_8
XFILLER_25_482 VPWR VGND sg13g2_decap_8
XFILLER_13_655 VPWR VGND sg13g2_decap_8
XFILLER_40_452 VPWR VGND sg13g2_decap_8
XFILLER_9_648 VPWR VGND sg13g2_decap_8
XFILLER_12_165 VPWR VGND sg13g2_decap_8
XFILLER_8_158 VPWR VGND sg13g2_decap_8
XFILLER_5_865 VPWR VGND sg13g2_decap_8
XFILLER_4_375 VPWR VGND sg13g2_decap_8
XFILLER_0_581 VPWR VGND sg13g2_decap_8
XFILLER_48_574 VPWR VGND sg13g2_decap_8
XFILLER_36_725 VPWR VGND sg13g2_decap_8
XFILLER_35_268 VPWR VGND sg13g2_decap_8
XFILLER_31_430 VPWR VGND sg13g2_decap_8
XFILLER_37_28 VPWR VGND sg13g2_decap_8
XFILLER_27_714 VPWR VGND sg13g2_decap_8
XFILLER_39_574 VPWR VGND sg13g2_decap_8
XFILLER_26_235 VPWR VGND sg13g2_decap_8
XFILLER_41_205 VPWR VGND sg13g2_decap_8
XFILLER_22_452 VPWR VGND sg13g2_decap_8
XFILLER_10_669 VPWR VGND sg13g2_decap_8
XFILLER_1_301 VPWR VGND sg13g2_decap_8
XFILLER_2_802 VPWR VGND sg13g2_decap_8
XFILLER_2_879 VPWR VGND sg13g2_decap_8
XFILLER_1_378 VPWR VGND sg13g2_decap_8
XFILLER_18_725 VPWR VGND sg13g2_decap_8
XFILLER_17_224 VPWR VGND sg13g2_decap_8
XFILLER_45_522 VPWR VGND sg13g2_decap_8
XFILLER_45_599 VPWR VGND sg13g2_decap_8
XFILLER_13_452 VPWR VGND sg13g2_decap_8
XFILLER_32_249 VPWR VGND sg13g2_decap_8
XFILLER_41_772 VPWR VGND sg13g2_decap_8
XFILLER_43_60 VPWR VGND sg13g2_decap_8
XFILLER_9_445 VPWR VGND sg13g2_decap_8
XFILLER_5_662 VPWR VGND sg13g2_decap_8
XFILLER_4_172 VPWR VGND sg13g2_decap_8
XFILLER_4_32 VPWR VGND sg13g2_decap_8
XFILLER_49_861 VPWR VGND sg13g2_decap_8
XFILLER_48_371 VPWR VGND sg13g2_decap_8
XFILLER_36_522 VPWR VGND sg13g2_decap_8
XFILLER_17_791 VPWR VGND sg13g2_decap_8
XFILLER_36_599 VPWR VGND sg13g2_decap_8
XFILLER_23_249 VPWR VGND sg13g2_decap_8
XFILLER_2_109 VPWR VGND sg13g2_decap_8
XFILLER_48_49 VPWR VGND sg13g2_decap_8
XFILLER_46_308 VPWR VGND sg13g2_decap_8
XFILLER_27_511 VPWR VGND sg13g2_decap_8
XFILLER_39_371 VPWR VGND sg13g2_decap_8
XFILLER_15_739 VPWR VGND sg13g2_decap_8
XFILLER_27_588 VPWR VGND sg13g2_decap_8
XFILLER_42_547 VPWR VGND sg13g2_decap_8
XFILLER_14_249 VPWR VGND sg13g2_decap_8
XFILLER_30_709 VPWR VGND sg13g2_decap_8
XFILLER_10_466 VPWR VGND sg13g2_decap_8
XFILLER_13_74 VPWR VGND sg13g2_decap_8
XFILLER_6_459 VPWR VGND sg13g2_decap_8
XFILLER_2_676 VPWR VGND sg13g2_decap_8
XFILLER_1_175 VPWR VGND sg13g2_decap_8
XFILLER_49_168 VPWR VGND sg13g2_decap_8
XFILLER_37_308 VPWR VGND sg13g2_decap_8
XFILLER_18_522 VPWR VGND sg13g2_decap_8
XFILLER_38_82 VPWR VGND sg13g2_decap_8
XFILLER_46_875 VPWR VGND sg13g2_decap_8
XFILLER_18_599 VPWR VGND sg13g2_decap_8
XFILLER_45_396 VPWR VGND sg13g2_decap_8
XFILLER_33_569 VPWR VGND sg13g2_decap_8
XFILLER_9_242 VPWR VGND sg13g2_decap_8
XFILLER_37_875 VPWR VGND sg13g2_decap_8
XFILLER_34_18 VPWR VGND sg13g2_decap_8
XFILLER_36_396 VPWR VGND sg13g2_decap_8
XFILLER_24_558 VPWR VGND sg13g2_decap_8
XFILLER_20_753 VPWR VGND sg13g2_decap_8
XFILLER_46_105 VPWR VGND sg13g2_decap_8
XFILLER_19_319 VPWR VGND sg13g2_decap_8
XFILLER_28_853 VPWR VGND sg13g2_decap_8
XFILLER_15_536 VPWR VGND sg13g2_decap_8
XFILLER_27_385 VPWR VGND sg13g2_decap_8
XFILLER_43_823 VPWR VGND sg13g2_decap_8
XFILLER_42_344 VPWR VGND sg13g2_decap_8
XFILLER_30_506 VPWR VGND sg13g2_decap_8
XFILLER_11_753 VPWR VGND sg13g2_decap_8
XFILLER_10_263 VPWR VGND sg13g2_decap_8
XFILLER_7_735 VPWR VGND sg13g2_decap_8
XFILLER_6_256 VPWR VGND sg13g2_decap_8
XFILLER_2_473 VPWR VGND sg13g2_decap_8
XFILLER_49_70 VPWR VGND sg13g2_decap_8
XFILLER_27_7 VPWR VGND sg13g2_decap_8
XFILLER_37_105 VPWR VGND sg13g2_decap_8
XFILLER_38_628 VPWR VGND sg13g2_decap_8
XFILLER_1_77 VPWR VGND sg13g2_decap_8
XFILLER_46_672 VPWR VGND sg13g2_decap_8
XFILLER_19_886 VPWR VGND sg13g2_decap_8
XFILLER_18_396 VPWR VGND sg13g2_decap_8
XFILLER_34_867 VPWR VGND sg13g2_decap_8
XFILLER_45_193 VPWR VGND sg13g2_decap_8
XFILLER_33_366 VPWR VGND sg13g2_decap_8
XFILLER_29_18 VPWR VGND sg13g2_decap_8
XFILLER_29_628 VPWR VGND sg13g2_decap_8
XFILLER_28_116 VPWR VGND sg13g2_fill_1
XFILLER_37_672 VPWR VGND sg13g2_decap_8
XFILLER_45_39 VPWR VGND sg13g2_decap_8
XFILLER_25_867 VPWR VGND sg13g2_decap_8
XFILLER_36_193 VPWR VGND sg13g2_decap_8
XFILLER_24_355 VPWR VGND sg13g2_decap_8
XFILLER_40_837 VPWR VGND sg13g2_decap_8
XFILLER_20_550 VPWR VGND sg13g2_decap_8
XFILLER_10_53 VPWR VGND sg13g2_decap_8
XFILLER_19_116 VPWR VGND sg13g2_decap_8
XFILLER_47_469 VPWR VGND sg13g2_decap_8
XFILLER_19_95 VPWR VGND sg13g2_decap_8
XFILLER_28_650 VPWR VGND sg13g2_decap_8
XFILLER_16_823 VPWR VGND sg13g2_decap_8
XFILLER_43_620 VPWR VGND sg13g2_decap_8
XFILLER_15_333 VPWR VGND sg13g2_decap_8
XFILLER_27_182 VPWR VGND sg13g2_decap_8
XFILLER_30_303 VPWR VGND sg13g2_decap_8
XFILLER_31_815 VPWR VGND sg13g2_decap_8
XFILLER_42_141 VPWR VGND sg13g2_decap_8
XFILLER_43_697 VPWR VGND sg13g2_decap_8
XFILLER_11_550 VPWR VGND sg13g2_decap_8
XFILLER_7_532 VPWR VGND sg13g2_decap_8
XFILLER_3_760 VPWR VGND sg13g2_decap_8
XFILLER_2_270 VPWR VGND sg13g2_decap_8
XFILLER_25_4 VPWR VGND sg13g2_decap_8
XFILLER_38_425 VPWR VGND sg13g2_decap_8
XFILLER_19_683 VPWR VGND sg13g2_decap_8
XFILLER_18_193 VPWR VGND sg13g2_decap_8
XFILLER_33_163 VPWR VGND sg13g2_decap_8
XFILLER_34_664 VPWR VGND sg13g2_decap_8
XFILLER_22_837 VPWR VGND sg13g2_decap_8
XFILLER_21_347 VPWR VGND sg13g2_decap_8
XFILLER_30_870 VPWR VGND sg13g2_decap_8
Xoutput19 net19 uo_out[2] VPWR VGND sg13g2_buf_1
XFILLER_29_425 VPWR VGND sg13g2_decap_8
XFILLER_45_907 VPWR VGND sg13g2_decap_8
XFILLER_17_609 VPWR VGND sg13g2_decap_8
XFILLER_44_417 VPWR VGND sg13g2_decap_8
XFILLER_24_152 VPWR VGND sg13g2_decap_8
XFILLER_25_664 VPWR VGND sg13g2_decap_8
XFILLER_13_837 VPWR VGND sg13g2_decap_8
XFILLER_40_634 VPWR VGND sg13g2_decap_8
XFILLER_12_347 VPWR VGND sg13g2_decap_8
XFILLER_4_557 VPWR VGND sg13g2_decap_8
XFILLER_21_74 VPWR VGND sg13g2_decap_8
XFILLER_0_763 VPWR VGND sg13g2_decap_8
XFILLER_48_756 VPWR VGND sg13g2_decap_8
XFILLER_36_907 VPWR VGND sg13g2_decap_8
XFILLER_47_266 VPWR VGND sg13g2_decap_8
XFILLER_16_620 VPWR VGND sg13g2_decap_8
XFILLER_15_130 VPWR VGND sg13g2_decap_8
XFILLER_16_697 VPWR VGND sg13g2_decap_8
XFILLER_31_612 VPWR VGND sg13g2_decap_8
XFILLER_43_494 VPWR VGND sg13g2_decap_8
XFILLER_8_830 VPWR VGND sg13g2_decap_8
XFILLER_7_21 VPWR VGND sg13g2_decap_8
XFILLER_30_177 VPWR VGND sg13g2_decap_8
XFILLER_31_689 VPWR VGND sg13g2_decap_8
XFILLER_7_98 VPWR VGND sg13g2_decap_8
XFILLER_38_222 VPWR VGND sg13g2_decap_8
XFILLER_39_756 VPWR VGND sg13g2_decap_8
XFILLER_26_417 VPWR VGND sg13g2_decap_8
XFILLER_19_480 VPWR VGND sg13g2_decap_8
XFILLER_38_299 VPWR VGND sg13g2_decap_8
XFILLER_34_461 VPWR VGND sg13g2_decap_8
XFILLER_22_634 VPWR VGND sg13g2_decap_8
XFILLER_21_144 VPWR VGND sg13g2_decap_8
XFILLER_42_18 VPWR VGND sg13g2_decap_8
XFILLER_18_907 VPWR VGND sg13g2_decap_8
XFILLER_29_222 VPWR VGND sg13g2_decap_8
XFILLER_45_704 VPWR VGND sg13g2_decap_8
XFILLER_17_406 VPWR VGND sg13g2_decap_8
XFILLER_44_214 VPWR VGND sg13g2_decap_8
XFILLER_29_299 VPWR VGND sg13g2_decap_8
XFILLER_25_461 VPWR VGND sg13g2_decap_8
XFILLER_13_634 VPWR VGND sg13g2_decap_8
XFILLER_16_74 VPWR VGND sg13g2_decap_8
XFILLER_12_144 VPWR VGND sg13g2_decap_8
XFILLER_40_431 VPWR VGND sg13g2_decap_8
XFILLER_9_627 VPWR VGND sg13g2_decap_8
XFILLER_8_137 VPWR VGND sg13g2_decap_8
XFILLER_32_95 VPWR VGND sg13g2_decap_8
XFILLER_5_844 VPWR VGND sg13g2_decap_8
XFILLER_4_354 VPWR VGND sg13g2_decap_8
XFILLER_0_560 VPWR VGND sg13g2_decap_8
XFILLER_48_553 VPWR VGND sg13g2_decap_8
XFILLER_36_704 VPWR VGND sg13g2_decap_8
XFILLER_35_247 VPWR VGND sg13g2_decap_8
XFILLER_16_494 VPWR VGND sg13g2_decap_8
XFILLER_32_921 VPWR VGND sg13g2_decap_4
XFILLER_44_781 VPWR VGND sg13g2_decap_8
XFILLER_43_291 VPWR VGND sg13g2_decap_8
XFILLER_31_486 VPWR VGND sg13g2_decap_8
XFILLER_39_553 VPWR VGND sg13g2_decap_8
XFILLER_26_214 VPWR VGND sg13g2_decap_8
XFILLER_42_729 VPWR VGND sg13g2_decap_8
XFILLER_23_921 VPWR VGND sg13g2_decap_4
XFILLER_22_431 VPWR VGND sg13g2_decap_8
XFILLER_10_648 VPWR VGND sg13g2_decap_8
XFILLER_2_858 VPWR VGND sg13g2_decap_8
XFILLER_1_357 VPWR VGND sg13g2_decap_8
XFILLER_17_203 VPWR VGND sg13g2_decap_8
XFILLER_18_704 VPWR VGND sg13g2_decap_8
XFILLER_45_501 VPWR VGND sg13g2_decap_8
XFILLER_27_84 VPWR VGND sg13g2_decap_8
XFILLER_45_578 VPWR VGND sg13g2_decap_8
XFILLER_14_921 VPWR VGND sg13g2_decap_4
XFILLER_26_781 VPWR VGND sg13g2_decap_8
XFILLER_32_228 VPWR VGND sg13g2_decap_8
XFILLER_13_431 VPWR VGND sg13g2_decap_8
XFILLER_41_751 VPWR VGND sg13g2_decap_8
XFILLER_9_424 VPWR VGND sg13g2_decap_8
XFILLER_5_641 VPWR VGND sg13g2_decap_8
XFILLER_4_151 VPWR VGND sg13g2_decap_8
XFILLER_4_11 VPWR VGND sg13g2_decap_8
XFILLER_4_88 VPWR VGND sg13g2_decap_8
XFILLER_49_840 VPWR VGND sg13g2_decap_8
XFILLER_48_350 VPWR VGND sg13g2_decap_8
XFILLER_36_501 VPWR VGND sg13g2_decap_8
XFILLER_36_578 VPWR VGND sg13g2_decap_8
XFILLER_17_770 VPWR VGND sg13g2_decap_8
XFILLER_23_228 VPWR VGND sg13g2_decap_8
XFILLER_16_291 VPWR VGND sg13g2_decap_8
XFILLER_31_283 VPWR VGND sg13g2_decap_8
XFILLER_32_795 VPWR VGND sg13g2_decap_8
XFILLER_48_28 VPWR VGND sg13g2_decap_8
XFILLER_39_350 VPWR VGND sg13g2_decap_8
XFILLER_15_718 VPWR VGND sg13g2_decap_8
XFILLER_27_567 VPWR VGND sg13g2_decap_8
XFILLER_14_228 VPWR VGND sg13g2_decap_8
XFILLER_42_526 VPWR VGND sg13g2_decap_8
XFILLER_7_917 VPWR VGND sg13g2_decap_8
XFILLER_23_795 VPWR VGND sg13g2_decap_8
XFILLER_10_445 VPWR VGND sg13g2_decap_8
XFILLER_13_53 VPWR VGND sg13g2_decap_8
XFILLER_6_438 VPWR VGND sg13g2_decap_8
XFILLER_2_655 VPWR VGND sg13g2_decap_8
XFILLER_1_154 VPWR VGND sg13g2_decap_8
XFILLER_49_147 VPWR VGND sg13g2_decap_8
XFILLER_18_501 VPWR VGND sg13g2_decap_8
XFILLER_38_61 VPWR VGND sg13g2_decap_8
XFILLER_46_854 VPWR VGND sg13g2_decap_8
XFILLER_18_578 VPWR VGND sg13g2_decap_8
XFILLER_45_375 VPWR VGND sg13g2_decap_8
XFILLER_33_548 VPWR VGND sg13g2_decap_8
XFILLER_9_221 VPWR VGND sg13g2_decap_8
XFILLER_14_795 VPWR VGND sg13g2_decap_8
XFILLER_9_298 VPWR VGND sg13g2_decap_8
XFILLER_37_854 VPWR VGND sg13g2_decap_8
XFILLER_24_537 VPWR VGND sg13g2_decap_8
XFILLER_36_375 VPWR VGND sg13g2_decap_8
XFILLER_20_732 VPWR VGND sg13g2_decap_8
XFILLER_32_592 VPWR VGND sg13g2_decap_8
XFILLER_28_832 VPWR VGND sg13g2_decap_8
XFILLER_43_802 VPWR VGND sg13g2_decap_8
XFILLER_15_515 VPWR VGND sg13g2_decap_8
XFILLER_27_364 VPWR VGND sg13g2_decap_8
XFILLER_42_323 VPWR VGND sg13g2_decap_8
XFILLER_43_879 VPWR VGND sg13g2_decap_8
XFILLER_11_732 VPWR VGND sg13g2_decap_8
XFILLER_23_592 VPWR VGND sg13g2_decap_8
XFILLER_24_74 VPWR VGND sg13g2_fill_2
XFILLER_10_242 VPWR VGND sg13g2_decap_8
XFILLER_7_714 VPWR VGND sg13g2_decap_8
XFILLER_24_96 VPWR VGND sg13g2_decap_8
XFILLER_6_235 VPWR VGND sg13g2_decap_8
XFILLER_40_95 VPWR VGND sg13g2_decap_8
XFILLER_2_452 VPWR VGND sg13g2_decap_8
XFILLER_38_607 VPWR VGND sg13g2_decap_8
XFILLER_1_56 VPWR VGND sg13g2_decap_8
XFILLER_46_651 VPWR VGND sg13g2_decap_8
XFILLER_19_865 VPWR VGND sg13g2_decap_8
XFILLER_18_375 VPWR VGND sg13g2_decap_8
XFILLER_45_172 VPWR VGND sg13g2_decap_8
XFILLER_33_345 VPWR VGND sg13g2_decap_8
XFILLER_34_846 VPWR VGND sg13g2_decap_8
XFILLER_14_592 VPWR VGND sg13g2_decap_8
XFILLER_21_529 VPWR VGND sg13g2_decap_8
XFILLER_42_890 VPWR VGND sg13g2_decap_8
XFILLER_46_0 VPWR VGND sg13g2_decap_8
XFILLER_29_607 VPWR VGND sg13g2_decap_8
XFILLER_28_106 VPWR VGND sg13g2_fill_2
XFILLER_28_139 VPWR VGND sg13g2_decap_8
XFILLER_37_651 VPWR VGND sg13g2_decap_8
XFILLER_45_18 VPWR VGND sg13g2_decap_8
XFILLER_43_109 VPWR VGND sg13g2_decap_8
XFILLER_24_334 VPWR VGND sg13g2_decap_8
XFILLER_25_846 VPWR VGND sg13g2_decap_8
XFILLER_36_172 VPWR VGND sg13g2_decap_8
XFILLER_40_816 VPWR VGND sg13g2_decap_8
XFILLER_12_529 VPWR VGND sg13g2_decap_8
XFILLER_4_739 VPWR VGND sg13g2_decap_8
XFILLER_10_32 VPWR VGND sg13g2_decap_8
XFILLER_3_249 VPWR VGND sg13g2_decap_8
XFILLER_19_74 VPWR VGND sg13g2_decap_8
XFILLER_47_448 VPWR VGND sg13g2_decap_8
XFILLER_16_802 VPWR VGND sg13g2_decap_8
XFILLER_27_161 VPWR VGND sg13g2_decap_8
XFILLER_15_312 VPWR VGND sg13g2_decap_8
XFILLER_42_120 VPWR VGND sg13g2_decap_8
XFILLER_16_879 VPWR VGND sg13g2_decap_8
XFILLER_43_676 VPWR VGND sg13g2_decap_8
XFILLER_15_389 VPWR VGND sg13g2_decap_8
XFILLER_35_95 VPWR VGND sg13g2_decap_8
XFILLER_42_197 VPWR VGND sg13g2_decap_8
XFILLER_30_359 VPWR VGND sg13g2_decap_8
XFILLER_7_511 VPWR VGND sg13g2_decap_8
XFILLER_7_588 VPWR VGND sg13g2_decap_8
XFILLER_38_404 VPWR VGND sg13g2_decap_8
XFILLER_18_4 VPWR VGND sg13g2_decap_8
XFILLER_19_662 VPWR VGND sg13g2_decap_8
XFILLER_18_172 VPWR VGND sg13g2_decap_8
XFILLER_34_643 VPWR VGND sg13g2_decap_8
XFILLER_22_816 VPWR VGND sg13g2_decap_8
XFILLER_33_142 VPWR VGND sg13g2_decap_8
XFILLER_21_326 VPWR VGND sg13g2_decap_8
XFILLER_29_404 VPWR VGND sg13g2_decap_8
XFILLER_16_109 VPWR VGND sg13g2_decap_8
XFILLER_25_643 VPWR VGND sg13g2_decap_8
XFILLER_13_816 VPWR VGND sg13g2_decap_8
XFILLER_24_131 VPWR VGND sg13g2_decap_8
XFILLER_9_809 VPWR VGND sg13g2_decap_8
XFILLER_12_326 VPWR VGND sg13g2_decap_8
XFILLER_40_613 VPWR VGND sg13g2_decap_8
XFILLER_8_319 VPWR VGND sg13g2_decap_8
XFILLER_21_893 VPWR VGND sg13g2_decap_8
XFILLER_21_53 VPWR VGND sg13g2_decap_8
XFILLER_4_536 VPWR VGND sg13g2_decap_8
XFILLER_0_742 VPWR VGND sg13g2_decap_8
XFILLER_48_735 VPWR VGND sg13g2_decap_8
XFILLER_47_245 VPWR VGND sg13g2_decap_8
XFILLER_35_429 VPWR VGND sg13g2_decap_8
XFILLER_16_676 VPWR VGND sg13g2_decap_8
XFILLER_15_186 VPWR VGND sg13g2_decap_8
XFILLER_43_473 VPWR VGND sg13g2_decap_8
XFILLER_31_668 VPWR VGND sg13g2_decap_8
XFILLER_30_156 VPWR VGND sg13g2_decap_8
XFILLER_12_893 VPWR VGND sg13g2_decap_8
XFILLER_8_886 VPWR VGND sg13g2_decap_8
XFILLER_7_77 VPWR VGND sg13g2_decap_8
XFILLER_7_385 VPWR VGND sg13g2_decap_8
XFILLER_38_201 VPWR VGND sg13g2_decap_8
XFILLER_39_735 VPWR VGND sg13g2_decap_8
XFILLER_38_278 VPWR VGND sg13g2_decap_8
XFILLER_34_440 VPWR VGND sg13g2_decap_8
XFILLER_22_613 VPWR VGND sg13g2_decap_8
XFILLER_21_123 VPWR VGND sg13g2_decap_8
XFILLER_1_539 VPWR VGND sg13g2_decap_8
XFILLER_29_201 VPWR VGND sg13g2_decap_8
XFILLER_29_278 VPWR VGND sg13g2_decap_8
XFILLER_16_53 VPWR VGND sg13g2_decap_8
XFILLER_25_440 VPWR VGND sg13g2_decap_8
XFILLER_13_613 VPWR VGND sg13g2_decap_8
XFILLER_40_410 VPWR VGND sg13g2_decap_8
XFILLER_9_606 VPWR VGND sg13g2_decap_8
XFILLER_12_123 VPWR VGND sg13g2_decap_8
XFILLER_8_116 VPWR VGND sg13g2_decap_8
XFILLER_40_487 VPWR VGND sg13g2_decap_8
XFILLER_21_690 VPWR VGND sg13g2_decap_8
XFILLER_32_74 VPWR VGND sg13g2_decap_8
XFILLER_5_823 VPWR VGND sg13g2_decap_8
XFILLER_4_333 VPWR VGND sg13g2_decap_8
XFILLER_48_532 VPWR VGND sg13g2_decap_8
XFILLER_35_226 VPWR VGND sg13g2_decap_8
XFILLER_32_900 VPWR VGND sg13g2_decap_8
XFILLER_44_760 VPWR VGND sg13g2_decap_8
XFILLER_16_473 VPWR VGND sg13g2_decap_8
XFILLER_43_270 VPWR VGND sg13g2_decap_8
XFILLER_31_465 VPWR VGND sg13g2_decap_8
XFILLER_12_690 VPWR VGND sg13g2_decap_8
XFILLER_8_683 VPWR VGND sg13g2_decap_8
XFILLER_7_182 VPWR VGND sg13g2_decap_8
XFILLER_39_532 VPWR VGND sg13g2_decap_8
XFILLER_27_749 VPWR VGND sg13g2_decap_8
XFILLER_23_900 VPWR VGND sg13g2_decap_8
XFILLER_42_708 VPWR VGND sg13g2_decap_8
XFILLER_22_410 VPWR VGND sg13g2_decap_8
XFILLER_35_793 VPWR VGND sg13g2_decap_8
XFILLER_10_627 VPWR VGND sg13g2_decap_8
XFILLER_22_487 VPWR VGND sg13g2_decap_8
XFILLER_2_837 VPWR VGND sg13g2_decap_8
XFILLER_1_336 VPWR VGND sg13g2_decap_8
XFILLER_49_329 VPWR VGND sg13g2_decap_8
XFILLER_27_63 VPWR VGND sg13g2_decap_8
XFILLER_14_900 VPWR VGND sg13g2_decap_8
XFILLER_17_259 VPWR VGND sg13g2_decap_8
XFILLER_45_557 VPWR VGND sg13g2_decap_8
XFILLER_13_410 VPWR VGND sg13g2_decap_8
XFILLER_26_760 VPWR VGND sg13g2_decap_8
XFILLER_32_207 VPWR VGND sg13g2_decap_8
XFILLER_41_730 VPWR VGND sg13g2_decap_8
XFILLER_9_403 VPWR VGND sg13g2_decap_8
XFILLER_13_487 VPWR VGND sg13g2_decap_8
XFILLER_40_284 VPWR VGND sg13g2_decap_8
XFILLER_43_95 VPWR VGND sg13g2_decap_8
XFILLER_5_620 VPWR VGND sg13g2_decap_8
XFILLER_4_130 VPWR VGND sg13g2_decap_8
XFILLER_5_697 VPWR VGND sg13g2_decap_8
XFILLER_4_67 VPWR VGND sg13g2_decap_8
XFILLER_49_896 VPWR VGND sg13g2_decap_8
XFILLER_24_719 VPWR VGND sg13g2_decap_8
XFILLER_36_557 VPWR VGND sg13g2_decap_8
XFILLER_23_207 VPWR VGND sg13g2_decap_8
XFILLER_16_270 VPWR VGND sg13g2_decap_8
XFILLER_20_914 VPWR VGND sg13g2_decap_8
XFILLER_31_262 VPWR VGND sg13g2_decap_8
XFILLER_32_774 VPWR VGND sg13g2_decap_8
XFILLER_8_480 VPWR VGND sg13g2_decap_8
XFILLER_27_546 VPWR VGND sg13g2_decap_8
XFILLER_14_207 VPWR VGND sg13g2_decap_8
XFILLER_42_505 VPWR VGND sg13g2_decap_8
XFILLER_35_590 VPWR VGND sg13g2_decap_8
XFILLER_11_914 VPWR VGND sg13g2_decap_8
XFILLER_23_774 VPWR VGND sg13g2_decap_8
XFILLER_10_424 VPWR VGND sg13g2_decap_8
XFILLER_13_32 VPWR VGND sg13g2_decap_8
XFILLER_22_284 VPWR VGND sg13g2_decap_8
XFILLER_6_417 VPWR VGND sg13g2_decap_8
XFILLER_1_133 VPWR VGND sg13g2_decap_8
XFILLER_2_634 VPWR VGND sg13g2_decap_8
XFILLER_49_126 VPWR VGND sg13g2_decap_8
XFILLER_38_40 VPWR VGND sg13g2_decap_8
XFILLER_46_833 VPWR VGND sg13g2_decap_8
XFILLER_18_557 VPWR VGND sg13g2_decap_8
XFILLER_45_354 VPWR VGND sg13g2_decap_8
XFILLER_33_527 VPWR VGND sg13g2_decap_8
XFILLER_9_200 VPWR VGND sg13g2_decap_8
XFILLER_14_774 VPWR VGND sg13g2_decap_8
XFILLER_13_284 VPWR VGND sg13g2_decap_8
XFILLER_9_277 VPWR VGND sg13g2_decap_8
XFILLER_5_494 VPWR VGND sg13g2_decap_8
XFILLER_49_693 VPWR VGND sg13g2_decap_8
XFILLER_37_833 VPWR VGND sg13g2_decap_8
XFILLER_36_354 VPWR VGND sg13g2_decap_8
XFILLER_24_516 VPWR VGND sg13g2_decap_8
XFILLER_20_711 VPWR VGND sg13g2_decap_8
XFILLER_32_571 VPWR VGND sg13g2_decap_8
XFILLER_20_788 VPWR VGND sg13g2_decap_8
XFILLER_28_811 VPWR VGND sg13g2_decap_8
XFILLER_27_343 VPWR VGND sg13g2_decap_8
XFILLER_28_888 VPWR VGND sg13g2_decap_8
XFILLER_42_302 VPWR VGND sg13g2_decap_8
XFILLER_43_858 VPWR VGND sg13g2_decap_8
XFILLER_42_379 VPWR VGND sg13g2_decap_8
XFILLER_11_711 VPWR VGND sg13g2_decap_8
XFILLER_23_571 VPWR VGND sg13g2_decap_8
XFILLER_24_53 VPWR VGND sg13g2_decap_8
XFILLER_10_221 VPWR VGND sg13g2_decap_8
XFILLER_6_214 VPWR VGND sg13g2_decap_8
XFILLER_11_788 VPWR VGND sg13g2_decap_8
XFILLER_10_298 VPWR VGND sg13g2_decap_8
XFILLER_3_921 VPWR VGND sg13g2_decap_4
XFILLER_40_74 VPWR VGND sg13g2_decap_8
XFILLER_2_431 VPWR VGND sg13g2_decap_8
XFILLER_1_35 VPWR VGND sg13g2_decap_8
XFILLER_46_630 VPWR VGND sg13g2_decap_8
XFILLER_19_844 VPWR VGND sg13g2_decap_8
XFILLER_18_354 VPWR VGND sg13g2_decap_8
XFILLER_34_825 VPWR VGND sg13g2_decap_8
XFILLER_45_151 VPWR VGND sg13g2_decap_8
XFILLER_33_324 VPWR VGND sg13g2_decap_8
XFILLER_21_508 VPWR VGND sg13g2_decap_8
XFILLER_14_571 VPWR VGND sg13g2_decap_8
XFILLER_6_781 VPWR VGND sg13g2_decap_8
XFILLER_5_291 VPWR VGND sg13g2_decap_8
Xinput1 ui_in[0] net1 VPWR VGND sg13g2_buf_1
XFILLER_49_490 VPWR VGND sg13g2_decap_8
XFILLER_37_630 VPWR VGND sg13g2_decap_8
XFILLER_25_825 VPWR VGND sg13g2_decap_8
XFILLER_36_151 VPWR VGND sg13g2_decap_8
XFILLER_24_313 VPWR VGND sg13g2_decap_8
XFILLER_12_508 VPWR VGND sg13g2_decap_8
XFILLER_33_891 VPWR VGND sg13g2_decap_8
XFILLER_20_585 VPWR VGND sg13g2_decap_8
XFILLER_10_11 VPWR VGND sg13g2_decap_8
XFILLER_4_718 VPWR VGND sg13g2_decap_8
XFILLER_3_228 VPWR VGND sg13g2_decap_8
XFILLER_10_88 VPWR VGND sg13g2_decap_8
XFILLER_0_924 VPWR VGND sg13g2_fill_1
XFILLER_48_917 VPWR VGND sg13g2_decap_8
XFILLER_47_427 VPWR VGND sg13g2_decap_8
XFILLER_19_53 VPWR VGND sg13g2_decap_8
XFILLER_27_140 VPWR VGND sg13g2_decap_8
XFILLER_28_685 VPWR VGND sg13g2_decap_8
XFILLER_16_858 VPWR VGND sg13g2_decap_8
XFILLER_15_368 VPWR VGND sg13g2_decap_8
XFILLER_35_74 VPWR VGND sg13g2_decap_8
XFILLER_43_655 VPWR VGND sg13g2_decap_8
XFILLER_24_880 VPWR VGND sg13g2_decap_8
XFILLER_42_176 VPWR VGND sg13g2_decap_8
XFILLER_30_338 VPWR VGND sg13g2_decap_8
XFILLER_11_585 VPWR VGND sg13g2_decap_8
XFILLER_7_567 VPWR VGND sg13g2_decap_8
XFILLER_3_795 VPWR VGND sg13g2_decap_8
XFILLER_39_917 VPWR VGND sg13g2_decap_8
XFILLER_19_641 VPWR VGND sg13g2_decap_8
XFILLER_18_151 VPWR VGND sg13g2_decap_8
XFILLER_34_622 VPWR VGND sg13g2_decap_8
XFILLER_33_121 VPWR VGND sg13g2_decap_8
XFILLER_21_305 VPWR VGND sg13g2_decap_8
XFILLER_34_699 VPWR VGND sg13g2_decap_8
XFILLER_33_198 VPWR VGND sg13g2_decap_8
XFILLER_24_110 VPWR VGND sg13g2_decap_8
XFILLER_25_622 VPWR VGND sg13g2_decap_8
XFILLER_12_305 VPWR VGND sg13g2_decap_8
XFILLER_24_187 VPWR VGND sg13g2_decap_8
XFILLER_25_699 VPWR VGND sg13g2_decap_8
XFILLER_40_669 VPWR VGND sg13g2_decap_8
XFILLER_21_872 VPWR VGND sg13g2_decap_8
XFILLER_20_382 VPWR VGND sg13g2_decap_8
XFILLER_4_515 VPWR VGND sg13g2_decap_8
XFILLER_21_32 VPWR VGND sg13g2_decap_8
XFILLER_0_721 VPWR VGND sg13g2_decap_8
XFILLER_48_714 VPWR VGND sg13g2_decap_8
XFILLER_0_798 VPWR VGND sg13g2_decap_8
XFILLER_47_224 VPWR VGND sg13g2_decap_8
XFILLER_35_408 VPWR VGND sg13g2_decap_8
XFILLER_46_84 VPWR VGND sg13g2_decap_8
XFILLER_28_482 VPWR VGND sg13g2_decap_8
XFILLER_16_655 VPWR VGND sg13g2_decap_8
XFILLER_43_452 VPWR VGND sg13g2_decap_8
XFILLER_15_165 VPWR VGND sg13g2_decap_8
XFILLER_30_135 VPWR VGND sg13g2_decap_8
XFILLER_31_647 VPWR VGND sg13g2_decap_8
XFILLER_12_872 VPWR VGND sg13g2_decap_8
XFILLER_11_382 VPWR VGND sg13g2_decap_8
XFILLER_8_865 VPWR VGND sg13g2_decap_8
XFILLER_7_364 VPWR VGND sg13g2_decap_8
XFILLER_7_56 VPWR VGND sg13g2_decap_8
XFILLER_3_592 VPWR VGND sg13g2_decap_8
XFILLER_30_4 VPWR VGND sg13g2_decap_8
XFILLER_39_714 VPWR VGND sg13g2_decap_8
XFILLER_38_257 VPWR VGND sg13g2_decap_8
XFILLER_47_791 VPWR VGND sg13g2_decap_8
XFILLER_21_102 VPWR VGND sg13g2_decap_8
XFILLER_10_809 VPWR VGND sg13g2_decap_8
XFILLER_22_669 VPWR VGND sg13g2_decap_8
XFILLER_34_496 VPWR VGND sg13g2_decap_8
XFILLER_21_179 VPWR VGND sg13g2_decap_8
XFILLER_1_518 VPWR VGND sg13g2_decap_8
XFILLER_29_257 VPWR VGND sg13g2_decap_8
XFILLER_45_739 VPWR VGND sg13g2_decap_8
XFILLER_16_32 VPWR VGND sg13g2_decap_8
XFILLER_44_249 VPWR VGND sg13g2_decap_8
XFILLER_12_102 VPWR VGND sg13g2_decap_8
XFILLER_41_912 VPWR VGND sg13g2_decap_8
XFILLER_41_923 VPWR VGND sg13g2_fill_2
XFILLER_25_496 VPWR VGND sg13g2_decap_8
XFILLER_13_669 VPWR VGND sg13g2_decap_8
XFILLER_40_466 VPWR VGND sg13g2_decap_8
XFILLER_12_179 VPWR VGND sg13g2_decap_8
XFILLER_32_53 VPWR VGND sg13g2_decap_8
XFILLER_5_802 VPWR VGND sg13g2_decap_8
XFILLER_4_312 VPWR VGND sg13g2_decap_8
XFILLER_5_879 VPWR VGND sg13g2_decap_8
XFILLER_4_389 VPWR VGND sg13g2_decap_8
XFILLER_48_511 VPWR VGND sg13g2_decap_8
XFILLER_0_595 VPWR VGND sg13g2_decap_8
XFILLER_48_588 VPWR VGND sg13g2_decap_8
XFILLER_35_205 VPWR VGND sg13g2_decap_8
XFILLER_36_739 VPWR VGND sg13g2_decap_8
XFILLER_16_452 VPWR VGND sg13g2_decap_8
XFILLER_31_444 VPWR VGND sg13g2_decap_8
XFILLER_8_662 VPWR VGND sg13g2_decap_8
XFILLER_7_161 VPWR VGND sg13g2_decap_8
XFILLER_39_511 VPWR VGND sg13g2_decap_8
XFILLER_27_728 VPWR VGND sg13g2_decap_8
XFILLER_39_588 VPWR VGND sg13g2_decap_8
XFILLER_26_249 VPWR VGND sg13g2_decap_8
XFILLER_35_772 VPWR VGND sg13g2_decap_8
XFILLER_41_219 VPWR VGND sg13g2_decap_8
XFILLER_34_293 VPWR VGND sg13g2_decap_8
XFILLER_10_606 VPWR VGND sg13g2_decap_8
XFILLER_22_466 VPWR VGND sg13g2_decap_8
XFILLER_5_109 VPWR VGND sg13g2_decap_8
XFILLER_2_816 VPWR VGND sg13g2_decap_8
XFILLER_1_315 VPWR VGND sg13g2_decap_8
XFILLER_49_308 VPWR VGND sg13g2_decap_8
XFILLER_18_739 VPWR VGND sg13g2_decap_8
XFILLER_27_42 VPWR VGND sg13g2_decap_8
XFILLER_45_536 VPWR VGND sg13g2_decap_8
XFILLER_17_238 VPWR VGND sg13g2_decap_8
XFILLER_33_709 VPWR VGND sg13g2_decap_8
XFILLER_25_293 VPWR VGND sg13g2_decap_8
XFILLER_13_466 VPWR VGND sg13g2_decap_8
XFILLER_41_786 VPWR VGND sg13g2_decap_8
XFILLER_43_74 VPWR VGND sg13g2_decap_8
XFILLER_9_459 VPWR VGND sg13g2_decap_8
XFILLER_40_263 VPWR VGND sg13g2_decap_8
XFILLER_5_676 VPWR VGND sg13g2_decap_8
XFILLER_4_186 VPWR VGND sg13g2_decap_8
XFILLER_4_46 VPWR VGND sg13g2_decap_8
XFILLER_1_882 VPWR VGND sg13g2_decap_8
XFILLER_49_875 VPWR VGND sg13g2_decap_8
XFILLER_0_392 VPWR VGND sg13g2_decap_8
XFILLER_48_385 VPWR VGND sg13g2_decap_8
XFILLER_36_536 VPWR VGND sg13g2_decap_8
XFILLER_31_241 VPWR VGND sg13g2_decap_8
XFILLER_32_753 VPWR VGND sg13g2_decap_8
XFILLER_27_525 VPWR VGND sg13g2_decap_8
XFILLER_39_385 VPWR VGND sg13g2_decap_8
XFILLER_23_753 VPWR VGND sg13g2_decap_8
XFILLER_10_403 VPWR VGND sg13g2_decap_8
XFILLER_13_11 VPWR VGND sg13g2_decap_8
XFILLER_22_263 VPWR VGND sg13g2_decap_8
XFILLER_13_88 VPWR VGND sg13g2_decap_8
XFILLER_2_613 VPWR VGND sg13g2_decap_8
XFILLER_8_4 VPWR VGND sg13g2_decap_8
XFILLER_1_112 VPWR VGND sg13g2_decap_8
XFILLER_49_105 VPWR VGND sg13g2_decap_8
XFILLER_1_189 VPWR VGND sg13g2_decap_8
XFILLER_46_812 VPWR VGND sg13g2_decap_8
XFILLER_38_96 VPWR VGND sg13g2_decap_8
XFILLER_18_536 VPWR VGND sg13g2_decap_8
XFILLER_45_333 VPWR VGND sg13g2_decap_8
XFILLER_46_889 VPWR VGND sg13g2_decap_8
XFILLER_33_506 VPWR VGND sg13g2_decap_8
XFILLER_14_753 VPWR VGND sg13g2_decap_8
XFILLER_13_263 VPWR VGND sg13g2_decap_8
XFILLER_41_583 VPWR VGND sg13g2_decap_8
XFILLER_9_256 VPWR VGND sg13g2_decap_8
XFILLER_5_473 VPWR VGND sg13g2_decap_8
XFILLER_49_672 VPWR VGND sg13g2_decap_8
XFILLER_37_812 VPWR VGND sg13g2_decap_8
XFILLER_48_182 VPWR VGND sg13g2_decap_8
XFILLER_36_333 VPWR VGND sg13g2_decap_8
XFILLER_37_889 VPWR VGND sg13g2_decap_8
XFILLER_32_550 VPWR VGND sg13g2_decap_8
XFILLER_20_767 VPWR VGND sg13g2_decap_8
XFILLER_47_609 VPWR VGND sg13g2_decap_8
XFILLER_46_119 VPWR VGND sg13g2_decap_8
XFILLER_27_322 VPWR VGND sg13g2_decap_8
XFILLER_28_867 VPWR VGND sg13g2_decap_8
XFILLER_39_182 VPWR VGND sg13g2_decap_8
XFILLER_27_399 VPWR VGND sg13g2_decap_8
XFILLER_43_837 VPWR VGND sg13g2_decap_8
XFILLER_23_550 VPWR VGND sg13g2_decap_8
XFILLER_24_32 VPWR VGND sg13g2_decap_8
XFILLER_42_358 VPWR VGND sg13g2_decap_8
XFILLER_10_200 VPWR VGND sg13g2_decap_8
XFILLER_24_76 VPWR VGND sg13g2_fill_1
XFILLER_11_767 VPWR VGND sg13g2_decap_8
XFILLER_10_277 VPWR VGND sg13g2_decap_8
XFILLER_7_749 VPWR VGND sg13g2_decap_8
XFILLER_40_53 VPWR VGND sg13g2_decap_8
XFILLER_3_900 VPWR VGND sg13g2_decap_8
XFILLER_2_410 VPWR VGND sg13g2_decap_8
XFILLER_2_487 VPWR VGND sg13g2_decap_8
XFILLER_49_84 VPWR VGND sg13g2_decap_8
XFILLER_1_14 VPWR VGND sg13g2_decap_8
XFILLER_19_823 VPWR VGND sg13g2_decap_8
XFILLER_37_119 VPWR VGND sg13g2_decap_8
XFILLER_18_333 VPWR VGND sg13g2_decap_8
XFILLER_46_686 VPWR VGND sg13g2_decap_8
XFILLER_33_303 VPWR VGND sg13g2_decap_8
XFILLER_34_804 VPWR VGND sg13g2_decap_8
XFILLER_45_130 VPWR VGND sg13g2_decap_8
XFILLER_14_550 VPWR VGND sg13g2_decap_8
XFILLER_41_380 VPWR VGND sg13g2_decap_8
XFILLER_6_760 VPWR VGND sg13g2_decap_8
XFILLER_5_270 VPWR VGND sg13g2_decap_8
Xinput2 ui_in[1] net2 VPWR VGND sg13g2_buf_1
XFILLER_25_804 VPWR VGND sg13g2_decap_8
XFILLER_36_130 VPWR VGND sg13g2_decap_8
XFILLER_37_686 VPWR VGND sg13g2_decap_8
XFILLER_24_369 VPWR VGND sg13g2_decap_8
XFILLER_33_870 VPWR VGND sg13g2_decap_8
XFILLER_20_564 VPWR VGND sg13g2_decap_8
XFILLER_3_207 VPWR VGND sg13g2_decap_8
XFILLER_10_67 VPWR VGND sg13g2_decap_8
XFILLER_0_903 VPWR VGND sg13g2_decap_8
XFILLER_47_406 VPWR VGND sg13g2_decap_8
XFILLER_19_32 VPWR VGND sg13g2_decap_8
XFILLER_28_664 VPWR VGND sg13g2_decap_8
XFILLER_16_837 VPWR VGND sg13g2_decap_8
XFILLER_43_634 VPWR VGND sg13g2_decap_8
XFILLER_15_347 VPWR VGND sg13g2_decap_8
XFILLER_27_196 VPWR VGND sg13g2_decap_8
XFILLER_35_53 VPWR VGND sg13g2_decap_8
XFILLER_30_317 VPWR VGND sg13g2_decap_8
XFILLER_31_829 VPWR VGND sg13g2_decap_8
XFILLER_42_155 VPWR VGND sg13g2_decap_8
XFILLER_11_564 VPWR VGND sg13g2_decap_8
XFILLER_7_546 VPWR VGND sg13g2_decap_8
XFILLER_3_774 VPWR VGND sg13g2_decap_8
XFILLER_2_284 VPWR VGND sg13g2_decap_8
XFILLER_19_620 VPWR VGND sg13g2_decap_8
XFILLER_38_439 VPWR VGND sg13g2_decap_8
XFILLER_18_130 VPWR VGND sg13g2_decap_8
XFILLER_34_601 VPWR VGND sg13g2_decap_8
XFILLER_46_483 VPWR VGND sg13g2_decap_8
XFILLER_19_697 VPWR VGND sg13g2_decap_8
XFILLER_33_100 VPWR VGND sg13g2_decap_8
XFILLER_34_678 VPWR VGND sg13g2_decap_8
XFILLER_33_177 VPWR VGND sg13g2_decap_8
XFILLER_30_884 VPWR VGND sg13g2_decap_8
XFILLER_29_439 VPWR VGND sg13g2_decap_8
XFILLER_25_601 VPWR VGND sg13g2_decap_8
XFILLER_37_483 VPWR VGND sg13g2_decap_8
XFILLER_24_166 VPWR VGND sg13g2_decap_8
XFILLER_25_678 VPWR VGND sg13g2_decap_8
XFILLER_40_648 VPWR VGND sg13g2_decap_8
XFILLER_21_851 VPWR VGND sg13g2_decap_8
XFILLER_20_361 VPWR VGND sg13g2_decap_8
XFILLER_21_11 VPWR VGND sg13g2_decap_8
XFILLER_21_88 VPWR VGND sg13g2_decap_8
XFILLER_0_700 VPWR VGND sg13g2_decap_8
XFILLER_47_203 VPWR VGND sg13g2_decap_8
XFILLER_0_777 VPWR VGND sg13g2_decap_8
XFILLER_46_63 VPWR VGND sg13g2_decap_8
XFILLER_16_634 VPWR VGND sg13g2_decap_8
XFILLER_28_461 VPWR VGND sg13g2_decap_8
XFILLER_44_921 VPWR VGND sg13g2_decap_4
XFILLER_15_144 VPWR VGND sg13g2_decap_8
XFILLER_43_431 VPWR VGND sg13g2_decap_8
XFILLER_30_103 VPWR VGND sg13g2_decap_8
XFILLER_31_626 VPWR VGND sg13g2_decap_8
XFILLER_30_114 VPWR VGND sg13g2_decap_8
XFILLER_12_851 VPWR VGND sg13g2_decap_8
XFILLER_11_361 VPWR VGND sg13g2_decap_8
XFILLER_8_844 VPWR VGND sg13g2_decap_8
XFILLER_7_35 VPWR VGND sg13g2_decap_8
XFILLER_7_343 VPWR VGND sg13g2_decap_8
XFILLER_3_571 VPWR VGND sg13g2_decap_8
XFILLER_23_4 VPWR VGND sg13g2_decap_8
XFILLER_38_236 VPWR VGND sg13g2_decap_8
XFILLER_47_770 VPWR VGND sg13g2_decap_8
XFILLER_46_280 VPWR VGND sg13g2_decap_8
XFILLER_19_494 VPWR VGND sg13g2_decap_8
XFILLER_34_475 VPWR VGND sg13g2_decap_8
XFILLER_22_648 VPWR VGND sg13g2_decap_8
XFILLER_21_158 VPWR VGND sg13g2_decap_8
XFILLER_30_681 VPWR VGND sg13g2_decap_8
XFILLER_29_236 VPWR VGND sg13g2_decap_8
XFILLER_45_718 VPWR VGND sg13g2_decap_8
XFILLER_16_11 VPWR VGND sg13g2_decap_8
XFILLER_26_921 VPWR VGND sg13g2_decap_4
XFILLER_44_228 VPWR VGND sg13g2_decap_8
XFILLER_37_280 VPWR VGND sg13g2_decap_8
XFILLER_25_475 VPWR VGND sg13g2_decap_8
XFILLER_13_648 VPWR VGND sg13g2_decap_8
XFILLER_16_88 VPWR VGND sg13g2_decap_8
XFILLER_40_445 VPWR VGND sg13g2_decap_8
XFILLER_12_158 VPWR VGND sg13g2_decap_8
XFILLER_32_32 VPWR VGND sg13g2_decap_8
XFILLER_5_858 VPWR VGND sg13g2_decap_8
XFILLER_4_368 VPWR VGND sg13g2_decap_8
XFILLER_0_574 VPWR VGND sg13g2_decap_8
XFILLER_48_567 VPWR VGND sg13g2_decap_8
XFILLER_36_718 VPWR VGND sg13g2_decap_8
XFILLER_17_910 VPWR VGND sg13g2_decap_8
XFILLER_16_431 VPWR VGND sg13g2_decap_8
XFILLER_31_423 VPWR VGND sg13g2_decap_8
XFILLER_44_795 VPWR VGND sg13g2_decap_8
XFILLER_8_641 VPWR VGND sg13g2_decap_8
XFILLER_7_140 VPWR VGND sg13g2_decap_8
XFILLER_27_707 VPWR VGND sg13g2_decap_8
XFILLER_39_567 VPWR VGND sg13g2_decap_8
XFILLER_26_228 VPWR VGND sg13g2_decap_8
XFILLER_19_291 VPWR VGND sg13g2_decap_8
XFILLER_35_751 VPWR VGND sg13g2_decap_8
XFILLER_34_272 VPWR VGND sg13g2_decap_8
XFILLER_22_445 VPWR VGND sg13g2_decap_8
XFILLER_18_718 VPWR VGND sg13g2_decap_8
XFILLER_17_217 VPWR VGND sg13g2_decap_8
XFILLER_27_21 VPWR VGND sg13g2_decap_8
XFILLER_45_515 VPWR VGND sg13g2_decap_8
XFILLER_27_98 VPWR VGND sg13g2_decap_8
XFILLER_25_272 VPWR VGND sg13g2_decap_8
XFILLER_26_795 VPWR VGND sg13g2_decap_8
XFILLER_13_445 VPWR VGND sg13g2_decap_8
XFILLER_40_242 VPWR VGND sg13g2_decap_8
XFILLER_41_765 VPWR VGND sg13g2_decap_8
XFILLER_43_53 VPWR VGND sg13g2_decap_8
XFILLER_9_438 VPWR VGND sg13g2_decap_8
XFILLER_5_655 VPWR VGND sg13g2_decap_8
XFILLER_4_165 VPWR VGND sg13g2_decap_8
XFILLER_4_25 VPWR VGND sg13g2_decap_8
XFILLER_1_861 VPWR VGND sg13g2_decap_8
XFILLER_0_371 VPWR VGND sg13g2_decap_8
XFILLER_49_854 VPWR VGND sg13g2_decap_8
XFILLER_48_364 VPWR VGND sg13g2_decap_8
XFILLER_36_515 VPWR VGND sg13g2_decap_8
XFILLER_17_784 VPWR VGND sg13g2_decap_8
XFILLER_32_732 VPWR VGND sg13g2_decap_8
XFILLER_44_592 VPWR VGND sg13g2_decap_8
XFILLER_31_220 VPWR VGND sg13g2_decap_8
XFILLER_31_297 VPWR VGND sg13g2_decap_8
XFILLER_27_504 VPWR VGND sg13g2_decap_8
XFILLER_39_364 VPWR VGND sg13g2_decap_8
XFILLER_23_732 VPWR VGND sg13g2_decap_8
XFILLER_22_242 VPWR VGND sg13g2_decap_8
XFILLER_10_459 VPWR VGND sg13g2_decap_8
XFILLER_13_67 VPWR VGND sg13g2_decap_8
XFILLER_2_669 VPWR VGND sg13g2_decap_8
XFILLER_1_168 VPWR VGND sg13g2_decap_8
XFILLER_18_515 VPWR VGND sg13g2_decap_8
XFILLER_38_75 VPWR VGND sg13g2_decap_8
XFILLER_45_312 VPWR VGND sg13g2_decap_8
XFILLER_46_868 VPWR VGND sg13g2_decap_8
XFILLER_14_732 VPWR VGND sg13g2_decap_8
XFILLER_26_592 VPWR VGND sg13g2_decap_8
XFILLER_45_389 VPWR VGND sg13g2_decap_8
XFILLER_13_242 VPWR VGND sg13g2_decap_8
XFILLER_41_562 VPWR VGND sg13g2_decap_8
XFILLER_9_235 VPWR VGND sg13g2_decap_8
XFILLER_5_452 VPWR VGND sg13g2_decap_8
XFILLER_49_651 VPWR VGND sg13g2_decap_8
XFILLER_48_161 VPWR VGND sg13g2_decap_8
XFILLER_36_312 VPWR VGND sg13g2_decap_8
XFILLER_37_868 VPWR VGND sg13g2_decap_8
XFILLER_17_581 VPWR VGND sg13g2_decap_8
XFILLER_36_389 VPWR VGND sg13g2_decap_8
XFILLER_20_746 VPWR VGND sg13g2_decap_8
XFILLER_27_301 VPWR VGND sg13g2_decap_8
XFILLER_39_161 VPWR VGND sg13g2_decap_8
XFILLER_28_846 VPWR VGND sg13g2_decap_8
XFILLER_27_378 VPWR VGND sg13g2_decap_8
XFILLER_43_816 VPWR VGND sg13g2_decap_8
XFILLER_15_529 VPWR VGND sg13g2_decap_8
XFILLER_42_337 VPWR VGND sg13g2_decap_8
XFILLER_24_11 VPWR VGND sg13g2_decap_8
XFILLER_11_746 VPWR VGND sg13g2_decap_8
XFILLER_10_256 VPWR VGND sg13g2_decap_8
XFILLER_7_728 VPWR VGND sg13g2_decap_8
XFILLER_6_249 VPWR VGND sg13g2_decap_8
XFILLER_40_32 VPWR VGND sg13g2_decap_8
XFILLER_2_466 VPWR VGND sg13g2_decap_8
XFILLER_49_63 VPWR VGND sg13g2_decap_8
XFILLER_19_802 VPWR VGND sg13g2_decap_8
XFILLER_18_312 VPWR VGND sg13g2_decap_8
XFILLER_46_665 VPWR VGND sg13g2_decap_8
XFILLER_19_879 VPWR VGND sg13g2_decap_8
XFILLER_18_389 VPWR VGND sg13g2_decap_8
XFILLER_45_186 VPWR VGND sg13g2_decap_8
XFILLER_33_359 VPWR VGND sg13g2_decap_8
Xinput3 ui_in[2] net3 VPWR VGND sg13g2_buf_1
XFILLER_37_665 VPWR VGND sg13g2_decap_8
XFILLER_36_186 VPWR VGND sg13g2_decap_8
XFILLER_24_348 VPWR VGND sg13g2_decap_8
XFILLER_20_543 VPWR VGND sg13g2_decap_8
XFILLER_10_46 VPWR VGND sg13g2_decap_8
XFILLER_19_11 VPWR VGND sg13g2_decap_8
XFILLER_19_109 VPWR VGND sg13g2_decap_8
XFILLER_19_88 VPWR VGND sg13g2_decap_8
XFILLER_28_643 VPWR VGND sg13g2_decap_8
XFILLER_16_816 VPWR VGND sg13g2_decap_8
XFILLER_15_326 VPWR VGND sg13g2_decap_8
XFILLER_27_175 VPWR VGND sg13g2_decap_8
XFILLER_35_32 VPWR VGND sg13g2_decap_8
XFILLER_43_613 VPWR VGND sg13g2_decap_8
XFILLER_31_808 VPWR VGND sg13g2_decap_8
XFILLER_42_134 VPWR VGND sg13g2_decap_8
XFILLER_11_543 VPWR VGND sg13g2_decap_8
XFILLER_7_525 VPWR VGND sg13g2_decap_8
XFILLER_3_753 VPWR VGND sg13g2_decap_8
XFILLER_2_263 VPWR VGND sg13g2_decap_8
XFILLER_38_418 VPWR VGND sg13g2_decap_8
XFILLER_19_676 VPWR VGND sg13g2_decap_8
XFILLER_46_462 VPWR VGND sg13g2_decap_8
XFILLER_18_186 VPWR VGND sg13g2_decap_8
XFILLER_34_657 VPWR VGND sg13g2_decap_8
XFILLER_33_156 VPWR VGND sg13g2_decap_8
XFILLER_15_893 VPWR VGND sg13g2_decap_8
XFILLER_30_863 VPWR VGND sg13g2_decap_8
XFILLER_29_418 VPWR VGND sg13g2_decap_8
XFILLER_37_462 VPWR VGND sg13g2_decap_8
XFILLER_25_657 VPWR VGND sg13g2_decap_8
XFILLER_24_145 VPWR VGND sg13g2_decap_8
XFILLER_40_627 VPWR VGND sg13g2_decap_8
XFILLER_21_830 VPWR VGND sg13g2_decap_8
XFILLER_20_340 VPWR VGND sg13g2_decap_8
XFILLER_21_67 VPWR VGND sg13g2_decap_8
XFILLER_0_756 VPWR VGND sg13g2_decap_8
XFILLER_48_749 VPWR VGND sg13g2_decap_8
XFILLER_47_259 VPWR VGND sg13g2_decap_8
XFILLER_46_42 VPWR VGND sg13g2_decap_8
XFILLER_28_440 VPWR VGND sg13g2_decap_8
XFILLER_44_900 VPWR VGND sg13g2_decap_8
XFILLER_16_613 VPWR VGND sg13g2_decap_8
XFILLER_43_410 VPWR VGND sg13g2_decap_8
XFILLER_15_123 VPWR VGND sg13g2_decap_8
XFILLER_31_605 VPWR VGND sg13g2_decap_8
XFILLER_43_487 VPWR VGND sg13g2_decap_8
XFILLER_12_830 VPWR VGND sg13g2_decap_8
XFILLER_11_340 VPWR VGND sg13g2_decap_8
XFILLER_8_823 VPWR VGND sg13g2_decap_8
XFILLER_7_322 VPWR VGND sg13g2_decap_8
XFILLER_7_14 VPWR VGND sg13g2_decap_8
XFILLER_7_399 VPWR VGND sg13g2_decap_8
XFILLER_3_550 VPWR VGND sg13g2_decap_8
XFILLER_16_4 VPWR VGND sg13g2_decap_8
XFILLER_38_215 VPWR VGND sg13g2_decap_8
XFILLER_39_749 VPWR VGND sg13g2_decap_8
XFILLER_19_473 VPWR VGND sg13g2_decap_8
XFILLER_34_454 VPWR VGND sg13g2_decap_8
XFILLER_15_690 VPWR VGND sg13g2_decap_8
XFILLER_22_627 VPWR VGND sg13g2_decap_8
XFILLER_21_137 VPWR VGND sg13g2_decap_8
XFILLER_30_660 VPWR VGND sg13g2_decap_8
XFILLER_29_215 VPWR VGND sg13g2_decap_8
XFILLER_26_900 VPWR VGND sg13g2_decap_8
XFILLER_38_782 VPWR VGND sg13g2_decap_8
XFILLER_44_207 VPWR VGND sg13g2_decap_8
XFILLER_16_67 VPWR VGND sg13g2_decap_8
XFILLER_25_454 VPWR VGND sg13g2_decap_8
XFILLER_13_627 VPWR VGND sg13g2_decap_8
XFILLER_40_424 VPWR VGND sg13g2_decap_8
XFILLER_12_137 VPWR VGND sg13g2_decap_8
XFILLER_32_11 VPWR VGND sg13g2_decap_8
XFILLER_32_88 VPWR VGND sg13g2_decap_8
XFILLER_5_837 VPWR VGND sg13g2_decap_8
XFILLER_4_347 VPWR VGND sg13g2_decap_8
XFILLER_0_553 VPWR VGND sg13g2_decap_8
XFILLER_48_546 VPWR VGND sg13g2_decap_8
XFILLER_29_782 VPWR VGND sg13g2_decap_8
XFILLER_16_410 VPWR VGND sg13g2_decap_8
XFILLER_31_402 VPWR VGND sg13g2_decap_8
XFILLER_32_914 VPWR VGND sg13g2_decap_8
XFILLER_44_774 VPWR VGND sg13g2_decap_8
XFILLER_16_487 VPWR VGND sg13g2_decap_8
XFILLER_43_284 VPWR VGND sg13g2_decap_8
XFILLER_8_620 VPWR VGND sg13g2_decap_8
XFILLER_31_479 VPWR VGND sg13g2_decap_8
XFILLER_8_697 VPWR VGND sg13g2_decap_8
XFILLER_7_196 VPWR VGND sg13g2_decap_8
XFILLER_39_546 VPWR VGND sg13g2_decap_8
XFILLER_26_207 VPWR VGND sg13g2_decap_8
XFILLER_19_270 VPWR VGND sg13g2_decap_8
XFILLER_35_730 VPWR VGND sg13g2_decap_8
XFILLER_23_914 VPWR VGND sg13g2_decap_8
XFILLER_34_251 VPWR VGND sg13g2_decap_8
XFILLER_22_424 VPWR VGND sg13g2_decap_8
XFILLER_27_77 VPWR VGND sg13g2_decap_8
XFILLER_14_914 VPWR VGND sg13g2_decap_8
XFILLER_25_251 VPWR VGND sg13g2_decap_8
XFILLER_26_774 VPWR VGND sg13g2_decap_8
XFILLER_13_424 VPWR VGND sg13g2_decap_8
XFILLER_43_32 VPWR VGND sg13g2_decap_8
XFILLER_9_417 VPWR VGND sg13g2_decap_8
XFILLER_40_221 VPWR VGND sg13g2_decap_8
XFILLER_41_744 VPWR VGND sg13g2_decap_8
XFILLER_40_298 VPWR VGND sg13g2_decap_8
XFILLER_5_634 VPWR VGND sg13g2_decap_8
XFILLER_4_144 VPWR VGND sg13g2_decap_8
XFILLER_1_840 VPWR VGND sg13g2_decap_8
XFILLER_49_833 VPWR VGND sg13g2_decap_8
XFILLER_0_350 VPWR VGND sg13g2_decap_8
XFILLER_48_343 VPWR VGND sg13g2_decap_8
XFILLER_17_763 VPWR VGND sg13g2_decap_8
XFILLER_16_284 VPWR VGND sg13g2_decap_8
XFILLER_32_711 VPWR VGND sg13g2_decap_8
XFILLER_44_571 VPWR VGND sg13g2_decap_8
XFILLER_31_276 VPWR VGND sg13g2_decap_8
XFILLER_32_788 VPWR VGND sg13g2_decap_8
XFILLER_8_494 VPWR VGND sg13g2_decap_8
XFILLER_39_343 VPWR VGND sg13g2_decap_8
XFILLER_42_519 VPWR VGND sg13g2_decap_8
XFILLER_23_711 VPWR VGND sg13g2_decap_8
XFILLER_22_221 VPWR VGND sg13g2_decap_8
XFILLER_23_788 VPWR VGND sg13g2_decap_8
XFILLER_10_438 VPWR VGND sg13g2_decap_8
XFILLER_13_46 VPWR VGND sg13g2_decap_8
XFILLER_22_298 VPWR VGND sg13g2_decap_8
XFILLER_2_648 VPWR VGND sg13g2_decap_8
XFILLER_1_147 VPWR VGND sg13g2_decap_8
XFILLER_38_54 VPWR VGND sg13g2_decap_8
XFILLER_46_847 VPWR VGND sg13g2_decap_8
XFILLER_45_368 VPWR VGND sg13g2_decap_8
XFILLER_14_711 VPWR VGND sg13g2_decap_8
XFILLER_26_571 VPWR VGND sg13g2_decap_8
XFILLER_13_221 VPWR VGND sg13g2_decap_8
XFILLER_41_541 VPWR VGND sg13g2_decap_8
XFILLER_9_214 VPWR VGND sg13g2_decap_8
XFILLER_14_788 VPWR VGND sg13g2_decap_8
XFILLER_13_298 VPWR VGND sg13g2_decap_8
XFILLER_6_921 VPWR VGND sg13g2_decap_4
XFILLER_5_431 VPWR VGND sg13g2_decap_8
XFILLER_48_7 VPWR VGND sg13g2_decap_8
XFILLER_49_630 VPWR VGND sg13g2_decap_8
XFILLER_48_140 VPWR VGND sg13g2_decap_8
XFILLER_37_847 VPWR VGND sg13g2_decap_8
XFILLER_36_368 VPWR VGND sg13g2_decap_8
XFILLER_17_560 VPWR VGND sg13g2_decap_8
XFILLER_20_725 VPWR VGND sg13g2_decap_8
XFILLER_32_585 VPWR VGND sg13g2_decap_8
XFILLER_9_781 VPWR VGND sg13g2_decap_8
XFILLER_8_291 VPWR VGND sg13g2_decap_8
XFILLER_28_825 VPWR VGND sg13g2_decap_8
XFILLER_39_140 VPWR VGND sg13g2_decap_8
XFILLER_15_508 VPWR VGND sg13g2_decap_8
XFILLER_27_357 VPWR VGND sg13g2_decap_8
XFILLER_42_316 VPWR VGND sg13g2_decap_8
XFILLER_11_725 VPWR VGND sg13g2_decap_8
XFILLER_24_67 VPWR VGND sg13g2_decap_8
XFILLER_7_707 VPWR VGND sg13g2_decap_8
XFILLER_23_585 VPWR VGND sg13g2_decap_8
XFILLER_24_89 VPWR VGND sg13g2_decap_8
XFILLER_10_235 VPWR VGND sg13g2_decap_8
XFILLER_40_11 VPWR VGND sg13g2_decap_8
XFILLER_6_228 VPWR VGND sg13g2_decap_8
XFILLER_40_88 VPWR VGND sg13g2_decap_8
XFILLER_2_445 VPWR VGND sg13g2_decap_8
XFILLER_49_42 VPWR VGND sg13g2_decap_8
XFILLER_46_644 VPWR VGND sg13g2_decap_8
XFILLER_1_49 VPWR VGND sg13g2_decap_8
XFILLER_19_858 VPWR VGND sg13g2_decap_8
XFILLER_18_368 VPWR VGND sg13g2_decap_8
XFILLER_34_839 VPWR VGND sg13g2_decap_8
XFILLER_45_165 VPWR VGND sg13g2_decap_8
XFILLER_33_338 VPWR VGND sg13g2_decap_8
XFILLER_42_883 VPWR VGND sg13g2_decap_8
XFILLER_14_585 VPWR VGND sg13g2_decap_8
XFILLER_6_795 VPWR VGND sg13g2_decap_8
Xinput4 ui_in[3] net4 VPWR VGND sg13g2_buf_1
XFILLER_37_644 VPWR VGND sg13g2_decap_8
XFILLER_24_327 VPWR VGND sg13g2_decap_8
XFILLER_25_839 VPWR VGND sg13g2_decap_8
XFILLER_36_165 VPWR VGND sg13g2_decap_8
XFILLER_40_809 VPWR VGND sg13g2_decap_8
XFILLER_20_522 VPWR VGND sg13g2_decap_8
XFILLER_32_382 VPWR VGND sg13g2_decap_8
XFILLER_20_599 VPWR VGND sg13g2_decap_8
XFILLER_10_25 VPWR VGND sg13g2_decap_8
XFILLER_19_67 VPWR VGND sg13g2_decap_8
XFILLER_28_622 VPWR VGND sg13g2_decap_8
XFILLER_15_305 VPWR VGND sg13g2_decap_8
XFILLER_27_154 VPWR VGND sg13g2_decap_8
XFILLER_28_699 VPWR VGND sg13g2_decap_8
XFILLER_35_11 VPWR VGND sg13g2_decap_8
XFILLER_42_113 VPWR VGND sg13g2_decap_8
XFILLER_43_669 VPWR VGND sg13g2_decap_8
XFILLER_35_88 VPWR VGND sg13g2_decap_8
XFILLER_11_522 VPWR VGND sg13g2_decap_8
XFILLER_23_382 VPWR VGND sg13g2_decap_8
XFILLER_24_894 VPWR VGND sg13g2_decap_8
XFILLER_7_504 VPWR VGND sg13g2_decap_8
XFILLER_11_599 VPWR VGND sg13g2_decap_8
XFILLER_3_732 VPWR VGND sg13g2_decap_8
XFILLER_2_242 VPWR VGND sg13g2_decap_8
XFILLER_46_441 VPWR VGND sg13g2_decap_8
XFILLER_19_655 VPWR VGND sg13g2_decap_8
XFILLER_18_165 VPWR VGND sg13g2_decap_8
XFILLER_22_809 VPWR VGND sg13g2_decap_8
XFILLER_33_135 VPWR VGND sg13g2_decap_8
XFILLER_34_636 VPWR VGND sg13g2_decap_8
XFILLER_15_872 VPWR VGND sg13g2_decap_8
XFILLER_21_319 VPWR VGND sg13g2_decap_8
XFILLER_14_382 VPWR VGND sg13g2_decap_8
XFILLER_42_680 VPWR VGND sg13g2_decap_8
XFILLER_30_842 VPWR VGND sg13g2_decap_8
XFILLER_6_592 VPWR VGND sg13g2_decap_8
XFILLER_37_0 VPWR VGND sg13g2_decap_8
XFILLER_2_81 VPWR VGND sg13g2_decap_8
XFILLER_37_441 VPWR VGND sg13g2_decap_8
XFILLER_24_124 VPWR VGND sg13g2_decap_8
XFILLER_25_636 VPWR VGND sg13g2_decap_8
XFILLER_13_809 VPWR VGND sg13g2_decap_8
XFILLER_40_606 VPWR VGND sg13g2_decap_8
XFILLER_12_319 VPWR VGND sg13g2_decap_8
XFILLER_21_886 VPWR VGND sg13g2_decap_8
XFILLER_20_396 VPWR VGND sg13g2_decap_8
XFILLER_21_46 VPWR VGND sg13g2_decap_8
XFILLER_4_529 VPWR VGND sg13g2_decap_8
XFILLER_0_735 VPWR VGND sg13g2_decap_8
XFILLER_48_728 VPWR VGND sg13g2_decap_8
XFILLER_47_238 VPWR VGND sg13g2_decap_8
XFILLER_46_21 VPWR VGND sg13g2_decap_8
XFILLER_46_98 VPWR VGND sg13g2_decap_8
XFILLER_15_102 VPWR VGND sg13g2_decap_8
XFILLER_28_496 VPWR VGND sg13g2_decap_8
XFILLER_16_669 VPWR VGND sg13g2_decap_8
XFILLER_43_466 VPWR VGND sg13g2_decap_8
XFILLER_15_179 VPWR VGND sg13g2_decap_8
XFILLER_24_691 VPWR VGND sg13g2_decap_8
XFILLER_8_802 VPWR VGND sg13g2_decap_8
XFILLER_30_149 VPWR VGND sg13g2_decap_8
XFILLER_7_301 VPWR VGND sg13g2_decap_8
XFILLER_12_886 VPWR VGND sg13g2_decap_8
XFILLER_11_396 VPWR VGND sg13g2_decap_8
XFILLER_8_879 VPWR VGND sg13g2_decap_8
XFILLER_7_378 VPWR VGND sg13g2_decap_8
XFILLER_39_728 VPWR VGND sg13g2_decap_8
XFILLER_19_452 VPWR VGND sg13g2_decap_8
XFILLER_35_912 VPWR VGND sg13g2_decap_8
XFILLER_35_923 VPWR VGND sg13g2_fill_2
XFILLER_34_433 VPWR VGND sg13g2_decap_8
XFILLER_22_606 VPWR VGND sg13g2_decap_8
XFILLER_21_116 VPWR VGND sg13g2_decap_8
XFILLER_38_761 VPWR VGND sg13g2_decap_8
XFILLER_25_433 VPWR VGND sg13g2_decap_8
XFILLER_13_606 VPWR VGND sg13g2_decap_8
XFILLER_16_46 VPWR VGND sg13g2_decap_8
XFILLER_12_116 VPWR VGND sg13g2_decap_8
XFILLER_40_403 VPWR VGND sg13g2_decap_8
XFILLER_8_109 VPWR VGND sg13g2_decap_8
XFILLER_21_683 VPWR VGND sg13g2_decap_8
XFILLER_20_193 VPWR VGND sg13g2_decap_8
XFILLER_32_67 VPWR VGND sg13g2_decap_8
XFILLER_5_816 VPWR VGND sg13g2_decap_8
XFILLER_4_326 VPWR VGND sg13g2_decap_8
XFILLER_0_532 VPWR VGND sg13g2_decap_8
XFILLER_48_525 VPWR VGND sg13g2_decap_8
XFILLER_29_761 VPWR VGND sg13g2_decap_8
XFILLER_35_219 VPWR VGND sg13g2_decap_8
XFILLER_28_293 VPWR VGND sg13g2_decap_8
XFILLER_16_466 VPWR VGND sg13g2_decap_8
XFILLER_44_753 VPWR VGND sg13g2_decap_8
XFILLER_43_263 VPWR VGND sg13g2_decap_8
XFILLER_31_458 VPWR VGND sg13g2_decap_8
XFILLER_12_683 VPWR VGND sg13g2_decap_8
XFILLER_11_193 VPWR VGND sg13g2_decap_8
XFILLER_8_676 VPWR VGND sg13g2_decap_8
XFILLER_7_175 VPWR VGND sg13g2_decap_8
XFILLER_4_893 VPWR VGND sg13g2_decap_8
XFILLER_39_525 VPWR VGND sg13g2_decap_8
XFILLER_34_230 VPWR VGND sg13g2_decap_8
XFILLER_22_403 VPWR VGND sg13g2_decap_8
XFILLER_35_786 VPWR VGND sg13g2_decap_8
XFILLER_1_329 VPWR VGND sg13g2_decap_8
XFILLER_27_56 VPWR VGND sg13g2_decap_8
XFILLER_25_230 VPWR VGND sg13g2_decap_8
XFILLER_26_753 VPWR VGND sg13g2_decap_8
XFILLER_13_403 VPWR VGND sg13g2_decap_8
XFILLER_40_200 VPWR VGND sg13g2_decap_8
XFILLER_41_723 VPWR VGND sg13g2_decap_8
XFILLER_43_11 VPWR VGND sg13g2_decap_8
XFILLER_40_277 VPWR VGND sg13g2_decap_8
XFILLER_43_88 VPWR VGND sg13g2_decap_8
XFILLER_21_480 VPWR VGND sg13g2_decap_8
XFILLER_5_613 VPWR VGND sg13g2_decap_8
XFILLER_4_123 VPWR VGND sg13g2_decap_8
XFILLER_49_812 VPWR VGND sg13g2_decap_8
XFILLER_1_896 VPWR VGND sg13g2_decap_8
XFILLER_48_322 VPWR VGND sg13g2_decap_8
XFILLER_49_889 VPWR VGND sg13g2_decap_8
XFILLER_48_399 VPWR VGND sg13g2_decap_8
XFILLER_17_742 VPWR VGND sg13g2_decap_8
XFILLER_44_550 VPWR VGND sg13g2_decap_8
XFILLER_16_263 VPWR VGND sg13g2_decap_8
XFILLER_20_907 VPWR VGND sg13g2_decap_8
XFILLER_32_767 VPWR VGND sg13g2_decap_8
XFILLER_31_255 VPWR VGND sg13g2_decap_8
XFILLER_12_480 VPWR VGND sg13g2_decap_8
XFILLER_8_473 VPWR VGND sg13g2_decap_8
XFILLER_4_690 VPWR VGND sg13g2_decap_8
XFILLER_39_322 VPWR VGND sg13g2_decap_8
XFILLER_27_539 VPWR VGND sg13g2_decap_8
XFILLER_39_399 VPWR VGND sg13g2_decap_8
XFILLER_22_200 VPWR VGND sg13g2_decap_8
XFILLER_35_583 VPWR VGND sg13g2_decap_8
XFILLER_11_907 VPWR VGND sg13g2_decap_8
XFILLER_23_767 VPWR VGND sg13g2_decap_8
XFILLER_10_417 VPWR VGND sg13g2_decap_8
XFILLER_22_277 VPWR VGND sg13g2_decap_8
XFILLER_13_25 VPWR VGND sg13g2_decap_8
XFILLER_2_627 VPWR VGND sg13g2_decap_8
XFILLER_1_126 VPWR VGND sg13g2_decap_8
XFILLER_49_119 VPWR VGND sg13g2_decap_8
XFILLER_38_11 VPWR VGND sg13g2_decap_4
XFILLER_38_33 VPWR VGND sg13g2_decap_8
XFILLER_46_826 VPWR VGND sg13g2_decap_8
XFILLER_26_550 VPWR VGND sg13g2_decap_8
XFILLER_45_347 VPWR VGND sg13g2_decap_8
XFILLER_13_200 VPWR VGND sg13g2_decap_8
XFILLER_41_520 VPWR VGND sg13g2_decap_8
XFILLER_14_767 VPWR VGND sg13g2_decap_8
XFILLER_13_277 VPWR VGND sg13g2_decap_8
XFILLER_41_597 VPWR VGND sg13g2_decap_8
XFILLER_6_900 VPWR VGND sg13g2_decap_8
XFILLER_5_410 VPWR VGND sg13g2_decap_8
XFILLER_5_487 VPWR VGND sg13g2_decap_8
XFILLER_1_693 VPWR VGND sg13g2_decap_8
XFILLER_37_826 VPWR VGND sg13g2_decap_8
XFILLER_49_686 VPWR VGND sg13g2_decap_8
XFILLER_48_196 VPWR VGND sg13g2_decap_8
XFILLER_24_509 VPWR VGND sg13g2_decap_8
XFILLER_36_347 VPWR VGND sg13g2_decap_8
XFILLER_20_704 VPWR VGND sg13g2_decap_8
XFILLER_32_564 VPWR VGND sg13g2_decap_8
XFILLER_9_760 VPWR VGND sg13g2_decap_8
XFILLER_8_270 VPWR VGND sg13g2_decap_8
XFILLER_5_81 VPWR VGND sg13g2_decap_8
XFILLER_28_804 VPWR VGND sg13g2_decap_8
XFILLER_27_336 VPWR VGND sg13g2_decap_8
XFILLER_39_196 VPWR VGND sg13g2_decap_8
XFILLER_35_380 VPWR VGND sg13g2_decap_8
XFILLER_11_704 VPWR VGND sg13g2_decap_8
XFILLER_23_564 VPWR VGND sg13g2_decap_8
XFILLER_24_46 VPWR VGND sg13g2_decap_8
XFILLER_10_214 VPWR VGND sg13g2_decap_8
XFILLER_6_207 VPWR VGND sg13g2_decap_8
XFILLER_40_67 VPWR VGND sg13g2_decap_8
XFILLER_3_914 VPWR VGND sg13g2_decap_8
XFILLER_49_21 VPWR VGND sg13g2_decap_8
XFILLER_6_4 VPWR VGND sg13g2_decap_8
XFILLER_2_424 VPWR VGND sg13g2_decap_8
XFILLER_49_98 VPWR VGND sg13g2_decap_8
XFILLER_1_28 VPWR VGND sg13g2_decap_8
XFILLER_46_623 VPWR VGND sg13g2_decap_8
XFILLER_19_837 VPWR VGND sg13g2_decap_8
XFILLER_18_347 VPWR VGND sg13g2_decap_8
XFILLER_34_818 VPWR VGND sg13g2_decap_8
XFILLER_45_144 VPWR VGND sg13g2_decap_8
XFILLER_33_317 VPWR VGND sg13g2_decap_8
XFILLER_14_564 VPWR VGND sg13g2_decap_8
XFILLER_42_862 VPWR VGND sg13g2_decap_8
XFILLER_41_394 VPWR VGND sg13g2_decap_8
XFILLER_10_781 VPWR VGND sg13g2_decap_8
XFILLER_6_774 VPWR VGND sg13g2_decap_8
XFILLER_5_284 VPWR VGND sg13g2_decap_8
XFILLER_39_4 VPWR VGND sg13g2_decap_8
XFILLER_1_490 VPWR VGND sg13g2_decap_8
XFILLER_49_483 VPWR VGND sg13g2_decap_8
Xinput5 ui_in[4] net5 VPWR VGND sg13g2_buf_1
XFILLER_37_623 VPWR VGND sg13g2_decap_8
XFILLER_36_144 VPWR VGND sg13g2_decap_8
XFILLER_24_306 VPWR VGND sg13g2_decap_8
XFILLER_25_818 VPWR VGND sg13g2_decap_8
XFILLER_20_501 VPWR VGND sg13g2_decap_8
XFILLER_32_361 VPWR VGND sg13g2_decap_8
XFILLER_33_884 VPWR VGND sg13g2_decap_8
XFILLER_20_578 VPWR VGND sg13g2_decap_8
XFILLER_0_917 VPWR VGND sg13g2_decap_8
XFILLER_19_46 VPWR VGND sg13g2_decap_8
XFILLER_28_601 VPWR VGND sg13g2_decap_8
XFILLER_27_133 VPWR VGND sg13g2_decap_8
XFILLER_28_678 VPWR VGND sg13g2_decap_8
XFILLER_35_67 VPWR VGND sg13g2_decap_8
XFILLER_43_648 VPWR VGND sg13g2_decap_8
XFILLER_24_873 VPWR VGND sg13g2_decap_8
XFILLER_42_169 VPWR VGND sg13g2_decap_8
XFILLER_11_501 VPWR VGND sg13g2_decap_8
XFILLER_23_361 VPWR VGND sg13g2_decap_8
XFILLER_11_578 VPWR VGND sg13g2_decap_8
XFILLER_3_711 VPWR VGND sg13g2_decap_8
XFILLER_2_221 VPWR VGND sg13g2_decap_8
XFILLER_3_788 VPWR VGND sg13g2_decap_8
XFILLER_2_298 VPWR VGND sg13g2_decap_8
XFILLER_47_910 VPWR VGND sg13g2_decap_8
XFILLER_46_420 VPWR VGND sg13g2_decap_8
XFILLER_19_634 VPWR VGND sg13g2_decap_8
XFILLER_18_144 VPWR VGND sg13g2_decap_8
XFILLER_34_615 VPWR VGND sg13g2_decap_8
XFILLER_46_497 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_40 VPWR VGND uio_out[7] sg13g2_tielo
XFILLER_33_114 VPWR VGND sg13g2_decap_8
XFILLER_15_851 VPWR VGND sg13g2_decap_8
XFILLER_14_361 VPWR VGND sg13g2_decap_8
XFILLER_30_821 VPWR VGND sg13g2_decap_8
XFILLER_41_191 VPWR VGND sg13g2_decap_8
XFILLER_30_898 VPWR VGND sg13g2_decap_8
XFILLER_6_571 VPWR VGND sg13g2_decap_8
XFILLER_2_60 VPWR VGND sg13g2_decap_8
XFILLER_49_280 VPWR VGND sg13g2_decap_8
XFILLER_37_420 VPWR VGND sg13g2_decap_8
XFILLER_25_615 VPWR VGND sg13g2_decap_8
X_59_ net7 net15 _25_ VPWR VGND sg13g2_nor2_1
XFILLER_24_103 VPWR VGND sg13g2_decap_8
XFILLER_37_497 VPWR VGND sg13g2_decap_8
XFILLER_33_681 VPWR VGND sg13g2_decap_8
XFILLER_21_865 VPWR VGND sg13g2_decap_8
XFILLER_20_375 VPWR VGND sg13g2_decap_8
XFILLER_21_25 VPWR VGND sg13g2_decap_8
XFILLER_4_508 VPWR VGND sg13g2_decap_8
XFILLER_0_714 VPWR VGND sg13g2_decap_8
XFILLER_48_707 VPWR VGND sg13g2_decap_8
XFILLER_47_217 VPWR VGND sg13g2_decap_8
XFILLER_46_77 VPWR VGND sg13g2_decap_8
XFILLER_28_475 VPWR VGND sg13g2_decap_8
XFILLER_16_648 VPWR VGND sg13g2_decap_8
XFILLER_15_158 VPWR VGND sg13g2_decap_8
XFILLER_43_445 VPWR VGND sg13g2_decap_8
XFILLER_24_670 VPWR VGND sg13g2_decap_8
XFILLER_30_128 VPWR VGND sg13g2_decap_8
XFILLER_12_865 VPWR VGND sg13g2_decap_8
XFILLER_11_375 VPWR VGND sg13g2_decap_8
XFILLER_8_858 VPWR VGND sg13g2_decap_8
XFILLER_7_357 VPWR VGND sg13g2_decap_8
XFILLER_7_49 VPWR VGND sg13g2_decap_8
XFILLER_3_585 VPWR VGND sg13g2_decap_8
XFILLER_39_707 VPWR VGND sg13g2_decap_8
XFILLER_19_431 VPWR VGND sg13g2_decap_8
XFILLER_47_784 VPWR VGND sg13g2_decap_8
XFILLER_46_294 VPWR VGND sg13g2_decap_8
XFILLER_34_412 VPWR VGND sg13g2_decap_8
XFILLER_34_489 VPWR VGND sg13g2_decap_8
XFILLER_30_695 VPWR VGND sg13g2_decap_8
XFILLER_38_740 VPWR VGND sg13g2_decap_8
XFILLER_16_25 VPWR VGND sg13g2_decap_8
XFILLER_25_412 VPWR VGND sg13g2_decap_8
XFILLER_37_294 VPWR VGND sg13g2_decap_8
XFILLER_41_905 VPWR VGND sg13g2_decap_8
XFILLER_25_489 VPWR VGND sg13g2_decap_8
XFILLER_40_459 VPWR VGND sg13g2_decap_8
XFILLER_21_662 VPWR VGND sg13g2_decap_8
XFILLER_32_46 VPWR VGND sg13g2_decap_8
XFILLER_20_172 VPWR VGND sg13g2_decap_8
XFILLER_4_305 VPWR VGND sg13g2_decap_8
XFILLER_0_511 VPWR VGND sg13g2_decap_8
XFILLER_48_504 VPWR VGND sg13g2_decap_8
XFILLER_0_588 VPWR VGND sg13g2_decap_8
XFILLER_29_740 VPWR VGND sg13g2_decap_8
XFILLER_17_924 VPWR VGND sg13g2_fill_1
XFILLER_28_272 VPWR VGND sg13g2_decap_8
XFILLER_44_732 VPWR VGND sg13g2_decap_8
XFILLER_16_445 VPWR VGND sg13g2_decap_8
XFILLER_43_242 VPWR VGND sg13g2_decap_8
XFILLER_31_437 VPWR VGND sg13g2_decap_8
XFILLER_12_662 VPWR VGND sg13g2_decap_8
XFILLER_11_172 VPWR VGND sg13g2_decap_8
XFILLER_8_655 VPWR VGND sg13g2_decap_8
XFILLER_7_154 VPWR VGND sg13g2_decap_8
XFILLER_4_872 VPWR VGND sg13g2_decap_8
XFILLER_3_382 VPWR VGND sg13g2_decap_8
XFILLER_21_4 VPWR VGND sg13g2_decap_8
XFILLER_39_504 VPWR VGND sg13g2_decap_8
XFILLER_47_581 VPWR VGND sg13g2_decap_8
XFILLER_35_765 VPWR VGND sg13g2_decap_8
XFILLER_22_459 VPWR VGND sg13g2_decap_8
XFILLER_34_286 VPWR VGND sg13g2_decap_8
XFILLER_30_492 VPWR VGND sg13g2_decap_8
XFILLER_8_81 VPWR VGND sg13g2_decap_8
XFILLER_2_809 VPWR VGND sg13g2_decap_8
XFILLER_1_308 VPWR VGND sg13g2_decap_8
XFILLER_27_35 VPWR VGND sg13g2_decap_8
XFILLER_26_732 VPWR VGND sg13g2_decap_8
XFILLER_45_529 VPWR VGND sg13g2_decap_8
XFILLER_41_702 VPWR VGND sg13g2_decap_8
XFILLER_13_459 VPWR VGND sg13g2_decap_8
XFILLER_25_286 VPWR VGND sg13g2_decap_8
XFILLER_40_256 VPWR VGND sg13g2_decap_8
XFILLER_41_779 VPWR VGND sg13g2_decap_8
XFILLER_43_67 VPWR VGND sg13g2_decap_8
XFILLER_4_102 VPWR VGND sg13g2_decap_8
XFILLER_5_669 VPWR VGND sg13g2_decap_8
XFILLER_4_179 VPWR VGND sg13g2_decap_8
XFILLER_4_39 VPWR VGND sg13g2_decap_8
XFILLER_48_301 VPWR VGND sg13g2_decap_8
XFILLER_1_875 VPWR VGND sg13g2_decap_8
XFILLER_49_868 VPWR VGND sg13g2_decap_8
XFILLER_0_385 VPWR VGND sg13g2_decap_8
XFILLER_48_378 VPWR VGND sg13g2_decap_8
XFILLER_17_721 VPWR VGND sg13g2_decap_8
XFILLER_36_529 VPWR VGND sg13g2_decap_8
XFILLER_16_242 VPWR VGND sg13g2_decap_8
XFILLER_17_798 VPWR VGND sg13g2_decap_8
XFILLER_31_234 VPWR VGND sg13g2_decap_8
XFILLER_32_746 VPWR VGND sg13g2_decap_8
XFILLER_8_452 VPWR VGND sg13g2_decap_8
XFILLER_39_301 VPWR VGND sg13g2_decap_8
XFILLER_27_518 VPWR VGND sg13g2_decap_8
XFILLER_39_378 VPWR VGND sg13g2_decap_8
XFILLER_35_562 VPWR VGND sg13g2_decap_8
XFILLER_23_746 VPWR VGND sg13g2_decap_8
XFILLER_22_256 VPWR VGND sg13g2_decap_8
XFILLER_2_606 VPWR VGND sg13g2_decap_8
XFILLER_1_105 VPWR VGND sg13g2_decap_8
XFILLER_46_805 VPWR VGND sg13g2_decap_8
XFILLER_18_529 VPWR VGND sg13g2_decap_8
XFILLER_38_89 VPWR VGND sg13g2_decap_8
XFILLER_45_326 VPWR VGND sg13g2_decap_8
XFILLER_14_746 VPWR VGND sg13g2_decap_8
XFILLER_13_256 VPWR VGND sg13g2_decap_8
XFILLER_41_576 VPWR VGND sg13g2_decap_8
XFILLER_9_249 VPWR VGND sg13g2_decap_8
XFILLER_5_466 VPWR VGND sg13g2_decap_8
XFILLER_1_672 VPWR VGND sg13g2_decap_8
XFILLER_49_665 VPWR VGND sg13g2_decap_8
XFILLER_0_182 VPWR VGND sg13g2_decap_8
XFILLER_37_805 VPWR VGND sg13g2_decap_8
XFILLER_48_175 VPWR VGND sg13g2_decap_8
XFILLER_36_326 VPWR VGND sg13g2_decap_8
XFILLER_45_893 VPWR VGND sg13g2_decap_8
XFILLER_17_595 VPWR VGND sg13g2_decap_8
XFILLER_32_543 VPWR VGND sg13g2_decap_8
XFILLER_5_60 VPWR VGND sg13g2_decap_8
XFILLER_27_315 VPWR VGND sg13g2_decap_8
XFILLER_39_175 VPWR VGND sg13g2_decap_8
XFILLER_36_893 VPWR VGND sg13g2_decap_8
XFILLER_23_543 VPWR VGND sg13g2_decap_8
XFILLER_24_25 VPWR VGND sg13g2_decap_8
XFILLER_40_46 VPWR VGND sg13g2_decap_8
XFILLER_2_403 VPWR VGND sg13g2_decap_8
XFILLER_49_77 VPWR VGND sg13g2_decap_8
XFILLER_19_816 VPWR VGND sg13g2_decap_8
XFILLER_46_602 VPWR VGND sg13g2_decap_8
XFILLER_18_326 VPWR VGND sg13g2_decap_8
XFILLER_45_123 VPWR VGND sg13g2_decap_8
XFILLER_46_679 VPWR VGND sg13g2_decap_8
XFILLER_27_882 VPWR VGND sg13g2_decap_8
XFILLER_42_841 VPWR VGND sg13g2_decap_8
XFILLER_14_543 VPWR VGND sg13g2_decap_8
XFILLER_41_373 VPWR VGND sg13g2_decap_8
XFILLER_10_760 VPWR VGND sg13g2_decap_8
XFILLER_6_753 VPWR VGND sg13g2_decap_8
XFILLER_5_263 VPWR VGND sg13g2_decap_8
XFILLER_49_462 VPWR VGND sg13g2_decap_8
Xinput6 ui_in[5] net6 VPWR VGND sg13g2_buf_1
XFILLER_37_602 VPWR VGND sg13g2_decap_8
XFILLER_36_123 VPWR VGND sg13g2_decap_8
XFILLER_37_679 VPWR VGND sg13g2_decap_8
XFILLER_18_893 VPWR VGND sg13g2_decap_8
XFILLER_45_690 VPWR VGND sg13g2_decap_8
XFILLER_17_392 VPWR VGND sg13g2_decap_8
XFILLER_32_340 VPWR VGND sg13g2_decap_8
XFILLER_33_863 VPWR VGND sg13g2_decap_8
XFILLER_20_557 VPWR VGND sg13g2_decap_8
XFILLER_19_25 VPWR VGND sg13g2_decap_8
XFILLER_27_112 VPWR VGND sg13g2_decap_8
XFILLER_28_657 VPWR VGND sg13g2_decap_8
XFILLER_27_189 VPWR VGND sg13g2_decap_8
XFILLER_35_46 VPWR VGND sg13g2_decap_8
XFILLER_36_690 VPWR VGND sg13g2_decap_8
XFILLER_43_627 VPWR VGND sg13g2_decap_8
XFILLER_23_340 VPWR VGND sg13g2_decap_8
XFILLER_24_852 VPWR VGND sg13g2_decap_8
XFILLER_42_148 VPWR VGND sg13g2_decap_8
XFILLER_11_557 VPWR VGND sg13g2_decap_8
XFILLER_7_539 VPWR VGND sg13g2_decap_8
XFILLER_2_200 VPWR VGND sg13g2_decap_8
XFILLER_3_767 VPWR VGND sg13g2_decap_8
XFILLER_2_277 VPWR VGND sg13g2_decap_8
XFILLER_19_613 VPWR VGND sg13g2_decap_8
XFILLER_18_123 VPWR VGND sg13g2_decap_8
XFILLER_46_476 VPWR VGND sg13g2_decap_8
XFILLER_15_830 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_30 VPWR VGND uio_oe[5] sg13g2_tielo
XFILLER_14_340 VPWR VGND sg13g2_decap_8
XFILLER_25_90 VPWR VGND sg13g2_decap_8
XFILLER_30_800 VPWR VGND sg13g2_decap_8
XFILLER_41_170 VPWR VGND sg13g2_decap_8
XFILLER_30_877 VPWR VGND sg13g2_decap_8
XFILLER_6_550 VPWR VGND sg13g2_decap_8
XFILLER_38_922 VPWR VGND sg13g2_fill_2
XFILLER_37_476 VPWR VGND sg13g2_decap_8
X_58_ _24_ net7 net15 VPWR VGND sg13g2_nand2_1
XFILLER_18_690 VPWR VGND sg13g2_decap_8
XFILLER_24_159 VPWR VGND sg13g2_decap_8
XFILLER_33_660 VPWR VGND sg13g2_decap_8
XFILLER_21_844 VPWR VGND sg13g2_decap_8
XFILLER_20_354 VPWR VGND sg13g2_decap_8
XFILLER_29_922 VPWR VGND sg13g2_fill_2
XFILLER_46_56 VPWR VGND sg13g2_decap_8
XFILLER_28_454 VPWR VGND sg13g2_decap_8
XFILLER_44_914 VPWR VGND sg13g2_decap_8
XFILLER_16_627 VPWR VGND sg13g2_decap_8
XFILLER_43_424 VPWR VGND sg13g2_decap_8
XFILLER_15_137 VPWR VGND sg13g2_decap_8
XFILLER_31_619 VPWR VGND sg13g2_decap_8
XFILLER_12_844 VPWR VGND sg13g2_decap_8
XFILLER_11_354 VPWR VGND sg13g2_decap_8
XFILLER_8_837 VPWR VGND sg13g2_decap_8
XFILLER_7_28 VPWR VGND sg13g2_decap_8
XFILLER_7_336 VPWR VGND sg13g2_decap_8
XFILLER_11_81 VPWR VGND sg13g2_decap_8
XFILLER_3_564 VPWR VGND sg13g2_decap_8
XFILLER_19_410 VPWR VGND sg13g2_decap_8
XFILLER_38_229 VPWR VGND sg13g2_decap_8
XFILLER_47_763 VPWR VGND sg13g2_decap_8
XFILLER_46_273 VPWR VGND sg13g2_decap_8
XFILLER_19_487 VPWR VGND sg13g2_decap_8
XFILLER_34_468 VPWR VGND sg13g2_decap_8
XFILLER_30_674 VPWR VGND sg13g2_decap_8
XFILLER_29_229 VPWR VGND sg13g2_decap_8
XFILLER_26_914 VPWR VGND sg13g2_decap_8
XFILLER_37_273 VPWR VGND sg13g2_decap_8
XFILLER_38_796 VPWR VGND sg13g2_decap_8
XFILLER_25_468 VPWR VGND sg13g2_decap_8
XFILLER_40_438 VPWR VGND sg13g2_decap_8
XFILLER_21_641 VPWR VGND sg13g2_decap_8
XFILLER_32_25 VPWR VGND sg13g2_decap_8
XFILLER_20_151 VPWR VGND sg13g2_decap_8
XFILLER_0_567 VPWR VGND sg13g2_decap_8
XFILLER_17_903 VPWR VGND sg13g2_decap_8
XFILLER_16_424 VPWR VGND sg13g2_decap_8
XFILLER_28_251 VPWR VGND sg13g2_decap_8
XFILLER_29_796 VPWR VGND sg13g2_decap_8
XFILLER_44_711 VPWR VGND sg13g2_decap_8
XFILLER_43_221 VPWR VGND sg13g2_decap_8
XFILLER_31_416 VPWR VGND sg13g2_decap_8
XFILLER_44_788 VPWR VGND sg13g2_decap_8
XFILLER_43_298 VPWR VGND sg13g2_decap_8
XFILLER_12_641 VPWR VGND sg13g2_decap_8
XFILLER_11_151 VPWR VGND sg13g2_decap_8
XFILLER_8_634 VPWR VGND sg13g2_decap_8
XFILLER_7_133 VPWR VGND sg13g2_decap_8
XFILLER_4_851 VPWR VGND sg13g2_decap_8
XFILLER_3_361 VPWR VGND sg13g2_decap_8
XFILLER_14_4 VPWR VGND sg13g2_decap_8
XFILLER_47_560 VPWR VGND sg13g2_decap_8
XFILLER_19_284 VPWR VGND sg13g2_decap_8
XFILLER_35_744 VPWR VGND sg13g2_decap_8
XFILLER_34_265 VPWR VGND sg13g2_decap_8
XFILLER_22_438 VPWR VGND sg13g2_decap_8
XFILLER_8_60 VPWR VGND sg13g2_decap_8
XFILLER_30_471 VPWR VGND sg13g2_decap_8
XFILLER_27_14 VPWR VGND sg13g2_decap_8
XFILLER_45_508 VPWR VGND sg13g2_decap_8
XFILLER_26_711 VPWR VGND sg13g2_decap_8
XFILLER_38_593 VPWR VGND sg13g2_decap_8
XFILLER_25_265 VPWR VGND sg13g2_decap_8
XFILLER_26_788 VPWR VGND sg13g2_decap_8
XFILLER_13_438 VPWR VGND sg13g2_decap_8
XFILLER_40_235 VPWR VGND sg13g2_decap_8
XFILLER_41_758 VPWR VGND sg13g2_decap_8
XFILLER_43_46 VPWR VGND sg13g2_decap_8
XFILLER_5_648 VPWR VGND sg13g2_decap_8
XFILLER_4_158 VPWR VGND sg13g2_decap_8
XFILLER_4_18 VPWR VGND sg13g2_decap_8
XFILLER_1_854 VPWR VGND sg13g2_decap_8
XFILLER_0_364 VPWR VGND sg13g2_decap_8
XFILLER_49_847 VPWR VGND sg13g2_decap_8
XFILLER_48_357 VPWR VGND sg13g2_decap_8
XFILLER_36_508 VPWR VGND sg13g2_decap_8
XFILLER_17_700 VPWR VGND sg13g2_decap_8
XFILLER_16_221 VPWR VGND sg13g2_decap_8
XFILLER_29_593 VPWR VGND sg13g2_decap_8
XFILLER_17_91 VPWR VGND sg13g2_decap_8
XFILLER_17_777 VPWR VGND sg13g2_decap_8
XFILLER_32_725 VPWR VGND sg13g2_decap_8
XFILLER_16_298 VPWR VGND sg13g2_decap_8
XFILLER_31_213 VPWR VGND sg13g2_decap_8
XFILLER_44_585 VPWR VGND sg13g2_decap_8
XFILLER_9_921 VPWR VGND sg13g2_decap_4
XFILLER_8_431 VPWR VGND sg13g2_decap_8
XFILLER_39_357 VPWR VGND sg13g2_decap_8
XFILLER_35_541 VPWR VGND sg13g2_decap_8
XFILLER_23_725 VPWR VGND sg13g2_decap_8
XFILLER_22_235 VPWR VGND sg13g2_decap_8
XFILLER_31_780 VPWR VGND sg13g2_decap_8
XFILLER_18_508 VPWR VGND sg13g2_decap_8
XFILLER_38_68 VPWR VGND sg13g2_decap_8
XFILLER_45_305 VPWR VGND sg13g2_decap_8
XFILLER_38_390 VPWR VGND sg13g2_decap_8
XFILLER_14_725 VPWR VGND sg13g2_decap_8
XFILLER_26_585 VPWR VGND sg13g2_decap_8
XFILLER_13_235 VPWR VGND sg13g2_decap_8
XFILLER_41_555 VPWR VGND sg13g2_decap_8
XFILLER_9_228 VPWR VGND sg13g2_decap_8
XFILLER_5_445 VPWR VGND sg13g2_decap_8
XFILLER_1_651 VPWR VGND sg13g2_decap_8
XFILLER_0_161 VPWR VGND sg13g2_decap_8
XFILLER_49_644 VPWR VGND sg13g2_decap_8
XFILLER_48_154 VPWR VGND sg13g2_decap_8
XFILLER_36_305 VPWR VGND sg13g2_decap_8
XFILLER_29_390 VPWR VGND sg13g2_decap_8
XFILLER_45_872 VPWR VGND sg13g2_decap_8
XFILLER_17_574 VPWR VGND sg13g2_decap_8
XFILLER_32_522 VPWR VGND sg13g2_decap_8
XFILLER_44_382 VPWR VGND sg13g2_decap_8
XFILLER_20_739 VPWR VGND sg13g2_decap_8
XFILLER_32_599 VPWR VGND sg13g2_decap_8
XFILLER_9_795 VPWR VGND sg13g2_decap_8
XFILLER_28_839 VPWR VGND sg13g2_decap_8
XFILLER_39_154 VPWR VGND sg13g2_decap_8
XFILLER_43_809 VPWR VGND sg13g2_decap_8
XFILLER_36_872 VPWR VGND sg13g2_decap_8
XFILLER_23_522 VPWR VGND sg13g2_decap_8
XFILLER_11_739 VPWR VGND sg13g2_decap_8
XFILLER_23_599 VPWR VGND sg13g2_decap_8
XFILLER_10_249 VPWR VGND sg13g2_decap_8
XFILLER_40_25 VPWR VGND sg13g2_decap_8
XFILLER_2_459 VPWR VGND sg13g2_decap_8
XFILLER_49_56 VPWR VGND sg13g2_decap_8
XFILLER_18_305 VPWR VGND sg13g2_decap_8
XFILLER_45_102 VPWR VGND sg13g2_decap_8
XFILLER_46_658 VPWR VGND sg13g2_decap_8
XFILLER_27_861 VPWR VGND sg13g2_decap_8
XFILLER_14_522 VPWR VGND sg13g2_decap_8
XFILLER_26_382 VPWR VGND sg13g2_decap_8
XFILLER_42_820 VPWR VGND sg13g2_decap_8
XFILLER_45_179 VPWR VGND sg13g2_decap_8
XFILLER_14_599 VPWR VGND sg13g2_decap_8
XFILLER_41_352 VPWR VGND sg13g2_decap_8
XFILLER_42_897 VPWR VGND sg13g2_decap_8
XFILLER_14_81 VPWR VGND sg13g2_decap_8
XFILLER_6_732 VPWR VGND sg13g2_decap_8
XFILLER_5_242 VPWR VGND sg13g2_decap_8
XFILLER_46_7 VPWR VGND sg13g2_decap_8
XFILLER_49_441 VPWR VGND sg13g2_decap_8
Xinput7 ui_in[6] net7 VPWR VGND sg13g2_buf_1
XFILLER_36_102 VPWR VGND sg13g2_decap_8
XFILLER_37_658 VPWR VGND sg13g2_decap_8
XFILLER_18_872 VPWR VGND sg13g2_decap_8
XFILLER_17_371 VPWR VGND sg13g2_decap_8
XFILLER_36_179 VPWR VGND sg13g2_decap_8
XFILLER_33_842 VPWR VGND sg13g2_decap_8
XFILLER_20_536 VPWR VGND sg13g2_decap_8
XFILLER_32_396 VPWR VGND sg13g2_decap_8
XFILLER_9_592 VPWR VGND sg13g2_decap_8
XFILLER_10_39 VPWR VGND sg13g2_decap_8
XFILLER_28_636 VPWR VGND sg13g2_decap_8
XFILLER_16_809 VPWR VGND sg13g2_decap_8
XFILLER_27_168 VPWR VGND sg13g2_decap_8
XFILLER_35_25 VPWR VGND sg13g2_decap_8
XFILLER_43_606 VPWR VGND sg13g2_decap_8
XFILLER_15_319 VPWR VGND sg13g2_decap_8
XFILLER_24_831 VPWR VGND sg13g2_decap_8
XFILLER_42_127 VPWR VGND sg13g2_decap_8
XFILLER_11_536 VPWR VGND sg13g2_decap_8
XFILLER_23_396 VPWR VGND sg13g2_decap_8
XFILLER_7_518 VPWR VGND sg13g2_decap_8
XFILLER_3_746 VPWR VGND sg13g2_decap_8
XFILLER_2_256 VPWR VGND sg13g2_decap_8
XFILLER_18_102 VPWR VGND sg13g2_decap_8
XFILLER_46_455 VPWR VGND sg13g2_decap_8
XFILLER_19_669 VPWR VGND sg13g2_decap_8
XFILLER_18_179 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_31 VPWR VGND uio_oe[6] sg13g2_tielo
XFILLER_33_149 VPWR VGND sg13g2_decap_8
XFILLER_15_886 VPWR VGND sg13g2_decap_8
XFILLER_14_396 VPWR VGND sg13g2_decap_8
XFILLER_30_856 VPWR VGND sg13g2_decap_8
XFILLER_42_694 VPWR VGND sg13g2_decap_8
XFILLER_44_4 VPWR VGND sg13g2_decap_8
XFILLER_38_901 VPWR VGND sg13g2_decap_8
XFILLER_2_95 VPWR VGND sg13g2_decap_8
X_57_ VPWR VGND _21_ _22_ _13_ net6 _23_ net14 sg13g2_a221oi_1
XFILLER_37_455 VPWR VGND sg13g2_decap_8
XFILLER_24_138 VPWR VGND sg13g2_decap_8
XFILLER_21_823 VPWR VGND sg13g2_decap_8
XFILLER_20_333 VPWR VGND sg13g2_decap_8
XFILLER_32_193 VPWR VGND sg13g2_decap_8
XFILLER_0_749 VPWR VGND sg13g2_decap_8
XFILLER_29_901 VPWR VGND sg13g2_decap_8
XFILLER_28_433 VPWR VGND sg13g2_decap_8
XFILLER_46_35 VPWR VGND sg13g2_decap_8
XFILLER_16_606 VPWR VGND sg13g2_decap_8
XFILLER_15_116 VPWR VGND sg13g2_decap_8
XFILLER_43_403 VPWR VGND sg13g2_decap_8
XFILLER_12_823 VPWR VGND sg13g2_decap_8
XFILLER_11_333 VPWR VGND sg13g2_decap_8
XFILLER_8_816 VPWR VGND sg13g2_decap_8
XFILLER_7_315 VPWR VGND sg13g2_decap_8
XFILLER_23_193 VPWR VGND sg13g2_decap_8
XFILLER_11_60 VPWR VGND sg13g2_decap_8
XFILLER_3_543 VPWR VGND sg13g2_decap_8
XFILLER_38_208 VPWR VGND sg13g2_decap_8
XFILLER_47_742 VPWR VGND sg13g2_decap_8
XFILLER_19_466 VPWR VGND sg13g2_decap_8
XFILLER_46_252 VPWR VGND sg13g2_decap_8
XFILLER_34_447 VPWR VGND sg13g2_decap_8
XFILLER_15_683 VPWR VGND sg13g2_decap_8
XFILLER_42_491 VPWR VGND sg13g2_decap_8
XFILLER_14_193 VPWR VGND sg13g2_decap_8
XFILLER_30_653 VPWR VGND sg13g2_decap_8
Xinput10 uio_in[1] net10 VPWR VGND sg13g2_buf_1
XFILLER_7_882 VPWR VGND sg13g2_decap_8
XFILLER_29_208 VPWR VGND sg13g2_decap_8
XFILLER_38_775 VPWR VGND sg13g2_decap_8
XFILLER_37_252 VPWR VGND sg13g2_decap_8
XFILLER_25_447 VPWR VGND sg13g2_decap_8
XFILLER_40_417 VPWR VGND sg13g2_decap_8
XFILLER_21_620 VPWR VGND sg13g2_decap_8
XFILLER_20_130 VPWR VGND sg13g2_decap_8
XFILLER_21_697 VPWR VGND sg13g2_decap_8
XFILLER_0_546 VPWR VGND sg13g2_decap_8
XFILLER_48_539 VPWR VGND sg13g2_decap_8
XFILLER_28_230 VPWR VGND sg13g2_decap_8
XFILLER_16_403 VPWR VGND sg13g2_decap_8
XFILLER_29_775 VPWR VGND sg13g2_decap_8
XFILLER_43_200 VPWR VGND sg13g2_decap_8
XFILLER_32_907 VPWR VGND sg13g2_decap_8
XFILLER_44_767 VPWR VGND sg13g2_decap_8
XFILLER_43_277 VPWR VGND sg13g2_decap_8
XFILLER_12_620 VPWR VGND sg13g2_decap_8
XFILLER_11_130 VPWR VGND sg13g2_decap_8
XFILLER_8_613 VPWR VGND sg13g2_decap_8
XFILLER_7_112 VPWR VGND sg13g2_decap_8
XFILLER_12_697 VPWR VGND sg13g2_decap_8
XFILLER_7_189 VPWR VGND sg13g2_decap_8
XFILLER_22_81 VPWR VGND sg13g2_decap_8
XFILLER_4_830 VPWR VGND sg13g2_decap_8
XFILLER_3_340 VPWR VGND sg13g2_decap_8
XFILLER_39_539 VPWR VGND sg13g2_decap_8
XFILLER_19_263 VPWR VGND sg13g2_decap_8
XFILLER_35_723 VPWR VGND sg13g2_decap_8
XFILLER_23_907 VPWR VGND sg13g2_decap_8
XFILLER_22_417 VPWR VGND sg13g2_decap_8
XFILLER_34_244 VPWR VGND sg13g2_decap_8
XFILLER_15_480 VPWR VGND sg13g2_decap_8
XFILLER_30_450 VPWR VGND sg13g2_decap_8
XFILLER_38_572 VPWR VGND sg13g2_decap_8
XFILLER_14_907 VPWR VGND sg13g2_decap_8
XFILLER_25_244 VPWR VGND sg13g2_decap_8
XFILLER_26_767 VPWR VGND sg13g2_decap_8
XFILLER_13_417 VPWR VGND sg13g2_decap_8
XFILLER_40_214 VPWR VGND sg13g2_decap_8
XFILLER_41_737 VPWR VGND sg13g2_decap_8
XFILLER_43_25 VPWR VGND sg13g2_decap_8
XFILLER_21_494 VPWR VGND sg13g2_decap_8
XFILLER_5_627 VPWR VGND sg13g2_decap_8
XFILLER_4_137 VPWR VGND sg13g2_decap_8
XFILLER_1_833 VPWR VGND sg13g2_decap_8
XFILLER_0_343 VPWR VGND sg13g2_decap_8
XFILLER_49_826 VPWR VGND sg13g2_decap_8
XFILLER_48_336 VPWR VGND sg13g2_decap_8
XFILLER_29_572 VPWR VGND sg13g2_decap_8
XFILLER_16_200 VPWR VGND sg13g2_decap_8
XFILLER_17_756 VPWR VGND sg13g2_decap_8
XFILLER_17_70 VPWR VGND sg13g2_decap_8
XFILLER_32_704 VPWR VGND sg13g2_decap_8
XFILLER_44_564 VPWR VGND sg13g2_decap_8
XFILLER_16_277 VPWR VGND sg13g2_decap_8
XFILLER_9_900 VPWR VGND sg13g2_decap_8
XFILLER_8_410 VPWR VGND sg13g2_decap_8
XFILLER_31_269 VPWR VGND sg13g2_decap_8
XFILLER_40_781 VPWR VGND sg13g2_decap_8
XFILLER_12_494 VPWR VGND sg13g2_decap_8
XFILLER_8_487 VPWR VGND sg13g2_decap_8
XFILLER_39_336 VPWR VGND sg13g2_decap_8
XFILLER_35_520 VPWR VGND sg13g2_decap_8
XFILLER_23_704 VPWR VGND sg13g2_decap_8
XFILLER_22_214 VPWR VGND sg13g2_decap_8
XFILLER_35_597 VPWR VGND sg13g2_decap_8
XFILLER_13_39 VPWR VGND sg13g2_decap_8
XFILLER_38_47 VPWR VGND sg13g2_decap_8
XFILLER_14_704 VPWR VGND sg13g2_decap_8
XFILLER_26_564 VPWR VGND sg13g2_decap_8
XFILLER_13_214 VPWR VGND sg13g2_decap_8
XFILLER_41_534 VPWR VGND sg13g2_decap_8
XFILLER_9_207 VPWR VGND sg13g2_decap_8
XFILLER_10_921 VPWR VGND sg13g2_decap_4
XFILLER_22_781 VPWR VGND sg13g2_decap_8
XFILLER_21_291 VPWR VGND sg13g2_decap_8
XFILLER_6_914 VPWR VGND sg13g2_decap_8
XFILLER_5_424 VPWR VGND sg13g2_decap_8
XFILLER_1_630 VPWR VGND sg13g2_decap_8
XFILLER_49_623 VPWR VGND sg13g2_decap_8
XFILLER_0_140 VPWR VGND sg13g2_decap_8
XFILLER_48_133 VPWR VGND sg13g2_decap_8
XFILLER_17_553 VPWR VGND sg13g2_decap_8
XFILLER_45_851 VPWR VGND sg13g2_decap_8
XFILLER_32_501 VPWR VGND sg13g2_decap_8
XFILLER_44_361 VPWR VGND sg13g2_decap_8
XFILLER_20_718 VPWR VGND sg13g2_decap_8
XFILLER_32_578 VPWR VGND sg13g2_decap_8
XFILLER_13_781 VPWR VGND sg13g2_decap_8
XFILLER_9_774 VPWR VGND sg13g2_decap_8
XFILLER_12_291 VPWR VGND sg13g2_decap_8
XFILLER_8_284 VPWR VGND sg13g2_decap_8
XFILLER_5_95 VPWR VGND sg13g2_decap_8
XFILLER_39_133 VPWR VGND sg13g2_decap_8
XFILLER_28_818 VPWR VGND sg13g2_decap_8
XFILLER_36_851 VPWR VGND sg13g2_decap_8
XFILLER_42_309 VPWR VGND sg13g2_decap_8
XFILLER_23_501 VPWR VGND sg13g2_decap_8
XFILLER_35_394 VPWR VGND sg13g2_decap_8
XFILLER_11_718 VPWR VGND sg13g2_decap_8
XFILLER_23_578 VPWR VGND sg13g2_decap_8
XFILLER_10_228 VPWR VGND sg13g2_decap_8
XFILLER_2_438 VPWR VGND sg13g2_decap_8
XFILLER_49_35 VPWR VGND sg13g2_decap_8
XFILLER_46_637 VPWR VGND sg13g2_decap_8
XFILLER_27_840 VPWR VGND sg13g2_decap_8
XFILLER_45_158 VPWR VGND sg13g2_decap_8
XFILLER_14_501 VPWR VGND sg13g2_decap_8
XFILLER_26_361 VPWR VGND sg13g2_decap_8
XFILLER_41_331 VPWR VGND sg13g2_decap_8
XFILLER_14_578 VPWR VGND sg13g2_decap_8
XFILLER_42_876 VPWR VGND sg13g2_decap_8
XFILLER_14_60 VPWR VGND sg13g2_decap_8
XFILLER_6_711 VPWR VGND sg13g2_decap_8
XFILLER_10_795 VPWR VGND sg13g2_decap_8
XFILLER_5_221 VPWR VGND sg13g2_decap_8
XFILLER_6_788 VPWR VGND sg13g2_decap_8
XFILLER_5_298 VPWR VGND sg13g2_decap_8
XFILLER_49_420 VPWR VGND sg13g2_decap_8
Xinput8 ui_in[7] net8 VPWR VGND sg13g2_buf_1
XFILLER_49_497 VPWR VGND sg13g2_decap_8
XFILLER_37_637 VPWR VGND sg13g2_decap_8
XFILLER_18_851 VPWR VGND sg13g2_decap_8
XFILLER_36_158 VPWR VGND sg13g2_decap_8
XFILLER_17_350 VPWR VGND sg13g2_decap_8
XFILLER_33_821 VPWR VGND sg13g2_decap_8
XFILLER_20_515 VPWR VGND sg13g2_decap_8
XFILLER_32_375 VPWR VGND sg13g2_decap_8
XFILLER_33_898 VPWR VGND sg13g2_decap_8
XFILLER_9_571 VPWR VGND sg13g2_decap_8
XFILLER_10_18 VPWR VGND sg13g2_decap_8
XFILLER_28_615 VPWR VGND sg13g2_decap_8
XFILLER_27_147 VPWR VGND sg13g2_decap_8
XFILLER_24_810 VPWR VGND sg13g2_decap_8
XFILLER_42_106 VPWR VGND sg13g2_decap_8
XFILLER_35_191 VPWR VGND sg13g2_decap_8
XFILLER_11_515 VPWR VGND sg13g2_decap_8
XFILLER_23_375 VPWR VGND sg13g2_decap_8
XFILLER_24_887 VPWR VGND sg13g2_decap_8
XFILLER_3_725 VPWR VGND sg13g2_decap_8
XFILLER_4_4 VPWR VGND sg13g2_decap_8
XFILLER_2_235 VPWR VGND sg13g2_decap_8
XFILLER_47_924 VPWR VGND sg13g2_fill_1
XFILLER_46_434 VPWR VGND sg13g2_decap_8
XFILLER_19_648 VPWR VGND sg13g2_decap_8
XFILLER_18_158 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_32 VPWR VGND uio_oe[7] sg13g2_tielo
XFILLER_34_629 VPWR VGND sg13g2_decap_8
XFILLER_33_128 VPWR VGND sg13g2_decap_8
XFILLER_15_865 VPWR VGND sg13g2_decap_8
XFILLER_42_673 VPWR VGND sg13g2_decap_8
XFILLER_14_375 VPWR VGND sg13g2_decap_8
XFILLER_30_835 VPWR VGND sg13g2_decap_8
XFILLER_10_592 VPWR VGND sg13g2_decap_8
XFILLER_6_585 VPWR VGND sg13g2_decap_8
XFILLER_38_924 VPWR VGND sg13g2_fill_1
XFILLER_2_74 VPWR VGND sg13g2_decap_8
XFILLER_37_434 VPWR VGND sg13g2_decap_8
XFILLER_49_294 VPWR VGND sg13g2_decap_8
X_56_ _14_ _18_ _22_ VPWR VGND sg13g2_nor2_1
XFILLER_24_117 VPWR VGND sg13g2_decap_8
XFILLER_25_629 VPWR VGND sg13g2_decap_8
XFILLER_21_802 VPWR VGND sg13g2_decap_8
XFILLER_20_312 VPWR VGND sg13g2_decap_8
XFILLER_32_172 VPWR VGND sg13g2_decap_8
XFILLER_33_695 VPWR VGND sg13g2_decap_8
XFILLER_21_879 VPWR VGND sg13g2_decap_8
XFILLER_20_389 VPWR VGND sg13g2_decap_8
XFILLER_21_39 VPWR VGND sg13g2_decap_8
XFILLER_0_728 VPWR VGND sg13g2_decap_8
XFILLER_46_14 VPWR VGND sg13g2_decap_8
XFILLER_28_412 VPWR VGND sg13g2_decap_8
XFILLER_29_924 VPWR VGND sg13g2_fill_1
XFILLER_28_489 VPWR VGND sg13g2_decap_8
XFILLER_43_459 VPWR VGND sg13g2_decap_8
XFILLER_12_802 VPWR VGND sg13g2_decap_8
XFILLER_11_312 VPWR VGND sg13g2_decap_8
XFILLER_23_172 VPWR VGND sg13g2_decap_8
XFILLER_24_684 VPWR VGND sg13g2_decap_8
XFILLER_12_879 VPWR VGND sg13g2_decap_8
XFILLER_11_389 VPWR VGND sg13g2_decap_8
XFILLER_3_522 VPWR VGND sg13g2_decap_8
XFILLER_3_599 VPWR VGND sg13g2_decap_8
XFILLER_47_721 VPWR VGND sg13g2_decap_8
XFILLER_46_231 VPWR VGND sg13g2_decap_8
XFILLER_19_445 VPWR VGND sg13g2_decap_8
XFILLER_35_905 VPWR VGND sg13g2_decap_8
XFILLER_47_798 VPWR VGND sg13g2_decap_8
XFILLER_34_426 VPWR VGND sg13g2_decap_8
XFILLER_15_662 VPWR VGND sg13g2_decap_8
XFILLER_21_109 VPWR VGND sg13g2_decap_8
XFILLER_14_172 VPWR VGND sg13g2_decap_8
XFILLER_30_632 VPWR VGND sg13g2_decap_8
XFILLER_42_470 VPWR VGND sg13g2_decap_8
Xinput11 uio_in[2] net11 VPWR VGND sg13g2_buf_1
XFILLER_7_861 VPWR VGND sg13g2_decap_8
XFILLER_6_382 VPWR VGND sg13g2_decap_8
XFILLER_37_231 VPWR VGND sg13g2_decap_8
XFILLER_38_754 VPWR VGND sg13g2_decap_8
X_39_ net4 net12 _08_ VPWR VGND sg13g2_and2_1
XFILLER_16_39 VPWR VGND sg13g2_decap_8
XFILLER_25_426 VPWR VGND sg13g2_decap_8
XFILLER_12_109 VPWR VGND sg13g2_decap_8
XFILLER_41_919 VPWR VGND sg13g2_decap_4
XFILLER_33_492 VPWR VGND sg13g2_decap_8
XFILLER_21_676 VPWR VGND sg13g2_decap_8
XFILLER_5_809 VPWR VGND sg13g2_decap_8
XFILLER_20_186 VPWR VGND sg13g2_decap_8
XFILLER_4_319 VPWR VGND sg13g2_decap_8
XFILLER_0_525 VPWR VGND sg13g2_decap_8
XFILLER_48_518 VPWR VGND sg13g2_decap_8
XFILLER_29_754 VPWR VGND sg13g2_decap_8
XFILLER_28_286 VPWR VGND sg13g2_decap_8
XFILLER_44_746 VPWR VGND sg13g2_decap_8
XFILLER_16_459 VPWR VGND sg13g2_decap_8
XFILLER_43_256 VPWR VGND sg13g2_decap_8
XFILLER_24_481 VPWR VGND sg13g2_decap_8
XFILLER_12_676 VPWR VGND sg13g2_decap_8
XFILLER_11_186 VPWR VGND sg13g2_decap_8
XFILLER_8_669 VPWR VGND sg13g2_decap_8
XFILLER_22_60 VPWR VGND sg13g2_decap_8
XFILLER_7_168 VPWR VGND sg13g2_decap_8
XFILLER_4_886 VPWR VGND sg13g2_decap_8
XFILLER_3_396 VPWR VGND sg13g2_decap_8
XFILLER_39_518 VPWR VGND sg13g2_decap_8
XFILLER_19_242 VPWR VGND sg13g2_decap_8
XFILLER_35_702 VPWR VGND sg13g2_decap_8
XFILLER_47_595 VPWR VGND sg13g2_decap_8
XFILLER_34_223 VPWR VGND sg13g2_decap_8
XFILLER_35_779 VPWR VGND sg13g2_decap_8
XFILLER_8_95 VPWR VGND sg13g2_decap_8
XFILLER_27_49 VPWR VGND sg13g2_decap_8
XFILLER_38_551 VPWR VGND sg13g2_decap_8
XFILLER_25_223 VPWR VGND sg13g2_decap_8
XFILLER_26_746 VPWR VGND sg13g2_decap_8
XFILLER_41_716 VPWR VGND sg13g2_decap_8
XFILLER_34_790 VPWR VGND sg13g2_decap_8
XFILLER_21_473 VPWR VGND sg13g2_decap_8
XFILLER_5_606 VPWR VGND sg13g2_decap_8
XFILLER_4_116 VPWR VGND sg13g2_decap_8
XFILLER_1_812 VPWR VGND sg13g2_decap_8
XFILLER_49_805 VPWR VGND sg13g2_decap_8
XFILLER_0_322 VPWR VGND sg13g2_decap_8
XFILLER_48_315 VPWR VGND sg13g2_decap_8
XFILLER_1_889 VPWR VGND sg13g2_decap_8
XFILLER_0_399 VPWR VGND sg13g2_decap_8
XFILLER_29_551 VPWR VGND sg13g2_decap_8
XFILLER_17_735 VPWR VGND sg13g2_decap_8
XFILLER_16_256 VPWR VGND sg13g2_decap_8
XFILLER_44_543 VPWR VGND sg13g2_decap_8
XFILLER_25_790 VPWR VGND sg13g2_decap_8
XFILLER_31_248 VPWR VGND sg13g2_decap_8
XFILLER_12_473 VPWR VGND sg13g2_decap_8
XFILLER_40_760 VPWR VGND sg13g2_decap_8
XFILLER_8_466 VPWR VGND sg13g2_decap_8
XFILLER_4_683 VPWR VGND sg13g2_decap_8
XFILLER_3_193 VPWR VGND sg13g2_decap_8
XFILLER_39_315 VPWR VGND sg13g2_decap_8
XFILLER_48_882 VPWR VGND sg13g2_decap_8
XFILLER_47_392 VPWR VGND sg13g2_decap_8
XFILLER_35_576 VPWR VGND sg13g2_decap_8
XFILLER_13_18 VPWR VGND sg13g2_decap_8
XFILLER_1_119 VPWR VGND sg13g2_decap_8
XFILLER_38_15 VPWR VGND sg13g2_fill_2
XFILLER_46_819 VPWR VGND sg13g2_decap_8
XFILLER_39_882 VPWR VGND sg13g2_decap_8
XFILLER_26_543 VPWR VGND sg13g2_decap_8
XFILLER_41_513 VPWR VGND sg13g2_decap_8
XFILLER_10_900 VPWR VGND sg13g2_decap_8
XFILLER_22_760 VPWR VGND sg13g2_decap_8
XFILLER_21_270 VPWR VGND sg13g2_decap_8
XFILLER_5_403 VPWR VGND sg13g2_decap_8
XFILLER_49_602 VPWR VGND sg13g2_decap_8
XFILLER_1_686 VPWR VGND sg13g2_decap_8
XFILLER_48_112 VPWR VGND sg13g2_decap_8
XFILLER_0_196 VPWR VGND sg13g2_decap_8
XFILLER_49_679 VPWR VGND sg13g2_decap_8
XFILLER_37_819 VPWR VGND sg13g2_decap_8
XFILLER_48_189 VPWR VGND sg13g2_decap_8
XFILLER_28_81 VPWR VGND sg13g2_decap_8
XFILLER_45_830 VPWR VGND sg13g2_decap_8
XFILLER_17_532 VPWR VGND sg13g2_decap_8
XFILLER_44_340 VPWR VGND sg13g2_decap_8
XFILLER_32_557 VPWR VGND sg13g2_decap_8
XFILLER_13_760 VPWR VGND sg13g2_decap_8
XFILLER_9_753 VPWR VGND sg13g2_decap_8
XFILLER_12_270 VPWR VGND sg13g2_decap_8
XFILLER_8_263 VPWR VGND sg13g2_decap_8
XFILLER_5_74 VPWR VGND sg13g2_decap_8
XFILLER_4_480 VPWR VGND sg13g2_decap_8
XFILLER_39_112 VPWR VGND sg13g2_decap_8
XFILLER_27_329 VPWR VGND sg13g2_decap_8
XFILLER_36_830 VPWR VGND sg13g2_decap_8
XFILLER_39_189 VPWR VGND sg13g2_decap_8
XFILLER_35_373 VPWR VGND sg13g2_decap_8
XFILLER_23_557 VPWR VGND sg13g2_decap_8
XFILLER_24_39 VPWR VGND sg13g2_decap_8
XFILLER_10_207 VPWR VGND sg13g2_decap_8
XFILLER_3_907 VPWR VGND sg13g2_decap_8
XFILLER_2_417 VPWR VGND sg13g2_decap_8
XFILLER_49_14 VPWR VGND sg13g2_decap_8
XFILLER_46_616 VPWR VGND sg13g2_decap_8
XFILLER_26_340 VPWR VGND sg13g2_decap_8
XFILLER_45_137 VPWR VGND sg13g2_decap_8
XFILLER_27_896 VPWR VGND sg13g2_decap_8
XFILLER_14_557 VPWR VGND sg13g2_decap_8
XFILLER_41_310 VPWR VGND sg13g2_decap_8
XFILLER_42_855 VPWR VGND sg13g2_decap_8
XFILLER_41_387 VPWR VGND sg13g2_decap_8
XFILLER_10_774 VPWR VGND sg13g2_decap_8
XFILLER_5_200 VPWR VGND sg13g2_decap_8
XFILLER_6_767 VPWR VGND sg13g2_decap_8
XFILLER_5_277 VPWR VGND sg13g2_decap_8
XFILLER_30_82 VPWR VGND sg13g2_decap_8
XFILLER_1_483 VPWR VGND sg13g2_decap_8
XFILLER_49_476 VPWR VGND sg13g2_decap_8
XFILLER_37_616 VPWR VGND sg13g2_decap_8
XFILLER_39_91 VPWR VGND sg13g2_decap_8
XFILLER_18_830 VPWR VGND sg13g2_decap_8
Xinput9 uio_in[0] net9 VPWR VGND sg13g2_buf_1
XFILLER_36_137 VPWR VGND sg13g2_decap_8
XFILLER_33_800 VPWR VGND sg13g2_decap_8
XFILLER_32_354 VPWR VGND sg13g2_decap_8
XFILLER_33_877 VPWR VGND sg13g2_decap_8
XFILLER_9_550 VPWR VGND sg13g2_decap_8
XFILLER_19_39 VPWR VGND sg13g2_decap_8
XFILLER_27_126 VPWR VGND sg13g2_decap_8
XFILLER_35_170 VPWR VGND sg13g2_decap_8
XFILLER_23_354 VPWR VGND sg13g2_decap_8
XFILLER_24_866 VPWR VGND sg13g2_decap_8
XFILLER_3_704 VPWR VGND sg13g2_decap_8
XFILLER_2_214 VPWR VGND sg13g2_decap_8
XFILLER_47_903 VPWR VGND sg13g2_decap_8
XFILLER_46_413 VPWR VGND sg13g2_decap_8
XFILLER_19_627 VPWR VGND sg13g2_decap_8
XFILLER_18_137 VPWR VGND sg13g2_decap_8
XFILLER_34_608 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_33 VPWR VGND uio_out[0] sg13g2_tielo
XFILLER_33_107 VPWR VGND sg13g2_fill_2
XFILLER_15_844 VPWR VGND sg13g2_decap_8
XFILLER_27_693 VPWR VGND sg13g2_decap_8
XFILLER_14_354 VPWR VGND sg13g2_decap_8
XFILLER_25_60 VPWR VGND sg13g2_decap_8
XFILLER_30_814 VPWR VGND sg13g2_decap_8
XFILLER_42_652 VPWR VGND sg13g2_decap_8
XFILLER_41_184 VPWR VGND sg13g2_decap_8
XFILLER_10_571 VPWR VGND sg13g2_decap_8
XFILLER_6_564 VPWR VGND sg13g2_decap_8
XFILLER_2_781 VPWR VGND sg13g2_decap_8
XFILLER_1_280 VPWR VGND sg13g2_decap_8
XFILLER_2_53 VPWR VGND sg13g2_decap_8
XFILLER_49_273 VPWR VGND sg13g2_decap_8
XFILLER_37_413 VPWR VGND sg13g2_decap_8
X_55_ _16_ _19_ _21_ VPWR VGND sg13g2_nor2_1
XFILLER_25_608 VPWR VGND sg13g2_decap_8
XFILLER_33_674 VPWR VGND sg13g2_decap_8
XFILLER_32_151 VPWR VGND sg13g2_decap_8
XFILLER_21_858 VPWR VGND sg13g2_decap_8
XFILLER_20_368 VPWR VGND sg13g2_decap_8
XFILLER_21_18 VPWR VGND sg13g2_decap_8
XFILLER_0_707 VPWR VGND sg13g2_decap_8
XFILLER_28_468 VPWR VGND sg13g2_decap_8
XFILLER_43_438 VPWR VGND sg13g2_decap_8
XFILLER_24_663 VPWR VGND sg13g2_decap_8
XFILLER_23_151 VPWR VGND sg13g2_decap_8
XFILLER_12_858 VPWR VGND sg13g2_decap_8
XFILLER_11_368 VPWR VGND sg13g2_decap_8
XFILLER_3_501 VPWR VGND sg13g2_decap_8
XFILLER_11_95 VPWR VGND sg13g2_decap_8
XFILLER_3_578 VPWR VGND sg13g2_decap_8
XFILLER_47_700 VPWR VGND sg13g2_decap_8
XFILLER_46_210 VPWR VGND sg13g2_decap_8
XFILLER_19_424 VPWR VGND sg13g2_decap_8
XFILLER_47_777 VPWR VGND sg13g2_decap_8
XFILLER_34_405 VPWR VGND sg13g2_decap_8
XFILLER_46_287 VPWR VGND sg13g2_decap_8
XFILLER_27_490 VPWR VGND sg13g2_decap_8
XFILLER_36_81 VPWR VGND sg13g2_decap_8
XFILLER_15_641 VPWR VGND sg13g2_decap_8
XFILLER_14_151 VPWR VGND sg13g2_decap_8
XFILLER_30_611 VPWR VGND sg13g2_decap_8
XFILLER_30_688 VPWR VGND sg13g2_decap_8
Xinput12 uio_in[3] net12 VPWR VGND sg13g2_buf_1
XFILLER_7_840 VPWR VGND sg13g2_decap_8
XFILLER_6_361 VPWR VGND sg13g2_decap_8
XFILLER_37_210 VPWR VGND sg13g2_decap_8
XFILLER_38_733 VPWR VGND sg13g2_decap_8
XFILLER_25_405 VPWR VGND sg13g2_decap_8
X_38_ VGND VPWR _07_ net12 net4 sg13g2_or2_1
XFILLER_16_18 VPWR VGND sg13g2_decap_8
XFILLER_37_287 VPWR VGND sg13g2_decap_8
XFILLER_33_471 VPWR VGND sg13g2_decap_8
XFILLER_21_655 VPWR VGND sg13g2_decap_8
XFILLER_20_165 VPWR VGND sg13g2_decap_8
XFILLER_32_39 VPWR VGND sg13g2_decap_8
XFILLER_0_504 VPWR VGND sg13g2_decap_8
XFILLER_29_733 VPWR VGND sg13g2_decap_8
XFILLER_17_917 VPWR VGND sg13g2_decap_8
XFILLER_28_265 VPWR VGND sg13g2_decap_8
XFILLER_16_438 VPWR VGND sg13g2_decap_8
XFILLER_44_725 VPWR VGND sg13g2_decap_8
XFILLER_43_235 VPWR VGND sg13g2_decap_8
XFILLER_24_460 VPWR VGND sg13g2_decap_8
XFILLER_12_655 VPWR VGND sg13g2_decap_8
XFILLER_11_165 VPWR VGND sg13g2_decap_8
XFILLER_8_648 VPWR VGND sg13g2_decap_8
XFILLER_7_147 VPWR VGND sg13g2_decap_8
XFILLER_4_865 VPWR VGND sg13g2_decap_8
XFILLER_3_375 VPWR VGND sg13g2_decap_8
XFILLER_19_221 VPWR VGND sg13g2_decap_8
XFILLER_47_574 VPWR VGND sg13g2_decap_8
XFILLER_47_91 VPWR VGND sg13g2_decap_8
XFILLER_19_298 VPWR VGND sg13g2_decap_8
XFILLER_34_202 VPWR VGND sg13g2_decap_8
XFILLER_35_758 VPWR VGND sg13g2_decap_8
XFILLER_31_920 VPWR VGND sg13g2_decap_4
XFILLER_34_279 VPWR VGND sg13g2_decap_8
XFILLER_8_74 VPWR VGND sg13g2_decap_8
XFILLER_30_485 VPWR VGND sg13g2_decap_8
XFILLER_38_530 VPWR VGND sg13g2_decap_8
XFILLER_27_28 VPWR VGND sg13g2_decap_8
XFILLER_25_202 VPWR VGND sg13g2_decap_8
XFILLER_26_725 VPWR VGND sg13g2_decap_8
XFILLER_25_279 VPWR VGND sg13g2_decap_8
XFILLER_40_249 VPWR VGND sg13g2_decap_8
XFILLER_21_452 VPWR VGND sg13g2_decap_8
XFILLER_0_301 VPWR VGND sg13g2_decap_8
XFILLER_1_868 VPWR VGND sg13g2_decap_8
XFILLER_0_378 VPWR VGND sg13g2_decap_8
XFILLER_29_530 VPWR VGND sg13g2_decap_8
XFILLER_17_714 VPWR VGND sg13g2_decap_8
XFILLER_44_522 VPWR VGND sg13g2_decap_8
XFILLER_16_235 VPWR VGND sg13g2_decap_8
XFILLER_32_739 VPWR VGND sg13g2_decap_8
XFILLER_44_599 VPWR VGND sg13g2_decap_8
XFILLER_31_227 VPWR VGND sg13g2_decap_8
XFILLER_12_452 VPWR VGND sg13g2_decap_8
XFILLER_8_445 VPWR VGND sg13g2_decap_8
XFILLER_33_93 VPWR VGND sg13g2_decap_8
XFILLER_4_662 VPWR VGND sg13g2_decap_8
XFILLER_3_172 VPWR VGND sg13g2_decap_8
XFILLER_12_4 VPWR VGND sg13g2_decap_8
XFILLER_48_861 VPWR VGND sg13g2_decap_8
XFILLER_47_371 VPWR VGND sg13g2_decap_8
XFILLER_35_555 VPWR VGND sg13g2_decap_8
XFILLER_23_739 VPWR VGND sg13g2_decap_8
XFILLER_22_249 VPWR VGND sg13g2_decap_8
XFILLER_30_282 VPWR VGND sg13g2_decap_8
XFILLER_31_794 VPWR VGND sg13g2_decap_8
XFILLER_39_861 VPWR VGND sg13g2_decap_8
XFILLER_26_522 VPWR VGND sg13g2_decap_8
XFILLER_45_319 VPWR VGND sg13g2_decap_8
XFILLER_14_739 VPWR VGND sg13g2_decap_8
XFILLER_26_599 VPWR VGND sg13g2_decap_8
XFILLER_13_249 VPWR VGND sg13g2_decap_8
XFILLER_41_569 VPWR VGND sg13g2_decap_8
XFILLER_5_459 VPWR VGND sg13g2_decap_8
XFILLER_1_665 VPWR VGND sg13g2_decap_8
XFILLER_49_658 VPWR VGND sg13g2_decap_8
XFILLER_0_175 VPWR VGND sg13g2_decap_8
XFILLER_48_168 VPWR VGND sg13g2_decap_8
XFILLER_17_511 VPWR VGND sg13g2_decap_8
XFILLER_28_60 VPWR VGND sg13g2_decap_8
XFILLER_36_319 VPWR VGND sg13g2_decap_8
XFILLER_45_886 VPWR VGND sg13g2_decap_8
XFILLER_17_588 VPWR VGND sg13g2_decap_8
XFILLER_32_536 VPWR VGND sg13g2_decap_8
XFILLER_44_396 VPWR VGND sg13g2_decap_8
XFILLER_44_81 VPWR VGND sg13g2_decap_8
XFILLER_9_732 VPWR VGND sg13g2_decap_8
XFILLER_8_242 VPWR VGND sg13g2_decap_8
XFILLER_5_53 VPWR VGND sg13g2_decap_8
XFILLER_27_308 VPWR VGND sg13g2_decap_8
XFILLER_39_168 VPWR VGND sg13g2_decap_8
XFILLER_35_352 VPWR VGND sg13g2_decap_8
XFILLER_36_886 VPWR VGND sg13g2_decap_8
XFILLER_23_536 VPWR VGND sg13g2_decap_8
XFILLER_24_18 VPWR VGND sg13g2_decap_8
XFILLER_31_591 VPWR VGND sg13g2_decap_8
XFILLER_40_39 VPWR VGND sg13g2_decap_8
XFILLER_19_809 VPWR VGND sg13g2_decap_8
XFILLER_18_319 VPWR VGND sg13g2_decap_8
XFILLER_45_116 VPWR VGND sg13g2_decap_8
XFILLER_27_875 VPWR VGND sg13g2_decap_8
XFILLER_14_536 VPWR VGND sg13g2_decap_8
XFILLER_26_396 VPWR VGND sg13g2_decap_8
XFILLER_42_834 VPWR VGND sg13g2_decap_8
XFILLER_41_366 VPWR VGND sg13g2_decap_8
XFILLER_10_753 VPWR VGND sg13g2_decap_8
XFILLER_14_95 VPWR VGND sg13g2_decap_8
XFILLER_6_746 VPWR VGND sg13g2_decap_8
XFILLER_5_256 VPWR VGND sg13g2_decap_8
XFILLER_30_61 VPWR VGND sg13g2_decap_8
XFILLER_1_462 VPWR VGND sg13g2_decap_8
XFILLER_49_455 VPWR VGND sg13g2_decap_8
XFILLER_39_70 VPWR VGND sg13g2_decap_8
XFILLER_36_116 VPWR VGND sg13g2_decap_8
XFILLER_18_886 VPWR VGND sg13g2_decap_8
XFILLER_17_385 VPWR VGND sg13g2_decap_8
XFILLER_33_856 VPWR VGND sg13g2_decap_8
XFILLER_45_683 VPWR VGND sg13g2_decap_8
XFILLER_32_333 VPWR VGND sg13g2_decap_8
XFILLER_44_193 VPWR VGND sg13g2_decap_8
XFILLER_19_18 VPWR VGND sg13g2_decap_8
XFILLER_27_105 VPWR VGND sg13g2_decap_8
XFILLER_35_39 VPWR VGND sg13g2_decap_8
XFILLER_24_845 VPWR VGND sg13g2_decap_8
XFILLER_36_683 VPWR VGND sg13g2_decap_8
XFILLER_23_333 VPWR VGND sg13g2_decap_8
XFILLER_19_606 VPWR VGND sg13g2_decap_8
XFILLER_18_116 VPWR VGND sg13g2_decap_8
XFILLER_46_469 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_34 VPWR VGND uio_out[1] sg13g2_tielo
XFILLER_27_672 VPWR VGND sg13g2_decap_8
XFILLER_15_823 VPWR VGND sg13g2_decap_8
XFILLER_42_631 VPWR VGND sg13g2_decap_8
XFILLER_14_333 VPWR VGND sg13g2_decap_8
XFILLER_26_193 VPWR VGND sg13g2_decap_8
XFILLER_41_163 VPWR VGND sg13g2_decap_8
XFILLER_10_550 VPWR VGND sg13g2_decap_8
XFILLER_6_543 VPWR VGND sg13g2_decap_8
XFILLER_41_93 VPWR VGND sg13g2_decap_8
XFILLER_2_760 VPWR VGND sg13g2_decap_8
XFILLER_2_32 VPWR VGND sg13g2_decap_8
XFILLER_38_915 VPWR VGND sg13g2_decap_8
XFILLER_49_252 VPWR VGND sg13g2_decap_8
X_54_ net22 _19_ _20_ VPWR VGND sg13g2_xnor2_1
XFILLER_37_469 VPWR VGND sg13g2_decap_8
XFILLER_17_182 VPWR VGND sg13g2_decap_8
XFILLER_18_683 VPWR VGND sg13g2_decap_8
XFILLER_45_480 VPWR VGND sg13g2_decap_8
XFILLER_32_130 VPWR VGND sg13g2_decap_8
XFILLER_33_653 VPWR VGND sg13g2_decap_8
XFILLER_21_837 VPWR VGND sg13g2_decap_8
XFILLER_20_347 VPWR VGND sg13g2_decap_8
XFILLER_29_915 VPWR VGND sg13g2_decap_8
XFILLER_46_49 VPWR VGND sg13g2_decap_8
XFILLER_28_447 VPWR VGND sg13g2_decap_8
XFILLER_44_907 VPWR VGND sg13g2_decap_8
XFILLER_43_417 VPWR VGND sg13g2_decap_8
XFILLER_36_480 VPWR VGND sg13g2_decap_8
XFILLER_23_130 VPWR VGND sg13g2_decap_8
XFILLER_24_642 VPWR VGND sg13g2_decap_8
XFILLER_12_837 VPWR VGND sg13g2_decap_8
XFILLER_11_347 VPWR VGND sg13g2_decap_8
XFILLER_7_329 VPWR VGND sg13g2_decap_8
XFILLER_11_74 VPWR VGND sg13g2_decap_8
XFILLER_3_557 VPWR VGND sg13g2_decap_8
XFILLER_19_403 VPWR VGND sg13g2_decap_8
XFILLER_47_756 VPWR VGND sg13g2_decap_8
XFILLER_46_266 VPWR VGND sg13g2_decap_8
XFILLER_15_620 VPWR VGND sg13g2_decap_8
XFILLER_36_60 VPWR VGND sg13g2_decap_8
XFILLER_14_130 VPWR VGND sg13g2_decap_8
XFILLER_15_697 VPWR VGND sg13g2_decap_8
XFILLER_30_667 VPWR VGND sg13g2_decap_8
Xinput13 uio_in[4] net13 VPWR VGND sg13g2_buf_1
XFILLER_6_340 VPWR VGND sg13g2_decap_8
XFILLER_7_896 VPWR VGND sg13g2_decap_8
XFILLER_42_4 VPWR VGND sg13g2_decap_8
XFILLER_38_712 VPWR VGND sg13g2_decap_8
XFILLER_26_907 VPWR VGND sg13g2_decap_8
X_37_ _05_ _03_ net19 VPWR VGND sg13g2_xor2_1
XFILLER_37_266 VPWR VGND sg13g2_decap_8
XFILLER_38_789 VPWR VGND sg13g2_decap_8
XFILLER_18_480 VPWR VGND sg13g2_decap_8
XFILLER_33_450 VPWR VGND sg13g2_decap_8
XFILLER_21_634 VPWR VGND sg13g2_decap_8
XFILLER_32_18 VPWR VGND sg13g2_decap_8
XFILLER_20_144 VPWR VGND sg13g2_decap_8
XFILLER_29_712 VPWR VGND sg13g2_decap_8
XFILLER_28_244 VPWR VGND sg13g2_decap_8
XFILLER_29_789 VPWR VGND sg13g2_decap_8
XFILLER_44_704 VPWR VGND sg13g2_decap_8
XFILLER_16_417 VPWR VGND sg13g2_decap_8
XFILLER_43_214 VPWR VGND sg13g2_decap_8
XFILLER_31_409 VPWR VGND sg13g2_decap_8
XFILLER_40_921 VPWR VGND sg13g2_decap_4
XFILLER_12_634 VPWR VGND sg13g2_decap_8
XFILLER_11_144 VPWR VGND sg13g2_decap_8
XFILLER_8_627 VPWR VGND sg13g2_decap_8
XFILLER_7_126 VPWR VGND sg13g2_decap_8
XFILLER_4_844 VPWR VGND sg13g2_decap_8
XFILLER_22_95 VPWR VGND sg13g2_decap_8
XFILLER_3_354 VPWR VGND sg13g2_decap_8
XFILLER_0_0 VPWR VGND sg13g2_decap_8
XFILLER_19_200 VPWR VGND sg13g2_decap_8
XFILLER_47_553 VPWR VGND sg13g2_decap_8
XFILLER_47_70 VPWR VGND sg13g2_decap_8
XFILLER_19_277 VPWR VGND sg13g2_decap_8
XFILLER_35_737 VPWR VGND sg13g2_decap_8
XFILLER_34_258 VPWR VGND sg13g2_decap_8
XFILLER_43_781 VPWR VGND sg13g2_decap_8
XFILLER_15_494 VPWR VGND sg13g2_decap_8
XFILLER_30_464 VPWR VGND sg13g2_decap_8
XFILLER_8_53 VPWR VGND sg13g2_decap_8
XFILLER_7_693 VPWR VGND sg13g2_decap_8
XFILLER_26_704 VPWR VGND sg13g2_decap_8
XFILLER_38_586 VPWR VGND sg13g2_decap_8
XFILLER_25_258 VPWR VGND sg13g2_decap_8
XFILLER_22_921 VPWR VGND sg13g2_decap_4
XFILLER_21_431 VPWR VGND sg13g2_decap_8
XFILLER_40_228 VPWR VGND sg13g2_decap_8
XFILLER_43_39 VPWR VGND sg13g2_decap_8
XFILLER_1_847 VPWR VGND sg13g2_decap_8
XFILLER_0_357 VPWR VGND sg13g2_decap_8
XFILLER_16_214 VPWR VGND sg13g2_decap_8
XFILLER_29_586 VPWR VGND sg13g2_decap_8
XFILLER_44_501 VPWR VGND sg13g2_decap_8
XFILLER_17_84 VPWR VGND sg13g2_decap_8
XFILLER_31_206 VPWR VGND sg13g2_decap_8
XFILLER_32_718 VPWR VGND sg13g2_decap_8
XFILLER_44_578 VPWR VGND sg13g2_decap_8
XFILLER_13_921 VPWR VGND sg13g2_decap_4
XFILLER_9_914 VPWR VGND sg13g2_decap_8
XFILLER_12_431 VPWR VGND sg13g2_decap_8
XFILLER_8_424 VPWR VGND sg13g2_decap_8
XFILLER_33_72 VPWR VGND sg13g2_decap_8
XFILLER_40_795 VPWR VGND sg13g2_decap_8
XFILLER_4_641 VPWR VGND sg13g2_decap_8
XFILLER_3_151 VPWR VGND sg13g2_decap_8
XFILLER_48_840 VPWR VGND sg13g2_decap_8
XFILLER_47_350 VPWR VGND sg13g2_decap_8
XFILLER_35_534 VPWR VGND sg13g2_decap_8
XFILLER_23_718 VPWR VGND sg13g2_decap_8
XFILLER_16_781 VPWR VGND sg13g2_decap_8
XFILLER_22_228 VPWR VGND sg13g2_decap_8
XFILLER_15_291 VPWR VGND sg13g2_decap_8
XFILLER_30_261 VPWR VGND sg13g2_decap_8
XFILLER_31_773 VPWR VGND sg13g2_decap_8
XFILLER_7_490 VPWR VGND sg13g2_decap_8
XFILLER_39_840 VPWR VGND sg13g2_decap_8
XFILLER_26_501 VPWR VGND sg13g2_decap_8
XFILLER_38_383 VPWR VGND sg13g2_decap_8
XFILLER_14_718 VPWR VGND sg13g2_decap_8
XFILLER_26_578 VPWR VGND sg13g2_decap_8
XFILLER_13_228 VPWR VGND sg13g2_decap_8
XFILLER_41_548 VPWR VGND sg13g2_decap_8
XFILLER_22_795 VPWR VGND sg13g2_decap_8
XFILLER_5_438 VPWR VGND sg13g2_decap_8
XFILLER_1_644 VPWR VGND sg13g2_decap_8
XFILLER_0_154 VPWR VGND sg13g2_decap_8
XFILLER_49_637 VPWR VGND sg13g2_decap_8
XFILLER_48_147 VPWR VGND sg13g2_decap_8
XFILLER_45_865 VPWR VGND sg13g2_decap_8
XFILLER_29_383 VPWR VGND sg13g2_decap_8
XFILLER_17_567 VPWR VGND sg13g2_decap_8
XFILLER_32_515 VPWR VGND sg13g2_decap_8
XFILLER_44_375 VPWR VGND sg13g2_decap_8
XFILLER_44_60 VPWR VGND sg13g2_decap_8
XFILLER_9_711 VPWR VGND sg13g2_decap_8
XFILLER_8_221 VPWR VGND sg13g2_decap_8
XFILLER_13_795 VPWR VGND sg13g2_decap_8
XFILLER_40_592 VPWR VGND sg13g2_decap_8
XFILLER_9_788 VPWR VGND sg13g2_decap_8
XFILLER_8_298 VPWR VGND sg13g2_decap_8
XFILLER_5_32 VPWR VGND sg13g2_decap_8
XFILLER_39_147 VPWR VGND sg13g2_decap_8
XFILLER_35_331 VPWR VGND sg13g2_decap_8
XFILLER_23_515 VPWR VGND sg13g2_decap_8
XFILLER_36_865 VPWR VGND sg13g2_decap_8
XFILLER_31_570 VPWR VGND sg13g2_decap_8
XFILLER_40_18 VPWR VGND sg13g2_decap_8
XFILLER_49_49 VPWR VGND sg13g2_decap_8
XFILLER_27_854 VPWR VGND sg13g2_decap_8
XFILLER_38_180 VPWR VGND sg13g2_decap_8
XFILLER_42_813 VPWR VGND sg13g2_decap_8
XFILLER_14_515 VPWR VGND sg13g2_decap_8
XFILLER_26_375 VPWR VGND sg13g2_decap_8
XFILLER_41_345 VPWR VGND sg13g2_decap_8
XFILLER_10_732 VPWR VGND sg13g2_decap_8
XFILLER_14_74 VPWR VGND sg13g2_decap_8
XFILLER_22_592 VPWR VGND sg13g2_decap_8
XFILLER_6_725 VPWR VGND sg13g2_decap_8
XFILLER_5_235 VPWR VGND sg13g2_decap_8
XFILLER_30_40 VPWR VGND sg13g2_decap_8
XFILLER_1_441 VPWR VGND sg13g2_decap_8
XFILLER_49_434 VPWR VGND sg13g2_decap_8
XFILLER_29_180 VPWR VGND sg13g2_decap_8
XFILLER_17_364 VPWR VGND sg13g2_decap_8
XFILLER_18_865 VPWR VGND sg13g2_decap_8
XFILLER_45_662 VPWR VGND sg13g2_decap_8
XFILLER_32_312 VPWR VGND sg13g2_decap_8
XFILLER_33_835 VPWR VGND sg13g2_decap_8
XFILLER_44_172 VPWR VGND sg13g2_decap_8
XFILLER_20_529 VPWR VGND sg13g2_decap_8
XFILLER_32_389 VPWR VGND sg13g2_decap_8
XFILLER_13_592 VPWR VGND sg13g2_decap_8
XFILLER_9_585 VPWR VGND sg13g2_decap_8
XFILLER_28_629 VPWR VGND sg13g2_decap_8
XFILLER_35_18 VPWR VGND sg13g2_decap_8
XFILLER_36_662 VPWR VGND sg13g2_decap_8
XFILLER_23_312 VPWR VGND sg13g2_decap_8
XFILLER_24_824 VPWR VGND sg13g2_decap_8
XFILLER_11_529 VPWR VGND sg13g2_decap_8
XFILLER_23_389 VPWR VGND sg13g2_decap_8
XFILLER_3_739 VPWR VGND sg13g2_decap_8
XFILLER_2_249 VPWR VGND sg13g2_decap_8
XFILLER_46_448 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_35 VPWR VGND uio_out[2] sg13g2_tielo
XFILLER_15_802 VPWR VGND sg13g2_decap_8
XFILLER_27_651 VPWR VGND sg13g2_decap_8
XFILLER_14_312 VPWR VGND sg13g2_decap_8
XFILLER_26_172 VPWR VGND sg13g2_decap_8
XFILLER_42_610 VPWR VGND sg13g2_decap_8
XFILLER_15_879 VPWR VGND sg13g2_decap_8
XFILLER_14_389 VPWR VGND sg13g2_decap_8
XFILLER_41_142 VPWR VGND sg13g2_decap_8
XFILLER_42_687 VPWR VGND sg13g2_decap_8
XFILLER_30_849 VPWR VGND sg13g2_decap_8
XFILLER_6_522 VPWR VGND sg13g2_decap_8
XFILLER_41_72 VPWR VGND sg13g2_decap_8
XFILLER_6_599 VPWR VGND sg13g2_decap_8
XFILLER_37_7 VPWR VGND sg13g2_decap_8
XFILLER_49_231 VPWR VGND sg13g2_decap_8
XFILLER_2_11 VPWR VGND sg13g2_decap_8
X_53_ _20_ _14_ _17_ VPWR VGND sg13g2_nand2_1
XFILLER_2_88 VPWR VGND sg13g2_decap_8
XFILLER_37_448 VPWR VGND sg13g2_decap_8
XFILLER_18_662 VPWR VGND sg13g2_decap_8
XFILLER_17_161 VPWR VGND sg13g2_decap_8
XFILLER_32_120 VPWR VGND sg13g2_fill_2
XFILLER_33_632 VPWR VGND sg13g2_decap_8
XFILLER_21_816 VPWR VGND sg13g2_decap_8
XFILLER_20_326 VPWR VGND sg13g2_decap_8
XFILLER_32_186 VPWR VGND sg13g2_decap_8
XFILLER_9_382 VPWR VGND sg13g2_decap_8
XFILLER_46_28 VPWR VGND sg13g2_decap_8
XFILLER_28_426 VPWR VGND sg13g2_decap_8
XFILLER_15_109 VPWR VGND sg13g2_decap_8
XFILLER_24_621 VPWR VGND sg13g2_decap_8
XFILLER_12_816 VPWR VGND sg13g2_decap_8
XFILLER_24_698 VPWR VGND sg13g2_decap_8
XFILLER_11_326 VPWR VGND sg13g2_decap_8
XFILLER_8_809 VPWR VGND sg13g2_decap_8
XFILLER_23_186 VPWR VGND sg13g2_decap_8
XFILLER_7_308 VPWR VGND sg13g2_decap_8
XFILLER_20_893 VPWR VGND sg13g2_decap_8
XFILLER_11_53 VPWR VGND sg13g2_decap_8
XFILLER_3_536 VPWR VGND sg13g2_decap_8
XFILLER_2_4 VPWR VGND sg13g2_decap_8
XFILLER_47_735 VPWR VGND sg13g2_decap_8
XFILLER_46_245 VPWR VGND sg13g2_decap_8
XFILLER_19_459 VPWR VGND sg13g2_decap_8
XFILLER_35_919 VPWR VGND sg13g2_decap_4
XFILLER_15_676 VPWR VGND sg13g2_decap_8
XFILLER_14_186 VPWR VGND sg13g2_decap_8
XFILLER_30_646 VPWR VGND sg13g2_decap_8
XFILLER_42_484 VPWR VGND sg13g2_decap_8
XFILLER_11_893 VPWR VGND sg13g2_decap_8
Xinput14 uio_in[5] net14 VPWR VGND sg13g2_buf_1
XFILLER_7_875 VPWR VGND sg13g2_decap_8
XFILLER_6_396 VPWR VGND sg13g2_decap_8
XFILLER_35_4 VPWR VGND sg13g2_decap_8
X_36_ _03_ _05_ _06_ VPWR VGND sg13g2_nor2_1
XFILLER_37_245 VPWR VGND sg13g2_decap_8
XFILLER_38_768 VPWR VGND sg13g2_decap_8
XFILLER_21_613 VPWR VGND sg13g2_decap_8
XFILLER_20_123 VPWR VGND sg13g2_decap_8
XFILLER_0_539 VPWR VGND sg13g2_decap_8
XFILLER_28_223 VPWR VGND sg13g2_decap_8
XFILLER_29_768 VPWR VGND sg13g2_decap_8
XFILLER_12_613 VPWR VGND sg13g2_decap_8
XFILLER_40_900 VPWR VGND sg13g2_decap_8
XFILLER_11_123 VPWR VGND sg13g2_decap_8
XFILLER_24_495 VPWR VGND sg13g2_decap_8
XFILLER_8_606 VPWR VGND sg13g2_decap_8
XFILLER_7_105 VPWR VGND sg13g2_decap_8
XFILLER_20_690 VPWR VGND sg13g2_decap_8
XFILLER_22_74 VPWR VGND sg13g2_decap_8
XFILLER_4_823 VPWR VGND sg13g2_decap_8
XFILLER_3_333 VPWR VGND sg13g2_decap_8
XFILLER_47_532 VPWR VGND sg13g2_decap_8
XFILLER_19_256 VPWR VGND sg13g2_decap_8
XFILLER_35_716 VPWR VGND sg13g2_decap_8
XFILLER_28_790 VPWR VGND sg13g2_decap_8
XFILLER_34_237 VPWR VGND sg13g2_decap_8
XFILLER_43_760 VPWR VGND sg13g2_decap_8
XFILLER_15_473 VPWR VGND sg13g2_decap_8
XFILLER_42_281 VPWR VGND sg13g2_decap_8
XFILLER_8_32 VPWR VGND sg13g2_decap_8
XFILLER_30_443 VPWR VGND sg13g2_decap_8
XFILLER_11_690 VPWR VGND sg13g2_decap_8
XFILLER_7_672 VPWR VGND sg13g2_decap_8
XFILLER_6_193 VPWR VGND sg13g2_decap_8
XFILLER_38_565 VPWR VGND sg13g2_decap_8
XFILLER_25_237 VPWR VGND sg13g2_decap_8
XFILLER_22_900 VPWR VGND sg13g2_decap_8
XFILLER_40_207 VPWR VGND sg13g2_decap_8
XFILLER_43_18 VPWR VGND sg13g2_decap_8
XFILLER_21_410 VPWR VGND sg13g2_decap_8
XFILLER_21_487 VPWR VGND sg13g2_decap_8
XFILLER_1_826 VPWR VGND sg13g2_decap_8
XFILLER_0_336 VPWR VGND sg13g2_decap_8
XFILLER_49_819 VPWR VGND sg13g2_decap_8
XFILLER_48_329 VPWR VGND sg13g2_decap_8
XFILLER_29_565 VPWR VGND sg13g2_decap_8
XFILLER_17_63 VPWR VGND sg13g2_decap_8
XFILLER_17_749 VPWR VGND sg13g2_decap_8
XFILLER_44_557 VPWR VGND sg13g2_decap_8
XFILLER_13_900 VPWR VGND sg13g2_decap_8
XFILLER_12_410 VPWR VGND sg13g2_decap_8
XFILLER_8_403 VPWR VGND sg13g2_decap_8
XFILLER_24_292 VPWR VGND sg13g2_decap_8
XFILLER_33_40 VPWR VGND sg13g2_decap_8
XFILLER_33_51 VPWR VGND sg13g2_decap_8
XFILLER_12_487 VPWR VGND sg13g2_decap_8
XFILLER_40_774 VPWR VGND sg13g2_decap_8
XFILLER_4_620 VPWR VGND sg13g2_decap_8
XFILLER_3_130 VPWR VGND sg13g2_decap_8
XFILLER_4_697 VPWR VGND sg13g2_decap_8
XFILLER_39_329 VPWR VGND sg13g2_decap_8
XFILLER_48_896 VPWR VGND sg13g2_decap_8
XFILLER_35_513 VPWR VGND sg13g2_decap_8
XFILLER_16_760 VPWR VGND sg13g2_decap_8
XFILLER_22_207 VPWR VGND sg13g2_decap_8
XFILLER_15_270 VPWR VGND sg13g2_decap_8
XFILLER_30_240 VPWR VGND sg13g2_decap_8
XFILLER_31_752 VPWR VGND sg13g2_decap_8
XFILLER_38_362 VPWR VGND sg13g2_decap_8
XFILLER_39_896 VPWR VGND sg13g2_decap_8
XFILLER_13_207 VPWR VGND sg13g2_decap_8
XFILLER_26_557 VPWR VGND sg13g2_decap_8
XFILLER_41_527 VPWR VGND sg13g2_decap_8
XFILLER_10_914 VPWR VGND sg13g2_decap_8
XFILLER_22_774 VPWR VGND sg13g2_decap_8
XFILLER_6_907 VPWR VGND sg13g2_decap_8
XFILLER_21_284 VPWR VGND sg13g2_decap_8
XFILLER_5_417 VPWR VGND sg13g2_decap_8
XFILLER_1_623 VPWR VGND sg13g2_decap_8
XFILLER_49_616 VPWR VGND sg13g2_decap_8
XFILLER_0_133 VPWR VGND sg13g2_decap_8
XFILLER_48_126 VPWR VGND sg13g2_decap_8
XFILLER_29_362 VPWR VGND sg13g2_decap_8
XFILLER_17_546 VPWR VGND sg13g2_decap_8
XFILLER_28_95 VPWR VGND sg13g2_decap_8
XFILLER_45_844 VPWR VGND sg13g2_decap_8
XFILLER_44_354 VPWR VGND sg13g2_decap_8
XFILLER_8_200 VPWR VGND sg13g2_decap_8
XFILLER_13_774 VPWR VGND sg13g2_decap_8
XFILLER_40_571 VPWR VGND sg13g2_decap_8
XFILLER_9_767 VPWR VGND sg13g2_decap_8
XFILLER_12_284 VPWR VGND sg13g2_decap_8
XFILLER_8_277 VPWR VGND sg13g2_decap_8
XFILLER_5_11 VPWR VGND sg13g2_decap_8
XFILLER_5_88 VPWR VGND sg13g2_decap_8
XFILLER_4_494 VPWR VGND sg13g2_decap_8
XFILLER_39_126 VPWR VGND sg13g2_decap_8
XFILLER_48_693 VPWR VGND sg13g2_decap_8
XFILLER_35_310 VPWR VGND sg13g2_decap_8
XFILLER_36_844 VPWR VGND sg13g2_decap_8
XFILLER_35_387 VPWR VGND sg13g2_decap_8
XFILLER_49_28 VPWR VGND sg13g2_decap_8
XFILLER_27_833 VPWR VGND sg13g2_decap_8
XFILLER_39_693 VPWR VGND sg13g2_decap_8
XFILLER_26_354 VPWR VGND sg13g2_decap_8
XFILLER_41_324 VPWR VGND sg13g2_decap_8
XFILLER_42_869 VPWR VGND sg13g2_decap_8
XFILLER_10_711 VPWR VGND sg13g2_decap_8
XFILLER_14_53 VPWR VGND sg13g2_decap_8
XFILLER_22_571 VPWR VGND sg13g2_decap_8
XFILLER_10_788 VPWR VGND sg13g2_decap_8
XFILLER_6_704 VPWR VGND sg13g2_decap_8
XFILLER_5_214 VPWR VGND sg13g2_decap_8
XFILLER_2_921 VPWR VGND sg13g2_decap_4
XFILLER_30_96 VPWR VGND sg13g2_decap_8
XFILLER_1_420 VPWR VGND sg13g2_decap_8
XFILLER_49_413 VPWR VGND sg13g2_decap_8
XFILLER_1_497 VPWR VGND sg13g2_decap_8
XFILLER_18_844 VPWR VGND sg13g2_decap_8
XFILLER_17_343 VPWR VGND sg13g2_decap_8
XFILLER_33_814 VPWR VGND sg13g2_decap_8
XFILLER_45_641 VPWR VGND sg13g2_decap_8
XFILLER_44_151 VPWR VGND sg13g2_decap_8
XFILLER_13_571 VPWR VGND sg13g2_decap_8
XFILLER_20_508 VPWR VGND sg13g2_decap_8
XFILLER_32_368 VPWR VGND sg13g2_decap_8
XFILLER_41_891 VPWR VGND sg13g2_decap_8
XFILLER_9_564 VPWR VGND sg13g2_decap_8
XFILLER_5_781 VPWR VGND sg13g2_decap_8
XFILLER_4_291 VPWR VGND sg13g2_decap_8
XFILLER_28_608 VPWR VGND sg13g2_decap_8
XFILLER_48_490 VPWR VGND sg13g2_decap_8
XFILLER_24_803 VPWR VGND sg13g2_decap_8
XFILLER_36_641 VPWR VGND sg13g2_decap_8
XFILLER_35_184 VPWR VGND sg13g2_decap_8
XFILLER_11_508 VPWR VGND sg13g2_decap_8
XFILLER_23_368 VPWR VGND sg13g2_decap_8
XFILLER_3_718 VPWR VGND sg13g2_decap_8
XFILLER_2_228 VPWR VGND sg13g2_decap_8
XFILLER_47_917 VPWR VGND sg13g2_decap_8
XFILLER_46_427 VPWR VGND sg13g2_decap_8
XFILLER_27_630 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_36 VPWR VGND uio_out[3] sg13g2_tielo
Xheichips25_example_small_25 VPWR VGND uio_oe[0] sg13g2_tielo
XFILLER_39_490 VPWR VGND sg13g2_decap_8
XFILLER_26_151 VPWR VGND sg13g2_decap_8
XFILLER_15_858 VPWR VGND sg13g2_decap_8
XFILLER_41_121 VPWR VGND sg13g2_decap_8
XFILLER_14_368 VPWR VGND sg13g2_decap_8
XFILLER_30_828 VPWR VGND sg13g2_decap_8
XFILLER_42_666 VPWR VGND sg13g2_decap_8
XFILLER_41_198 VPWR VGND sg13g2_decap_8
XFILLER_6_501 VPWR VGND sg13g2_decap_8
XFILLER_10_585 VPWR VGND sg13g2_decap_8
XFILLER_41_51 VPWR VGND sg13g2_decap_8
XFILLER_6_578 VPWR VGND sg13g2_decap_8
XFILLER_49_210 VPWR VGND sg13g2_decap_8
XFILLER_1_294 VPWR VGND sg13g2_decap_8
XFILLER_2_795 VPWR VGND sg13g2_decap_8
XFILLER_2_67 VPWR VGND sg13g2_decap_8
X_52_ _19_ net6 net14 VPWR VGND sg13g2_xnor2_1
XFILLER_49_287 VPWR VGND sg13g2_decap_8
XFILLER_37_427 VPWR VGND sg13g2_decap_8
XFILLER_18_641 VPWR VGND sg13g2_decap_8
XFILLER_17_140 VPWR VGND sg13g2_decap_8
XFILLER_33_611 VPWR VGND sg13g2_decap_8
XFILLER_20_305 VPWR VGND sg13g2_decap_8
XFILLER_32_165 VPWR VGND sg13g2_decap_8
XFILLER_33_688 VPWR VGND sg13g2_decap_8
XFILLER_9_361 VPWR VGND sg13g2_decap_8
XFILLER_28_405 VPWR VGND sg13g2_decap_8
XFILLER_24_600 VPWR VGND sg13g2_decap_8
XFILLER_11_305 VPWR VGND sg13g2_decap_8
XFILLER_23_165 VPWR VGND sg13g2_decap_8
XFILLER_24_677 VPWR VGND sg13g2_decap_8
XFILLER_20_872 VPWR VGND sg13g2_decap_8
XFILLER_11_32 VPWR VGND sg13g2_decap_8
XFILLER_3_515 VPWR VGND sg13g2_decap_8
XFILLER_47_714 VPWR VGND sg13g2_decap_8
XFILLER_46_224 VPWR VGND sg13g2_decap_8
XFILLER_19_438 VPWR VGND sg13g2_decap_8
XFILLER_34_419 VPWR VGND sg13g2_decap_8
XFILLER_36_95 VPWR VGND sg13g2_decap_8
XFILLER_15_655 VPWR VGND sg13g2_decap_8
XFILLER_42_463 VPWR VGND sg13g2_decap_8
XFILLER_14_165 VPWR VGND sg13g2_decap_8
XFILLER_30_625 VPWR VGND sg13g2_decap_8
XFILLER_11_872 VPWR VGND sg13g2_decap_8
Xinput15 uio_in[6] net15 VPWR VGND sg13g2_buf_1
XFILLER_10_382 VPWR VGND sg13g2_decap_8
XFILLER_7_854 VPWR VGND sg13g2_decap_8
XFILLER_6_375 VPWR VGND sg13g2_decap_8
XFILLER_2_592 VPWR VGND sg13g2_decap_8
XFILLER_28_4 VPWR VGND sg13g2_decap_8
XFILLER_37_224 VPWR VGND sg13g2_decap_8
XFILLER_38_747 VPWR VGND sg13g2_decap_8
X_35_ _05_ net3 net11 VPWR VGND sg13g2_xnor2_1
XFILLER_25_419 VPWR VGND sg13g2_decap_8
XFILLER_46_791 VPWR VGND sg13g2_decap_8
XFILLER_20_102 VPWR VGND sg13g2_decap_8
XFILLER_33_485 VPWR VGND sg13g2_decap_8
XFILLER_21_669 VPWR VGND sg13g2_decap_8
XFILLER_20_179 VPWR VGND sg13g2_decap_8
XFILLER_0_518 VPWR VGND sg13g2_decap_8
XFILLER_28_202 VPWR VGND sg13g2_decap_8
XFILLER_29_747 VPWR VGND sg13g2_decap_8
XFILLER_28_279 VPWR VGND sg13g2_decap_8
XFILLER_44_739 VPWR VGND sg13g2_decap_8
XFILLER_37_791 VPWR VGND sg13g2_decap_8
XFILLER_43_249 VPWR VGND sg13g2_decap_8
XFILLER_11_102 VPWR VGND sg13g2_decap_8
XFILLER_24_474 VPWR VGND sg13g2_decap_8
XFILLER_12_669 VPWR VGND sg13g2_decap_8
XFILLER_11_179 VPWR VGND sg13g2_decap_8
XFILLER_4_802 VPWR VGND sg13g2_decap_8
XFILLER_22_53 VPWR VGND sg13g2_decap_8
XFILLER_3_312 VPWR VGND sg13g2_decap_8
XFILLER_4_879 VPWR VGND sg13g2_decap_8
XFILLER_3_389 VPWR VGND sg13g2_decap_8
XFILLER_47_511 VPWR VGND sg13g2_decap_8
XFILLER_19_235 VPWR VGND sg13g2_decap_8
XFILLER_47_588 VPWR VGND sg13g2_decap_8
XFILLER_34_216 VPWR VGND sg13g2_decap_8
XFILLER_15_452 VPWR VGND sg13g2_decap_8
XFILLER_30_422 VPWR VGND sg13g2_decap_8
XFILLER_42_260 VPWR VGND sg13g2_decap_8
XFILLER_8_11 VPWR VGND sg13g2_decap_8
XFILLER_8_88 VPWR VGND sg13g2_decap_8
XFILLER_7_651 VPWR VGND sg13g2_decap_8
XFILLER_30_499 VPWR VGND sg13g2_decap_8
XFILLER_6_172 VPWR VGND sg13g2_decap_8
XFILLER_38_544 VPWR VGND sg13g2_decap_8
XFILLER_26_739 VPWR VGND sg13g2_decap_8
XFILLER_25_216 VPWR VGND sg13g2_decap_8
XFILLER_41_709 VPWR VGND sg13g2_decap_8
XFILLER_34_783 VPWR VGND sg13g2_decap_8
XFILLER_33_282 VPWR VGND sg13g2_decap_8
XFILLER_21_466 VPWR VGND sg13g2_decap_8
XFILLER_4_109 VPWR VGND sg13g2_decap_8
XFILLER_1_805 VPWR VGND sg13g2_decap_8
XFILLER_0_315 VPWR VGND sg13g2_decap_8
XFILLER_48_308 VPWR VGND sg13g2_decap_8
XFILLER_29_544 VPWR VGND sg13g2_decap_8
XFILLER_17_728 VPWR VGND sg13g2_decap_8
XFILLER_17_42 VPWR VGND sg13g2_decap_8
XFILLER_44_536 VPWR VGND sg13g2_decap_8
XFILLER_16_249 VPWR VGND sg13g2_decap_8
XFILLER_24_271 VPWR VGND sg13g2_decap_8
XFILLER_25_783 VPWR VGND sg13g2_decap_8
XFILLER_40_753 VPWR VGND sg13g2_decap_8
XFILLER_12_466 VPWR VGND sg13g2_decap_8
XFILLER_8_459 VPWR VGND sg13g2_decap_8
XFILLER_4_676 VPWR VGND sg13g2_decap_8
XFILLER_3_186 VPWR VGND sg13g2_decap_8
XFILLER_39_308 VPWR VGND sg13g2_decap_8
XFILLER_0_882 VPWR VGND sg13g2_decap_8
XFILLER_48_875 VPWR VGND sg13g2_decap_8
XFILLER_47_385 VPWR VGND sg13g2_decap_8
XFILLER_35_569 VPWR VGND sg13g2_decap_8
XFILLER_31_731 VPWR VGND sg13g2_decap_8
XFILLER_30_296 VPWR VGND sg13g2_decap_8
XFILLER_38_341 VPWR VGND sg13g2_decap_8
XFILLER_39_875 VPWR VGND sg13g2_decap_8
XFILLER_26_536 VPWR VGND sg13g2_decap_8
XFILLER_41_506 VPWR VGND sg13g2_decap_8
XFILLER_34_580 VPWR VGND sg13g2_decap_8
XFILLER_22_753 VPWR VGND sg13g2_decap_8
XFILLER_21_263 VPWR VGND sg13g2_decap_8
XFILLER_1_602 VPWR VGND sg13g2_decap_8
XFILLER_0_112 VPWR VGND sg13g2_decap_8
XFILLER_48_105 VPWR VGND sg13g2_decap_8
XFILLER_1_679 VPWR VGND sg13g2_decap_8
XFILLER_0_189 VPWR VGND sg13g2_decap_8
XFILLER_28_74 VPWR VGND sg13g2_decap_8
XFILLER_29_341 VPWR VGND sg13g2_decap_8
XFILLER_17_525 VPWR VGND sg13g2_decap_8
XFILLER_45_823 VPWR VGND sg13g2_decap_8
XFILLER_44_333 VPWR VGND sg13g2_decap_8
XFILLER_13_753 VPWR VGND sg13g2_decap_8
XFILLER_25_580 VPWR VGND sg13g2_decap_8
XFILLER_44_95 VPWR VGND sg13g2_decap_8
XFILLER_12_263 VPWR VGND sg13g2_decap_8
XFILLER_40_550 VPWR VGND sg13g2_decap_8
XFILLER_9_746 VPWR VGND sg13g2_decap_8
XFILLER_8_256 VPWR VGND sg13g2_decap_8
XFILLER_5_67 VPWR VGND sg13g2_decap_8
XFILLER_4_473 VPWR VGND sg13g2_decap_8
XFILLER_39_105 VPWR VGND sg13g2_decap_8
XFILLER_48_672 VPWR VGND sg13g2_decap_8
XFILLER_10_4 VPWR VGND sg13g2_decap_8
XFILLER_47_182 VPWR VGND sg13g2_decap_8
XFILLER_36_823 VPWR VGND sg13g2_decap_8
XFILLER_35_366 VPWR VGND sg13g2_decap_8
XFILLER_46_609 VPWR VGND sg13g2_decap_8
XFILLER_27_812 VPWR VGND sg13g2_decap_8
XFILLER_39_672 VPWR VGND sg13g2_decap_8
XFILLER_26_333 VPWR VGND sg13g2_decap_8
XFILLER_27_889 VPWR VGND sg13g2_decap_8
XFILLER_41_303 VPWR VGND sg13g2_decap_8
XFILLER_42_848 VPWR VGND sg13g2_decap_8
XFILLER_14_32 VPWR VGND sg13g2_decap_8
XFILLER_22_550 VPWR VGND sg13g2_decap_8
XFILLER_10_767 VPWR VGND sg13g2_decap_8
XFILLER_30_31 VPWR VGND sg13g2_decap_4
XFILLER_2_900 VPWR VGND sg13g2_decap_8
XFILLER_30_75 VPWR VGND sg13g2_decap_8
XFILLER_1_476 VPWR VGND sg13g2_decap_8
XFILLER_39_84 VPWR VGND sg13g2_decap_8
XFILLER_49_469 VPWR VGND sg13g2_decap_8
XFILLER_37_609 VPWR VGND sg13g2_decap_8
XFILLER_17_322 VPWR VGND sg13g2_decap_8
XFILLER_18_823 VPWR VGND sg13g2_decap_8
XFILLER_45_620 VPWR VGND sg13g2_decap_8
XFILLER_44_130 VPWR VGND sg13g2_decap_8
XFILLER_45_697 VPWR VGND sg13g2_decap_8
XFILLER_17_399 VPWR VGND sg13g2_decap_8
XFILLER_32_347 VPWR VGND sg13g2_decap_8
XFILLER_13_550 VPWR VGND sg13g2_decap_8
XFILLER_41_870 VPWR VGND sg13g2_decap_8
XFILLER_9_543 VPWR VGND sg13g2_decap_8
XFILLER_5_760 VPWR VGND sg13g2_decap_8
XFILLER_4_270 VPWR VGND sg13g2_decap_8
XFILLER_27_119 VPWR VGND sg13g2_decap_8
XFILLER_36_620 VPWR VGND sg13g2_decap_8
XFILLER_35_163 VPWR VGND sg13g2_decap_8
XFILLER_36_697 VPWR VGND sg13g2_decap_8
XFILLER_23_347 VPWR VGND sg13g2_decap_8
XFILLER_24_859 VPWR VGND sg13g2_decap_8
XFILLER_2_207 VPWR VGND sg13g2_decap_8
XFILLER_46_406 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_26 VPWR VGND uio_oe[1] sg13g2_tielo
XFILLER_26_130 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_37 VPWR VGND uio_out[4] sg13g2_tielo
XFILLER_15_837 VPWR VGND sg13g2_decap_8
XFILLER_27_686 VPWR VGND sg13g2_decap_8
XFILLER_14_347 VPWR VGND sg13g2_decap_8
XFILLER_25_53 VPWR VGND sg13g2_decap_8
XFILLER_41_100 VPWR VGND sg13g2_decap_8
XFILLER_42_645 VPWR VGND sg13g2_decap_8
XFILLER_25_97 VPWR VGND sg13g2_decap_8
XFILLER_30_807 VPWR VGND sg13g2_decap_8
XFILLER_41_177 VPWR VGND sg13g2_decap_8
XFILLER_10_564 VPWR VGND sg13g2_decap_8
XFILLER_6_557 VPWR VGND sg13g2_decap_8
XFILLER_2_774 VPWR VGND sg13g2_decap_8
XFILLER_1_273 VPWR VGND sg13g2_decap_8
XFILLER_49_266 VPWR VGND sg13g2_decap_8
XFILLER_2_46 VPWR VGND sg13g2_decap_8
X_51_ net6 net14 _18_ VPWR VGND sg13g2_nor2_1
XFILLER_37_406 VPWR VGND sg13g2_decap_8
XFILLER_18_620 VPWR VGND sg13g2_decap_8
XFILLER_17_196 VPWR VGND sg13g2_decap_8
XFILLER_18_697 VPWR VGND sg13g2_decap_8
XFILLER_45_494 VPWR VGND sg13g2_decap_8
XFILLER_32_144 VPWR VGND sg13g2_decap_8
XFILLER_33_667 VPWR VGND sg13g2_decap_8
XFILLER_9_340 VPWR VGND sg13g2_decap_8
XFILLER_49_0 VPWR VGND sg13g2_decap_8
XFILLER_36_494 VPWR VGND sg13g2_decap_8
XFILLER_23_144 VPWR VGND sg13g2_decap_8
XFILLER_24_656 VPWR VGND sg13g2_decap_8
XFILLER_20_851 VPWR VGND sg13g2_decap_8
XFILLER_11_11 VPWR VGND sg13g2_decap_8
XFILLER_11_88 VPWR VGND sg13g2_decap_8
XFILLER_46_203 VPWR VGND sg13g2_decap_8
XFILLER_19_417 VPWR VGND sg13g2_decap_8
XFILLER_43_921 VPWR VGND sg13g2_decap_4
XFILLER_15_634 VPWR VGND sg13g2_decap_8
XFILLER_27_483 VPWR VGND sg13g2_decap_8
XFILLER_36_74 VPWR VGND sg13g2_decap_8
XFILLER_14_144 VPWR VGND sg13g2_decap_8
XFILLER_30_604 VPWR VGND sg13g2_decap_8
XFILLER_42_442 VPWR VGND sg13g2_decap_8
XFILLER_11_851 VPWR VGND sg13g2_decap_8
XFILLER_10_361 VPWR VGND sg13g2_decap_8
XFILLER_7_833 VPWR VGND sg13g2_decap_8
Xinput16 uio_in[7] net16 VPWR VGND sg13g2_buf_1
XFILLER_6_354 VPWR VGND sg13g2_decap_8
XFILLER_2_571 VPWR VGND sg13g2_decap_8
XFILLER_37_203 VPWR VGND sg13g2_decap_8
XFILLER_38_726 VPWR VGND sg13g2_decap_8
X_34_ net3 net11 _04_ VPWR VGND sg13g2_and2_1
XFILLER_46_770 VPWR VGND sg13g2_decap_8
XFILLER_18_494 VPWR VGND sg13g2_decap_8
XFILLER_33_464 VPWR VGND sg13g2_decap_8
XFILLER_45_291 VPWR VGND sg13g2_decap_8
XFILLER_21_648 VPWR VGND sg13g2_decap_8
XFILLER_20_158 VPWR VGND sg13g2_decap_8
XFILLER_29_726 VPWR VGND sg13g2_decap_8
XFILLER_28_258 VPWR VGND sg13g2_decap_8
XFILLER_37_770 VPWR VGND sg13g2_decap_8
XFILLER_44_718 VPWR VGND sg13g2_decap_8
XFILLER_43_228 VPWR VGND sg13g2_decap_8
XFILLER_24_453 VPWR VGND sg13g2_decap_8
XFILLER_36_291 VPWR VGND sg13g2_decap_8
XFILLER_12_648 VPWR VGND sg13g2_decap_8
XFILLER_11_158 VPWR VGND sg13g2_decap_8
XFILLER_22_32 VPWR VGND sg13g2_decap_8
XFILLER_4_858 VPWR VGND sg13g2_decap_8
XFILLER_3_368 VPWR VGND sg13g2_decap_8
XFILLER_19_214 VPWR VGND sg13g2_decap_8
XFILLER_47_567 VPWR VGND sg13g2_decap_8
XFILLER_47_84 VPWR VGND sg13g2_decap_8
XFILLER_16_921 VPWR VGND sg13g2_decap_4
XFILLER_27_280 VPWR VGND sg13g2_decap_8
XFILLER_15_431 VPWR VGND sg13g2_decap_8
XFILLER_30_401 VPWR VGND sg13g2_decap_8
XFILLER_31_913 VPWR VGND sg13g2_decap_8
XFILLER_31_924 VPWR VGND sg13g2_fill_1
XFILLER_43_795 VPWR VGND sg13g2_decap_8
XFILLER_8_67 VPWR VGND sg13g2_decap_8
XFILLER_30_478 VPWR VGND sg13g2_decap_8
XFILLER_7_630 VPWR VGND sg13g2_decap_8
XFILLER_6_151 VPWR VGND sg13g2_decap_8
XFILLER_40_4 VPWR VGND sg13g2_decap_8
XFILLER_38_523 VPWR VGND sg13g2_decap_8
XFILLER_26_718 VPWR VGND sg13g2_decap_8
XFILLER_19_781 VPWR VGND sg13g2_decap_8
XFILLER_18_291 VPWR VGND sg13g2_decap_8
XFILLER_34_762 VPWR VGND sg13g2_decap_8
XFILLER_33_261 VPWR VGND sg13g2_decap_8
XFILLER_21_445 VPWR VGND sg13g2_decap_8
XFILLER_29_523 VPWR VGND sg13g2_decap_8
XFILLER_17_21 VPWR VGND sg13g2_decap_8
XFILLER_17_707 VPWR VGND sg13g2_decap_8
XFILLER_44_515 VPWR VGND sg13g2_decap_8
XFILLER_16_228 VPWR VGND sg13g2_decap_8
XFILLER_17_98 VPWR VGND sg13g2_decap_8
XFILLER_25_762 VPWR VGND sg13g2_decap_8
XFILLER_24_250 VPWR VGND sg13g2_decap_8
XFILLER_12_445 VPWR VGND sg13g2_decap_8
XFILLER_40_732 VPWR VGND sg13g2_decap_8
XFILLER_33_86 VPWR VGND sg13g2_decap_8
XFILLER_8_438 VPWR VGND sg13g2_decap_8
XFILLER_4_655 VPWR VGND sg13g2_decap_8
XFILLER_3_165 VPWR VGND sg13g2_decap_8
XFILLER_0_861 VPWR VGND sg13g2_decap_8
XFILLER_48_854 VPWR VGND sg13g2_decap_8
XFILLER_47_364 VPWR VGND sg13g2_decap_8
XFILLER_35_548 VPWR VGND sg13g2_decap_8
XFILLER_16_795 VPWR VGND sg13g2_decap_8
XFILLER_31_710 VPWR VGND sg13g2_decap_8
XFILLER_43_592 VPWR VGND sg13g2_decap_8
XFILLER_31_787 VPWR VGND sg13g2_decap_8
XFILLER_30_275 VPWR VGND sg13g2_decap_8
XFILLER_38_320 VPWR VGND sg13g2_decap_8
XFILLER_39_854 VPWR VGND sg13g2_decap_8
XFILLER_26_515 VPWR VGND sg13g2_decap_8
XFILLER_38_397 VPWR VGND sg13g2_decap_8
XFILLER_22_732 VPWR VGND sg13g2_decap_8
XFILLER_21_242 VPWR VGND sg13g2_decap_8
XFILLER_1_658 VPWR VGND sg13g2_decap_8
XFILLER_0_168 VPWR VGND sg13g2_decap_8
XFILLER_29_320 VPWR VGND sg13g2_decap_8
XFILLER_17_504 VPWR VGND sg13g2_decap_8
XFILLER_28_53 VPWR VGND sg13g2_decap_8
XFILLER_45_802 VPWR VGND sg13g2_decap_8
XFILLER_29_397 VPWR VGND sg13g2_decap_8
XFILLER_44_312 VPWR VGND sg13g2_decap_8
XFILLER_45_879 VPWR VGND sg13g2_decap_8
XFILLER_32_529 VPWR VGND sg13g2_decap_8
XFILLER_44_389 VPWR VGND sg13g2_decap_8
XFILLER_13_732 VPWR VGND sg13g2_decap_8
XFILLER_44_74 VPWR VGND sg13g2_decap_8
XFILLER_9_725 VPWR VGND sg13g2_decap_8
XFILLER_12_242 VPWR VGND sg13g2_decap_8
XFILLER_8_235 VPWR VGND sg13g2_decap_8
XFILLER_5_46 VPWR VGND sg13g2_decap_8
XFILLER_4_452 VPWR VGND sg13g2_decap_8
XFILLER_48_651 VPWR VGND sg13g2_decap_8
XFILLER_36_802 VPWR VGND sg13g2_decap_8
XFILLER_47_161 VPWR VGND sg13g2_decap_8
XFILLER_35_345 VPWR VGND sg13g2_decap_8
XFILLER_36_879 VPWR VGND sg13g2_decap_8
XFILLER_23_529 VPWR VGND sg13g2_decap_8
XFILLER_16_592 VPWR VGND sg13g2_decap_8
XFILLER_31_584 VPWR VGND sg13g2_decap_8
XFILLER_39_651 VPWR VGND sg13g2_decap_8
XFILLER_26_312 VPWR VGND sg13g2_decap_8
XFILLER_45_109 VPWR VGND sg13g2_decap_8
XFILLER_27_868 VPWR VGND sg13g2_decap_8
XFILLER_38_194 VPWR VGND sg13g2_decap_8
XFILLER_14_529 VPWR VGND sg13g2_decap_8
XFILLER_26_389 VPWR VGND sg13g2_decap_8
XFILLER_42_827 VPWR VGND sg13g2_decap_8
XFILLER_14_11 VPWR VGND sg13g2_decap_8
XFILLER_41_359 VPWR VGND sg13g2_decap_8
XFILLER_10_746 VPWR VGND sg13g2_decap_8
XFILLER_14_88 VPWR VGND sg13g2_decap_8
XFILLER_6_739 VPWR VGND sg13g2_decap_8
XFILLER_5_249 VPWR VGND sg13g2_decap_8
XFILLER_30_54 VPWR VGND sg13g2_decap_8
XFILLER_1_455 VPWR VGND sg13g2_decap_8
XFILLER_49_448 VPWR VGND sg13g2_decap_8
XFILLER_39_63 VPWR VGND sg13g2_decap_8
XFILLER_18_802 VPWR VGND sg13g2_decap_8
XFILLER_17_301 VPWR VGND sg13g2_decap_8
XFILLER_36_109 VPWR VGND sg13g2_decap_8
XFILLER_18_879 VPWR VGND sg13g2_decap_8
XFILLER_29_194 VPWR VGND sg13g2_decap_8
XFILLER_17_378 VPWR VGND sg13g2_decap_8
XFILLER_45_676 VPWR VGND sg13g2_decap_8
XFILLER_32_326 VPWR VGND sg13g2_decap_8
XFILLER_33_849 VPWR VGND sg13g2_decap_8
XFILLER_44_186 VPWR VGND sg13g2_decap_8
XFILLER_9_522 VPWR VGND sg13g2_decap_8
XFILLER_9_599 VPWR VGND sg13g2_decap_8
XFILLER_24_838 VPWR VGND sg13g2_decap_8
XFILLER_35_142 VPWR VGND sg13g2_decap_8
XFILLER_36_676 VPWR VGND sg13g2_decap_8
XFILLER_23_326 VPWR VGND sg13g2_decap_8
XFILLER_32_893 VPWR VGND sg13g2_decap_8
XFILLER_31_381 VPWR VGND sg13g2_decap_8
XFILLER_18_109 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_27 VPWR VGND uio_oe[2] sg13g2_tielo
XFILLER_15_816 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_38 VPWR VGND uio_out[5] sg13g2_tielo
XFILLER_27_665 VPWR VGND sg13g2_decap_8
XFILLER_14_326 VPWR VGND sg13g2_decap_8
XFILLER_25_32 VPWR VGND sg13g2_decap_8
XFILLER_26_186 VPWR VGND sg13g2_decap_8
XFILLER_42_624 VPWR VGND sg13g2_decap_8
XFILLER_41_156 VPWR VGND sg13g2_decap_8
XFILLER_23_893 VPWR VGND sg13g2_decap_8
XFILLER_10_543 VPWR VGND sg13g2_decap_8
XFILLER_6_536 VPWR VGND sg13g2_decap_8
XFILLER_41_86 VPWR VGND sg13g2_decap_8
XFILLER_1_252 VPWR VGND sg13g2_decap_8
XFILLER_2_753 VPWR VGND sg13g2_decap_8
XFILLER_2_25 VPWR VGND sg13g2_decap_8
XFILLER_49_245 VPWR VGND sg13g2_decap_8
X_50_ net21 _13_ _16_ VPWR VGND sg13g2_xnor2_1
XFILLER_38_908 VPWR VGND sg13g2_decap_8
XFILLER_18_676 VPWR VGND sg13g2_decap_8
XFILLER_45_473 VPWR VGND sg13g2_decap_8
XFILLER_17_175 VPWR VGND sg13g2_decap_8
XFILLER_33_646 VPWR VGND sg13g2_decap_8
XFILLER_14_893 VPWR VGND sg13g2_decap_8
XFILLER_9_396 VPWR VGND sg13g2_decap_8
XFILLER_29_908 VPWR VGND sg13g2_decap_8
XFILLER_24_635 VPWR VGND sg13g2_decap_8
XFILLER_36_473 VPWR VGND sg13g2_decap_8
XFILLER_23_123 VPWR VGND sg13g2_decap_8
XFILLER_20_830 VPWR VGND sg13g2_decap_8
XFILLER_32_690 VPWR VGND sg13g2_decap_8
XFILLER_11_67 VPWR VGND sg13g2_decap_8
XFILLER_47_749 VPWR VGND sg13g2_decap_8
XFILLER_46_259 VPWR VGND sg13g2_decap_8
XFILLER_27_462 VPWR VGND sg13g2_decap_8
XFILLER_36_53 VPWR VGND sg13g2_decap_8
XFILLER_43_900 VPWR VGND sg13g2_decap_8
XFILLER_15_613 VPWR VGND sg13g2_decap_8
XFILLER_42_421 VPWR VGND sg13g2_decap_8
XFILLER_14_123 VPWR VGND sg13g2_decap_8
XFILLER_42_498 VPWR VGND sg13g2_decap_8
XFILLER_11_830 VPWR VGND sg13g2_decap_8
XFILLER_23_690 VPWR VGND sg13g2_decap_8
XFILLER_10_340 VPWR VGND sg13g2_decap_8
XFILLER_7_812 VPWR VGND sg13g2_decap_8
XFILLER_6_333 VPWR VGND sg13g2_decap_8
XFILLER_7_889 VPWR VGND sg13g2_decap_8
XFILLER_2_550 VPWR VGND sg13g2_decap_8
XFILLER_38_705 VPWR VGND sg13g2_decap_8
X_33_ VGND VPWR _01_ _03_ _02_ _00_ sg13g2_a21oi_2
XFILLER_37_259 VPWR VGND sg13g2_decap_8
XFILLER_18_473 VPWR VGND sg13g2_decap_8
XFILLER_45_270 VPWR VGND sg13g2_decap_8
XFILLER_33_443 VPWR VGND sg13g2_decap_8
XFILLER_21_627 VPWR VGND sg13g2_decap_8
XFILLER_14_690 VPWR VGND sg13g2_decap_8
XFILLER_20_137 VPWR VGND sg13g2_decap_8
XFILLER_9_193 VPWR VGND sg13g2_decap_8
XFILLER_29_705 VPWR VGND sg13g2_decap_8
XFILLER_28_237 VPWR VGND sg13g2_decap_8
XFILLER_43_207 VPWR VGND sg13g2_decap_8
XFILLER_36_270 VPWR VGND sg13g2_decap_8
XFILLER_24_432 VPWR VGND sg13g2_decap_8
XFILLER_12_627 VPWR VGND sg13g2_decap_8
XFILLER_40_914 VPWR VGND sg13g2_decap_8
XFILLER_11_137 VPWR VGND sg13g2_decap_8
XFILLER_7_119 VPWR VGND sg13g2_decap_8
XFILLER_22_11 VPWR VGND sg13g2_decap_8
XFILLER_22_88 VPWR VGND sg13g2_decap_8
XFILLER_4_837 VPWR VGND sg13g2_decap_8
XFILLER_3_347 VPWR VGND sg13g2_decap_8
XFILLER_47_546 VPWR VGND sg13g2_decap_8
XFILLER_47_63 VPWR VGND sg13g2_decap_8
XFILLER_16_900 VPWR VGND sg13g2_decap_8
XFILLER_15_410 VPWR VGND sg13g2_decap_8
XFILLER_15_487 VPWR VGND sg13g2_decap_8
XFILLER_43_774 VPWR VGND sg13g2_decap_8
XFILLER_42_295 VPWR VGND sg13g2_decap_8
XFILLER_8_46 VPWR VGND sg13g2_decap_8
XFILLER_30_457 VPWR VGND sg13g2_decap_8
XFILLER_6_130 VPWR VGND sg13g2_decap_8
XFILLER_7_686 VPWR VGND sg13g2_decap_8
XFILLER_33_4 VPWR VGND sg13g2_decap_8
XFILLER_38_502 VPWR VGND sg13g2_decap_8
XFILLER_19_760 VPWR VGND sg13g2_decap_8
XFILLER_38_579 VPWR VGND sg13g2_decap_8
XFILLER_18_270 VPWR VGND sg13g2_decap_8
XFILLER_34_741 VPWR VGND sg13g2_decap_8
XFILLER_22_914 VPWR VGND sg13g2_decap_8
XFILLER_33_240 VPWR VGND sg13g2_decap_8
XFILLER_21_424 VPWR VGND sg13g2_decap_8
XFILLER_29_502 VPWR VGND sg13g2_decap_8
XFILLER_29_579 VPWR VGND sg13g2_decap_8
XFILLER_16_207 VPWR VGND sg13g2_decap_8
XFILLER_17_77 VPWR VGND sg13g2_decap_8
XFILLER_25_741 VPWR VGND sg13g2_decap_8
XFILLER_13_914 VPWR VGND sg13g2_decap_8
XFILLER_40_711 VPWR VGND sg13g2_decap_8
XFILLER_9_907 VPWR VGND sg13g2_decap_8
XFILLER_12_424 VPWR VGND sg13g2_decap_8
XFILLER_8_417 VPWR VGND sg13g2_decap_8
XFILLER_33_65 VPWR VGND sg13g2_decap_8
XFILLER_40_788 VPWR VGND sg13g2_decap_8
XFILLER_4_634 VPWR VGND sg13g2_decap_8
XFILLER_3_144 VPWR VGND sg13g2_decap_8
XFILLER_0_840 VPWR VGND sg13g2_decap_8
XFILLER_48_833 VPWR VGND sg13g2_decap_8
XFILLER_47_343 VPWR VGND sg13g2_decap_8
XFILLER_35_527 VPWR VGND sg13g2_decap_8
XFILLER_16_774 VPWR VGND sg13g2_decap_8
XFILLER_43_571 VPWR VGND sg13g2_decap_8
XFILLER_15_284 VPWR VGND sg13g2_decap_8
XFILLER_30_254 VPWR VGND sg13g2_decap_8
XFILLER_31_766 VPWR VGND sg13g2_decap_8
XFILLER_7_483 VPWR VGND sg13g2_decap_8
XFILLER_39_833 VPWR VGND sg13g2_decap_8
XFILLER_38_376 VPWR VGND sg13g2_decap_8
XFILLER_0_91 VPWR VGND sg13g2_decap_8
XFILLER_22_711 VPWR VGND sg13g2_decap_8
XFILLER_21_221 VPWR VGND sg13g2_decap_8
XFILLER_22_788 VPWR VGND sg13g2_decap_8
XFILLER_21_298 VPWR VGND sg13g2_decap_8
XFILLER_1_637 VPWR VGND sg13g2_decap_8
XFILLER_0_147 VPWR VGND sg13g2_decap_8
XFILLER_28_32 VPWR VGND sg13g2_decap_8
XFILLER_29_376 VPWR VGND sg13g2_decap_8
XFILLER_45_858 VPWR VGND sg13g2_decap_8
XFILLER_13_711 VPWR VGND sg13g2_decap_8
XFILLER_32_508 VPWR VGND sg13g2_decap_8
XFILLER_44_53 VPWR VGND sg13g2_decap_8
XFILLER_44_368 VPWR VGND sg13g2_decap_8
XFILLER_12_221 VPWR VGND sg13g2_decap_8
XFILLER_9_704 VPWR VGND sg13g2_decap_8
XFILLER_8_214 VPWR VGND sg13g2_decap_8
XFILLER_13_788 VPWR VGND sg13g2_decap_8
XFILLER_40_585 VPWR VGND sg13g2_decap_8
XFILLER_12_298 VPWR VGND sg13g2_decap_8
XFILLER_5_921 VPWR VGND sg13g2_decap_4
XFILLER_5_25 VPWR VGND sg13g2_decap_8
XFILLER_4_431 VPWR VGND sg13g2_decap_8
XFILLER_48_630 VPWR VGND sg13g2_decap_8
XFILLER_47_140 VPWR VGND sg13g2_decap_8
XFILLER_35_324 VPWR VGND sg13g2_decap_8
XFILLER_36_858 VPWR VGND sg13g2_decap_8
XFILLER_23_508 VPWR VGND sg13g2_decap_8
XFILLER_16_571 VPWR VGND sg13g2_decap_8
XFILLER_31_563 VPWR VGND sg13g2_decap_8
XFILLER_8_781 VPWR VGND sg13g2_decap_8
XFILLER_7_280 VPWR VGND sg13g2_decap_8
XFILLER_39_630 VPWR VGND sg13g2_decap_8
XFILLER_38_173 VPWR VGND sg13g2_decap_8
XFILLER_27_847 VPWR VGND sg13g2_decap_8
XFILLER_14_508 VPWR VGND sg13g2_decap_8
XFILLER_26_368 VPWR VGND sg13g2_decap_8
XFILLER_42_806 VPWR VGND sg13g2_decap_8
XFILLER_35_891 VPWR VGND sg13g2_decap_8
XFILLER_41_338 VPWR VGND sg13g2_decap_8
XFILLER_10_725 VPWR VGND sg13g2_decap_8
XFILLER_14_67 VPWR VGND sg13g2_decap_8
XFILLER_22_585 VPWR VGND sg13g2_decap_8
XFILLER_6_718 VPWR VGND sg13g2_decap_8
XFILLER_5_228 VPWR VGND sg13g2_decap_8
XFILLER_30_11 VPWR VGND sg13g2_fill_1
XFILLER_1_434 VPWR VGND sg13g2_decap_8
XFILLER_39_20 VPWR VGND sg13g2_fill_1
XFILLER_39_42 VPWR VGND sg13g2_decap_8
XFILLER_49_427 VPWR VGND sg13g2_decap_8
XFILLER_18_858 VPWR VGND sg13g2_decap_8
XFILLER_29_173 VPWR VGND sg13g2_decap_8
XFILLER_45_655 VPWR VGND sg13g2_decap_8
XFILLER_17_357 VPWR VGND sg13g2_decap_8
XFILLER_32_305 VPWR VGND sg13g2_decap_8
XFILLER_33_828 VPWR VGND sg13g2_decap_8
XFILLER_44_165 VPWR VGND sg13g2_decap_8
XFILLER_9_501 VPWR VGND sg13g2_decap_8
XFILLER_13_585 VPWR VGND sg13g2_decap_8
XFILLER_9_578 VPWR VGND sg13g2_decap_8
XFILLER_40_382 VPWR VGND sg13g2_decap_8
XFILLER_5_795 VPWR VGND sg13g2_decap_8
XFILLER_35_121 VPWR VGND sg13g2_decap_8
XFILLER_36_655 VPWR VGND sg13g2_decap_8
XFILLER_23_305 VPWR VGND sg13g2_decap_8
XFILLER_24_817 VPWR VGND sg13g2_decap_8
XFILLER_35_198 VPWR VGND sg13g2_decap_8
XFILLER_31_360 VPWR VGND sg13g2_decap_8
XFILLER_32_872 VPWR VGND sg13g2_decap_8
XFILLER_27_644 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_39 VPWR VGND uio_out[6] sg13g2_tielo
Xheichips25_example_small_28 VPWR VGND uio_oe[3] sg13g2_tielo
XFILLER_25_11 VPWR VGND sg13g2_decap_8
XFILLER_42_603 VPWR VGND sg13g2_decap_8
XFILLER_14_305 VPWR VGND sg13g2_decap_8
XFILLER_26_165 VPWR VGND sg13g2_decap_8
XFILLER_41_135 VPWR VGND sg13g2_decap_8
XFILLER_23_872 VPWR VGND sg13g2_decap_8
XFILLER_10_522 VPWR VGND sg13g2_decap_8
XFILLER_22_382 VPWR VGND sg13g2_decap_8
XFILLER_41_32 VPWR VGND sg13g2_decap_4
XFILLER_6_515 VPWR VGND sg13g2_decap_8
XFILLER_41_65 VPWR VGND sg13g2_decap_8
XFILLER_10_599 VPWR VGND sg13g2_decap_8
XFILLER_2_732 VPWR VGND sg13g2_decap_8
XFILLER_1_231 VPWR VGND sg13g2_decap_8
XFILLER_49_224 VPWR VGND sg13g2_decap_8
XFILLER_17_154 VPWR VGND sg13g2_decap_8
XFILLER_18_655 VPWR VGND sg13g2_decap_8
XFILLER_45_452 VPWR VGND sg13g2_decap_8
XFILLER_32_102 VPWR VGND sg13g2_decap_8
XFILLER_33_625 VPWR VGND sg13g2_decap_8
XFILLER_21_809 VPWR VGND sg13g2_decap_8
XFILLER_14_872 VPWR VGND sg13g2_decap_8
XFILLER_20_319 VPWR VGND sg13g2_decap_8
XFILLER_32_179 VPWR VGND sg13g2_decap_8
XFILLER_13_382 VPWR VGND sg13g2_decap_8
XFILLER_9_375 VPWR VGND sg13g2_decap_8
XFILLER_5_592 VPWR VGND sg13g2_decap_8
XFILLER_28_419 VPWR VGND sg13g2_decap_8
XFILLER_49_791 VPWR VGND sg13g2_decap_8
XFILLER_36_452 VPWR VGND sg13g2_decap_8
XFILLER_23_102 VPWR VGND sg13g2_decap_8
XFILLER_24_614 VPWR VGND sg13g2_decap_8
XFILLER_12_809 VPWR VGND sg13g2_decap_8
XFILLER_11_319 VPWR VGND sg13g2_decap_8
XFILLER_23_179 VPWR VGND sg13g2_decap_8
XFILLER_20_886 VPWR VGND sg13g2_decap_8
XFILLER_11_46 VPWR VGND sg13g2_decap_8
XFILLER_3_529 VPWR VGND sg13g2_decap_8
XFILLER_47_728 VPWR VGND sg13g2_decap_8
XFILLER_46_238 VPWR VGND sg13g2_decap_8
XFILLER_27_441 VPWR VGND sg13g2_decap_8
XFILLER_36_32 VPWR VGND sg13g2_decap_8
XFILLER_14_102 VPWR VGND sg13g2_decap_8
XFILLER_42_400 VPWR VGND sg13g2_decap_8
XFILLER_15_669 VPWR VGND sg13g2_decap_8
XFILLER_14_179 VPWR VGND sg13g2_decap_8
XFILLER_42_477 VPWR VGND sg13g2_decap_8
XFILLER_30_639 VPWR VGND sg13g2_decap_8
XFILLER_11_886 VPWR VGND sg13g2_decap_8
XFILLER_7_868 VPWR VGND sg13g2_decap_8
XFILLER_6_312 VPWR VGND sg13g2_decap_8
XFILLER_10_396 VPWR VGND sg13g2_decap_8
XFILLER_6_389 VPWR VGND sg13g2_decap_8
X_32_ _02_ _00_ net18 VPWR VGND sg13g2_xor2_1
XFILLER_37_238 VPWR VGND sg13g2_decap_8
XFILLER_18_452 VPWR VGND sg13g2_decap_8
XFILLER_34_923 VPWR VGND sg13g2_fill_2
XFILLER_33_422 VPWR VGND sg13g2_decap_8
XFILLER_21_606 VPWR VGND sg13g2_decap_8
XFILLER_20_116 VPWR VGND sg13g2_decap_8
XFILLER_33_499 VPWR VGND sg13g2_decap_8
XFILLER_9_172 VPWR VGND sg13g2_decap_8
XFILLER_28_216 VPWR VGND sg13g2_decap_8
XFILLER_24_411 VPWR VGND sg13g2_decap_8
XFILLER_25_923 VPWR VGND sg13g2_fill_2
XFILLER_12_606 VPWR VGND sg13g2_decap_8
XFILLER_24_488 VPWR VGND sg13g2_decap_8
XFILLER_11_116 VPWR VGND sg13g2_decap_8
XFILLER_20_683 VPWR VGND sg13g2_decap_8
XFILLER_22_67 VPWR VGND sg13g2_decap_8
XFILLER_4_816 VPWR VGND sg13g2_decap_8
XFILLER_3_326 VPWR VGND sg13g2_decap_8
XFILLER_47_525 VPWR VGND sg13g2_decap_8
XFILLER_47_42 VPWR VGND sg13g2_decap_8
XFILLER_19_249 VPWR VGND sg13g2_decap_8
XFILLER_35_709 VPWR VGND sg13g2_decap_8
XFILLER_28_783 VPWR VGND sg13g2_decap_8
XFILLER_43_753 VPWR VGND sg13g2_decap_8
XFILLER_15_466 VPWR VGND sg13g2_decap_8
XFILLER_30_436 VPWR VGND sg13g2_decap_8
XFILLER_42_274 VPWR VGND sg13g2_decap_8
XFILLER_8_25 VPWR VGND sg13g2_decap_8
XFILLER_11_683 VPWR VGND sg13g2_decap_8
XFILLER_10_193 VPWR VGND sg13g2_decap_8
XFILLER_7_665 VPWR VGND sg13g2_decap_8
XFILLER_6_186 VPWR VGND sg13g2_decap_8
XFILLER_3_893 VPWR VGND sg13g2_decap_8
XFILLER_26_4 VPWR VGND sg13g2_decap_8
XFILLER_38_558 VPWR VGND sg13g2_decap_8
XFILLER_34_720 VPWR VGND sg13g2_decap_8
XFILLER_21_403 VPWR VGND sg13g2_decap_8
XFILLER_33_296 VPWR VGND sg13g2_decap_8
XFILLER_34_797 VPWR VGND sg13g2_decap_8
XFILLER_1_819 VPWR VGND sg13g2_decap_8
XFILLER_0_329 VPWR VGND sg13g2_decap_8
XFILLER_29_558 VPWR VGND sg13g2_decap_8
XFILLER_17_56 VPWR VGND sg13g2_decap_8
XFILLER_25_720 VPWR VGND sg13g2_decap_8
XFILLER_12_403 VPWR VGND sg13g2_decap_8
XFILLER_24_285 VPWR VGND sg13g2_decap_8
XFILLER_25_797 VPWR VGND sg13g2_decap_8
XFILLER_33_11 VPWR VGND sg13g2_decap_8
XFILLER_33_33 VPWR VGND sg13g2_decap_8
XFILLER_40_767 VPWR VGND sg13g2_decap_8
XFILLER_20_480 VPWR VGND sg13g2_decap_8
XFILLER_4_613 VPWR VGND sg13g2_decap_8
XFILLER_3_123 VPWR VGND sg13g2_decap_8
XFILLER_48_812 VPWR VGND sg13g2_decap_8
XFILLER_47_322 VPWR VGND sg13g2_decap_8
XFILLER_0_896 VPWR VGND sg13g2_decap_8
XFILLER_48_889 VPWR VGND sg13g2_decap_8
XFILLER_35_506 VPWR VGND sg13g2_decap_8
XFILLER_47_399 VPWR VGND sg13g2_decap_8
XFILLER_28_580 VPWR VGND sg13g2_decap_8
XFILLER_16_753 VPWR VGND sg13g2_decap_8
XFILLER_43_550 VPWR VGND sg13g2_decap_8
XFILLER_15_263 VPWR VGND sg13g2_decap_8
XFILLER_31_745 VPWR VGND sg13g2_decap_8
XFILLER_30_233 VPWR VGND sg13g2_decap_8
XFILLER_11_480 VPWR VGND sg13g2_decap_8
XFILLER_7_462 VPWR VGND sg13g2_decap_8
XFILLER_3_690 VPWR VGND sg13g2_decap_8
XFILLER_39_812 VPWR VGND sg13g2_decap_8
XFILLER_17_0 VPWR VGND sg13g2_decap_8
XFILLER_38_355 VPWR VGND sg13g2_decap_8
XFILLER_39_889 VPWR VGND sg13g2_decap_8
XFILLER_0_70 VPWR VGND sg13g2_decap_8
XFILLER_21_200 VPWR VGND sg13g2_decap_8
XFILLER_34_594 VPWR VGND sg13g2_decap_8
XFILLER_10_907 VPWR VGND sg13g2_decap_8
XFILLER_22_767 VPWR VGND sg13g2_decap_8
XFILLER_21_277 VPWR VGND sg13g2_decap_8
XFILLER_1_616 VPWR VGND sg13g2_decap_8
XFILLER_0_126 VPWR VGND sg13g2_decap_8
XFILLER_49_609 VPWR VGND sg13g2_decap_8
XFILLER_48_119 VPWR VGND sg13g2_decap_8
XFILLER_28_11 VPWR VGND sg13g2_decap_8
XFILLER_29_355 VPWR VGND sg13g2_decap_8
XFILLER_28_88 VPWR VGND sg13g2_decap_8
XFILLER_45_837 VPWR VGND sg13g2_decap_8
XFILLER_17_539 VPWR VGND sg13g2_decap_8
XFILLER_44_347 VPWR VGND sg13g2_decap_8
XFILLER_44_32 VPWR VGND sg13g2_decap_8
XFILLER_12_200 VPWR VGND sg13g2_decap_8
XFILLER_25_594 VPWR VGND sg13g2_decap_8
XFILLER_13_767 VPWR VGND sg13g2_decap_8
XFILLER_12_277 VPWR VGND sg13g2_decap_8
XFILLER_40_564 VPWR VGND sg13g2_decap_8
XFILLER_5_900 VPWR VGND sg13g2_decap_8
XFILLER_4_410 VPWR VGND sg13g2_decap_8
XFILLER_4_487 VPWR VGND sg13g2_decap_8
XFILLER_39_119 VPWR VGND sg13g2_decap_8
XFILLER_0_693 VPWR VGND sg13g2_decap_8
XFILLER_48_686 VPWR VGND sg13g2_decap_8
XFILLER_35_303 VPWR VGND sg13g2_decap_8
XFILLER_36_837 VPWR VGND sg13g2_decap_8
XFILLER_47_196 VPWR VGND sg13g2_decap_8
XFILLER_16_550 VPWR VGND sg13g2_decap_8
XFILLER_31_542 VPWR VGND sg13g2_decap_8
XFILLER_8_760 VPWR VGND sg13g2_decap_8
XFILLER_27_826 VPWR VGND sg13g2_decap_8
XFILLER_38_152 VPWR VGND sg13g2_decap_8
XFILLER_39_686 VPWR VGND sg13g2_decap_8
XFILLER_26_347 VPWR VGND sg13g2_decap_8
XFILLER_35_870 VPWR VGND sg13g2_decap_8
XFILLER_41_317 VPWR VGND sg13g2_decap_8
XFILLER_34_391 VPWR VGND sg13g2_decap_8
XFILLER_10_704 VPWR VGND sg13g2_decap_8
XFILLER_14_46 VPWR VGND sg13g2_decap_8
XFILLER_22_564 VPWR VGND sg13g2_decap_8
XFILLER_5_207 VPWR VGND sg13g2_decap_8
XFILLER_2_914 VPWR VGND sg13g2_decap_8
XFILLER_30_89 VPWR VGND sg13g2_decap_8
XFILLER_1_413 VPWR VGND sg13g2_decap_8
XFILLER_49_406 VPWR VGND sg13g2_decap_8
XFILLER_39_98 VPWR VGND sg13g2_decap_8
XFILLER_29_152 VPWR VGND sg13g2_decap_8
XFILLER_17_336 VPWR VGND sg13g2_decap_8
XFILLER_18_837 VPWR VGND sg13g2_decap_8
XFILLER_45_634 VPWR VGND sg13g2_decap_8
XFILLER_33_807 VPWR VGND sg13g2_decap_8
XFILLER_44_144 VPWR VGND sg13g2_decap_8
XFILLER_25_391 VPWR VGND sg13g2_decap_8
XFILLER_13_564 VPWR VGND sg13g2_decap_8
XFILLER_40_361 VPWR VGND sg13g2_decap_8
XFILLER_41_884 VPWR VGND sg13g2_decap_8
XFILLER_9_557 VPWR VGND sg13g2_decap_8
XFILLER_5_774 VPWR VGND sg13g2_decap_8
XFILLER_4_284 VPWR VGND sg13g2_decap_8
XFILLER_0_490 VPWR VGND sg13g2_decap_8
XFILLER_48_483 VPWR VGND sg13g2_decap_8
XFILLER_36_634 VPWR VGND sg13g2_decap_8
XFILLER_35_177 VPWR VGND sg13g2_decap_8
XFILLER_32_851 VPWR VGND sg13g2_decap_8
XFILLER_27_623 VPWR VGND sg13g2_decap_8
XFILLER_39_483 VPWR VGND sg13g2_decap_8
Xheichips25_example_small_29 VPWR VGND uio_oe[4] sg13g2_tielo
XFILLER_26_144 VPWR VGND sg13g2_decap_8
XFILLER_41_114 VPWR VGND sg13g2_decap_8
XFILLER_23_851 VPWR VGND sg13g2_decap_8
XFILLER_25_67 VPWR VGND sg13g2_decap_8
XFILLER_42_659 VPWR VGND sg13g2_decap_8
XFILLER_10_501 VPWR VGND sg13g2_decap_8
XFILLER_22_361 VPWR VGND sg13g2_decap_8
XFILLER_41_11 VPWR VGND sg13g2_decap_8
XFILLER_10_578 VPWR VGND sg13g2_decap_8
XFILLER_41_44 VPWR VGND sg13g2_decap_8
XFILLER_1_210 VPWR VGND sg13g2_decap_8
XFILLER_2_711 VPWR VGND sg13g2_decap_8
XFILLER_49_203 VPWR VGND sg13g2_decap_8
XFILLER_2_788 VPWR VGND sg13g2_decap_8
XFILLER_1_287 VPWR VGND sg13g2_decap_8
XFILLER_46_910 VPWR VGND sg13g2_decap_8
XFILLER_18_634 VPWR VGND sg13g2_decap_8
XFILLER_17_133 VPWR VGND sg13g2_decap_8
XFILLER_33_604 VPWR VGND sg13g2_decap_8
XFILLER_45_431 VPWR VGND sg13g2_decap_8
XFILLER_14_851 VPWR VGND sg13g2_decap_8
XFILLER_13_361 VPWR VGND sg13g2_decap_8
XFILLER_32_158 VPWR VGND sg13g2_decap_8
XFILLER_41_681 VPWR VGND sg13g2_decap_8
XFILLER_9_354 VPWR VGND sg13g2_decap_8
XFILLER_5_571 VPWR VGND sg13g2_decap_8
XFILLER_49_770 VPWR VGND sg13g2_decap_8
XFILLER_37_910 VPWR VGND sg13g2_decap_8
XFILLER_48_280 VPWR VGND sg13g2_decap_8
XFILLER_36_431 VPWR VGND sg13g2_decap_8
XFILLER_23_158 VPWR VGND sg13g2_decap_8
XFILLER_20_865 VPWR VGND sg13g2_decap_8
XFILLER_11_25 VPWR VGND sg13g2_decap_8
XFILLER_3_508 VPWR VGND sg13g2_decap_8
XFILLER_47_707 VPWR VGND sg13g2_decap_8
XFILLER_46_217 VPWR VGND sg13g2_decap_8
XFILLER_27_420 VPWR VGND sg13g2_decap_8
XFILLER_36_11 VPWR VGND sg13g2_decap_8
XFILLER_39_280 VPWR VGND sg13g2_decap_8
XFILLER_36_88 VPWR VGND sg13g2_decap_8
XFILLER_15_648 VPWR VGND sg13g2_decap_8
XFILLER_27_497 VPWR VGND sg13g2_decap_8
XFILLER_14_158 VPWR VGND sg13g2_decap_8
XFILLER_30_618 VPWR VGND sg13g2_decap_8
XFILLER_42_456 VPWR VGND sg13g2_decap_8
XFILLER_11_865 VPWR VGND sg13g2_decap_8
XFILLER_10_375 VPWR VGND sg13g2_decap_8
XFILLER_7_847 VPWR VGND sg13g2_decap_8
XFILLER_6_368 VPWR VGND sg13g2_decap_8
XFILLER_2_585 VPWR VGND sg13g2_decap_8
X_31_ net10 net2 _02_ VPWR VGND sg13g2_xor2_1
XFILLER_19_921 VPWR VGND sg13g2_decap_4
XFILLER_37_217 VPWR VGND sg13g2_decap_8
XFILLER_18_431 VPWR VGND sg13g2_decap_8
XFILLER_34_902 VPWR VGND sg13g2_decap_8
XFILLER_46_784 VPWR VGND sg13g2_decap_8
XFILLER_33_401 VPWR VGND sg13g2_decap_8
XFILLER_33_478 VPWR VGND sg13g2_decap_8
XFILLER_9_151 VPWR VGND sg13g2_decap_8
XFILLER_47_0 VPWR VGND sg13g2_decap_8
XFILLER_3_81 VPWR VGND sg13g2_decap_8
XFILLER_25_902 VPWR VGND sg13g2_decap_8
XFILLER_37_784 VPWR VGND sg13g2_decap_8
XFILLER_24_467 VPWR VGND sg13g2_decap_8
XFILLER_20_662 VPWR VGND sg13g2_decap_8
XFILLER_22_46 VPWR VGND sg13g2_decap_8
XFILLER_3_305 VPWR VGND sg13g2_decap_8
XFILLER_47_504 VPWR VGND sg13g2_decap_8
XFILLER_47_21 VPWR VGND sg13g2_decap_8
XFILLER_19_228 VPWR VGND sg13g2_decap_8
XFILLER_47_98 VPWR VGND sg13g2_decap_8
XFILLER_28_762 VPWR VGND sg13g2_decap_8
XFILLER_34_209 VPWR VGND sg13g2_decap_8
XFILLER_15_445 VPWR VGND sg13g2_decap_8
XFILLER_27_294 VPWR VGND sg13g2_decap_8
XFILLER_43_732 VPWR VGND sg13g2_decap_8
XFILLER_42_253 VPWR VGND sg13g2_decap_8
XFILLER_30_415 VPWR VGND sg13g2_decap_8
XFILLER_11_662 VPWR VGND sg13g2_decap_8
XFILLER_10_172 VPWR VGND sg13g2_decap_8
XFILLER_7_644 VPWR VGND sg13g2_decap_8
XFILLER_6_165 VPWR VGND sg13g2_decap_8
XFILLER_3_872 VPWR VGND sg13g2_decap_8
XFILLER_2_382 VPWR VGND sg13g2_decap_8
XFILLER_19_4 VPWR VGND sg13g2_decap_8
XFILLER_38_537 VPWR VGND sg13g2_decap_8
XFILLER_25_209 VPWR VGND sg13g2_decap_8
XFILLER_46_581 VPWR VGND sg13g2_decap_8
XFILLER_19_795 VPWR VGND sg13g2_decap_8
XFILLER_34_776 VPWR VGND sg13g2_decap_8
XFILLER_33_275 VPWR VGND sg13g2_decap_8
XFILLER_21_459 VPWR VGND sg13g2_decap_8
XFILLER_0_308 VPWR VGND sg13g2_decap_8
XFILLER_29_537 VPWR VGND sg13g2_decap_8
XFILLER_17_35 VPWR VGND sg13g2_decap_8
XFILLER_44_529 VPWR VGND sg13g2_decap_8
XFILLER_37_581 VPWR VGND sg13g2_decap_8
XFILLER_25_776 VPWR VGND sg13g2_decap_8
XFILLER_24_264 VPWR VGND sg13g2_decap_8
XFILLER_40_746 VPWR VGND sg13g2_decap_8
XFILLER_12_459 VPWR VGND sg13g2_decap_8
XFILLER_3_102 VPWR VGND sg13g2_decap_8
XFILLER_4_669 VPWR VGND sg13g2_decap_8
XFILLER_3_179 VPWR VGND sg13g2_decap_8
XFILLER_0_875 VPWR VGND sg13g2_decap_8
XFILLER_47_301 VPWR VGND sg13g2_decap_8
XFILLER_48_868 VPWR VGND sg13g2_decap_8
XFILLER_47_378 VPWR VGND sg13g2_decap_8
XFILLER_16_732 VPWR VGND sg13g2_decap_8
XFILLER_15_242 VPWR VGND sg13g2_decap_8
XFILLER_30_212 VPWR VGND sg13g2_decap_8
XFILLER_31_724 VPWR VGND sg13g2_decap_8
XFILLER_30_289 VPWR VGND sg13g2_decap_8
XFILLER_7_441 VPWR VGND sg13g2_decap_8
XFILLER_38_334 VPWR VGND sg13g2_decap_8
XFILLER_39_868 VPWR VGND sg13g2_decap_8
XFILLER_26_529 VPWR VGND sg13g2_decap_8
XFILLER_19_592 VPWR VGND sg13g2_decap_8
XFILLER_34_573 VPWR VGND sg13g2_decap_8
XFILLER_22_746 VPWR VGND sg13g2_decap_8
XFILLER_21_256 VPWR VGND sg13g2_decap_8
XFILLER_0_105 VPWR VGND sg13g2_decap_8
XFILLER_29_334 VPWR VGND sg13g2_decap_8
XFILLER_17_518 VPWR VGND sg13g2_decap_8
XFILLER_28_67 VPWR VGND sg13g2_decap_8
XFILLER_45_816 VPWR VGND sg13g2_decap_8
XFILLER_44_326 VPWR VGND sg13g2_decap_8
XFILLER_44_11 VPWR VGND sg13g2_decap_8
XFILLER_25_573 VPWR VGND sg13g2_decap_8
XFILLER_13_746 VPWR VGND sg13g2_decap_8
XFILLER_40_543 VPWR VGND sg13g2_decap_8
XFILLER_44_88 VPWR VGND sg13g2_decap_8
XFILLER_9_739 VPWR VGND sg13g2_decap_8
XFILLER_12_256 VPWR VGND sg13g2_decap_8
XFILLER_8_249 VPWR VGND sg13g2_decap_8
XFILLER_4_466 VPWR VGND sg13g2_decap_8
XFILLER_0_672 VPWR VGND sg13g2_decap_8
XFILLER_48_665 VPWR VGND sg13g2_decap_8
XFILLER_36_816 VPWR VGND sg13g2_decap_8
XFILLER_47_175 VPWR VGND sg13g2_decap_8
XFILLER_35_359 VPWR VGND sg13g2_decap_8
XFILLER_44_893 VPWR VGND sg13g2_decap_8
XFILLER_31_521 VPWR VGND sg13g2_decap_8
XFILLER_31_598 VPWR VGND sg13g2_decap_8
XFILLER_27_805 VPWR VGND sg13g2_decap_8
XFILLER_38_131 VPWR VGND sg13g2_decap_8
XFILLER_39_665 VPWR VGND sg13g2_decap_8
XFILLER_26_326 VPWR VGND sg13g2_decap_8
XFILLER_34_370 VPWR VGND sg13g2_decap_8
XFILLER_14_25 VPWR VGND sg13g2_decap_8
XFILLER_22_543 VPWR VGND sg13g2_decap_8
XFILLER_30_24 VPWR VGND sg13g2_decap_8
XFILLER_30_35 VPWR VGND sg13g2_fill_1
XFILLER_30_68 VPWR VGND sg13g2_decap_8
XFILLER_39_11 VPWR VGND sg13g2_decap_8
XFILLER_1_469 VPWR VGND sg13g2_decap_8
XFILLER_39_77 VPWR VGND sg13g2_decap_8
XFILLER_18_816 VPWR VGND sg13g2_decap_8
XFILLER_29_131 VPWR VGND sg13g2_decap_8
XFILLER_45_613 VPWR VGND sg13g2_decap_8
XFILLER_17_315 VPWR VGND sg13g2_decap_8
XFILLER_44_123 VPWR VGND sg13g2_decap_8
XFILLER_25_370 VPWR VGND sg13g2_decap_8
XFILLER_26_893 VPWR VGND sg13g2_decap_8
XFILLER_13_543 VPWR VGND sg13g2_decap_8
XFILLER_40_340 VPWR VGND sg13g2_decap_8
XFILLER_41_863 VPWR VGND sg13g2_decap_8
XFILLER_9_536 VPWR VGND sg13g2_decap_8
XFILLER_5_753 VPWR VGND sg13g2_decap_8
XFILLER_4_263 VPWR VGND sg13g2_decap_8
XFILLER_48_462 VPWR VGND sg13g2_decap_8
XFILLER_36_613 VPWR VGND sg13g2_decap_8
XFILLER_35_156 VPWR VGND sg13g2_decap_8
XFILLER_17_882 VPWR VGND sg13g2_decap_8
XFILLER_32_830 VPWR VGND sg13g2_decap_8
XFILLER_44_690 VPWR VGND sg13g2_decap_8
XFILLER_31_395 VPWR VGND sg13g2_decap_8
XFILLER_6_81 VPWR VGND sg13g2_decap_8
XFILLER_27_602 VPWR VGND sg13g2_decap_8
XFILLER_39_462 VPWR VGND sg13g2_decap_8
XFILLER_26_123 VPWR VGND sg13g2_decap_8
XFILLER_27_679 VPWR VGND sg13g2_decap_8
XFILLER_42_638 VPWR VGND sg13g2_decap_8
XFILLER_23_830 VPWR VGND sg13g2_decap_8
XFILLER_25_46 VPWR VGND sg13g2_decap_8
XFILLER_22_340 VPWR VGND sg13g2_decap_8
XFILLER_10_557 VPWR VGND sg13g2_decap_8
XFILLER_2_767 VPWR VGND sg13g2_decap_8
XFILLER_1_266 VPWR VGND sg13g2_decap_8
XFILLER_2_39 VPWR VGND sg13g2_decap_8
XFILLER_49_259 VPWR VGND sg13g2_decap_8
XFILLER_17_112 VPWR VGND sg13g2_decap_8
XFILLER_18_613 VPWR VGND sg13g2_decap_8
XFILLER_45_410 VPWR VGND sg13g2_decap_8
XFILLER_45_487 VPWR VGND sg13g2_decap_8
XFILLER_14_830 VPWR VGND sg13g2_decap_8
XFILLER_17_189 VPWR VGND sg13g2_decap_8
XFILLER_26_690 VPWR VGND sg13g2_decap_8
XFILLER_32_137 VPWR VGND sg13g2_decap_8
XFILLER_13_340 VPWR VGND sg13g2_decap_8
XFILLER_41_660 VPWR VGND sg13g2_decap_8
XFILLER_9_333 VPWR VGND sg13g2_decap_8
XFILLER_5_550 VPWR VGND sg13g2_decap_8
XFILLER_36_410 VPWR VGND sg13g2_decap_8
XFILLER_36_487 VPWR VGND sg13g2_decap_8
XFILLER_23_137 VPWR VGND sg13g2_decap_8
XFILLER_24_649 VPWR VGND sg13g2_decap_8
XFILLER_20_844 VPWR VGND sg13g2_decap_8
XFILLER_31_192 VPWR VGND sg13g2_decap_8
XFILLER_15_627 VPWR VGND sg13g2_decap_8
XFILLER_27_476 VPWR VGND sg13g2_decap_8
XFILLER_36_67 VPWR VGND sg13g2_decap_8
XFILLER_43_914 VPWR VGND sg13g2_decap_8
XFILLER_14_137 VPWR VGND sg13g2_decap_8
XFILLER_42_435 VPWR VGND sg13g2_decap_8
XFILLER_11_844 VPWR VGND sg13g2_decap_8
XFILLER_10_354 VPWR VGND sg13g2_decap_8
XFILLER_7_826 VPWR VGND sg13g2_decap_8
XFILLER_6_347 VPWR VGND sg13g2_decap_8
XFILLER_7_0 VPWR VGND sg13g2_decap_8
XFILLER_2_564 VPWR VGND sg13g2_decap_8
XFILLER_19_900 VPWR VGND sg13g2_decap_8
X_30_ net2 net10 _01_ VPWR VGND sg13g2_and2_1
XFILLER_38_719 VPWR VGND sg13g2_decap_8
XFILLER_18_410 VPWR VGND sg13g2_decap_8
XFILLER_46_763 VPWR VGND sg13g2_decap_8
XFILLER_18_487 VPWR VGND sg13g2_decap_8
XFILLER_45_284 VPWR VGND sg13g2_decap_8
XFILLER_33_457 VPWR VGND sg13g2_decap_8
XFILLER_9_130 VPWR VGND sg13g2_decap_8
XFILLER_3_60 VPWR VGND sg13g2_decap_8
XFILLER_29_719 VPWR VGND sg13g2_decap_8
XFILLER_37_763 VPWR VGND sg13g2_decap_8
XFILLER_36_284 VPWR VGND sg13g2_decap_8
XFILLER_24_446 VPWR VGND sg13g2_decap_8
XFILLER_20_641 VPWR VGND sg13g2_decap_8
XFILLER_22_25 VPWR VGND sg13g2_decap_8
XFILLER_0_7 VPWR VGND sg13g2_decap_8
XFILLER_19_207 VPWR VGND sg13g2_decap_8
XFILLER_47_77 VPWR VGND sg13g2_decap_8
XFILLER_28_741 VPWR VGND sg13g2_decap_8
XFILLER_16_914 VPWR VGND sg13g2_decap_8
XFILLER_43_711 VPWR VGND sg13g2_decap_8
XFILLER_15_424 VPWR VGND sg13g2_decap_8
XFILLER_27_273 VPWR VGND sg13g2_decap_8
XFILLER_31_906 VPWR VGND sg13g2_decap_8
XFILLER_42_232 VPWR VGND sg13g2_decap_8
XFILLER_43_788 VPWR VGND sg13g2_decap_8
XFILLER_11_641 VPWR VGND sg13g2_decap_8
XFILLER_10_151 VPWR VGND sg13g2_decap_8
XFILLER_7_623 VPWR VGND sg13g2_decap_8
XFILLER_6_144 VPWR VGND sg13g2_decap_8
XFILLER_3_851 VPWR VGND sg13g2_decap_8
XFILLER_2_361 VPWR VGND sg13g2_decap_8
XFILLER_38_516 VPWR VGND sg13g2_decap_8
XFILLER_46_560 VPWR VGND sg13g2_decap_8
XFILLER_19_774 VPWR VGND sg13g2_decap_8
XFILLER_18_284 VPWR VGND sg13g2_decap_8
XFILLER_33_254 VPWR VGND sg13g2_decap_8
XFILLER_34_755 VPWR VGND sg13g2_decap_8
XFILLER_21_438 VPWR VGND sg13g2_decap_8
XFILLER_29_516 VPWR VGND sg13g2_decap_8
XFILLER_17_14 VPWR VGND sg13g2_decap_8
XFILLER_37_560 VPWR VGND sg13g2_decap_8
XFILLER_44_508 VPWR VGND sg13g2_decap_8
XFILLER_24_243 VPWR VGND sg13g2_decap_8
XFILLER_25_755 VPWR VGND sg13g2_decap_8
XFILLER_40_725 VPWR VGND sg13g2_decap_8
XFILLER_12_438 VPWR VGND sg13g2_decap_8
XFILLER_33_79 VPWR VGND sg13g2_decap_8
XFILLER_4_648 VPWR VGND sg13g2_decap_8
XFILLER_3_158 VPWR VGND sg13g2_decap_8
XFILLER_0_854 VPWR VGND sg13g2_decap_8
XFILLER_48_847 VPWR VGND sg13g2_decap_8
XFILLER_47_357 VPWR VGND sg13g2_decap_8
XFILLER_16_711 VPWR VGND sg13g2_decap_8
XFILLER_15_221 VPWR VGND sg13g2_decap_8
XFILLER_31_703 VPWR VGND sg13g2_decap_8
XFILLER_16_788 VPWR VGND sg13g2_decap_8
XFILLER_43_585 VPWR VGND sg13g2_decap_8
XFILLER_15_298 VPWR VGND sg13g2_decap_8
XFILLER_8_921 VPWR VGND sg13g2_decap_4
XFILLER_30_268 VPWR VGND sg13g2_decap_8
XFILLER_7_420 VPWR VGND sg13g2_decap_8
XFILLER_7_497 VPWR VGND sg13g2_decap_8
XFILLER_31_4 VPWR VGND sg13g2_decap_8
XFILLER_38_313 VPWR VGND sg13g2_decap_8
XFILLER_39_847 VPWR VGND sg13g2_decap_8
XFILLER_26_508 VPWR VGND sg13g2_decap_8
XFILLER_19_571 VPWR VGND sg13g2_decap_8
XFILLER_34_552 VPWR VGND sg13g2_decap_8
XFILLER_22_725 VPWR VGND sg13g2_decap_8
XFILLER_21_235 VPWR VGND sg13g2_decap_8
XFILLER_9_81 VPWR VGND sg13g2_decap_8
XFILLER_28_46 VPWR VGND sg13g2_decap_8
XFILLER_29_313 VPWR VGND sg13g2_decap_8
XFILLER_44_305 VPWR VGND sg13g2_decap_8
XFILLER_38_880 VPWR VGND sg13g2_decap_8
XFILLER_25_552 VPWR VGND sg13g2_decap_8
XFILLER_13_725 VPWR VGND sg13g2_decap_8
XFILLER_44_67 VPWR VGND sg13g2_decap_8
XFILLER_9_718 VPWR VGND sg13g2_decap_8
XFILLER_12_235 VPWR VGND sg13g2_decap_8
XFILLER_40_522 VPWR VGND sg13g2_decap_8
XFILLER_8_228 VPWR VGND sg13g2_decap_8
XFILLER_40_599 VPWR VGND sg13g2_decap_8
XFILLER_5_39 VPWR VGND sg13g2_decap_8
XFILLER_4_445 VPWR VGND sg13g2_decap_8
XFILLER_0_651 VPWR VGND sg13g2_decap_8
XFILLER_48_644 VPWR VGND sg13g2_decap_8
XFILLER_47_154 VPWR VGND sg13g2_decap_8
XFILLER_29_880 VPWR VGND sg13g2_decap_8
XFILLER_35_338 VPWR VGND sg13g2_decap_8
XFILLER_16_585 VPWR VGND sg13g2_decap_8
XFILLER_31_500 VPWR VGND sg13g2_decap_8
XFILLER_44_872 VPWR VGND sg13g2_decap_8
XFILLER_43_382 VPWR VGND sg13g2_decap_8
XFILLER_31_577 VPWR VGND sg13g2_decap_8
XFILLER_8_795 VPWR VGND sg13g2_decap_8
XFILLER_7_294 VPWR VGND sg13g2_decap_8
XFILLER_38_110 VPWR VGND sg13g2_decap_8
XFILLER_39_644 VPWR VGND sg13g2_decap_8
XFILLER_26_305 VPWR VGND sg13g2_decap_8
XFILLER_38_187 VPWR VGND sg13g2_decap_8
XFILLER_22_522 VPWR VGND sg13g2_decap_8
XFILLER_10_739 VPWR VGND sg13g2_decap_8
XFILLER_22_599 VPWR VGND sg13g2_decap_8
XFILLER_30_47 VPWR VGND sg13g2_decap_8
XFILLER_1_448 VPWR VGND sg13g2_decap_8
XFILLER_39_56 VPWR VGND sg13g2_decap_8
XFILLER_29_187 VPWR VGND sg13g2_decap_8
XFILLER_44_102 VPWR VGND sg13g2_decap_8
XFILLER_45_669 VPWR VGND sg13g2_decap_8
XFILLER_26_872 VPWR VGND sg13g2_decap_8
XFILLER_32_319 VPWR VGND sg13g2_decap_8
XFILLER_44_179 VPWR VGND sg13g2_decap_8
XFILLER_13_522 VPWR VGND sg13g2_decap_8
XFILLER_41_842 VPWR VGND sg13g2_decap_8
XFILLER_9_515 VPWR VGND sg13g2_decap_8
XFILLER_13_599 VPWR VGND sg13g2_decap_8
XFILLER_40_396 VPWR VGND sg13g2_decap_8
XFILLER_5_732 VPWR VGND sg13g2_decap_8
XFILLER_4_242 VPWR VGND sg13g2_decap_8
XFILLER_48_441 VPWR VGND sg13g2_decap_8
XFILLER_35_102 VPWR VGND sg13g2_decap_8
XFILLER_35_135 VPWR VGND sg13g2_decap_8
XFILLER_36_669 VPWR VGND sg13g2_decap_8
XFILLER_17_861 VPWR VGND sg13g2_decap_8
XFILLER_23_319 VPWR VGND sg13g2_decap_8
XFILLER_16_382 VPWR VGND sg13g2_decap_8
XFILLER_32_886 VPWR VGND sg13g2_decap_8
XFILLER_31_374 VPWR VGND sg13g2_decap_8
XFILLER_8_592 VPWR VGND sg13g2_decap_8
XFILLER_6_60 VPWR VGND sg13g2_decap_8
XFILLER_39_441 VPWR VGND sg13g2_decap_8
XFILLER_26_102 VPWR VGND sg13g2_decap_8
XFILLER_15_809 VPWR VGND sg13g2_decap_8
XFILLER_27_658 VPWR VGND sg13g2_decap_8
XFILLER_14_319 VPWR VGND sg13g2_decap_8
XFILLER_25_25 VPWR VGND sg13g2_decap_8
XFILLER_26_179 VPWR VGND sg13g2_decap_8
XFILLER_42_617 VPWR VGND sg13g2_decap_8
XFILLER_41_149 VPWR VGND sg13g2_decap_8
XFILLER_23_886 VPWR VGND sg13g2_decap_8
XFILLER_10_536 VPWR VGND sg13g2_decap_8
XFILLER_22_396 VPWR VGND sg13g2_decap_8
XFILLER_6_529 VPWR VGND sg13g2_decap_8
XFILLER_41_79 VPWR VGND sg13g2_decap_8
XFILLER_9_4 VPWR VGND sg13g2_decap_8
XFILLER_2_746 VPWR VGND sg13g2_decap_8
XFILLER_1_245 VPWR VGND sg13g2_decap_8
XFILLER_49_238 VPWR VGND sg13g2_decap_8
XFILLER_2_18 VPWR VGND sg13g2_decap_8
XFILLER_18_669 VPWR VGND sg13g2_decap_8
XFILLER_17_168 VPWR VGND sg13g2_decap_8
XFILLER_45_466 VPWR VGND sg13g2_decap_8
XFILLER_32_116 VPWR VGND sg13g2_decap_4
XFILLER_33_639 VPWR VGND sg13g2_decap_8
XFILLER_9_312 VPWR VGND sg13g2_decap_8
XFILLER_14_886 VPWR VGND sg13g2_decap_8
XFILLER_13_396 VPWR VGND sg13g2_decap_8
XFILLER_40_193 VPWR VGND sg13g2_decap_8
XFILLER_9_389 VPWR VGND sg13g2_decap_8
XFILLER_24_628 VPWR VGND sg13g2_decap_8
XFILLER_36_466 VPWR VGND sg13g2_decap_8
XFILLER_23_116 VPWR VGND sg13g2_decap_8
XFILLER_20_823 VPWR VGND sg13g2_decap_8
XFILLER_32_683 VPWR VGND sg13g2_decap_8
XFILLER_31_171 VPWR VGND sg13g2_decap_8
XFILLER_28_923 VPWR VGND sg13g2_fill_2
XFILLER_36_46 VPWR VGND sg13g2_decap_8
XFILLER_15_606 VPWR VGND sg13g2_decap_8
XFILLER_27_455 VPWR VGND sg13g2_decap_8
XFILLER_14_116 VPWR VGND sg13g2_decap_8
XFILLER_42_414 VPWR VGND sg13g2_decap_8
XFILLER_11_823 VPWR VGND sg13g2_decap_8
XFILLER_23_683 VPWR VGND sg13g2_decap_8
XFILLER_10_333 VPWR VGND sg13g2_decap_8
XFILLER_7_805 VPWR VGND sg13g2_decap_8
XFILLER_22_193 VPWR VGND sg13g2_decap_8
XFILLER_6_326 VPWR VGND sg13g2_decap_8
XFILLER_2_543 VPWR VGND sg13g2_decap_8
XFILLER_46_742 VPWR VGND sg13g2_decap_8
XFILLER_18_466 VPWR VGND sg13g2_decap_8
XFILLER_45_263 VPWR VGND sg13g2_decap_8
XFILLER_33_436 VPWR VGND sg13g2_decap_8
XFILLER_14_683 VPWR VGND sg13g2_decap_8
XFILLER_13_193 VPWR VGND sg13g2_decap_8
XFILLER_9_186 VPWR VGND sg13g2_decap_8
XFILLER_6_893 VPWR VGND sg13g2_decap_8
XFILLER_37_742 VPWR VGND sg13g2_decap_8
XFILLER_24_425 VPWR VGND sg13g2_decap_8
XFILLER_36_263 VPWR VGND sg13g2_decap_8
XFILLER_40_907 VPWR VGND sg13g2_decap_8
XFILLER_20_620 VPWR VGND sg13g2_decap_8
XFILLER_32_480 VPWR VGND sg13g2_decap_8
XFILLER_20_697 VPWR VGND sg13g2_decap_8
XFILLER_47_539 VPWR VGND sg13g2_decap_8
XFILLER_47_56 VPWR VGND sg13g2_decap_8
XFILLER_28_720 VPWR VGND sg13g2_decap_8
XFILLER_27_252 VPWR VGND sg13g2_decap_8
XFILLER_15_403 VPWR VGND sg13g2_decap_8
XFILLER_28_797 VPWR VGND sg13g2_decap_8
XFILLER_42_211 VPWR VGND sg13g2_decap_8
XFILLER_43_767 VPWR VGND sg13g2_decap_8
XFILLER_42_288 VPWR VGND sg13g2_decap_8
XFILLER_8_39 VPWR VGND sg13g2_decap_8
XFILLER_11_620 VPWR VGND sg13g2_decap_8
XFILLER_23_480 VPWR VGND sg13g2_decap_8
XFILLER_10_130 VPWR VGND sg13g2_decap_8
XFILLER_7_602 VPWR VGND sg13g2_decap_8
XFILLER_6_123 VPWR VGND sg13g2_decap_8
XFILLER_11_697 VPWR VGND sg13g2_decap_8
XFILLER_7_679 VPWR VGND sg13g2_decap_8
XFILLER_12_81 VPWR VGND sg13g2_decap_8
XFILLER_3_830 VPWR VGND sg13g2_decap_8
XFILLER_2_340 VPWR VGND sg13g2_decap_8
XFILLER_19_753 VPWR VGND sg13g2_decap_8
XFILLER_18_263 VPWR VGND sg13g2_decap_8
XFILLER_34_734 VPWR VGND sg13g2_decap_8
XFILLER_22_907 VPWR VGND sg13g2_decap_8
XFILLER_33_233 VPWR VGND sg13g2_decap_8
XFILLER_21_417 VPWR VGND sg13g2_decap_8
XFILLER_14_480 VPWR VGND sg13g2_decap_8
XFILLER_6_690 VPWR VGND sg13g2_decap_8
XFILLER_25_734 VPWR VGND sg13g2_decap_8
XFILLER_13_907 VPWR VGND sg13g2_decap_8
XFILLER_24_222 VPWR VGND sg13g2_decap_8
XFILLER_12_417 VPWR VGND sg13g2_decap_8
XFILLER_33_25 VPWR VGND sg13g2_decap_4
XFILLER_40_704 VPWR VGND sg13g2_decap_8
XFILLER_24_299 VPWR VGND sg13g2_decap_8
XFILLER_33_58 VPWR VGND sg13g2_decap_8
XFILLER_20_494 VPWR VGND sg13g2_decap_8
XFILLER_4_627 VPWR VGND sg13g2_decap_8
XFILLER_3_137 VPWR VGND sg13g2_decap_8
XFILLER_0_833 VPWR VGND sg13g2_decap_8
XFILLER_48_826 VPWR VGND sg13g2_decap_8
XFILLER_47_336 VPWR VGND sg13g2_decap_8
XFILLER_15_200 VPWR VGND sg13g2_decap_8
XFILLER_28_594 VPWR VGND sg13g2_decap_8
XFILLER_16_767 VPWR VGND sg13g2_decap_8
XFILLER_15_277 VPWR VGND sg13g2_decap_8
XFILLER_43_564 VPWR VGND sg13g2_decap_8
XFILLER_31_759 VPWR VGND sg13g2_decap_8
XFILLER_8_900 VPWR VGND sg13g2_decap_8
XFILLER_30_247 VPWR VGND sg13g2_decap_8
XFILLER_11_494 VPWR VGND sg13g2_decap_8
XFILLER_7_476 VPWR VGND sg13g2_decap_8
XFILLER_24_4 VPWR VGND sg13g2_decap_8
XFILLER_39_826 VPWR VGND sg13g2_decap_8
XFILLER_19_550 VPWR VGND sg13g2_decap_8
XFILLER_38_369 VPWR VGND sg13g2_decap_8
XFILLER_0_84 VPWR VGND sg13g2_decap_8
XFILLER_34_531 VPWR VGND sg13g2_decap_8
XFILLER_22_704 VPWR VGND sg13g2_decap_8
XFILLER_21_214 VPWR VGND sg13g2_decap_8
XFILLER_9_60 VPWR VGND sg13g2_decap_8
XFILLER_28_25 VPWR VGND sg13g2_decap_8
XFILLER_29_369 VPWR VGND sg13g2_decap_8
XFILLER_25_531 VPWR VGND sg13g2_decap_8
XFILLER_13_704 VPWR VGND sg13g2_decap_8
XFILLER_40_501 VPWR VGND sg13g2_decap_8
XFILLER_44_46 VPWR VGND sg13g2_decap_8
XFILLER_12_214 VPWR VGND sg13g2_decap_8
XFILLER_8_207 VPWR VGND sg13g2_decap_8
XFILLER_40_578 VPWR VGND sg13g2_decap_8
XFILLER_21_781 VPWR VGND sg13g2_decap_8
XFILLER_5_914 VPWR VGND sg13g2_decap_8
XFILLER_20_291 VPWR VGND sg13g2_decap_8
XFILLER_5_18 VPWR VGND sg13g2_decap_8
XFILLER_4_424 VPWR VGND sg13g2_decap_8
XFILLER_0_630 VPWR VGND sg13g2_decap_8
XFILLER_48_623 VPWR VGND sg13g2_decap_8
XFILLER_47_133 VPWR VGND sg13g2_decap_8
XFILLER_35_317 VPWR VGND sg13g2_decap_8
XFILLER_28_391 VPWR VGND sg13g2_decap_8
XFILLER_44_851 VPWR VGND sg13g2_decap_8
XFILLER_16_564 VPWR VGND sg13g2_decap_8
XFILLER_43_361 VPWR VGND sg13g2_decap_8
XFILLER_31_556 VPWR VGND sg13g2_decap_8
XFILLER_12_781 VPWR VGND sg13g2_decap_8
XFILLER_11_291 VPWR VGND sg13g2_decap_8
XFILLER_8_774 VPWR VGND sg13g2_decap_8
XFILLER_7_273 VPWR VGND sg13g2_decap_8
XFILLER_39_623 VPWR VGND sg13g2_decap_8
XFILLER_38_166 VPWR VGND sg13g2_decap_8
XFILLER_22_501 VPWR VGND sg13g2_decap_8
XFILLER_35_884 VPWR VGND sg13g2_decap_8
XFILLER_10_718 VPWR VGND sg13g2_decap_8
XFILLER_22_578 VPWR VGND sg13g2_decap_8
XFILLER_1_427 VPWR VGND sg13g2_decap_8
XFILLER_39_35 VPWR VGND sg13g2_decap_8
XFILLER_29_166 VPWR VGND sg13g2_decap_8
XFILLER_26_851 VPWR VGND sg13g2_decap_8
XFILLER_45_648 VPWR VGND sg13g2_decap_8
XFILLER_13_501 VPWR VGND sg13g2_decap_8
XFILLER_44_158 VPWR VGND sg13g2_decap_8
XFILLER_41_821 VPWR VGND sg13g2_decap_8
XFILLER_13_578 VPWR VGND sg13g2_decap_8
XFILLER_40_375 VPWR VGND sg13g2_decap_8
XFILLER_41_898 VPWR VGND sg13g2_decap_8
XFILLER_5_711 VPWR VGND sg13g2_decap_8
XFILLER_4_221 VPWR VGND sg13g2_decap_8
XFILLER_5_788 VPWR VGND sg13g2_decap_8
XFILLER_4_298 VPWR VGND sg13g2_decap_8
XFILLER_20_81 VPWR VGND sg13g2_decap_8
XFILLER_49_910 VPWR VGND sg13g2_decap_8
XFILLER_48_420 VPWR VGND sg13g2_decap_8
XFILLER_48_497 VPWR VGND sg13g2_decap_8
XFILLER_17_840 VPWR VGND sg13g2_decap_8
XFILLER_35_114 VPWR VGND sg13g2_decap_8
XFILLER_36_648 VPWR VGND sg13g2_decap_8
XFILLER_16_361 VPWR VGND sg13g2_decap_8
XFILLER_31_353 VPWR VGND sg13g2_decap_8
XFILLER_32_865 VPWR VGND sg13g2_decap_8
XFILLER_8_571 VPWR VGND sg13g2_decap_8
XFILLER_39_420 VPWR VGND sg13g2_decap_8
XFILLER_27_637 VPWR VGND sg13g2_decap_8
XFILLER_39_497 VPWR VGND sg13g2_decap_8
XFILLER_26_158 VPWR VGND sg13g2_decap_8
XFILLER_35_681 VPWR VGND sg13g2_decap_8
XFILLER_41_128 VPWR VGND sg13g2_decap_8
XFILLER_23_865 VPWR VGND sg13g2_decap_8
XFILLER_10_515 VPWR VGND sg13g2_decap_8
XFILLER_22_375 VPWR VGND sg13g2_decap_8
XFILLER_6_508 VPWR VGND sg13g2_decap_8
XFILLER_41_25 VPWR VGND sg13g2_decap_8
XFILLER_41_58 VPWR VGND sg13g2_decap_8
XFILLER_1_224 VPWR VGND sg13g2_decap_8
XFILLER_2_725 VPWR VGND sg13g2_decap_8
XFILLER_49_217 VPWR VGND sg13g2_decap_8
XFILLER_46_924 VPWR VGND sg13g2_fill_1
XFILLER_18_648 VPWR VGND sg13g2_decap_8
XFILLER_45_445 VPWR VGND sg13g2_decap_8
XFILLER_17_147 VPWR VGND sg13g2_decap_8
XFILLER_33_618 VPWR VGND sg13g2_decap_8
XFILLER_14_865 VPWR VGND sg13g2_decap_8
XFILLER_13_375 VPWR VGND sg13g2_decap_8
XFILLER_15_81 VPWR VGND sg13g2_decap_8
XFILLER_41_695 VPWR VGND sg13g2_decap_8
XFILLER_9_368 VPWR VGND sg13g2_decap_8
XFILLER_40_172 VPWR VGND sg13g2_decap_8
XFILLER_5_585 VPWR VGND sg13g2_decap_8
XFILLER_1_791 VPWR VGND sg13g2_decap_8
XFILLER_49_784 VPWR VGND sg13g2_decap_8
XFILLER_37_924 VPWR VGND sg13g2_fill_1
XFILLER_48_294 VPWR VGND sg13g2_decap_8
XFILLER_36_445 VPWR VGND sg13g2_decap_8
XFILLER_24_607 VPWR VGND sg13g2_decap_8
XFILLER_20_802 VPWR VGND sg13g2_decap_8
XFILLER_31_150 VPWR VGND sg13g2_decap_8
XFILLER_32_662 VPWR VGND sg13g2_decap_8
XFILLER_20_879 VPWR VGND sg13g2_decap_8
XFILLER_11_39 VPWR VGND sg13g2_decap_8
XFILLER_28_902 VPWR VGND sg13g2_decap_8
XFILLER_27_434 VPWR VGND sg13g2_decap_8
XFILLER_36_25 VPWR VGND sg13g2_decap_8
XFILLER_39_294 VPWR VGND sg13g2_decap_8
XFILLER_11_802 VPWR VGND sg13g2_decap_8
XFILLER_23_662 VPWR VGND sg13g2_decap_8
XFILLER_10_312 VPWR VGND sg13g2_decap_8
XFILLER_22_172 VPWR VGND sg13g2_decap_8
XFILLER_6_305 VPWR VGND sg13g2_decap_8
XFILLER_11_879 VPWR VGND sg13g2_decap_8
XFILLER_10_389 VPWR VGND sg13g2_decap_8
XFILLER_2_522 VPWR VGND sg13g2_decap_8
XFILLER_2_599 VPWR VGND sg13g2_decap_8
XFILLER_46_721 VPWR VGND sg13g2_decap_8
XFILLER_18_445 VPWR VGND sg13g2_decap_8
XFILLER_34_916 VPWR VGND sg13g2_decap_8
XFILLER_45_242 VPWR VGND sg13g2_decap_8
XFILLER_46_798 VPWR VGND sg13g2_decap_8
XFILLER_33_415 VPWR VGND sg13g2_decap_8
XFILLER_14_662 VPWR VGND sg13g2_decap_8
XFILLER_20_109 VPWR VGND sg13g2_decap_8
XFILLER_13_172 VPWR VGND sg13g2_decap_8
XFILLER_41_492 VPWR VGND sg13g2_decap_8
XFILLER_9_165 VPWR VGND sg13g2_decap_8
XFILLER_6_872 VPWR VGND sg13g2_decap_8
XFILLER_5_382 VPWR VGND sg13g2_decap_8
XFILLER_3_95 VPWR VGND sg13g2_decap_8
XFILLER_28_209 VPWR VGND sg13g2_decap_8
XFILLER_49_581 VPWR VGND sg13g2_decap_8
XFILLER_37_721 VPWR VGND sg13g2_decap_8
XFILLER_25_916 VPWR VGND sg13g2_decap_8
XFILLER_36_242 VPWR VGND sg13g2_decap_8
XFILLER_24_404 VPWR VGND sg13g2_decap_8
XFILLER_37_798 VPWR VGND sg13g2_decap_8
XFILLER_11_109 VPWR VGND sg13g2_decap_8
XFILLER_20_676 VPWR VGND sg13g2_decap_8
XFILLER_4_809 VPWR VGND sg13g2_decap_8
XFILLER_3_319 VPWR VGND sg13g2_decap_8
XFILLER_47_518 VPWR VGND sg13g2_decap_8
XFILLER_47_35 VPWR VGND sg13g2_decap_8
XFILLER_27_231 VPWR VGND sg13g2_decap_8
XFILLER_28_776 VPWR VGND sg13g2_decap_8
XFILLER_15_459 VPWR VGND sg13g2_decap_8
XFILLER_43_746 VPWR VGND sg13g2_decap_8
XFILLER_30_429 VPWR VGND sg13g2_decap_8
XFILLER_42_267 VPWR VGND sg13g2_decap_8
XFILLER_8_18 VPWR VGND sg13g2_decap_8
XFILLER_11_676 VPWR VGND sg13g2_decap_8
XFILLER_10_186 VPWR VGND sg13g2_decap_8
XFILLER_7_658 VPWR VGND sg13g2_decap_8
XFILLER_6_102 VPWR VGND sg13g2_decap_8
XFILLER_12_60 VPWR VGND sg13g2_decap_8
XFILLER_6_179 VPWR VGND sg13g2_decap_8
XFILLER_3_886 VPWR VGND sg13g2_decap_8
XFILLER_2_396 VPWR VGND sg13g2_decap_8
XFILLER_19_732 VPWR VGND sg13g2_decap_8
XFILLER_18_242 VPWR VGND sg13g2_decap_8
XFILLER_46_595 VPWR VGND sg13g2_decap_8
XFILLER_33_212 VPWR VGND sg13g2_decap_8
XFILLER_34_713 VPWR VGND sg13g2_decap_8
XFILLER_33_289 VPWR VGND sg13g2_decap_8
XFILLER_17_49 VPWR VGND sg13g2_decap_8
XFILLER_24_201 VPWR VGND sg13g2_decap_8
XFILLER_25_713 VPWR VGND sg13g2_decap_8
XFILLER_37_595 VPWR VGND sg13g2_decap_8
XFILLER_24_278 VPWR VGND sg13g2_decap_8
XFILLER_20_473 VPWR VGND sg13g2_decap_8
XFILLER_4_606 VPWR VGND sg13g2_decap_8
XFILLER_3_116 VPWR VGND sg13g2_decap_8
XFILLER_0_812 VPWR VGND sg13g2_decap_8
XFILLER_48_805 VPWR VGND sg13g2_decap_8
XFILLER_0_889 VPWR VGND sg13g2_decap_8
XFILLER_47_315 VPWR VGND sg13g2_decap_8
XFILLER_28_573 VPWR VGND sg13g2_decap_8
XFILLER_16_746 VPWR VGND sg13g2_decap_8
XFILLER_43_543 VPWR VGND sg13g2_decap_8
XFILLER_15_256 VPWR VGND sg13g2_decap_8
XFILLER_30_226 VPWR VGND sg13g2_decap_8
XFILLER_31_738 VPWR VGND sg13g2_decap_8
XFILLER_11_473 VPWR VGND sg13g2_decap_8
XFILLER_23_81 VPWR VGND sg13g2_decap_8
XFILLER_7_455 VPWR VGND sg13g2_decap_8
XFILLER_3_683 VPWR VGND sg13g2_decap_8
XFILLER_2_193 VPWR VGND sg13g2_decap_8
XFILLER_39_805 VPWR VGND sg13g2_decap_8
XFILLER_38_348 VPWR VGND sg13g2_decap_8
XFILLER_47_882 VPWR VGND sg13g2_decap_8
XFILLER_34_510 VPWR VGND sg13g2_decap_8
XFILLER_46_392 VPWR VGND sg13g2_decap_8
XFILLER_0_63 VPWR VGND sg13g2_decap_8
XFILLER_34_587 VPWR VGND sg13g2_decap_8
XFILLER_30_793 VPWR VGND sg13g2_decap_8
XFILLER_1_609 VPWR VGND sg13g2_decap_8
XFILLER_0_119 VPWR VGND sg13g2_decap_8
XFILLER_29_348 VPWR VGND sg13g2_decap_8
XFILLER_25_510 VPWR VGND sg13g2_decap_8
XFILLER_37_392 VPWR VGND sg13g2_decap_8
XFILLER_44_25 VPWR VGND sg13g2_decap_8
XFILLER_25_587 VPWR VGND sg13g2_decap_8
XFILLER_40_557 VPWR VGND sg13g2_decap_8
XFILLER_21_760 VPWR VGND sg13g2_decap_8
XFILLER_20_270 VPWR VGND sg13g2_decap_8
XFILLER_4_403 VPWR VGND sg13g2_decap_8
XFILLER_48_602 VPWR VGND sg13g2_decap_8
XFILLER_47_112 VPWR VGND sg13g2_decap_8
XFILLER_0_686 VPWR VGND sg13g2_decap_8
XFILLER_48_679 VPWR VGND sg13g2_decap_8
XFILLER_47_189 VPWR VGND sg13g2_decap_8
XFILLER_16_543 VPWR VGND sg13g2_decap_8
XFILLER_18_81 VPWR VGND sg13g2_decap_8
XFILLER_28_370 VPWR VGND sg13g2_decap_8
XFILLER_44_830 VPWR VGND sg13g2_decap_8
XFILLER_43_340 VPWR VGND sg13g2_decap_8
XFILLER_31_535 VPWR VGND sg13g2_decap_8
XFILLER_34_91 VPWR VGND sg13g2_decap_8
XFILLER_12_760 VPWR VGND sg13g2_decap_8
XFILLER_11_270 VPWR VGND sg13g2_decap_8
XFILLER_8_753 VPWR VGND sg13g2_decap_8
XFILLER_7_252 VPWR VGND sg13g2_decap_8
XFILLER_3_480 VPWR VGND sg13g2_decap_8
XFILLER_39_602 VPWR VGND sg13g2_decap_8
XFILLER_27_819 VPWR VGND sg13g2_decap_8
XFILLER_38_145 VPWR VGND sg13g2_decap_8
XFILLER_39_679 VPWR VGND sg13g2_decap_8
XFILLER_35_863 VPWR VGND sg13g2_decap_8
XFILLER_34_384 VPWR VGND sg13g2_decap_8
XFILLER_14_39 VPWR VGND sg13g2_decap_8
XFILLER_22_557 VPWR VGND sg13g2_decap_8
XFILLER_30_590 VPWR VGND sg13g2_decap_8
XFILLER_2_907 VPWR VGND sg13g2_decap_8
XFILLER_1_406 VPWR VGND sg13g2_decap_8
XFILLER_29_145 VPWR VGND sg13g2_decap_8
XFILLER_45_627 VPWR VGND sg13g2_decap_8
XFILLER_17_329 VPWR VGND sg13g2_decap_8
XFILLER_26_830 VPWR VGND sg13g2_decap_8
XFILLER_44_137 VPWR VGND sg13g2_decap_8
XFILLER_41_800 VPWR VGND sg13g2_decap_8
XFILLER_25_384 VPWR VGND sg13g2_decap_8
XFILLER_13_557 VPWR VGND sg13g2_decap_8
XFILLER_41_877 VPWR VGND sg13g2_decap_8
XFILLER_40_354 VPWR VGND sg13g2_decap_8
XFILLER_4_200 VPWR VGND sg13g2_decap_8
XFILLER_5_767 VPWR VGND sg13g2_decap_8
XFILLER_20_60 VPWR VGND sg13g2_decap_8
XFILLER_4_277 VPWR VGND sg13g2_decap_8
XFILLER_0_483 VPWR VGND sg13g2_decap_8
XFILLER_48_476 VPWR VGND sg13g2_decap_8
XFILLER_36_627 VPWR VGND sg13g2_decap_8
XFILLER_16_340 VPWR VGND sg13g2_decap_8
XFILLER_17_896 VPWR VGND sg13g2_decap_8
XFILLER_31_332 VPWR VGND sg13g2_decap_8
XFILLER_32_844 VPWR VGND sg13g2_decap_8
XFILLER_8_550 VPWR VGND sg13g2_decap_8
XFILLER_6_95 VPWR VGND sg13g2_decap_8
XFILLER_27_616 VPWR VGND sg13g2_decap_8
XFILLER_39_476 VPWR VGND sg13g2_decap_8
XFILLER_26_137 VPWR VGND sg13g2_decap_8
XFILLER_35_660 VPWR VGND sg13g2_decap_8
XFILLER_41_107 VPWR VGND sg13g2_decap_8
XFILLER_23_844 VPWR VGND sg13g2_decap_8
XFILLER_34_181 VPWR VGND sg13g2_decap_8
XFILLER_22_354 VPWR VGND sg13g2_decap_8
XFILLER_2_704 VPWR VGND sg13g2_decap_8
XFILLER_1_203 VPWR VGND sg13g2_decap_8
XFILLER_46_903 VPWR VGND sg13g2_decap_8
XFILLER_18_627 VPWR VGND sg13g2_decap_8
XFILLER_17_126 VPWR VGND sg13g2_decap_8
XFILLER_45_424 VPWR VGND sg13g2_decap_8
XFILLER_14_844 VPWR VGND sg13g2_decap_8
XFILLER_25_181 VPWR VGND sg13g2_decap_8
XFILLER_13_354 VPWR VGND sg13g2_decap_8
XFILLER_15_60 VPWR VGND sg13g2_decap_8
XFILLER_40_151 VPWR VGND sg13g2_decap_8
XFILLER_41_674 VPWR VGND sg13g2_decap_8
XFILLER_9_347 VPWR VGND sg13g2_decap_8
XFILLER_5_564 VPWR VGND sg13g2_decap_8
XFILLER_31_81 VPWR VGND sg13g2_decap_8
XFILLER_49_7 VPWR VGND sg13g2_decap_8
XFILLER_1_770 VPWR VGND sg13g2_decap_8
XFILLER_0_280 VPWR VGND sg13g2_decap_8
XFILLER_49_763 VPWR VGND sg13g2_decap_8
XFILLER_37_903 VPWR VGND sg13g2_decap_8
XFILLER_48_273 VPWR VGND sg13g2_decap_8
XFILLER_36_424 VPWR VGND sg13g2_decap_8
XFILLER_17_693 VPWR VGND sg13g2_decap_8
XFILLER_32_641 VPWR VGND sg13g2_decap_8
XFILLER_20_858 VPWR VGND sg13g2_decap_8
XFILLER_11_18 VPWR VGND sg13g2_decap_8
XFILLER_27_413 VPWR VGND sg13g2_decap_8
XFILLER_39_273 VPWR VGND sg13g2_decap_8
XFILLER_23_641 VPWR VGND sg13g2_decap_8
XFILLER_42_449 VPWR VGND sg13g2_decap_8
XFILLER_22_151 VPWR VGND sg13g2_decap_8
XFILLER_11_858 VPWR VGND sg13g2_decap_8
XFILLER_10_368 VPWR VGND sg13g2_decap_8
XFILLER_2_501 VPWR VGND sg13g2_decap_8
XFILLER_2_578 VPWR VGND sg13g2_decap_8
XFILLER_46_700 VPWR VGND sg13g2_decap_8
XFILLER_19_914 VPWR VGND sg13g2_decap_8
XFILLER_18_424 VPWR VGND sg13g2_decap_8
XFILLER_46_777 VPWR VGND sg13g2_decap_8
XFILLER_45_221 VPWR VGND sg13g2_decap_8
XFILLER_14_641 VPWR VGND sg13g2_decap_8
XFILLER_45_298 VPWR VGND sg13g2_decap_8
XFILLER_13_151 VPWR VGND sg13g2_decap_8
XFILLER_41_471 VPWR VGND sg13g2_decap_8
XFILLER_9_144 VPWR VGND sg13g2_decap_8
XFILLER_6_851 VPWR VGND sg13g2_decap_8
XFILLER_5_361 VPWR VGND sg13g2_decap_8
XFILLER_3_74 VPWR VGND sg13g2_decap_8
XFILLER_49_560 VPWR VGND sg13g2_decap_8
XFILLER_37_700 VPWR VGND sg13g2_decap_8
XFILLER_36_221 VPWR VGND sg13g2_decap_8
XFILLER_37_777 VPWR VGND sg13g2_decap_8
XFILLER_17_490 VPWR VGND sg13g2_decap_8
XFILLER_36_298 VPWR VGND sg13g2_decap_8
XFILLER_20_655 VPWR VGND sg13g2_decap_8
XFILLER_22_39 VPWR VGND sg13g2_decap_8
XFILLER_47_14 VPWR VGND sg13g2_decap_8
XFILLER_27_210 VPWR VGND sg13g2_decap_8
XFILLER_28_755 VPWR VGND sg13g2_decap_8
XFILLER_43_725 VPWR VGND sg13g2_decap_8
XFILLER_15_438 VPWR VGND sg13g2_decap_8
XFILLER_27_287 VPWR VGND sg13g2_decap_8
XFILLER_42_246 VPWR VGND sg13g2_decap_8
XFILLER_30_408 VPWR VGND sg13g2_decap_8
XFILLER_11_655 VPWR VGND sg13g2_decap_8
XFILLER_10_165 VPWR VGND sg13g2_decap_8
XFILLER_7_637 VPWR VGND sg13g2_decap_8
XFILLER_6_158 VPWR VGND sg13g2_decap_8
XFILLER_3_865 VPWR VGND sg13g2_decap_8
XFILLER_2_375 VPWR VGND sg13g2_decap_8
XFILLER_19_711 VPWR VGND sg13g2_decap_8
XFILLER_18_221 VPWR VGND sg13g2_decap_8
XFILLER_46_574 VPWR VGND sg13g2_decap_8
XFILLER_19_788 VPWR VGND sg13g2_decap_8
XFILLER_37_91 VPWR VGND sg13g2_decap_8
XFILLER_18_298 VPWR VGND sg13g2_decap_8
XFILLER_34_769 VPWR VGND sg13g2_decap_8
XFILLER_33_268 VPWR VGND sg13g2_decap_8
XFILLER_17_28 VPWR VGND sg13g2_decap_8
XFILLER_37_574 VPWR VGND sg13g2_decap_8
XFILLER_24_257 VPWR VGND sg13g2_decap_8
XFILLER_25_769 VPWR VGND sg13g2_decap_8
XFILLER_40_739 VPWR VGND sg13g2_decap_8
XFILLER_20_452 VPWR VGND sg13g2_decap_8
XFILLER_0_868 VPWR VGND sg13g2_decap_8
XFILLER_16_725 VPWR VGND sg13g2_decap_8
XFILLER_28_552 VPWR VGND sg13g2_decap_8
XFILLER_15_235 VPWR VGND sg13g2_decap_8
XFILLER_43_522 VPWR VGND sg13g2_decap_8
XFILLER_31_717 VPWR VGND sg13g2_decap_8
XFILLER_30_205 VPWR VGND sg13g2_decap_8
XFILLER_43_599 VPWR VGND sg13g2_decap_8
XFILLER_11_452 VPWR VGND sg13g2_decap_8
XFILLER_23_60 VPWR VGND sg13g2_decap_8
XFILLER_7_434 VPWR VGND sg13g2_decap_8
XFILLER_3_662 VPWR VGND sg13g2_decap_8
XFILLER_2_172 VPWR VGND sg13g2_decap_8
XFILLER_38_327 VPWR VGND sg13g2_decap_8
XFILLER_47_861 VPWR VGND sg13g2_decap_8
XFILLER_0_42 VPWR VGND sg13g2_decap_8
XFILLER_46_371 VPWR VGND sg13g2_decap_8
XFILLER_19_585 VPWR VGND sg13g2_decap_8
XFILLER_34_566 VPWR VGND sg13g2_decap_8
XFILLER_22_739 VPWR VGND sg13g2_decap_8
XFILLER_21_249 VPWR VGND sg13g2_decap_8
XFILLER_9_95 VPWR VGND sg13g2_decap_8
XFILLER_30_772 VPWR VGND sg13g2_decap_8
XFILLER_29_327 VPWR VGND sg13g2_decap_8
XFILLER_45_809 VPWR VGND sg13g2_decap_8
XFILLER_44_319 VPWR VGND sg13g2_decap_8
XFILLER_37_371 VPWR VGND sg13g2_decap_8
XFILLER_38_894 VPWR VGND sg13g2_decap_8
XFILLER_25_566 VPWR VGND sg13g2_decap_8
XFILLER_13_739 VPWR VGND sg13g2_decap_8
XFILLER_40_536 VPWR VGND sg13g2_decap_8
XFILLER_12_249 VPWR VGND sg13g2_decap_8
XFILLER_4_459 VPWR VGND sg13g2_decap_8
XFILLER_0_665 VPWR VGND sg13g2_decap_8
XFILLER_48_658 VPWR VGND sg13g2_decap_8
XFILLER_36_809 VPWR VGND sg13g2_decap_8
XFILLER_47_168 VPWR VGND sg13g2_decap_8
XFILLER_18_60 VPWR VGND sg13g2_decap_8
XFILLER_16_522 VPWR VGND sg13g2_decap_8
XFILLER_29_894 VPWR VGND sg13g2_decap_8
XFILLER_16_599 VPWR VGND sg13g2_decap_8
XFILLER_31_514 VPWR VGND sg13g2_decap_8
XFILLER_44_886 VPWR VGND sg13g2_decap_8
XFILLER_34_70 VPWR VGND sg13g2_decap_8
XFILLER_43_396 VPWR VGND sg13g2_decap_8
XFILLER_8_732 VPWR VGND sg13g2_decap_8
XFILLER_7_231 VPWR VGND sg13g2_decap_8
XFILLER_38_124 VPWR VGND sg13g2_decap_8
XFILLER_39_658 VPWR VGND sg13g2_decap_8
XFILLER_26_319 VPWR VGND sg13g2_decap_8
XFILLER_19_382 VPWR VGND sg13g2_decap_8
XFILLER_35_842 VPWR VGND sg13g2_decap_8
XFILLER_14_18 VPWR VGND sg13g2_decap_8
XFILLER_34_363 VPWR VGND sg13g2_decap_8
XFILLER_22_536 VPWR VGND sg13g2_decap_8
XFILLER_29_102 VPWR VGND sg13g2_decap_8
XFILLER_18_809 VPWR VGND sg13g2_decap_8
XFILLER_29_124 VPWR VGND sg13g2_decap_8
XFILLER_17_308 VPWR VGND sg13g2_decap_8
XFILLER_45_606 VPWR VGND sg13g2_decap_8
XFILLER_38_691 VPWR VGND sg13g2_decap_8
XFILLER_44_116 VPWR VGND sg13g2_decap_8
XFILLER_25_363 VPWR VGND sg13g2_decap_8
XFILLER_26_886 VPWR VGND sg13g2_decap_8
XFILLER_13_536 VPWR VGND sg13g2_decap_8
XFILLER_40_333 VPWR VGND sg13g2_decap_8
XFILLER_41_856 VPWR VGND sg13g2_decap_8
XFILLER_9_529 VPWR VGND sg13g2_decap_8
XFILLER_5_746 VPWR VGND sg13g2_decap_8
XFILLER_4_256 VPWR VGND sg13g2_decap_8
XFILLER_0_462 VPWR VGND sg13g2_decap_8
XFILLER_48_455 VPWR VGND sg13g2_decap_8
XFILLER_29_81 VPWR VGND sg13g2_decap_8
XFILLER_36_606 VPWR VGND sg13g2_decap_8
XFILLER_29_691 VPWR VGND sg13g2_decap_8
XFILLER_17_875 VPWR VGND sg13g2_decap_8
XFILLER_35_149 VPWR VGND sg13g2_decap_8
XFILLER_32_823 VPWR VGND sg13g2_decap_8
XFILLER_44_683 VPWR VGND sg13g2_decap_8
XFILLER_16_396 VPWR VGND sg13g2_decap_8
XFILLER_31_311 VPWR VGND sg13g2_decap_8
XFILLER_43_193 VPWR VGND sg13g2_decap_8
XFILLER_31_388 VPWR VGND sg13g2_decap_8
XFILLER_6_74 VPWR VGND sg13g2_decap_8
XFILLER_39_455 VPWR VGND sg13g2_decap_8
XFILLER_26_116 VPWR VGND sg13g2_decap_8
XFILLER_23_823 VPWR VGND sg13g2_decap_8
XFILLER_25_39 VPWR VGND sg13g2_decap_8
XFILLER_34_160 VPWR VGND sg13g2_decap_8
XFILLER_22_333 VPWR VGND sg13g2_decap_8
XFILLER_1_259 VPWR VGND sg13g2_decap_8
XFILLER_18_606 VPWR VGND sg13g2_decap_8
XFILLER_45_403 VPWR VGND sg13g2_decap_8
XFILLER_17_105 VPWR VGND sg13g2_decap_8
XFILLER_14_823 VPWR VGND sg13g2_decap_8
XFILLER_25_160 VPWR VGND sg13g2_decap_8
XFILLER_26_683 VPWR VGND sg13g2_decap_8
XFILLER_13_333 VPWR VGND sg13g2_decap_8
XFILLER_40_130 VPWR VGND sg13g2_decap_8
XFILLER_41_653 VPWR VGND sg13g2_decap_8
XFILLER_9_326 VPWR VGND sg13g2_decap_8
XFILLER_5_543 VPWR VGND sg13g2_decap_8
XFILLER_49_742 VPWR VGND sg13g2_decap_8
XFILLER_48_252 VPWR VGND sg13g2_decap_8
XFILLER_36_403 VPWR VGND sg13g2_decap_8
XFILLER_17_672 VPWR VGND sg13g2_decap_8
XFILLER_16_193 VPWR VGND sg13g2_decap_8
XFILLER_32_620 VPWR VGND sg13g2_decap_8
XFILLER_44_480 VPWR VGND sg13g2_decap_8
XFILLER_20_837 VPWR VGND sg13g2_decap_8
XFILLER_31_185 VPWR VGND sg13g2_decap_8
XFILLER_32_697 VPWR VGND sg13g2_decap_8
XFILLER_9_893 VPWR VGND sg13g2_decap_8
XFILLER_39_252 VPWR VGND sg13g2_decap_8
XFILLER_27_469 VPWR VGND sg13g2_decap_8
XFILLER_43_907 VPWR VGND sg13g2_decap_8
XFILLER_42_428 VPWR VGND sg13g2_decap_8
XFILLER_23_620 VPWR VGND sg13g2_decap_8
XFILLER_22_130 VPWR VGND sg13g2_decap_8
XFILLER_11_837 VPWR VGND sg13g2_decap_8
XFILLER_23_697 VPWR VGND sg13g2_decap_8
XFILLER_10_347 VPWR VGND sg13g2_decap_8
XFILLER_7_819 VPWR VGND sg13g2_decap_8
XFILLER_2_557 VPWR VGND sg13g2_decap_8
XFILLER_18_403 VPWR VGND sg13g2_decap_8
XFILLER_45_200 VPWR VGND sg13g2_decap_8
XFILLER_46_756 VPWR VGND sg13g2_decap_8
XFILLER_45_277 VPWR VGND sg13g2_decap_8
XFILLER_14_620 VPWR VGND sg13g2_decap_8
XFILLER_26_480 VPWR VGND sg13g2_decap_8
XFILLER_13_130 VPWR VGND sg13g2_decap_8
XFILLER_41_450 VPWR VGND sg13g2_decap_8
XFILLER_9_123 VPWR VGND sg13g2_decap_8
XFILLER_14_697 VPWR VGND sg13g2_decap_8
XFILLER_6_830 VPWR VGND sg13g2_decap_8
XFILLER_42_92 VPWR VGND sg13g2_decap_8
XFILLER_5_340 VPWR VGND sg13g2_decap_8
XFILLER_3_53 VPWR VGND sg13g2_decap_8
XFILLER_36_200 VPWR VGND sg13g2_decap_8
XFILLER_37_756 VPWR VGND sg13g2_decap_8
XFILLER_36_277 VPWR VGND sg13g2_decap_8
XFILLER_24_439 VPWR VGND sg13g2_decap_8
XFILLER_20_634 VPWR VGND sg13g2_decap_8
XFILLER_22_18 VPWR VGND sg13g2_decap_8
XFILLER_32_494 VPWR VGND sg13g2_decap_8
XFILLER_9_690 VPWR VGND sg13g2_decap_8
XFILLER_28_734 VPWR VGND sg13g2_decap_8
XFILLER_16_907 VPWR VGND sg13g2_decap_8
XFILLER_15_417 VPWR VGND sg13g2_decap_8
XFILLER_27_266 VPWR VGND sg13g2_decap_8
XFILLER_43_704 VPWR VGND sg13g2_decap_8
XFILLER_42_225 VPWR VGND sg13g2_decap_8
XFILLER_7_616 VPWR VGND sg13g2_decap_8
XFILLER_11_634 VPWR VGND sg13g2_decap_8
XFILLER_23_494 VPWR VGND sg13g2_decap_8
XFILLER_10_144 VPWR VGND sg13g2_decap_8
XFILLER_6_137 VPWR VGND sg13g2_decap_8
XFILLER_12_95 VPWR VGND sg13g2_decap_8
XFILLER_3_844 VPWR VGND sg13g2_decap_8
XFILLER_2_354 VPWR VGND sg13g2_decap_8
XFILLER_38_509 VPWR VGND sg13g2_decap_8
XFILLER_18_200 VPWR VGND sg13g2_decap_8
XFILLER_19_767 VPWR VGND sg13g2_decap_8
XFILLER_46_553 VPWR VGND sg13g2_decap_8
XFILLER_18_277 VPWR VGND sg13g2_decap_8
XFILLER_37_70 VPWR VGND sg13g2_decap_8
XFILLER_34_748 VPWR VGND sg13g2_decap_8
XFILLER_33_247 VPWR VGND sg13g2_decap_8
XFILLER_42_792 VPWR VGND sg13g2_decap_8
XFILLER_14_494 VPWR VGND sg13g2_decap_8
XFILLER_29_509 VPWR VGND sg13g2_decap_8
XFILLER_37_553 VPWR VGND sg13g2_decap_8
XFILLER_24_236 VPWR VGND sg13g2_decap_8
XFILLER_25_748 VPWR VGND sg13g2_decap_8
XFILLER_40_718 VPWR VGND sg13g2_decap_8
XFILLER_21_921 VPWR VGND sg13g2_decap_4
XFILLER_20_431 VPWR VGND sg13g2_decap_8
XFILLER_32_291 VPWR VGND sg13g2_decap_8
XFILLER_0_847 VPWR VGND sg13g2_decap_8
XFILLER_28_531 VPWR VGND sg13g2_decap_8
XFILLER_16_704 VPWR VGND sg13g2_decap_8
XFILLER_43_501 VPWR VGND sg13g2_decap_8
XFILLER_15_214 VPWR VGND sg13g2_decap_8
XFILLER_43_578 VPWR VGND sg13g2_decap_8
XFILLER_12_921 VPWR VGND sg13g2_decap_4
XFILLER_11_431 VPWR VGND sg13g2_decap_8
XFILLER_8_914 VPWR VGND sg13g2_decap_8
XFILLER_23_291 VPWR VGND sg13g2_decap_8
XFILLER_7_413 VPWR VGND sg13g2_decap_8
XFILLER_3_641 VPWR VGND sg13g2_decap_8
XFILLER_2_151 VPWR VGND sg13g2_decap_8
XFILLER_38_306 VPWR VGND sg13g2_decap_8
XFILLER_47_840 VPWR VGND sg13g2_decap_8
XFILLER_48_91 VPWR VGND sg13g2_decap_8
XFILLER_46_350 VPWR VGND sg13g2_decap_8
XFILLER_0_21 VPWR VGND sg13g2_decap_8
XFILLER_19_564 VPWR VGND sg13g2_decap_8
XFILLER_0_98 VPWR VGND sg13g2_decap_8
XFILLER_22_718 VPWR VGND sg13g2_decap_8
XFILLER_34_545 VPWR VGND sg13g2_decap_8
XFILLER_15_781 VPWR VGND sg13g2_decap_8
XFILLER_21_228 VPWR VGND sg13g2_decap_8
XFILLER_14_291 VPWR VGND sg13g2_decap_8
XFILLER_9_74 VPWR VGND sg13g2_decap_8
XFILLER_30_751 VPWR VGND sg13g2_decap_8
XFILLER_28_39 VPWR VGND sg13g2_decap_8
XFILLER_29_306 VPWR VGND sg13g2_decap_8
XFILLER_37_350 VPWR VGND sg13g2_decap_8
XFILLER_38_873 VPWR VGND sg13g2_decap_8
XFILLER_25_545 VPWR VGND sg13g2_decap_8
XFILLER_13_718 VPWR VGND sg13g2_decap_8
XFILLER_40_515 VPWR VGND sg13g2_decap_8
XFILLER_12_228 VPWR VGND sg13g2_decap_8
XFILLER_21_795 VPWR VGND sg13g2_decap_8
XFILLER_4_438 VPWR VGND sg13g2_decap_8
XFILLER_0_644 VPWR VGND sg13g2_decap_8
XFILLER_48_637 VPWR VGND sg13g2_decap_8
XFILLER_47_147 VPWR VGND sg13g2_decap_8
XFILLER_29_873 VPWR VGND sg13g2_decap_8
XFILLER_16_501 VPWR VGND sg13g2_decap_8
XFILLER_44_865 VPWR VGND sg13g2_decap_8
XFILLER_16_578 VPWR VGND sg13g2_decap_8
XFILLER_43_375 VPWR VGND sg13g2_decap_8
XFILLER_8_711 VPWR VGND sg13g2_decap_8
XFILLER_7_210 VPWR VGND sg13g2_decap_8
XFILLER_12_795 VPWR VGND sg13g2_decap_8
XFILLER_8_788 VPWR VGND sg13g2_decap_8
XFILLER_7_287 VPWR VGND sg13g2_decap_8
XFILLER_22_4 VPWR VGND sg13g2_decap_8
XFILLER_38_103 VPWR VGND sg13g2_decap_8
XFILLER_39_637 VPWR VGND sg13g2_decap_8
XFILLER_19_361 VPWR VGND sg13g2_decap_8
XFILLER_35_821 VPWR VGND sg13g2_decap_8
XFILLER_34_342 VPWR VGND sg13g2_decap_8
XFILLER_22_515 VPWR VGND sg13g2_decap_8
XFILLER_35_898 VPWR VGND sg13g2_decap_8
XFILLER_39_49 VPWR VGND sg13g2_decap_8
XFILLER_38_670 VPWR VGND sg13g2_decap_8
XFILLER_25_342 VPWR VGND sg13g2_decap_8
XFILLER_26_865 VPWR VGND sg13g2_decap_8
XFILLER_13_515 VPWR VGND sg13g2_decap_8
XFILLER_41_835 VPWR VGND sg13g2_decap_8
XFILLER_9_508 VPWR VGND sg13g2_decap_8
XFILLER_40_312 VPWR VGND sg13g2_decap_8
XFILLER_21_592 VPWR VGND sg13g2_decap_8
XFILLER_40_389 VPWR VGND sg13g2_decap_8
XFILLER_5_725 VPWR VGND sg13g2_decap_8
XFILLER_4_235 VPWR VGND sg13g2_decap_8
XFILLER_20_95 VPWR VGND sg13g2_decap_8
XFILLER_49_924 VPWR VGND sg13g2_fill_1
XFILLER_0_441 VPWR VGND sg13g2_decap_8
XFILLER_48_434 VPWR VGND sg13g2_decap_8
XFILLER_29_60 VPWR VGND sg13g2_decap_8
XFILLER_29_670 VPWR VGND sg13g2_decap_8
XFILLER_35_128 VPWR VGND sg13g2_decap_8
XFILLER_17_854 VPWR VGND sg13g2_decap_8
XFILLER_16_375 VPWR VGND sg13g2_decap_8
XFILLER_32_802 VPWR VGND sg13g2_decap_8
XFILLER_44_662 VPWR VGND sg13g2_decap_8
XFILLER_45_81 VPWR VGND sg13g2_decap_8
XFILLER_43_172 VPWR VGND sg13g2_decap_8
XFILLER_31_367 VPWR VGND sg13g2_decap_8
XFILLER_32_879 VPWR VGND sg13g2_decap_8
XFILLER_12_592 VPWR VGND sg13g2_decap_8
XFILLER_8_585 VPWR VGND sg13g2_decap_8
XFILLER_6_53 VPWR VGND sg13g2_decap_8
XFILLER_39_434 VPWR VGND sg13g2_decap_8
XFILLER_25_18 VPWR VGND sg13g2_decap_8
XFILLER_23_802 VPWR VGND sg13g2_decap_8
XFILLER_22_312 VPWR VGND sg13g2_decap_8
XFILLER_35_695 VPWR VGND sg13g2_decap_8
XFILLER_23_879 VPWR VGND sg13g2_decap_8
XFILLER_10_529 VPWR VGND sg13g2_decap_8
XFILLER_22_389 VPWR VGND sg13g2_decap_8
XFILLER_2_739 VPWR VGND sg13g2_decap_8
XFILLER_1_238 VPWR VGND sg13g2_decap_8
XFILLER_45_459 VPWR VGND sg13g2_decap_8
XFILLER_14_802 VPWR VGND sg13g2_decap_8
XFILLER_26_662 VPWR VGND sg13g2_decap_8
XFILLER_32_109 VPWR VGND sg13g2_decap_8
XFILLER_13_312 VPWR VGND sg13g2_decap_8
XFILLER_41_632 VPWR VGND sg13g2_decap_8
XFILLER_9_305 VPWR VGND sg13g2_decap_8
XFILLER_14_879 VPWR VGND sg13g2_decap_8
XFILLER_13_389 VPWR VGND sg13g2_decap_8
XFILLER_15_95 VPWR VGND sg13g2_decap_8
XFILLER_40_186 VPWR VGND sg13g2_decap_8
XFILLER_5_522 VPWR VGND sg13g2_decap_8
XFILLER_5_599 VPWR VGND sg13g2_decap_8
XFILLER_49_721 VPWR VGND sg13g2_decap_8
XFILLER_48_231 VPWR VGND sg13g2_decap_8
XFILLER_49_798 VPWR VGND sg13g2_decap_8
XFILLER_36_459 VPWR VGND sg13g2_decap_8
XFILLER_17_651 VPWR VGND sg13g2_decap_8
XFILLER_23_109 VPWR VGND sg13g2_decap_8
XFILLER_16_172 VPWR VGND sg13g2_decap_8
XFILLER_20_816 VPWR VGND sg13g2_decap_8
XFILLER_32_676 VPWR VGND sg13g2_decap_8
XFILLER_31_164 VPWR VGND sg13g2_decap_8
XFILLER_9_872 VPWR VGND sg13g2_decap_8
XFILLER_8_382 VPWR VGND sg13g2_decap_8
XFILLER_28_916 VPWR VGND sg13g2_decap_8
XFILLER_39_231 VPWR VGND sg13g2_decap_8
XFILLER_27_448 VPWR VGND sg13g2_decap_8
XFILLER_36_39 VPWR VGND sg13g2_decap_8
XFILLER_14_109 VPWR VGND sg13g2_decap_8
XFILLER_42_407 VPWR VGND sg13g2_decap_8
XFILLER_35_492 VPWR VGND sg13g2_decap_8
XFILLER_11_816 VPWR VGND sg13g2_decap_8
XFILLER_23_676 VPWR VGND sg13g2_decap_8
XFILLER_10_326 VPWR VGND sg13g2_decap_8
XFILLER_22_186 VPWR VGND sg13g2_decap_8
XFILLER_6_319 VPWR VGND sg13g2_decap_8
XFILLER_2_536 VPWR VGND sg13g2_decap_8
XFILLER_46_735 VPWR VGND sg13g2_decap_8
XFILLER_18_459 VPWR VGND sg13g2_decap_8
XFILLER_45_256 VPWR VGND sg13g2_decap_8
XFILLER_26_61 VPWR VGND sg13g2_decap_8
XFILLER_33_429 VPWR VGND sg13g2_decap_8
XFILLER_9_102 VPWR VGND sg13g2_decap_8
XFILLER_14_676 VPWR VGND sg13g2_decap_8
XFILLER_13_186 VPWR VGND sg13g2_decap_8
XFILLER_42_71 VPWR VGND sg13g2_decap_8
XFILLER_9_179 VPWR VGND sg13g2_decap_8
XFILLER_10_893 VPWR VGND sg13g2_decap_8
XFILLER_6_886 VPWR VGND sg13g2_decap_8
XFILLER_5_396 VPWR VGND sg13g2_decap_8
XFILLER_3_32 VPWR VGND sg13g2_decap_8
XFILLER_49_595 VPWR VGND sg13g2_decap_8
XFILLER_37_735 VPWR VGND sg13g2_decap_8
XFILLER_24_418 VPWR VGND sg13g2_decap_8
XFILLER_36_256 VPWR VGND sg13g2_decap_8
XFILLER_20_613 VPWR VGND sg13g2_decap_8
XFILLER_32_473 VPWR VGND sg13g2_decap_8
XFILLER_47_49 VPWR VGND sg13g2_decap_8
XFILLER_28_713 VPWR VGND sg13g2_decap_8
XFILLER_27_245 VPWR VGND sg13g2_decap_8
XFILLER_42_204 VPWR VGND sg13g2_decap_8
XFILLER_11_613 VPWR VGND sg13g2_decap_8
XFILLER_23_473 VPWR VGND sg13g2_decap_8
XFILLER_10_123 VPWR VGND sg13g2_decap_8
XFILLER_6_116 VPWR VGND sg13g2_decap_8
XFILLER_12_74 VPWR VGND sg13g2_decap_8
XFILLER_3_823 VPWR VGND sg13g2_decap_8
XFILLER_2_333 VPWR VGND sg13g2_decap_8
XFILLER_46_532 VPWR VGND sg13g2_decap_8
XFILLER_19_746 VPWR VGND sg13g2_decap_8
XFILLER_18_256 VPWR VGND sg13g2_decap_8
XFILLER_33_226 VPWR VGND sg13g2_decap_8
XFILLER_34_727 VPWR VGND sg13g2_decap_8
XFILLER_14_473 VPWR VGND sg13g2_decap_8
XFILLER_42_771 VPWR VGND sg13g2_decap_8
XFILLER_10_690 VPWR VGND sg13g2_decap_8
XFILLER_6_683 VPWR VGND sg13g2_decap_8
XFILLER_5_193 VPWR VGND sg13g2_decap_8
XFILLER_49_392 VPWR VGND sg13g2_decap_8
XFILLER_37_532 VPWR VGND sg13g2_decap_8
XFILLER_24_215 VPWR VGND sg13g2_decap_8
XFILLER_25_727 VPWR VGND sg13g2_decap_8
XFILLER_21_900 VPWR VGND sg13g2_decap_8
XFILLER_33_18 VPWR VGND sg13g2_decap_8
XFILLER_20_410 VPWR VGND sg13g2_decap_8
XFILLER_32_270 VPWR VGND sg13g2_decap_8
XFILLER_33_793 VPWR VGND sg13g2_decap_8
XFILLER_20_487 VPWR VGND sg13g2_decap_8
XFILLER_0_826 VPWR VGND sg13g2_decap_8
XFILLER_48_819 VPWR VGND sg13g2_decap_8
XFILLER_47_329 VPWR VGND sg13g2_decap_8
XFILLER_28_510 VPWR VGND sg13g2_decap_8
XFILLER_28_587 VPWR VGND sg13g2_decap_8
XFILLER_43_557 VPWR VGND sg13g2_decap_8
XFILLER_12_900 VPWR VGND sg13g2_decap_8
XFILLER_24_782 VPWR VGND sg13g2_decap_8
XFILLER_11_410 VPWR VGND sg13g2_decap_8
XFILLER_23_270 VPWR VGND sg13g2_decap_8
XFILLER_11_487 VPWR VGND sg13g2_decap_8
XFILLER_23_95 VPWR VGND sg13g2_decap_8
XFILLER_7_469 VPWR VGND sg13g2_decap_8
XFILLER_3_620 VPWR VGND sg13g2_decap_8
XFILLER_2_130 VPWR VGND sg13g2_decap_8
XFILLER_3_697 VPWR VGND sg13g2_decap_8
XFILLER_48_70 VPWR VGND sg13g2_decap_8
XFILLER_39_819 VPWR VGND sg13g2_decap_8
XFILLER_17_7 VPWR VGND sg13g2_decap_8
XFILLER_19_543 VPWR VGND sg13g2_decap_8
XFILLER_47_896 VPWR VGND sg13g2_decap_8
XFILLER_0_77 VPWR VGND sg13g2_decap_8
XFILLER_34_524 VPWR VGND sg13g2_decap_8
XFILLER_15_760 VPWR VGND sg13g2_decap_8
XFILLER_21_207 VPWR VGND sg13g2_decap_8
XFILLER_9_53 VPWR VGND sg13g2_decap_8
XFILLER_14_270 VPWR VGND sg13g2_decap_8
XFILLER_30_730 VPWR VGND sg13g2_decap_8
XFILLER_6_480 VPWR VGND sg13g2_decap_8
XFILLER_28_18 VPWR VGND sg13g2_decap_8
XFILLER_38_852 VPWR VGND sg13g2_decap_8
XFILLER_25_524 VPWR VGND sg13g2_decap_8
XFILLER_44_39 VPWR VGND sg13g2_decap_8
XFILLER_12_207 VPWR VGND sg13g2_decap_8
XFILLER_33_590 VPWR VGND sg13g2_decap_8
XFILLER_21_774 VPWR VGND sg13g2_decap_8
XFILLER_20_284 VPWR VGND sg13g2_decap_8
XFILLER_5_907 VPWR VGND sg13g2_decap_8
XFILLER_4_417 VPWR VGND sg13g2_decap_8
XFILLER_0_623 VPWR VGND sg13g2_decap_8
XFILLER_48_616 VPWR VGND sg13g2_decap_8
XFILLER_47_126 VPWR VGND sg13g2_decap_8
XFILLER_29_852 VPWR VGND sg13g2_decap_8
XFILLER_18_95 VPWR VGND sg13g2_decap_8
XFILLER_28_384 VPWR VGND sg13g2_decap_8
XFILLER_16_557 VPWR VGND sg13g2_decap_8
XFILLER_44_844 VPWR VGND sg13g2_decap_8
XFILLER_43_354 VPWR VGND sg13g2_decap_8
XFILLER_31_549 VPWR VGND sg13g2_decap_8
XFILLER_12_774 VPWR VGND sg13g2_decap_8
XFILLER_11_284 VPWR VGND sg13g2_decap_8
XFILLER_8_767 VPWR VGND sg13g2_decap_8
XFILLER_7_266 VPWR VGND sg13g2_decap_8
XFILLER_3_494 VPWR VGND sg13g2_decap_8
XFILLER_39_616 VPWR VGND sg13g2_decap_8
XFILLER_15_4 VPWR VGND sg13g2_decap_8
XFILLER_19_340 VPWR VGND sg13g2_decap_8
XFILLER_35_800 VPWR VGND sg13g2_decap_8
XFILLER_38_159 VPWR VGND sg13g2_decap_8
XFILLER_47_693 VPWR VGND sg13g2_decap_8
XFILLER_34_321 VPWR VGND sg13g2_decap_8
XFILLER_35_877 VPWR VGND sg13g2_decap_8
XFILLER_34_398 VPWR VGND sg13g2_decap_8
XFILLER_29_159 VPWR VGND sg13g2_decap_8
XFILLER_25_321 VPWR VGND sg13g2_decap_8
XFILLER_26_844 VPWR VGND sg13g2_decap_8
XFILLER_41_814 VPWR VGND sg13g2_decap_8
XFILLER_25_398 VPWR VGND sg13g2_decap_8
XFILLER_40_368 VPWR VGND sg13g2_decap_8
XFILLER_21_571 VPWR VGND sg13g2_decap_8
XFILLER_5_704 VPWR VGND sg13g2_decap_8
XFILLER_4_214 VPWR VGND sg13g2_decap_8
XFILLER_1_910 VPWR VGND sg13g2_decap_8
XFILLER_20_74 VPWR VGND sg13g2_decap_8
XFILLER_0_420 VPWR VGND sg13g2_decap_8
XFILLER_49_903 VPWR VGND sg13g2_decap_8
XFILLER_48_413 VPWR VGND sg13g2_decap_8
XFILLER_0_497 VPWR VGND sg13g2_decap_8
XFILLER_17_833 VPWR VGND sg13g2_decap_8
XFILLER_28_181 VPWR VGND sg13g2_decap_8
XFILLER_44_641 VPWR VGND sg13g2_decap_8
XFILLER_16_354 VPWR VGND sg13g2_decap_8
XFILLER_43_151 VPWR VGND sg13g2_decap_8
XFILLER_45_60 VPWR VGND sg13g2_decap_8
XFILLER_32_858 VPWR VGND sg13g2_decap_8
XFILLER_31_346 VPWR VGND sg13g2_decap_8
XFILLER_12_571 VPWR VGND sg13g2_decap_8
XFILLER_8_564 VPWR VGND sg13g2_decap_8
XFILLER_6_32 VPWR VGND sg13g2_decap_8
XFILLER_4_781 VPWR VGND sg13g2_decap_8
XFILLER_3_291 VPWR VGND sg13g2_decap_8
XFILLER_39_413 VPWR VGND sg13g2_decap_8
XFILLER_47_490 VPWR VGND sg13g2_decap_8
XFILLER_35_674 VPWR VGND sg13g2_decap_8
XFILLER_23_858 VPWR VGND sg13g2_decap_8
XFILLER_10_508 VPWR VGND sg13g2_decap_8
XFILLER_22_368 VPWR VGND sg13g2_decap_8
XFILLER_34_195 VPWR VGND sg13g2_decap_8
XFILLER_41_18 VPWR VGND sg13g2_decap_8
XFILLER_2_718 VPWR VGND sg13g2_decap_8
XFILLER_1_217 VPWR VGND sg13g2_decap_8
XFILLER_46_917 VPWR VGND sg13g2_decap_8
XFILLER_26_641 VPWR VGND sg13g2_decap_8
XFILLER_45_438 VPWR VGND sg13g2_decap_8
XFILLER_14_858 VPWR VGND sg13g2_decap_8
XFILLER_41_611 VPWR VGND sg13g2_decap_8
XFILLER_13_368 VPWR VGND sg13g2_decap_8
XFILLER_15_74 VPWR VGND sg13g2_decap_8
XFILLER_25_195 VPWR VGND sg13g2_decap_8
XFILLER_40_165 VPWR VGND sg13g2_decap_8
XFILLER_41_688 VPWR VGND sg13g2_decap_8
XFILLER_5_501 VPWR VGND sg13g2_decap_8
XFILLER_31_40 VPWR VGND sg13g2_fill_2
XFILLER_5_578 VPWR VGND sg13g2_decap_8
XFILLER_49_700 VPWR VGND sg13g2_decap_8
XFILLER_48_210 VPWR VGND sg13g2_decap_8
XFILLER_1_784 VPWR VGND sg13g2_decap_8
XFILLER_49_777 VPWR VGND sg13g2_decap_8
XFILLER_0_294 VPWR VGND sg13g2_decap_8
XFILLER_37_917 VPWR VGND sg13g2_decap_8
XFILLER_48_287 VPWR VGND sg13g2_decap_8
XFILLER_17_630 VPWR VGND sg13g2_decap_8
XFILLER_36_438 VPWR VGND sg13g2_decap_8
XFILLER_16_151 VPWR VGND sg13g2_decap_8
XFILLER_31_143 VPWR VGND sg13g2_decap_8
XFILLER_32_655 VPWR VGND sg13g2_decap_8
XFILLER_9_851 VPWR VGND sg13g2_decap_8
XFILLER_8_361 VPWR VGND sg13g2_decap_8
XFILLER_39_210 VPWR VGND sg13g2_decap_8
XFILLER_36_18 VPWR VGND sg13g2_decap_8
XFILLER_27_427 VPWR VGND sg13g2_decap_8
XFILLER_39_287 VPWR VGND sg13g2_decap_8
XFILLER_35_471 VPWR VGND sg13g2_decap_8
XFILLER_23_655 VPWR VGND sg13g2_decap_8
XFILLER_10_305 VPWR VGND sg13g2_decap_8
XFILLER_22_165 VPWR VGND sg13g2_decap_8
XFILLER_2_515 VPWR VGND sg13g2_decap_8
XFILLER_46_714 VPWR VGND sg13g2_decap_8
XFILLER_18_438 VPWR VGND sg13g2_decap_8
XFILLER_34_909 VPWR VGND sg13g2_decap_8
XFILLER_45_235 VPWR VGND sg13g2_decap_8
XFILLER_26_40 VPWR VGND sg13g2_decap_8
XFILLER_33_408 VPWR VGND sg13g2_decap_8
XFILLER_14_655 VPWR VGND sg13g2_decap_8
XFILLER_26_95 VPWR VGND sg13g2_decap_8
XFILLER_13_165 VPWR VGND sg13g2_decap_8
XFILLER_41_485 VPWR VGND sg13g2_decap_8
XFILLER_9_158 VPWR VGND sg13g2_decap_8
XFILLER_42_50 VPWR VGND sg13g2_decap_8
XFILLER_10_872 VPWR VGND sg13g2_decap_8
XFILLER_6_865 VPWR VGND sg13g2_decap_8
XFILLER_47_7 VPWR VGND sg13g2_decap_8
XFILLER_5_375 VPWR VGND sg13g2_decap_8
XFILLER_3_11 VPWR VGND sg13g2_decap_8
XFILLER_3_88 VPWR VGND sg13g2_decap_8
XFILLER_1_581 VPWR VGND sg13g2_decap_8
XFILLER_49_574 VPWR VGND sg13g2_decap_8
XFILLER_37_714 VPWR VGND sg13g2_decap_8
XFILLER_36_235 VPWR VGND sg13g2_decap_8
XFILLER_25_909 VPWR VGND sg13g2_decap_8
XFILLER_32_452 VPWR VGND sg13g2_decap_8
XFILLER_20_669 VPWR VGND sg13g2_decap_8
XFILLER_47_28 VPWR VGND sg13g2_decap_8
XFILLER_27_224 VPWR VGND sg13g2_decap_8
XFILLER_28_769 VPWR VGND sg13g2_decap_8
XFILLER_43_739 VPWR VGND sg13g2_decap_8
XFILLER_23_452 VPWR VGND sg13g2_decap_8
XFILLER_10_102 VPWR VGND sg13g2_decap_8
XFILLER_11_669 VPWR VGND sg13g2_decap_8
XFILLER_10_179 VPWR VGND sg13g2_decap_8
XFILLER_12_53 VPWR VGND sg13g2_decap_8
XFILLER_3_802 VPWR VGND sg13g2_decap_8
XFILLER_2_312 VPWR VGND sg13g2_decap_8
XFILLER_3_879 VPWR VGND sg13g2_decap_8
XFILLER_2_389 VPWR VGND sg13g2_decap_8
XFILLER_46_511 VPWR VGND sg13g2_decap_8
XFILLER_19_725 VPWR VGND sg13g2_decap_8
XFILLER_18_235 VPWR VGND sg13g2_decap_8
XFILLER_34_706 VPWR VGND sg13g2_decap_8
XFILLER_46_588 VPWR VGND sg13g2_decap_8
XFILLER_27_791 VPWR VGND sg13g2_decap_8
XFILLER_33_205 VPWR VGND sg13g2_decap_8
XFILLER_42_750 VPWR VGND sg13g2_decap_8
XFILLER_14_452 VPWR VGND sg13g2_decap_8
XFILLER_30_912 VPWR VGND sg13g2_decap_8
XFILLER_30_923 VPWR VGND sg13g2_fill_2
XFILLER_41_282 VPWR VGND sg13g2_decap_8
XFILLER_6_662 VPWR VGND sg13g2_decap_8
XFILLER_5_172 VPWR VGND sg13g2_decap_8
XFILLER_45_4 VPWR VGND sg13g2_decap_8
XFILLER_49_371 VPWR VGND sg13g2_decap_8
XFILLER_37_511 VPWR VGND sg13g2_decap_8
XFILLER_25_706 VPWR VGND sg13g2_decap_8
XFILLER_37_588 VPWR VGND sg13g2_decap_8
XFILLER_33_772 VPWR VGND sg13g2_decap_8
XFILLER_20_466 VPWR VGND sg13g2_decap_8
XFILLER_3_109 VPWR VGND sg13g2_decap_8
XFILLER_0_805 VPWR VGND sg13g2_decap_8
XFILLER_47_308 VPWR VGND sg13g2_decap_8
XFILLER_28_566 VPWR VGND sg13g2_decap_8
XFILLER_16_739 VPWR VGND sg13g2_decap_8
XFILLER_15_249 VPWR VGND sg13g2_decap_8
XFILLER_43_536 VPWR VGND sg13g2_decap_8
XFILLER_24_761 VPWR VGND sg13g2_decap_8
XFILLER_30_219 VPWR VGND sg13g2_decap_8
XFILLER_11_466 VPWR VGND sg13g2_decap_8
XFILLER_7_448 VPWR VGND sg13g2_decap_8
XFILLER_23_74 VPWR VGND sg13g2_decap_8
XFILLER_3_676 VPWR VGND sg13g2_decap_8
XFILLER_2_186 VPWR VGND sg13g2_decap_8
XFILLER_19_522 VPWR VGND sg13g2_decap_8
XFILLER_47_875 VPWR VGND sg13g2_decap_8
XFILLER_46_385 VPWR VGND sg13g2_decap_8
XFILLER_0_56 VPWR VGND sg13g2_decap_8
XFILLER_19_599 VPWR VGND sg13g2_decap_8
XFILLER_34_503 VPWR VGND sg13g2_decap_8
XFILLER_9_32 VPWR VGND sg13g2_decap_8
XFILLER_30_786 VPWR VGND sg13g2_decap_8
XFILLER_38_831 VPWR VGND sg13g2_decap_8
XFILLER_25_503 VPWR VGND sg13g2_decap_8
XFILLER_37_385 VPWR VGND sg13g2_decap_8
XFILLER_44_18 VPWR VGND sg13g2_decap_8
XFILLER_21_753 VPWR VGND sg13g2_decap_8
XFILLER_20_263 VPWR VGND sg13g2_decap_8
XFILLER_0_602 VPWR VGND sg13g2_decap_8
XFILLER_0_679 VPWR VGND sg13g2_decap_8
XFILLER_47_105 VPWR VGND sg13g2_decap_8
XFILLER_29_831 VPWR VGND sg13g2_decap_8
XFILLER_18_74 VPWR VGND sg13g2_decap_8
XFILLER_28_363 VPWR VGND sg13g2_decap_8
XFILLER_44_823 VPWR VGND sg13g2_decap_8
XFILLER_16_536 VPWR VGND sg13g2_decap_8
XFILLER_43_333 VPWR VGND sg13g2_decap_8
XFILLER_31_528 VPWR VGND sg13g2_decap_8
XFILLER_12_753 VPWR VGND sg13g2_decap_8
XFILLER_34_84 VPWR VGND sg13g2_decap_8
XFILLER_11_263 VPWR VGND sg13g2_decap_8
XFILLER_8_746 VPWR VGND sg13g2_decap_8
XFILLER_7_245 VPWR VGND sg13g2_decap_8
XFILLER_3_473 VPWR VGND sg13g2_decap_8
XFILLER_38_138 VPWR VGND sg13g2_decap_8
XFILLER_47_672 VPWR VGND sg13g2_decap_8
XFILLER_34_300 VPWR VGND sg13g2_decap_8
XFILLER_46_182 VPWR VGND sg13g2_decap_8
XFILLER_19_396 VPWR VGND sg13g2_decap_8
XFILLER_35_856 VPWR VGND sg13g2_decap_8
XFILLER_34_377 VPWR VGND sg13g2_decap_8
XFILLER_30_583 VPWR VGND sg13g2_decap_8
XFILLER_39_18 VPWR VGND sg13g2_fill_2
XFILLER_39_29 VPWR VGND sg13g2_fill_1
XFILLER_29_116 VPWR VGND sg13g2_fill_2
XFILLER_29_138 VPWR VGND sg13g2_decap_8
XFILLER_25_300 VPWR VGND sg13g2_decap_8
XFILLER_26_823 VPWR VGND sg13g2_decap_8
XFILLER_37_182 VPWR VGND sg13g2_decap_8
XFILLER_25_377 VPWR VGND sg13g2_decap_8
XFILLER_40_347 VPWR VGND sg13g2_decap_8
XFILLER_21_550 VPWR VGND sg13g2_decap_8
XFILLER_20_53 VPWR VGND sg13g2_decap_8
XFILLER_0_476 VPWR VGND sg13g2_decap_8
XFILLER_48_469 VPWR VGND sg13g2_decap_8
XFILLER_29_95 VPWR VGND sg13g2_decap_8
XFILLER_17_812 VPWR VGND sg13g2_decap_8
XFILLER_16_333 VPWR VGND sg13g2_decap_8
XFILLER_28_160 VPWR VGND sg13g2_decap_8
XFILLER_44_620 VPWR VGND sg13g2_decap_8
XFILLER_17_889 VPWR VGND sg13g2_decap_8
XFILLER_43_130 VPWR VGND sg13g2_decap_8
XFILLER_31_325 VPWR VGND sg13g2_decap_8
XFILLER_32_837 VPWR VGND sg13g2_decap_8
XFILLER_44_697 VPWR VGND sg13g2_decap_8
XFILLER_12_550 VPWR VGND sg13g2_decap_8
XFILLER_8_543 VPWR VGND sg13g2_decap_8
XFILLER_6_11 VPWR VGND sg13g2_decap_8
XFILLER_6_88 VPWR VGND sg13g2_decap_8
XFILLER_4_760 VPWR VGND sg13g2_decap_8
XFILLER_3_270 VPWR VGND sg13g2_decap_8
XFILLER_27_609 VPWR VGND sg13g2_decap_8
XFILLER_39_469 VPWR VGND sg13g2_decap_8
XFILLER_19_193 VPWR VGND sg13g2_decap_8
XFILLER_35_653 VPWR VGND sg13g2_decap_8
XFILLER_23_837 VPWR VGND sg13g2_decap_8
XFILLER_34_174 VPWR VGND sg13g2_decap_8
XFILLER_22_347 VPWR VGND sg13g2_decap_8
XFILLER_30_380 VPWR VGND sg13g2_decap_8
XFILLER_31_892 VPWR VGND sg13g2_decap_8
XFILLER_45_417 VPWR VGND sg13g2_decap_8
XFILLER_17_119 VPWR VGND sg13g2_decap_8
XFILLER_26_620 VPWR VGND sg13g2_decap_8
XFILLER_14_837 VPWR VGND sg13g2_decap_8
XFILLER_25_174 VPWR VGND sg13g2_decap_8
XFILLER_26_697 VPWR VGND sg13g2_decap_8
XFILLER_13_347 VPWR VGND sg13g2_decap_8
XFILLER_15_53 VPWR VGND sg13g2_decap_8
XFILLER_40_144 VPWR VGND sg13g2_decap_8
XFILLER_41_667 VPWR VGND sg13g2_decap_8
XFILLER_31_74 VPWR VGND sg13g2_decap_8
XFILLER_5_557 VPWR VGND sg13g2_decap_8
XFILLER_1_763 VPWR VGND sg13g2_decap_8
XFILLER_0_273 VPWR VGND sg13g2_decap_8
XFILLER_49_756 VPWR VGND sg13g2_decap_8
XFILLER_48_266 VPWR VGND sg13g2_decap_8
XFILLER_36_417 VPWR VGND sg13g2_decap_8
XFILLER_16_130 VPWR VGND sg13g2_decap_8
XFILLER_17_686 VPWR VGND sg13g2_decap_8
XFILLER_31_100 VPWR VGND sg13g2_decap_4
XFILLER_31_111 VPWR VGND sg13g2_decap_8
XFILLER_31_122 VPWR VGND sg13g2_decap_8
XFILLER_32_634 VPWR VGND sg13g2_decap_8
XFILLER_44_494 VPWR VGND sg13g2_decap_8
XFILLER_9_830 VPWR VGND sg13g2_decap_8
XFILLER_31_199 VPWR VGND sg13g2_decap_8
XFILLER_8_340 VPWR VGND sg13g2_decap_8
.ends

