module NE_term (UserCLK,
    UserCLKo,
    FrameData,
    FrameData_O,
    FrameStrobe,
    FrameStrobe_O,
    N1END,
    N2END,
    N2MID,
    N4END,
    S1BEG,
    S2BEG,
    S2BEGb,
    S4BEG);
 input UserCLK;
 output UserCLKo;
 input [31:0] FrameData;
 output [31:0] FrameData_O;
 input [19:0] FrameStrobe;
 output [19:0] FrameStrobe_O;
 input [3:0] N1END;
 input [7:0] N2END;
 input [7:0] N2MID;
 input [15:0] N4END;
 output [3:0] S1BEG;
 output [7:0] S2BEG;
 output [7:0] S2BEGb;
 output [15:0] S4BEG;


 sg13g2_buf_1 _00_ (.A(FrameData[0]),
    .X(FrameData_O[0]));
 sg13g2_buf_1 _01_ (.A(FrameData[1]),
    .X(FrameData_O[1]));
 sg13g2_buf_1 _02_ (.A(FrameData[2]),
    .X(FrameData_O[2]));
 sg13g2_buf_1 _03_ (.A(FrameData[3]),
    .X(FrameData_O[3]));
 sg13g2_buf_1 _04_ (.A(FrameData[4]),
    .X(FrameData_O[4]));
 sg13g2_buf_1 _05_ (.A(FrameData[5]),
    .X(FrameData_O[5]));
 sg13g2_buf_1 _06_ (.A(FrameData[6]),
    .X(FrameData_O[6]));
 sg13g2_buf_1 _07_ (.A(FrameData[7]),
    .X(FrameData_O[7]));
 sg13g2_buf_1 _08_ (.A(FrameData[8]),
    .X(FrameData_O[8]));
 sg13g2_buf_1 _09_ (.A(FrameData[9]),
    .X(FrameData_O[9]));
 sg13g2_buf_1 _10_ (.A(FrameData[10]),
    .X(FrameData_O[10]));
 sg13g2_buf_1 _11_ (.A(FrameData[11]),
    .X(FrameData_O[11]));
 sg13g2_buf_1 _12_ (.A(FrameData[12]),
    .X(FrameData_O[12]));
 sg13g2_buf_1 _13_ (.A(FrameData[13]),
    .X(FrameData_O[13]));
 sg13g2_buf_1 _14_ (.A(FrameData[14]),
    .X(FrameData_O[14]));
 sg13g2_buf_1 _15_ (.A(FrameData[15]),
    .X(FrameData_O[15]));
 sg13g2_buf_1 _16_ (.A(FrameData[16]),
    .X(FrameData_O[16]));
 sg13g2_buf_1 _17_ (.A(FrameData[17]),
    .X(FrameData_O[17]));
 sg13g2_buf_1 _18_ (.A(FrameData[18]),
    .X(FrameData_O[18]));
 sg13g2_buf_1 _19_ (.A(FrameData[19]),
    .X(FrameData_O[19]));
 sg13g2_buf_1 _20_ (.A(FrameData[20]),
    .X(FrameData_O[20]));
 sg13g2_buf_1 _21_ (.A(FrameData[21]),
    .X(FrameData_O[21]));
 sg13g2_buf_1 _22_ (.A(FrameData[22]),
    .X(FrameData_O[22]));
 sg13g2_buf_1 _23_ (.A(FrameData[23]),
    .X(FrameData_O[23]));
 sg13g2_buf_1 _24_ (.A(FrameData[24]),
    .X(FrameData_O[24]));
 sg13g2_buf_1 _25_ (.A(FrameData[25]),
    .X(FrameData_O[25]));
 sg13g2_buf_1 _26_ (.A(FrameData[26]),
    .X(FrameData_O[26]));
 sg13g2_buf_1 _27_ (.A(FrameData[27]),
    .X(FrameData_O[27]));
 sg13g2_buf_1 _28_ (.A(FrameData[28]),
    .X(FrameData_O[28]));
 sg13g2_buf_1 _29_ (.A(FrameData[29]),
    .X(FrameData_O[29]));
 sg13g2_buf_1 _30_ (.A(FrameData[30]),
    .X(FrameData_O[30]));
 sg13g2_buf_1 _31_ (.A(FrameData[31]),
    .X(FrameData_O[31]));
 sg13g2_buf_1 _32_ (.A(FrameStrobe[0]),
    .X(FrameStrobe_O[0]));
 sg13g2_buf_1 _33_ (.A(FrameStrobe[1]),
    .X(FrameStrobe_O[1]));
 sg13g2_buf_1 _34_ (.A(FrameStrobe[2]),
    .X(FrameStrobe_O[2]));
 sg13g2_buf_1 _35_ (.A(FrameStrobe[3]),
    .X(FrameStrobe_O[3]));
 sg13g2_buf_1 _36_ (.A(FrameStrobe[4]),
    .X(FrameStrobe_O[4]));
 sg13g2_buf_1 _37_ (.A(FrameStrobe[5]),
    .X(FrameStrobe_O[5]));
 sg13g2_buf_1 _38_ (.A(FrameStrobe[6]),
    .X(FrameStrobe_O[6]));
 sg13g2_buf_1 _39_ (.A(FrameStrobe[7]),
    .X(FrameStrobe_O[7]));
 sg13g2_buf_1 _40_ (.A(FrameStrobe[8]),
    .X(FrameStrobe_O[8]));
 sg13g2_buf_1 _41_ (.A(FrameStrobe[9]),
    .X(FrameStrobe_O[9]));
 sg13g2_buf_1 _42_ (.A(FrameStrobe[10]),
    .X(FrameStrobe_O[10]));
 sg13g2_buf_1 _43_ (.A(FrameStrobe[11]),
    .X(FrameStrobe_O[11]));
 sg13g2_buf_1 _44_ (.A(FrameStrobe[12]),
    .X(FrameStrobe_O[12]));
 sg13g2_buf_1 _45_ (.A(FrameStrobe[13]),
    .X(FrameStrobe_O[13]));
 sg13g2_buf_1 _46_ (.A(FrameStrobe[14]),
    .X(FrameStrobe_O[14]));
 sg13g2_buf_1 _47_ (.A(FrameStrobe[15]),
    .X(FrameStrobe_O[15]));
 sg13g2_buf_1 _48_ (.A(FrameStrobe[16]),
    .X(FrameStrobe_O[16]));
 sg13g2_buf_1 _49_ (.A(FrameStrobe[17]),
    .X(FrameStrobe_O[17]));
 sg13g2_buf_1 _50_ (.A(FrameStrobe[18]),
    .X(FrameStrobe_O[18]));
 sg13g2_buf_1 _51_ (.A(FrameStrobe[19]),
    .X(FrameStrobe_O[19]));
 sg13g2_buf_1 _52_ (.A(N1END[3]),
    .X(S1BEG[0]));
 sg13g2_buf_1 _53_ (.A(N1END[2]),
    .X(S1BEG[1]));
 sg13g2_buf_1 _54_ (.A(N1END[1]),
    .X(S1BEG[2]));
 sg13g2_buf_1 _55_ (.A(N1END[0]),
    .X(S1BEG[3]));
 sg13g2_buf_1 _56_ (.A(N2MID[7]),
    .X(S2BEG[0]));
 sg13g2_buf_1 _57_ (.A(N2MID[6]),
    .X(S2BEG[1]));
 sg13g2_buf_1 _58_ (.A(N2MID[5]),
    .X(S2BEG[2]));
 sg13g2_buf_1 _59_ (.A(N2MID[4]),
    .X(S2BEG[3]));
 sg13g2_buf_1 _60_ (.A(N2MID[3]),
    .X(S2BEG[4]));
 sg13g2_buf_1 _61_ (.A(N2MID[2]),
    .X(S2BEG[5]));
 sg13g2_buf_1 _62_ (.A(N2MID[1]),
    .X(S2BEG[6]));
 sg13g2_buf_1 _63_ (.A(N2MID[0]),
    .X(S2BEG[7]));
 sg13g2_buf_1 _64_ (.A(N2END[7]),
    .X(S2BEGb[0]));
 sg13g2_buf_1 _65_ (.A(N2END[6]),
    .X(S2BEGb[1]));
 sg13g2_buf_1 _66_ (.A(N2END[5]),
    .X(S2BEGb[2]));
 sg13g2_buf_1 _67_ (.A(N2END[4]),
    .X(S2BEGb[3]));
 sg13g2_buf_1 _68_ (.A(N2END[3]),
    .X(S2BEGb[4]));
 sg13g2_buf_1 _69_ (.A(N2END[2]),
    .X(S2BEGb[5]));
 sg13g2_buf_1 _70_ (.A(N2END[1]),
    .X(S2BEGb[6]));
 sg13g2_buf_1 _71_ (.A(N2END[0]),
    .X(S2BEGb[7]));
 sg13g2_buf_1 _72_ (.A(N4END[15]),
    .X(S4BEG[0]));
 sg13g2_buf_1 _73_ (.A(N4END[14]),
    .X(S4BEG[1]));
 sg13g2_buf_1 _74_ (.A(N4END[13]),
    .X(S4BEG[2]));
 sg13g2_buf_1 _75_ (.A(N4END[12]),
    .X(S4BEG[3]));
 sg13g2_buf_1 _76_ (.A(N4END[11]),
    .X(S4BEG[4]));
 sg13g2_buf_1 _77_ (.A(N4END[10]),
    .X(S4BEG[5]));
 sg13g2_buf_1 _78_ (.A(N4END[9]),
    .X(S4BEG[6]));
 sg13g2_buf_1 _79_ (.A(N4END[8]),
    .X(S4BEG[7]));
 sg13g2_buf_1 _80_ (.A(N4END[7]),
    .X(S4BEG[8]));
 sg13g2_buf_1 _81_ (.A(N4END[6]),
    .X(S4BEG[9]));
 sg13g2_buf_1 _82_ (.A(N4END[5]),
    .X(S4BEG[10]));
 sg13g2_buf_1 _83_ (.A(N4END[4]),
    .X(S4BEG[11]));
 sg13g2_buf_1 _84_ (.A(N4END[3]),
    .X(S4BEG[12]));
 sg13g2_buf_1 _85_ (.A(N4END[2]),
    .X(S4BEG[13]));
 sg13g2_buf_1 _86_ (.A(N4END[1]),
    .X(S4BEG[14]));
 sg13g2_buf_1 _87_ (.A(N4END[0]),
    .X(S4BEG[15]));
 sg13g2_buf_1 _88_ (.A(UserCLK),
    .X(UserCLKo));
 sg13g2_decap_8 FILLER_0_0 ();
 sg13g2_decap_8 FILLER_0_7 ();
 sg13g2_decap_8 FILLER_0_14 ();
 sg13g2_decap_8 FILLER_0_21 ();
 sg13g2_decap_8 FILLER_0_28 ();
 sg13g2_decap_8 FILLER_0_35 ();
 sg13g2_decap_8 FILLER_0_42 ();
 sg13g2_decap_8 FILLER_0_49 ();
 sg13g2_decap_8 FILLER_0_56 ();
 sg13g2_decap_8 FILLER_0_63 ();
 sg13g2_decap_8 FILLER_0_70 ();
 sg13g2_decap_8 FILLER_0_77 ();
 sg13g2_decap_8 FILLER_0_84 ();
 sg13g2_decap_8 FILLER_0_91 ();
 sg13g2_decap_8 FILLER_0_98 ();
 sg13g2_decap_8 FILLER_0_105 ();
 sg13g2_decap_8 FILLER_0_112 ();
 sg13g2_decap_8 FILLER_0_119 ();
 sg13g2_decap_8 FILLER_0_126 ();
 sg13g2_decap_8 FILLER_0_133 ();
 sg13g2_decap_8 FILLER_0_140 ();
 sg13g2_decap_8 FILLER_0_147 ();
 sg13g2_decap_8 FILLER_0_154 ();
 sg13g2_decap_8 FILLER_0_161 ();
 sg13g2_decap_8 FILLER_0_172 ();
 sg13g2_decap_8 FILLER_0_179 ();
 sg13g2_decap_8 FILLER_0_186 ();
 sg13g2_decap_8 FILLER_0_193 ();
 sg13g2_decap_8 FILLER_1_0 ();
 sg13g2_decap_8 FILLER_1_19 ();
 sg13g2_fill_2 FILLER_1_38 ();
 sg13g2_fill_1 FILLER_1_40 ();
 sg13g2_fill_1 FILLER_1_45 ();
 sg13g2_fill_1 FILLER_1_50 ();
 sg13g2_decap_4 FILLER_1_55 ();
 sg13g2_decap_8 FILLER_1_79 ();
 sg13g2_decap_4 FILLER_1_86 ();
 sg13g2_fill_1 FILLER_1_90 ();
 sg13g2_fill_1 FILLER_1_99 ();
 sg13g2_decap_4 FILLER_1_116 ();
 sg13g2_fill_1 FILLER_1_120 ();
 sg13g2_fill_2 FILLER_1_137 ();
 sg13g2_decap_8 FILLER_1_143 ();
 sg13g2_fill_2 FILLER_1_150 ();
 sg13g2_fill_1 FILLER_1_152 ();
 sg13g2_decap_8 FILLER_1_157 ();
 sg13g2_decap_8 FILLER_1_176 ();
 sg13g2_fill_2 FILLER_1_183 ();
 sg13g2_fill_2 FILLER_1_197 ();
 sg13g2_fill_1 FILLER_1_199 ();
 sg13g2_decap_8 FILLER_2_0 ();
 sg13g2_decap_4 FILLER_2_11 ();
 sg13g2_fill_1 FILLER_2_15 ();
 sg13g2_decap_4 FILLER_2_20 ();
 sg13g2_decap_8 FILLER_2_28 ();
 sg13g2_decap_8 FILLER_2_35 ();
 sg13g2_decap_8 FILLER_2_42 ();
 sg13g2_decap_8 FILLER_2_49 ();
 sg13g2_fill_1 FILLER_2_56 ();
 sg13g2_decap_8 FILLER_2_61 ();
 sg13g2_decap_8 FILLER_2_68 ();
 sg13g2_fill_2 FILLER_2_75 ();
 sg13g2_fill_1 FILLER_2_77 ();
 sg13g2_decap_4 FILLER_2_82 ();
 sg13g2_fill_2 FILLER_2_86 ();
 sg13g2_decap_8 FILLER_2_92 ();
 sg13g2_decap_8 FILLER_2_99 ();
 sg13g2_decap_8 FILLER_2_106 ();
 sg13g2_decap_8 FILLER_2_113 ();
 sg13g2_decap_8 FILLER_2_120 ();
 sg13g2_decap_8 FILLER_2_127 ();
 sg13g2_decap_8 FILLER_2_134 ();
 sg13g2_fill_2 FILLER_2_141 ();
 sg13g2_fill_2 FILLER_2_151 ();
 sg13g2_decap_8 FILLER_2_157 ();
 sg13g2_decap_4 FILLER_2_164 ();
 sg13g2_decap_8 FILLER_2_172 ();
 sg13g2_decap_8 FILLER_2_179 ();
 sg13g2_decap_8 FILLER_2_186 ();
 sg13g2_decap_8 FILLER_2_193 ();
 sg13g2_decap_8 FILLER_3_0 ();
 sg13g2_decap_8 FILLER_3_11 ();
 sg13g2_decap_8 FILLER_3_18 ();
 sg13g2_decap_8 FILLER_3_25 ();
 sg13g2_decap_8 FILLER_3_32 ();
 sg13g2_decap_8 FILLER_3_39 ();
 sg13g2_decap_8 FILLER_3_46 ();
 sg13g2_decap_8 FILLER_3_53 ();
 sg13g2_decap_8 FILLER_3_60 ();
 sg13g2_decap_8 FILLER_3_67 ();
 sg13g2_decap_8 FILLER_3_74 ();
 sg13g2_decap_8 FILLER_3_81 ();
 sg13g2_decap_8 FILLER_3_88 ();
 sg13g2_decap_8 FILLER_3_95 ();
 sg13g2_decap_8 FILLER_3_102 ();
 sg13g2_decap_8 FILLER_3_109 ();
 sg13g2_decap_8 FILLER_3_116 ();
 sg13g2_decap_8 FILLER_3_123 ();
 sg13g2_decap_8 FILLER_3_130 ();
 sg13g2_decap_8 FILLER_3_137 ();
 sg13g2_decap_8 FILLER_3_144 ();
 sg13g2_decap_8 FILLER_3_151 ();
 sg13g2_decap_8 FILLER_3_158 ();
 sg13g2_decap_8 FILLER_3_165 ();
 sg13g2_decap_8 FILLER_3_172 ();
 sg13g2_decap_8 FILLER_3_179 ();
 sg13g2_fill_2 FILLER_3_186 ();
 sg13g2_decap_8 FILLER_3_192 ();
 sg13g2_fill_1 FILLER_3_199 ();
 sg13g2_decap_8 FILLER_4_0 ();
 sg13g2_decap_8 FILLER_4_11 ();
 sg13g2_decap_8 FILLER_4_18 ();
 sg13g2_decap_8 FILLER_4_25 ();
 sg13g2_decap_8 FILLER_4_32 ();
 sg13g2_decap_8 FILLER_4_39 ();
 sg13g2_decap_8 FILLER_4_46 ();
 sg13g2_decap_8 FILLER_4_53 ();
 sg13g2_decap_8 FILLER_4_60 ();
 sg13g2_decap_8 FILLER_4_67 ();
 sg13g2_decap_8 FILLER_4_74 ();
 sg13g2_decap_8 FILLER_4_81 ();
 sg13g2_decap_8 FILLER_4_88 ();
 sg13g2_decap_8 FILLER_4_95 ();
 sg13g2_decap_8 FILLER_4_102 ();
 sg13g2_decap_8 FILLER_4_109 ();
 sg13g2_decap_8 FILLER_4_116 ();
 sg13g2_decap_8 FILLER_4_123 ();
 sg13g2_decap_8 FILLER_4_130 ();
 sg13g2_decap_8 FILLER_4_137 ();
 sg13g2_decap_8 FILLER_4_144 ();
 sg13g2_decap_8 FILLER_4_151 ();
 sg13g2_decap_8 FILLER_4_158 ();
 sg13g2_decap_8 FILLER_4_165 ();
 sg13g2_decap_8 FILLER_4_172 ();
 sg13g2_decap_4 FILLER_4_179 ();
 sg13g2_decap_4 FILLER_4_195 ();
 sg13g2_fill_1 FILLER_4_199 ();
 sg13g2_decap_8 FILLER_5_0 ();
 sg13g2_decap_8 FILLER_5_11 ();
 sg13g2_decap_8 FILLER_5_18 ();
 sg13g2_decap_8 FILLER_5_25 ();
 sg13g2_decap_8 FILLER_5_32 ();
 sg13g2_decap_8 FILLER_5_39 ();
 sg13g2_decap_8 FILLER_5_46 ();
 sg13g2_decap_8 FILLER_5_53 ();
 sg13g2_decap_8 FILLER_5_60 ();
 sg13g2_decap_8 FILLER_5_67 ();
 sg13g2_decap_8 FILLER_5_74 ();
 sg13g2_decap_8 FILLER_5_81 ();
 sg13g2_decap_8 FILLER_5_88 ();
 sg13g2_decap_8 FILLER_5_95 ();
 sg13g2_decap_8 FILLER_5_102 ();
 sg13g2_decap_8 FILLER_5_109 ();
 sg13g2_decap_8 FILLER_5_116 ();
 sg13g2_decap_8 FILLER_5_123 ();
 sg13g2_decap_8 FILLER_5_130 ();
 sg13g2_decap_8 FILLER_5_137 ();
 sg13g2_decap_8 FILLER_5_144 ();
 sg13g2_decap_8 FILLER_5_151 ();
 sg13g2_fill_2 FILLER_5_158 ();
 sg13g2_fill_1 FILLER_5_160 ();
 sg13g2_fill_2 FILLER_5_165 ();
 sg13g2_decap_8 FILLER_5_171 ();
 sg13g2_decap_8 FILLER_5_178 ();
 sg13g2_decap_8 FILLER_5_185 ();
 sg13g2_decap_8 FILLER_5_192 ();
 sg13g2_fill_1 FILLER_5_199 ();
 sg13g2_decap_8 FILLER_6_0 ();
 sg13g2_decap_8 FILLER_6_11 ();
 sg13g2_decap_8 FILLER_6_18 ();
 sg13g2_decap_8 FILLER_6_25 ();
 sg13g2_decap_8 FILLER_6_32 ();
 sg13g2_decap_8 FILLER_6_39 ();
 sg13g2_decap_8 FILLER_6_46 ();
 sg13g2_decap_8 FILLER_6_53 ();
 sg13g2_decap_8 FILLER_6_60 ();
 sg13g2_decap_8 FILLER_6_67 ();
 sg13g2_decap_8 FILLER_6_74 ();
 sg13g2_decap_8 FILLER_6_81 ();
 sg13g2_decap_8 FILLER_6_88 ();
 sg13g2_decap_8 FILLER_6_95 ();
 sg13g2_decap_8 FILLER_6_102 ();
 sg13g2_decap_8 FILLER_6_109 ();
 sg13g2_decap_8 FILLER_6_116 ();
 sg13g2_decap_8 FILLER_6_123 ();
 sg13g2_decap_8 FILLER_6_130 ();
 sg13g2_decap_8 FILLER_6_137 ();
 sg13g2_decap_8 FILLER_6_144 ();
 sg13g2_decap_8 FILLER_6_151 ();
 sg13g2_decap_8 FILLER_6_158 ();
 sg13g2_decap_8 FILLER_6_165 ();
 sg13g2_decap_8 FILLER_6_172 ();
 sg13g2_decap_8 FILLER_6_179 ();
 sg13g2_fill_1 FILLER_6_186 ();
 sg13g2_decap_8 FILLER_6_191 ();
 sg13g2_fill_2 FILLER_6_198 ();
 sg13g2_decap_4 FILLER_7_0 ();
 sg13g2_fill_2 FILLER_7_4 ();
 sg13g2_decap_8 FILLER_7_18 ();
 sg13g2_decap_8 FILLER_7_25 ();
 sg13g2_decap_8 FILLER_7_32 ();
 sg13g2_decap_8 FILLER_7_39 ();
 sg13g2_decap_8 FILLER_7_46 ();
 sg13g2_decap_8 FILLER_7_53 ();
 sg13g2_decap_8 FILLER_7_60 ();
 sg13g2_decap_8 FILLER_7_67 ();
 sg13g2_decap_8 FILLER_7_74 ();
 sg13g2_decap_8 FILLER_7_81 ();
 sg13g2_decap_8 FILLER_7_88 ();
 sg13g2_decap_8 FILLER_7_95 ();
 sg13g2_decap_8 FILLER_7_102 ();
 sg13g2_decap_8 FILLER_7_109 ();
 sg13g2_decap_8 FILLER_7_116 ();
 sg13g2_decap_8 FILLER_7_123 ();
 sg13g2_decap_8 FILLER_7_130 ();
 sg13g2_decap_8 FILLER_7_137 ();
 sg13g2_decap_8 FILLER_7_144 ();
 sg13g2_decap_8 FILLER_7_151 ();
 sg13g2_decap_8 FILLER_7_158 ();
 sg13g2_decap_8 FILLER_7_165 ();
 sg13g2_fill_2 FILLER_7_172 ();
 sg13g2_decap_8 FILLER_7_178 ();
 sg13g2_fill_2 FILLER_7_185 ();
 sg13g2_fill_1 FILLER_7_187 ();
 sg13g2_decap_4 FILLER_7_196 ();
 sg13g2_decap_8 FILLER_8_0 ();
 sg13g2_decap_8 FILLER_8_7 ();
 sg13g2_decap_8 FILLER_8_14 ();
 sg13g2_decap_8 FILLER_8_21 ();
 sg13g2_decap_8 FILLER_8_28 ();
 sg13g2_decap_8 FILLER_8_35 ();
 sg13g2_decap_8 FILLER_8_42 ();
 sg13g2_decap_8 FILLER_8_49 ();
 sg13g2_decap_8 FILLER_8_56 ();
 sg13g2_decap_8 FILLER_8_63 ();
 sg13g2_decap_8 FILLER_8_70 ();
 sg13g2_decap_8 FILLER_8_77 ();
 sg13g2_decap_8 FILLER_8_84 ();
 sg13g2_decap_8 FILLER_8_91 ();
 sg13g2_decap_8 FILLER_8_98 ();
 sg13g2_decap_8 FILLER_8_105 ();
 sg13g2_decap_8 FILLER_8_112 ();
 sg13g2_decap_8 FILLER_8_119 ();
 sg13g2_decap_8 FILLER_8_126 ();
 sg13g2_decap_8 FILLER_8_133 ();
 sg13g2_decap_8 FILLER_8_140 ();
 sg13g2_decap_8 FILLER_8_147 ();
 sg13g2_decap_8 FILLER_8_154 ();
 sg13g2_decap_8 FILLER_8_161 ();
 sg13g2_decap_8 FILLER_8_168 ();
 sg13g2_decap_8 FILLER_8_175 ();
 sg13g2_decap_4 FILLER_8_182 ();
 sg13g2_fill_2 FILLER_8_186 ();
 sg13g2_decap_8 FILLER_8_192 ();
 sg13g2_fill_1 FILLER_8_199 ();
 sg13g2_decap_8 FILLER_9_0 ();
 sg13g2_fill_2 FILLER_9_7 ();
 sg13g2_fill_1 FILLER_9_9 ();
 sg13g2_decap_8 FILLER_9_14 ();
 sg13g2_decap_8 FILLER_9_21 ();
 sg13g2_decap_8 FILLER_9_28 ();
 sg13g2_decap_8 FILLER_9_35 ();
 sg13g2_decap_8 FILLER_9_42 ();
 sg13g2_decap_8 FILLER_9_49 ();
 sg13g2_decap_8 FILLER_9_56 ();
 sg13g2_decap_8 FILLER_9_63 ();
 sg13g2_decap_8 FILLER_9_70 ();
 sg13g2_decap_8 FILLER_9_77 ();
 sg13g2_decap_8 FILLER_9_84 ();
 sg13g2_decap_8 FILLER_9_91 ();
 sg13g2_decap_8 FILLER_9_98 ();
 sg13g2_decap_8 FILLER_9_105 ();
 sg13g2_decap_8 FILLER_9_112 ();
 sg13g2_decap_8 FILLER_9_119 ();
 sg13g2_fill_2 FILLER_9_126 ();
 sg13g2_fill_1 FILLER_9_128 ();
 sg13g2_decap_8 FILLER_9_133 ();
 sg13g2_decap_8 FILLER_9_140 ();
 sg13g2_decap_8 FILLER_9_147 ();
 sg13g2_decap_8 FILLER_9_154 ();
 sg13g2_decap_8 FILLER_9_161 ();
 sg13g2_decap_8 FILLER_9_168 ();
 sg13g2_decap_8 FILLER_9_175 ();
 sg13g2_decap_8 FILLER_9_182 ();
 sg13g2_decap_8 FILLER_9_189 ();
 sg13g2_decap_4 FILLER_9_196 ();
 sg13g2_fill_2 FILLER_10_0 ();
 sg13g2_fill_1 FILLER_10_2 ();
 sg13g2_decap_8 FILLER_10_15 ();
 sg13g2_fill_1 FILLER_10_22 ();
 sg13g2_decap_4 FILLER_10_31 ();
 sg13g2_fill_2 FILLER_10_35 ();
 sg13g2_decap_4 FILLER_10_41 ();
 sg13g2_fill_2 FILLER_10_45 ();
 sg13g2_decap_4 FILLER_10_51 ();
 sg13g2_fill_1 FILLER_10_55 ();
 sg13g2_decap_8 FILLER_10_60 ();
 sg13g2_fill_2 FILLER_10_67 ();
 sg13g2_decap_4 FILLER_10_73 ();
 sg13g2_fill_2 FILLER_10_77 ();
 sg13g2_fill_2 FILLER_10_83 ();
 sg13g2_decap_8 FILLER_10_89 ();
 sg13g2_decap_4 FILLER_10_100 ();
 sg13g2_decap_8 FILLER_10_116 ();
 sg13g2_decap_8 FILLER_10_127 ();
 sg13g2_decap_8 FILLER_10_138 ();
 sg13g2_fill_2 FILLER_10_145 ();
 sg13g2_fill_1 FILLER_10_147 ();
 sg13g2_fill_2 FILLER_10_152 ();
 sg13g2_fill_1 FILLER_10_154 ();
 sg13g2_decap_4 FILLER_10_167 ();
 sg13g2_fill_2 FILLER_10_175 ();
 sg13g2_decap_4 FILLER_10_181 ();
 sg13g2_fill_2 FILLER_10_197 ();
 sg13g2_fill_1 FILLER_10_199 ();
 sg13g2_decap_8 FILLER_11_0 ();
 sg13g2_decap_8 FILLER_11_7 ();
 sg13g2_decap_8 FILLER_11_14 ();
 sg13g2_decap_8 FILLER_11_21 ();
 sg13g2_decap_8 FILLER_11_28 ();
 sg13g2_decap_8 FILLER_11_35 ();
 sg13g2_decap_8 FILLER_11_42 ();
 sg13g2_decap_8 FILLER_11_49 ();
 sg13g2_decap_8 FILLER_11_56 ();
 sg13g2_decap_8 FILLER_11_63 ();
 sg13g2_decap_8 FILLER_11_70 ();
 sg13g2_decap_8 FILLER_11_77 ();
 sg13g2_decap_8 FILLER_11_84 ();
 sg13g2_decap_8 FILLER_11_91 ();
 sg13g2_decap_8 FILLER_11_98 ();
 sg13g2_decap_8 FILLER_11_105 ();
 sg13g2_decap_8 FILLER_11_112 ();
 sg13g2_decap_8 FILLER_11_119 ();
 sg13g2_decap_8 FILLER_11_126 ();
 sg13g2_decap_8 FILLER_11_133 ();
 sg13g2_decap_8 FILLER_11_140 ();
 sg13g2_decap_8 FILLER_11_147 ();
 sg13g2_decap_8 FILLER_11_154 ();
 sg13g2_decap_8 FILLER_11_161 ();
 sg13g2_decap_8 FILLER_11_168 ();
 sg13g2_decap_8 FILLER_11_175 ();
 sg13g2_decap_8 FILLER_11_182 ();
 sg13g2_decap_8 FILLER_11_189 ();
 sg13g2_decap_4 FILLER_11_196 ();
endmodule
