* NGSPICE file created from N_IO4.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

.subckt N_IO4 A_I_top A_O_top A_T_top B_I_top B_O_top B_T_top C_I_top C_O_top C_T_top
+ Ci D_I_top D_O_top D_T_top FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1END[0] N1END[1]
+ N1END[2] N1END[3] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4] N2END[5] N2END[6]
+ N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3] S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7]
+ S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4] S2BEGb[5] S2BEGb[6] S2BEGb[7]
+ S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1] S4BEG[2]
+ S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] SS4BEG[0] SS4BEG[10]
+ SS4BEG[11] SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3]
+ SS4BEG[4] SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] UserCLK UserCLKo VGND
+ VPWR
X_294_ FrameData[4] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
X_432_ Inst_N_IO4_switch_matrix.S2BEGb6 S2BEGb[6] VPWR VGND sg13g2_buf_1
X_363_ FrameData[1] FrameData_O[1] VPWR VGND sg13g2_buf_1
XFILLER_5_332 VPWR VGND sg13g2_fill_1
X_346_ FrameData[24] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_415_ Inst_N_IO4_switch_matrix.S1BEG1 S1BEG[1] VPWR VGND sg13g2_buf_1
X_277_ FrameData[19] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_11_423 VPWR VGND sg13g2_fill_1
X_131_ Inst_N_IO4_ConfigMem.Inst_frame0_bit28.Q VPWR _034_ VGND _026_ _029_ sg13g2_o21ai_1
X_200_ Inst_N_IO4_ConfigMem.Inst_frame2_bit26.Q N4END[8] NN4END[8] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_D_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame2_bit27.Q
+ Inst_N_IO4_switch_matrix.S4BEG11 VPWR VGND sg13g2_mux4_1
X_329_ FrameData[7] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
X_114_ _018_ VPWR C_T_top VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit24.Q _015_ sg13g2_o21ai_1
XFILLER_0_411 VPWR VGND sg13g2_fill_2
XFILLER_4_238 VPWR VGND sg13g2_fill_1
XFILLER_8_385 VPWR VGND sg13g2_fill_2
XFILLER_11_0 VPWR VGND sg13g2_fill_2
X_362_ FrameData[0] FrameData_O[0] VPWR VGND sg13g2_buf_1
X_293_ FrameData[3] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_3_79 VPWR VGND sg13g2_fill_2
X_431_ Inst_N_IO4_switch_matrix.S2BEGb5 S2BEGb[5] VPWR VGND sg13g2_buf_1
X_345_ FrameData[23] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_276_ FrameData[18] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_414_ Inst_N_IO4_switch_matrix.S1BEG0 S1BEG[0] VPWR VGND sg13g2_buf_1
X_130_ VPWR VGND _032_ Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q _031_ Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q
+ _033_ _030_ sg13g2_a221oi_1
X_259_ FrameData[1] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
X_328_ FrameData[6] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
X_113_ _018_ _016_ _017_ VPWR VGND sg13g2_nand2b_1
XFILLER_0_423 VPWR VGND sg13g2_fill_1
X_292_ FrameData[2] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
X_430_ Inst_N_IO4_switch_matrix.S2BEGb4 S2BEGb[4] VPWR VGND sg13g2_buf_1
X_361_ VPWR VGND _082_ sg13g2_tiehi
XFILLER_2_348 VPWR VGND sg13g2_fill_2
X_413_ FrameStrobe[19] FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_275_ FrameData[17] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_344_ FrameData[22] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_2_178 VPWR VGND sg13g2_decap_8
X_189_ Inst_N_IO4_ConfigMem.Inst_frame1_bit17.Q N2MID[2] N2MID[6] N2MID[4] C_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit16.Q Inst_N_IO4_switch_matrix.SS4BEG6 VPWR VGND
+ sg13g2_mux4_1
X_327_ FrameData[5] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_258_ FrameData[0] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
X_112_ Inst_N_IO4_ConfigMem.Inst_frame0_bit24.Q VPWR _017_ VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q
+ _014_ sg13g2_o21ai_1
XFILLER_1_0 VPWR VGND sg13g2_fill_1
XFILLER_3_421 VPWR VGND sg13g2_fill_2
XFILLER_8_387 VPWR VGND sg13g2_fill_1
X_360_ VPWR VGND _081_ sg13g2_tiehi
X_291_ FrameData[1] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
X_412_ FrameStrobe[18] FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_343_ FrameData[21] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_274_ FrameData[16] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_187 VPWR VGND sg13g2_decap_8
XFILLER_2_157 VPWR VGND sg13g2_decap_8
XFILLER_9_36 VPWR VGND sg13g2_fill_2
X_326_ FrameData[4] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
X_257_ FrameData[31] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_188_ Inst_N_IO4_ConfigMem.Inst_frame1_bit18.Q N2MID[3] N2MID[5] N2MID[7] D_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit19.Q Inst_N_IO4_switch_matrix.SS4BEG7 VPWR VGND
+ sg13g2_mux4_1
X_309_ FrameData[19] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_111_ Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q VPWR _016_ VGND N2END[6] Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q
+ sg13g2_o21ai_1
XFILLER_0_200 VPWR VGND sg13g2_fill_2
X_290_ FrameData[0] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_5_358 VPWR VGND sg13g2_fill_1
X_411_ FrameStrobe[17] FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_273_ FrameData[15] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_342_ FrameData[20] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_187_ Inst_N_IO4_ConfigMem.Inst_frame1_bit20.Q N4END[6] N4END[8] N4END[10] Inst_C_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit21.Q Inst_N_IO4_switch_matrix.SS4BEG8 VPWR VGND
+ sg13g2_mux4_1
X_325_ FrameData[3] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
X_256_ FrameData[30] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_110_ Inst_N_IO4_ConfigMem.Inst_frame0_bit22.Q N2MID[6] N2MID[7] N2END[0] N2END[4]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q _015_ VPWR VGND sg13g2_mux4_1
XFILLER_3_423 VPWR VGND sg13g2_fill_1
X_308_ FrameData[18] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_239_ FrameData[13] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_410_ FrameStrobe[16] FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
X_272_ FrameData[14] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_341_ FrameData[19] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_4_71 VPWR VGND sg13g2_fill_2
X_255_ FrameData[29] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_324_ FrameData[2] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_6_421 VPWR VGND sg13g2_fill_2
X_186_ Inst_N_IO4_ConfigMem.Inst_frame1_bit22.Q N4END[3] N4END[5] N4END[7] Inst_D_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit23.Q Inst_N_IO4_switch_matrix.SS4BEG9 VPWR VGND
+ sg13g2_mux4_1
X_307_ FrameData[17] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_1_61 VPWR VGND sg13g2_fill_2
X_169_ Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q VPWR _069_ VGND N2END[6] Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q
+ sg13g2_o21ai_1
X_238_ FrameData[12] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_0_202 VPWR VGND sg13g2_fill_1
X_340_ FrameData[18] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_271_ FrameData[13] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_135 VPWR VGND sg13g2_decap_8
XFILLER_4_190 VPWR VGND sg13g2_decap_4
X_254_ FrameData[28] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_323_ FrameData[1] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
X_185_ Inst_N_IO4_ConfigMem.Inst_frame1_bit24.Q N4END[0] N4END[2] N4END[4] A_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit25.Q Inst_N_IO4_switch_matrix.SS4BEG10 VPWR
+ VGND sg13g2_mux4_1
X_306_ FrameData[16] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_168_ N2END[7] Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q _068_ VPWR VGND sg13g2_nor2b_1
X_237_ FrameData[11] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_099_ Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q
+ _006_ VPWR VGND sg13g2_nor2_1
XFILLER_6_274 VPWR VGND sg13g2_fill_1
XFILLER_3_222 VPWR VGND sg13g2_fill_2
XFILLER_3_277 VPWR VGND sg13g2_fill_2
X_270_ FrameData[12] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_399_ FrameStrobe[5] FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
X_322_ FrameData[0] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
X_253_ FrameData[27] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_184_ Inst_N_IO4_ConfigMem.Inst_frame1_bit26.Q N4END[6] N4END[8] N4END[10] B_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit27.Q Inst_N_IO4_switch_matrix.SS4BEG11 VPWR
+ VGND sg13g2_mux4_1
XFILLER_6_423 VPWR VGND sg13g2_fill_1
XFILLER_11_227 VPWR VGND sg13g2_fill_2
X_098_ Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q VPWR _005_ VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q
+ N2END[4] sg13g2_o21ai_1
X_167_ VPWR VGND _066_ Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q _065_ Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q
+ _067_ _064_ sg13g2_a221oi_1
X_236_ FrameData[10] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_305_ FrameData[15] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_6_231 VPWR VGND sg13g2_decap_4
XFILLER_10_50 VPWR VGND sg13g2_fill_1
XFILLER_3_245 VPWR VGND sg13g2_fill_2
X_219_ Inst_N_IO4_ConfigMem.Inst_frame3_bit21.Q N2END[7] NN4END[7] N4END[7] NN4END[15]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit20.Q Inst_N_IO4_switch_matrix.S2BEGb0 VPWR VGND
+ sg13g2_mux4_1
XFILLER_1_343 VPWR VGND sg13g2_fill_1
X_398_ FrameStrobe[4] FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
X_252_ FrameData[26] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_183_ Inst_N_IO4_ConfigMem.Inst_frame1_bit29.Q N4END[1] N4END[5] N4END[3] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit28.Q Inst_N_IO4_switch_matrix.SS4BEG12 VPWR
+ VGND sg13g2_mux4_1
X_321_ FrameData[31] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_6_402 VPWR VGND sg13g2_fill_1
X_235_ FrameData[9] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
X_304_ FrameData[14] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_166_ VGND VPWR _000_ Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q _066_ Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q
+ sg13g2_a21oi_1
X_097_ Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q N2MID[7] N2END[0] N2END[1] N2END[2]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q _004_ VPWR VGND sg13g2_mux4_1
XFILLER_6_265 VPWR VGND sg13g2_decap_4
XFILLER_3_279 VPWR VGND sg13g2_fill_1
X_149_ N2MID[4] N2MID[5] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q _051_ VPWR VGND
+ sg13g2_mux2_1
X_218_ Inst_N_IO4_ConfigMem.Inst_frame3_bit23.Q N2END[6] NN4END[6] N4END[6] NN4END[14]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit22.Q Inst_N_IO4_switch_matrix.S2BEGb1 VPWR VGND
+ sg13g2_mux4_1
XFILLER_7_393 VPWR VGND sg13g2_fill_2
X_466_ clknet_1_0__leaf_UserCLK UserCLKo VPWR VGND sg13g2_buf_1
X_397_ FrameStrobe[3] FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
X_251_ FrameData[25] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_10_421 VPWR VGND sg13g2_fill_2
XFILLER_1_196 VPWR VGND sg13g2_decap_8
XFILLER_1_130 VPWR VGND sg13g2_fill_1
X_182_ Inst_N_IO4_ConfigMem.Inst_frame1_bit30.Q N4END[7] N4END[9] N4END[11] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit31.Q Inst_N_IO4_switch_matrix.SS4BEG13 VPWR
+ VGND sg13g2_mux4_1
X_320_ FrameData[30] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_449_ Inst_N_IO4_switch_matrix.S4BEG15 S4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_10_273 VPWR VGND sg13g2_fill_2
X_165_ VGND VPWR _065_ Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q N2END[0] sg13g2_or2_1
X_096_ Inst_N_IO4_ConfigMem.Inst_frame4_bit29.Q N1END[2] A_O_top N1END[3] C_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame4_bit28.Q Inst_N_IO4_switch_matrix.S1BEG0 VPWR VGND
+ sg13g2_mux4_1
X_234_ FrameData[8] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
X_303_ FrameData[13] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_6_222 VPWR VGND sg13g2_fill_1
X_217_ Inst_N_IO4_ConfigMem.Inst_frame3_bit25.Q N2END[5] NN4END[5] N4END[5] NN4END[13]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit24.Q Inst_N_IO4_switch_matrix.S2BEGb2 VPWR VGND
+ sg13g2_mux4_1
XFILLER_10_85 VPWR VGND sg13g2_fill_1
X_148_ N2MID[6] N2MID[7] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q _050_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_3_247 VPWR VGND sg13g2_fill_1
XFILLER_8_328 VPWR VGND sg13g2_fill_2
XFILLER_7_86 VPWR VGND sg13g2_fill_1
XFILLER_9_423 VPWR VGND sg13g2_fill_1
X_396_ FrameStrobe[2] FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
X_465_ Inst_N_IO4_switch_matrix.SS4BEG15 SS4BEG[15] VPWR VGND sg13g2_buf_1
XFILLER_4_194 VPWR VGND sg13g2_fill_2
X_250_ FrameData[24] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_181_ Inst_N_IO4_ConfigMem.Inst_frame0_bit0.Q N2MID[0] N2MID[2] N2MID[4] C_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit1.Q Inst_N_IO4_switch_matrix.SS4BEG14 VPWR VGND
+ sg13g2_mux4_1
X_448_ Inst_N_IO4_switch_matrix.S4BEG14 S4BEG[14] VPWR VGND sg13g2_buf_1
X_379_ FrameData[17] FrameData_O[17] VPWR VGND sg13g2_buf_1
X_164_ N2END[2] N2END[3] Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q _064_ VPWR VGND sg13g2_mux2_1
X_233_ FrameData[7] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
X_095_ Inst_N_IO4_ConfigMem.Inst_frame4_bit30.Q N1END[1] N1END[2] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_C_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame4_bit31.Q
+ Inst_N_IO4_switch_matrix.S1BEG1 VPWR VGND sg13g2_mux4_1
X_302_ FrameData[12] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_147_ N2MID[0] N2MID[1] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q _049_ VPWR VGND
+ sg13g2_mux2_1
X_216_ Inst_N_IO4_ConfigMem.Inst_frame3_bit27.Q N2END[4] NN4END[4] N4END[4] NN4END[12]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit26.Q Inst_N_IO4_switch_matrix.S2BEGb3 VPWR VGND
+ sg13g2_mux4_1
XFILLER_7_54 VPWR VGND sg13g2_fill_1
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_0__leaf_UserCLK_regs VPWR
+ VGND sg13g2_buf_8
X_464_ Inst_N_IO4_switch_matrix.SS4BEG14 SS4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_4_162 VPWR VGND sg13g2_decap_8
X_395_ FrameStrobe[1] FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
XFILLER_10_423 VPWR VGND sg13g2_fill_1
XFILLER_10_412 VPWR VGND sg13g2_fill_1
X_180_ Inst_N_IO4_ConfigMem.Inst_frame0_bit3.Q N2MID[1] N2MID[5] N2MID[3] D_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit2.Q Inst_N_IO4_switch_matrix.SS4BEG15 VPWR VGND
+ sg13g2_mux4_1
XFILLER_9_287 VPWR VGND sg13g2_fill_2
X_447_ Inst_N_IO4_switch_matrix.S4BEG13 S4BEG[13] VPWR VGND sg13g2_buf_1
X_378_ FrameData[16] FrameData_O[16] VPWR VGND sg13g2_buf_1
X_094_ Inst_N_IO4_ConfigMem.Inst_frame3_bit0.Q N1END[0] N1END[1] B_O_top D_O_top Inst_N_IO4_ConfigMem.Inst_frame3_bit1.Q
+ Inst_N_IO4_switch_matrix.S1BEG2 VPWR VGND sg13g2_mux4_1
X_301_ FrameData[11] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_232_ FrameData[6] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
X_163_ _063_ VPWR B_I_top VGND _058_ _059_ sg13g2_o21ai_1
XFILLER_6_235 VPWR VGND sg13g2_fill_1
X_215_ Inst_N_IO4_ConfigMem.Inst_frame3_bit29.Q N2END[3] NN4END[3] N4END[3] NN4END[11]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit28.Q Inst_N_IO4_switch_matrix.S2BEGb4 VPWR VGND
+ sg13g2_mux4_1
X_146_ N2MID[2] N2MID[3] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q _048_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_7_22 VPWR VGND sg13g2_fill_2
XFILLER_7_374 VPWR VGND sg13g2_fill_2
X_129_ VGND VPWR _000_ Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q _032_ Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q
+ sg13g2_a21oi_1
X_463_ Inst_N_IO4_switch_matrix.SS4BEG13 SS4BEG[13] VPWR VGND sg13g2_buf_1
X_394_ FrameStrobe[0] FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
X_446_ Inst_N_IO4_switch_matrix.S4BEG12 S4BEG[12] VPWR VGND sg13g2_buf_1
X_377_ FrameData[15] FrameData_O[15] VPWR VGND sg13g2_buf_1
X_231_ FrameData[5] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_093_ Inst_N_IO4_ConfigMem.Inst_frame3_bit2.Q N1END[0] N1END[3] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_D_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame3_bit3.Q
+ Inst_N_IO4_switch_matrix.S1BEG3 VPWR VGND sg13g2_mux4_1
X_300_ FrameData[10] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_162_ _063_ _062_ Inst_N_IO4_ConfigMem.Inst_frame0_bit14.Q VPWR VGND sg13g2_nand2b_1
XFILLER_6_269 VPWR VGND sg13g2_fill_1
XFILLER_5_291 VPWR VGND sg13g2_fill_1
X_429_ Inst_N_IO4_switch_matrix.S2BEGb3 S2BEGb[3] VPWR VGND sg13g2_buf_1
X_145_ VPWR VGND _046_ _002_ _044_ _041_ _047_ _042_ sg13g2_a221oi_1
X_214_ Inst_N_IO4_ConfigMem.Inst_frame3_bit30.Q N2END[2] N4END[2] NN4END[2] NN4END[10]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit31.Q Inst_N_IO4_switch_matrix.S2BEGb5 VPWR VGND
+ sg13g2_mux4_1
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK clknet_1_0__leaf_UserCLK VPWR VGND sg13g2_buf_8
X_128_ VGND VPWR _031_ Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q N2END[0] sg13g2_or2_1
XFILLER_7_172 VPWR VGND sg13g2_fill_2
X_393_ FrameData[31] FrameData_O[31] VPWR VGND sg13g2_buf_1
X_462_ Inst_N_IO4_switch_matrix.SS4BEG12 SS4BEG[12] VPWR VGND sg13g2_buf_1
XFILLER_1_156 VPWR VGND sg13g2_fill_2
XFILLER_6_407 VPWR VGND sg13g2_fill_2
X_376_ FrameData[14] FrameData_O[14] VPWR VGND sg13g2_buf_1
X_445_ Inst_N_IO4_switch_matrix.S4BEG11 S4BEG[11] VPWR VGND sg13g2_buf_1
XFILLER_10_200 VPWR VGND sg13g2_fill_1
X_230_ FrameData[4] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
X_161_ _060_ _061_ Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q _062_ VPWR VGND sg13g2_mux2_1
X_428_ Inst_N_IO4_switch_matrix.S2BEGb2 S2BEGb[2] VPWR VGND sg13g2_buf_1
X_092_ Inst_N_IO4_ConfigMem.Inst_frame3_bit4.Q N2MID[7] N4END[7] NN4END[7] NN4END[15]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit5.Q Inst_N_IO4_switch_matrix.S2BEG0 VPWR VGND
+ sg13g2_mux4_1
X_359_ VPWR VGND _080_ sg13g2_tiehi
XFILLER_3_218 VPWR VGND sg13g2_decap_4
X_213_ Inst_N_IO4_ConfigMem.Inst_frame2_bit0.Q N2END[1] N4END[1] NN4END[1] NN4END[9]
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit1.Q Inst_N_IO4_switch_matrix.S2BEGb6 VPWR VGND
+ sg13g2_mux4_1
X_144_ VGND VPWR Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q _045_ _046_ _001_ sg13g2_a21oi_1
X_127_ N2END[2] N2END[3] Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q _030_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_8_107 VPWR VGND sg13g2_decap_4
XFILLER_4_379 VPWR VGND sg13g2_fill_2
X_392_ FrameData[30] FrameData_O[30] VPWR VGND sg13g2_buf_1
X_461_ Inst_N_IO4_switch_matrix.SS4BEG11 SS4BEG[11] VPWR VGND sg13g2_buf_1
X_444_ Inst_N_IO4_switch_matrix.S4BEG10 S4BEG[10] VPWR VGND sg13g2_buf_1
X_375_ FrameData[13] FrameData_O[13] VPWR VGND sg13g2_buf_1
X_358_ VPWR VGND _079_ sg13g2_tiehi
Xclkbuf_regs_0_UserCLK UserCLK UserCLK_regs VPWR VGND sg13g2_buf_8
X_160_ Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q _061_ VPWR VGND sg13g2_mux4_1
X_091_ Inst_N_IO4_ConfigMem.Inst_frame3_bit6.Q N2MID[6] N4END[6] NN4END[6] NN4END[14]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit7.Q Inst_N_IO4_switch_matrix.S2BEG1 VPWR VGND
+ sg13g2_mux4_1
X_427_ Inst_N_IO4_switch_matrix.S2BEGb1 S2BEGb[1] VPWR VGND sg13g2_buf_1
XFILLER_5_260 VPWR VGND sg13g2_decap_4
X_289_ FrameData[31] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_212_ Inst_N_IO4_ConfigMem.Inst_frame2_bit2.Q N2END[0] N4END[0] NN4END[0] NN4END[8]
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit3.Q Inst_N_IO4_switch_matrix.S2BEGb7 VPWR VGND
+ sg13g2_mux4_1
X_143_ N2END[6] N2END[7] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q _045_ VPWR VGND
+ sg13g2_mux2_1
X_126_ Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q VPWR _029_ VGND _027_ _028_ sg13g2_o21ai_1
X_109_ _014_ N2END[5] Inst_N_IO4_ConfigMem.Inst_frame0_bit23.Q VPWR VGND sg13g2_nand2b_1
XFILLER_7_174 VPWR VGND sg13g2_fill_1
X_391_ FrameData[29] FrameData_O[29] VPWR VGND sg13g2_buf_1
XFILLER_1_317 VPWR VGND sg13g2_fill_1
X_460_ Inst_N_IO4_switch_matrix.SS4BEG10 SS4BEG[10] VPWR VGND sg13g2_buf_1
XFILLER_4_155 VPWR VGND sg13g2_decap_8
XFILLER_9_225 VPWR VGND sg13g2_decap_8
X_374_ FrameData[12] FrameData_O[12] VPWR VGND sg13g2_buf_1
X_443_ Inst_N_IO4_switch_matrix.S4BEG9 S4BEG[9] VPWR VGND sg13g2_buf_1
Xclkbuf_0_UserCLK_regs UserCLK_regs clknet_0_UserCLK_regs VPWR VGND sg13g2_buf_8
XFILLER_2_423 VPWR VGND sg13g2_fill_1
X_090_ Inst_N_IO4_ConfigMem.Inst_frame3_bit8.Q N2MID[5] N4END[5] NN4END[5] NN4END[13]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit9.Q Inst_N_IO4_switch_matrix.S2BEG2 VPWR VGND
+ sg13g2_mux4_1
X_357_ _080_ VGND VPWR D_O_top Inst_D_IO_1_bidirectional_frame_config_pass.Q clknet_1_1__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_426_ Inst_N_IO4_switch_matrix.S2BEGb0 S2BEGb[0] VPWR VGND sg13g2_buf_1
X_288_ FrameData[30] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_142_ _044_ _043_ Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q VPWR VGND sg13g2_nand2b_1
X_211_ Inst_N_IO4_ConfigMem.Inst_frame2_bit5.Q N4END[15] A_O_top NN4END[15] C_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit4.Q Inst_N_IO4_switch_matrix.S4BEG0 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_0 VPWR VGND sg13g2_fill_2
X_409_ FrameStrobe[15] FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_125_ Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q VPWR _028_ VGND N2END[6] Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q
+ sg13g2_o21ai_1
XFILLER_4_348 VPWR VGND sg13g2_fill_2
X_108_ _013_ VPWR B_T_top VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit17.Q _009_ sg13g2_o21ai_1
X_390_ FrameData[28] FrameData_O[28] VPWR VGND sg13g2_buf_1
X_373_ FrameData[11] FrameData_O[11] VPWR VGND sg13g2_buf_1
XFILLER_5_421 VPWR VGND sg13g2_fill_2
X_442_ Inst_N_IO4_switch_matrix.S4BEG8 S4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_10_247 VPWR VGND sg13g2_fill_1
X_287_ FrameData[29] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_356_ _079_ VGND VPWR C_O_top Inst_C_IO_1_bidirectional_frame_config_pass.Q clknet_1_0__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_425_ Inst_N_IO4_switch_matrix.S2BEG7 S2BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_10_48 VPWR VGND sg13g2_fill_2
X_408_ FrameStrobe[14] FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
X_141_ N2END[4] N2END[5] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q _043_ VPWR VGND
+ sg13g2_mux2_1
X_210_ Inst_N_IO4_ConfigMem.Inst_frame2_bit7.Q N4END[14] B_O_top NN4END[14] D_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit6.Q Inst_N_IO4_switch_matrix.S4BEG1 VPWR VGND
+ sg13g2_mux4_1
X_339_ FrameData[17] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_124_ N2END[7] Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q _027_ VPWR VGND sg13g2_nor2b_1
X_107_ _010_ _012_ Inst_N_IO4_ConfigMem.Inst_frame0_bit17.Q _013_ VPWR VGND sg13g2_nand3_1
XFILLER_3_371 VPWR VGND sg13g2_fill_1
X_372_ FrameData[10] FrameData_O[10] VPWR VGND sg13g2_buf_1
X_441_ Inst_N_IO4_switch_matrix.S4BEG7 S4BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_0_193 VPWR VGND sg13g2_decap_8
XFILLER_0_160 VPWR VGND sg13g2_decap_8
X_286_ FrameData[28] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_355_ _082_ VGND VPWR B_O_top Inst_B_IO_1_bidirectional_frame_config_pass.Q clknet_1_1__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_424_ Inst_N_IO4_switch_matrix.S2BEG6 S2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_5_241 VPWR VGND sg13g2_fill_2
X_140_ VGND VPWR Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q _039_ _042_ Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q
+ sg13g2_a21oi_1
X_338_ FrameData[16] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_269_ FrameData[11] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_1__leaf_UserCLK_regs VPWR
+ VGND sg13g2_buf_8
X_407_ FrameStrobe[13] FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
X_123_ VGND VPWR _024_ _025_ _026_ Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q sg13g2_a21oi_1
XFILLER_4_317 VPWR VGND sg13g2_fill_2
X_106_ _012_ N2END[5] _011_ VPWR VGND sg13g2_nand2_1
X_440_ Inst_N_IO4_switch_matrix.S4BEG6 S4BEG[6] VPWR VGND sg13g2_buf_1
X_371_ FrameData[9] FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_5_423 VPWR VGND sg13g2_fill_1
X_285_ FrameData[27] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_354_ _081_ VGND VPWR A_O_top Inst_A_IO_1_bidirectional_frame_config_pass.Q clknet_1_0__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_423_ Inst_N_IO4_switch_matrix.S2BEG5 S2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_10_39 VPWR VGND sg13g2_fill_2
X_406_ FrameStrobe[12] FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
X_199_ Inst_N_IO4_ConfigMem.Inst_frame2_bit28.Q N4END[5] NN4END[5] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_C_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame2_bit29.Q
+ Inst_N_IO4_switch_matrix.S4BEG12 VPWR VGND sg13g2_mux4_1
X_337_ FrameData[15] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_268_ FrameData[10] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_122_ _025_ N2END[4] Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q VPWR VGND sg13g2_nand2b_1
XFILLER_2_0 VPWR VGND sg13g2_fill_1
XFILLER_6_370 VPWR VGND sg13g2_fill_2
X_105_ Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q
+ _011_ VPWR VGND sg13g2_nor2_1
XFILLER_8_421 VPWR VGND sg13g2_fill_2
X_370_ FrameData[8] FrameData_O[8] VPWR VGND sg13g2_buf_1
XFILLER_5_95 VPWR VGND sg13g2_fill_1
X_284_ FrameData[26] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_353_ FrameData[31] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_422_ Inst_N_IO4_switch_matrix.S2BEG4 S2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_5_210 VPWR VGND sg13g2_decap_8
XFILLER_2_213 VPWR VGND sg13g2_fill_2
XFILLER_2_257 VPWR VGND sg13g2_fill_2
X_267_ FrameData[9] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
X_405_ FrameStrobe[11] FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
X_336_ FrameData[14] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_198_ Inst_N_IO4_ConfigMem.Inst_frame2_bit30.Q N4END[4] NN4END[4] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_D_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame2_bit31.Q
+ Inst_N_IO4_switch_matrix.S4BEG13 VPWR VGND sg13g2_mux4_1
X_121_ _024_ N2END[5] Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q VPWR VGND sg13g2_nand2_1
X_319_ FrameData[29] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_11_175 VPWR VGND sg13g2_fill_1
X_104_ Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q VPWR _010_ VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q
+ N2END[6] sg13g2_o21ai_1
XFILLER_3_330 VPWR VGND sg13g2_fill_1
XFILLER_0_174 VPWR VGND sg13g2_fill_2
XFILLER_10_0 VPWR VGND sg13g2_fill_1
X_421_ Inst_N_IO4_switch_matrix.S2BEG3 S2BEG[3] VPWR VGND sg13g2_buf_1
X_283_ FrameData[25] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_352_ FrameData[30] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_404_ FrameStrobe[10] FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
X_266_ FrameData[8] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
X_197_ Inst_N_IO4_ConfigMem.Inst_frame1_bit0.Q N4END[1] NN4END[1] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_C_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame1_bit1.Q
+ Inst_N_IO4_switch_matrix.S4BEG14 VPWR VGND sg13g2_mux4_1
X_335_ FrameData[13] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_120_ _023_ VPWR D_T_top VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit31.Q _020_ sg13g2_o21ai_1
XFILLER_7_306 VPWR VGND sg13g2_fill_1
X_318_ FrameData[28] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_6_372 VPWR VGND sg13g2_fill_1
X_249_ FrameData[23] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_103_ Inst_N_IO4_ConfigMem.Inst_frame0_bit15.Q N2MID[6] N2MID[7] N2END[0] N2END[4]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit16.Q _009_ VPWR VGND sg13g2_mux4_1
XFILLER_8_423 VPWR VGND sg13g2_fill_1
XFILLER_0_153 VPWR VGND sg13g2_decap_8
X_351_ FrameData[29] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_282_ FrameData[24] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_420_ Inst_N_IO4_switch_matrix.S2BEG2 S2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_5_234 VPWR VGND sg13g2_decap_8
XFILLER_5_289 VPWR VGND sg13g2_fill_2
X_403_ FrameStrobe[9] FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
X_334_ FrameData[12] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_265_ FrameData[7] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
X_196_ Inst_N_IO4_ConfigMem.Inst_frame1_bit2.Q N4END[0] NN4END[0] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_D_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame1_bit3.Q
+ Inst_N_IO4_switch_matrix.S4BEG15 VPWR VGND sg13g2_mux4_1
X_317_ FrameData[27] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_248_ FrameData[22] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_179_ _078_ VPWR A_I_top VGND _067_ _074_ sg13g2_o21ai_1
XFILLER_0_0 VPWR VGND sg13g2_fill_1
X_102_ _008_ VPWR A_T_top VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit10.Q _004_ sg13g2_o21ai_1
XFILLER_7_104 VPWR VGND sg13g2_fill_2
XFILLER_3_151 VPWR VGND sg13g2_fill_2
X_350_ FrameData[28] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_202 VPWR VGND sg13g2_decap_4
X_281_ FrameData[23] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_402_ FrameStrobe[8] FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_195_ Inst_N_IO4_ConfigMem.Inst_frame1_bit4.Q N4END[0] N4END[2] N4END[4] A_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit5.Q Inst_N_IO4_switch_matrix.SS4BEG0 VPWR VGND
+ sg13g2_mux4_1
X_264_ FrameData[6] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
X_333_ FrameData[11] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_316_ FrameData[26] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_247_ FrameData[21] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_178_ _078_ _077_ Inst_N_IO4_ConfigMem.Inst_frame0_bit7.Q VPWR VGND sg13g2_nand2b_1
X_101_ _005_ _007_ Inst_N_IO4_ConfigMem.Inst_frame0_bit10.Q _008_ VPWR VGND sg13g2_nand3_1
XFILLER_7_149 VPWR VGND sg13g2_fill_2
XFILLER_5_406 VPWR VGND sg13g2_fill_2
X_280_ FrameData[22] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_401_ FrameStrobe[7] FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
X_194_ Inst_N_IO4_ConfigMem.Inst_frame1_bit6.Q N4END[6] N4END[8] N4END[10] B_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit7.Q Inst_N_IO4_switch_matrix.SS4BEG1 VPWR VGND
+ sg13g2_mux4_1
X_263_ FrameData[5] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_332_ FrameData[10] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_11_327 VPWR VGND sg13g2_fill_2
XFILLER_11_87 VPWR VGND sg13g2_fill_2
X_315_ FrameData[25] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_10_393 VPWR VGND sg13g2_fill_2
X_246_ FrameData[20] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_177_ _075_ _076_ Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q _077_ VPWR VGND sg13g2_mux2_1
X_100_ _007_ N2END[3] _006_ VPWR VGND sg13g2_nand2_1
X_229_ FrameData[3] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_3_301 VPWR VGND sg13g2_fill_2
XFILLER_6_194 VPWR VGND sg13g2_decap_8
XFILLER_3_153 VPWR VGND sg13g2_fill_1
XFILLER_0_167 VPWR VGND sg13g2_decap_8
XFILLER_8_256 VPWR VGND sg13g2_fill_1
XFILLER_5_34 VPWR VGND sg13g2_fill_1
X_262_ FrameData[4] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit4.Q VPWR VGND
+ sg13g2_dlhq_1
X_331_ FrameData[9] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
X_193_ Inst_N_IO4_ConfigMem.Inst_frame1_bit8.Q N2END[6] N2END[7] N4END[1] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit9.Q Inst_N_IO4_switch_matrix.SS4BEG2 VPWR VGND
+ sg13g2_mux4_1
X_400_ FrameStrobe[6] FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
XFILLER_9_340 VPWR VGND sg13g2_fill_1
X_314_ FrameData[24] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_176_ Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q _076_ VPWR VGND sg13g2_mux4_1
XFILLER_6_321 VPWR VGND sg13g2_fill_2
X_245_ FrameData[19] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_6_398 VPWR VGND sg13g2_decap_4
X_228_ FrameData[2] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
X_159_ Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q N2MID[0] N2MID[1] N2MID[2] N2MID[3]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q _060_ VPWR VGND sg13g2_mux4_1
XFILLER_5_408 VPWR VGND sg13g2_fill_1
X_261_ FrameData[3] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit3.Q VPWR VGND
+ sg13g2_dlhq_1
X_192_ Inst_N_IO4_ConfigMem.Inst_frame1_bit10.Q N4END[7] N4END[9] N4END[11] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit11.Q Inst_N_IO4_switch_matrix.SS4BEG3 VPWR VGND
+ sg13g2_mux4_1
X_330_ FrameData[8] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_9_0 VPWR VGND sg13g2_fill_2
XFILLER_1_285 VPWR VGND sg13g2_fill_2
X_459_ Inst_N_IO4_switch_matrix.SS4BEG9 SS4BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_11_329 VPWR VGND sg13g2_fill_1
XFILLER_11_89 VPWR VGND sg13g2_fill_1
X_313_ FrameData[23] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_175_ Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q N2MID[0] N2MID[1] N2MID[2] N2MID[3]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q _075_ VPWR VGND sg13g2_mux4_1
X_244_ FrameData[18] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_3_369 VPWR VGND sg13g2_fill_2
X_227_ FrameData[1] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit1.Q VPWR VGND
+ sg13g2_dlhq_1
X_089_ Inst_N_IO4_ConfigMem.Inst_frame3_bit10.Q N2MID[4] N4END[4] NN4END[4] NN4END[12]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit11.Q Inst_N_IO4_switch_matrix.S2BEG3 VPWR VGND
+ sg13g2_mux4_1
X_158_ Inst_N_IO4_ConfigMem.Inst_frame0_bit14.Q VPWR _059_ VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q
+ _053_ sg13g2_o21ai_1
XFILLER_3_144 VPWR VGND sg13g2_decap_8
XFILLER_3_188 VPWR VGND sg13g2_decap_8
XFILLER_3_199 VPWR VGND sg13g2_fill_2
XFILLER_0_125 VPWR VGND sg13g2_fill_2
XFILLER_1_423 VPWR VGND sg13g2_fill_1
X_260_ FrameData[2] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit2.Q VPWR VGND
+ sg13g2_dlhq_1
X_191_ Inst_N_IO4_ConfigMem.Inst_frame1_bit12.Q N2END[0] N2END[2] N2END[4] Inst_C_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit13.Q Inst_N_IO4_switch_matrix.SS4BEG4 VPWR VGND
+ sg13g2_mux4_1
X_389_ FrameData[27] FrameData_O[27] VPWR VGND sg13g2_buf_1
X_458_ Inst_N_IO4_switch_matrix.SS4BEG8 SS4BEG[8] VPWR VGND sg13g2_buf_1
X_243_ FrameData[17] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_312_ FrameData[22] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_174_ Inst_N_IO4_ConfigMem.Inst_frame0_bit7.Q VPWR _074_ VGND _072_ _073_ sg13g2_o21ai_1
X_226_ FrameData[0] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit0.Q VPWR VGND
+ sg13g2_dlhq_1
X_088_ Inst_N_IO4_ConfigMem.Inst_frame3_bit12.Q N2MID[3] N4END[3] NN4END[3] NN4END[11]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit13.Q Inst_N_IO4_switch_matrix.S2BEG4 VPWR VGND
+ sg13g2_mux4_1
X_157_ VGND VPWR _003_ _054_ _058_ _057_ sg13g2_a21oi_1
XFILLER_6_153 VPWR VGND sg13g2_fill_2
X_209_ Inst_N_IO4_ConfigMem.Inst_frame2_bit9.Q N4END[11] A_O_top NN4END[11] C_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit8.Q Inst_N_IO4_switch_matrix.S4BEG2 VPWR VGND
+ sg13g2_mux4_1
XFILLER_4_421 VPWR VGND sg13g2_fill_2
XFILLER_1_287 VPWR VGND sg13g2_fill_1
X_190_ Inst_N_IO4_ConfigMem.Inst_frame1_bit14.Q N2END[1] N2END[3] N2END[5] Inst_D_IO_1_bidirectional_frame_config_pass.Q
+ Inst_N_IO4_ConfigMem.Inst_frame1_bit15.Q Inst_N_IO4_switch_matrix.SS4BEG5 VPWR VGND
+ sg13g2_mux4_1
X_457_ Inst_N_IO4_switch_matrix.SS4BEG7 SS4BEG[7] VPWR VGND sg13g2_buf_1
X_388_ FrameData[26] FrameData_O[26] VPWR VGND sg13g2_buf_1
X_242_ FrameData[16] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_173_ Inst_N_IO4_ConfigMem.Inst_frame0_bit6.Q VPWR _073_ VGND _068_ _069_ sg13g2_o21ai_1
X_311_ FrameData[21] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_10_194 VPWR VGND sg13g2_fill_2
XFILLER_8_59 VPWR VGND sg13g2_fill_1
X_156_ Inst_N_IO4_ConfigMem.Inst_frame0_bit13.Q VPWR _057_ VGND _055_ _056_ sg13g2_o21ai_1
X_225_ FrameData[31] FrameStrobe[4] Inst_N_IO4_ConfigMem.Inst_frame4_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_087_ Inst_N_IO4_ConfigMem.Inst_frame3_bit14.Q N2MID[2] N4END[2] NN4END[2] NN4END[10]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit15.Q Inst_N_IO4_switch_matrix.S2BEG5 VPWR VGND
+ sg13g2_mux4_1
X_208_ Inst_N_IO4_ConfigMem.Inst_frame2_bit11.Q N4END[10] B_O_top NN4END[10] D_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit10.Q Inst_N_IO4_switch_matrix.S4BEG3 VPWR VGND
+ sg13g2_mux4_1
X_139_ _041_ _040_ Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q VPWR VGND sg13g2_nand2b_1
XFILLER_4_411 VPWR VGND sg13g2_fill_2
X_387_ FrameData[25] FrameData_O[25] VPWR VGND sg13g2_buf_1
X_456_ Inst_N_IO4_switch_matrix.SS4BEG6 SS4BEG[6] VPWR VGND sg13g2_buf_1
X_310_ FrameData[20] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_10_343 VPWR VGND sg13g2_fill_2
X_172_ VGND VPWR _070_ _071_ _072_ Inst_N_IO4_ConfigMem.Inst_frame0_bit5.Q sg13g2_a21oi_1
X_241_ FrameData[15] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_439_ Inst_N_IO4_switch_matrix.S4BEG5 S4BEG[5] VPWR VGND sg13g2_buf_1
X_155_ Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q VPWR _056_ VGND N2END[6] Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q
+ sg13g2_o21ai_1
X_224_ FrameData[30] FrameStrobe[4] Inst_N_IO4_ConfigMem.Inst_frame4_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_3_328 VPWR VGND sg13g2_fill_2
XFILLER_6_100 VPWR VGND sg13g2_fill_1
X_086_ VPWR _003_ Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q VGND sg13g2_inv_1
XFILLER_6_155 VPWR VGND sg13g2_fill_1
XFILLER_2_350 VPWR VGND sg13g2_fill_1
X_207_ Inst_N_IO4_ConfigMem.Inst_frame2_bit12.Q N4END[7] NN4END[7] A_O_top C_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit13.Q Inst_N_IO4_switch_matrix.S4BEG4 VPWR VGND
+ sg13g2_mux4_1
X_138_ N2END[0] N2END[1] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q _040_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_8_206 VPWR VGND sg13g2_decap_4
XFILLER_4_423 VPWR VGND sg13g2_fill_1
XFILLER_6_71 VPWR VGND sg13g2_fill_1
X_386_ FrameData[24] FrameData_O[24] VPWR VGND sg13g2_buf_1
XFILLER_9_389 VPWR VGND sg13g2_fill_1
X_455_ Inst_N_IO4_switch_matrix.SS4BEG5 SS4BEG[5] VPWR VGND sg13g2_buf_1
X_171_ _071_ N2END[4] Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q VPWR VGND sg13g2_nand2b_1
X_240_ FrameData[14] FrameStrobe[3] Inst_N_IO4_ConfigMem.Inst_frame3_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_6_348 VPWR VGND sg13g2_fill_1
XFILLER_9_197 VPWR VGND sg13g2_fill_2
X_369_ FrameData[7] FrameData_O[7] VPWR VGND sg13g2_buf_1
X_438_ Inst_N_IO4_switch_matrix.S4BEG4 S4BEG[4] VPWR VGND sg13g2_buf_1
X_223_ FrameData[29] FrameStrobe[4] Inst_N_IO4_ConfigMem.Inst_frame4_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_085_ VPWR _002_ Inst_N_IO4_ConfigMem.Inst_frame0_bit21.Q VGND sg13g2_inv_1
X_154_ N2END[7] Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q _055_ VPWR VGND sg13g2_nor2b_1
XFILLER_2_192 VPWR VGND sg13g2_decap_4
X_206_ Inst_N_IO4_ConfigMem.Inst_frame2_bit14.Q N4END[6] NN4END[6] B_O_top D_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit15.Q Inst_N_IO4_switch_matrix.S4BEG5 VPWR VGND
+ sg13g2_mux4_1
X_137_ N2END[2] N2END[3] Inst_N_IO4_ConfigMem.Inst_frame0_bit18.Q _039_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_7_421 VPWR VGND sg13g2_fill_2
XFILLER_4_402 VPWR VGND sg13g2_fill_1
XFILLER_5_18 VPWR VGND sg13g2_fill_1
X_385_ FrameData[23] FrameData_O[23] VPWR VGND sg13g2_buf_1
X_454_ Inst_N_IO4_switch_matrix.SS4BEG4 SS4BEG[4] VPWR VGND sg13g2_buf_1
X_170_ _070_ N2END[5] Inst_N_IO4_ConfigMem.Inst_frame0_bit4.Q VPWR VGND sg13g2_nand2_1
X_368_ FrameData[6] FrameData_O[6] VPWR VGND sg13g2_buf_1
X_437_ Inst_N_IO4_switch_matrix.S4BEG3 S4BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_3_51 VPWR VGND sg13g2_fill_1
X_299_ FrameData[9] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit9.Q VPWR VGND
+ sg13g2_dlhq_1
XFILLER_10_153 VPWR VGND sg13g2_fill_2
X_084_ VPWR _001_ Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q VGND sg13g2_inv_1
X_153_ N2END[4] N2END[5] Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q _054_ VPWR VGND
+ sg13g2_mux2_1
X_222_ FrameData[28] FrameStrobe[4] Inst_N_IO4_ConfigMem.Inst_frame4_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_6_146 VPWR VGND sg13g2_decap_8
X_136_ _038_ VPWR D_I_top VGND _033_ _034_ sg13g2_o21ai_1
X_205_ Inst_N_IO4_ConfigMem.Inst_frame2_bit16.Q N4END[3] NN4END[3] A_O_top C_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit17.Q Inst_N_IO4_switch_matrix.S4BEG6 VPWR VGND
+ sg13g2_mux4_1
XFILLER_2_171 VPWR VGND sg13g2_decap_8
X_119_ _023_ _021_ _022_ VPWR VGND sg13g2_nand2b_1
XFILLER_4_277 VPWR VGND sg13g2_fill_2
X_384_ FrameData[22] FrameData_O[22] VPWR VGND sg13g2_buf_1
XFILLER_1_203 VPWR VGND sg13g2_fill_2
X_453_ Inst_N_IO4_switch_matrix.SS4BEG3 SS4BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_11_29 VPWR VGND sg13g2_fill_2
XFILLER_9_199 VPWR VGND sg13g2_fill_1
X_367_ FrameData[5] FrameData_O[5] VPWR VGND sg13g2_buf_1
X_436_ Inst_N_IO4_switch_matrix.S4BEG2 S4BEG[2] VPWR VGND sg13g2_buf_1
X_298_ FrameData[8] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit8.Q VPWR VGND
+ sg13g2_dlhq_1
X_083_ VPWR _000_ N2END[1] VGND sg13g2_inv_1
X_221_ Inst_N_IO4_ConfigMem.Inst_frame3_bit16.Q N2MID[1] N4END[1] NN4END[1] NN4END[9]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit17.Q Inst_N_IO4_switch_matrix.S2BEG6 VPWR VGND
+ sg13g2_mux4_1
XFILLER_5_0 VPWR VGND sg13g2_fill_1
X_152_ Inst_N_IO4_ConfigMem.Inst_frame0_bit12.Q N2END[0] N2END[2] N2END[1] N2END[3]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit11.Q _053_ VPWR VGND sg13g2_mux4_1
X_419_ Inst_N_IO4_switch_matrix.S2BEG1 S2BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_5_180 VPWR VGND sg13g2_decap_8
X_204_ Inst_N_IO4_ConfigMem.Inst_frame2_bit19.Q N4END[2] B_O_top NN4END[2] D_O_top
+ Inst_N_IO4_ConfigMem.Inst_frame2_bit18.Q Inst_N_IO4_switch_matrix.S4BEG7 VPWR VGND
+ sg13g2_mux4_1
X_135_ _038_ _037_ Inst_N_IO4_ConfigMem.Inst_frame0_bit28.Q VPWR VGND sg13g2_nand2b_1
XFILLER_7_412 VPWR VGND sg13g2_fill_1
XFILLER_7_423 VPWR VGND sg13g2_fill_1
X_118_ Inst_N_IO4_ConfigMem.Inst_frame0_bit31.Q VPWR _022_ VGND Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q
+ _019_ sg13g2_o21ai_1
XFILLER_7_264 VPWR VGND sg13g2_decap_4
XFILLER_4_234 VPWR VGND sg13g2_decap_4
X_383_ FrameData[21] FrameData_O[21] VPWR VGND sg13g2_buf_1
X_452_ Inst_N_IO4_switch_matrix.SS4BEG2 SS4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_9_112 VPWR VGND sg13g2_fill_2
X_297_ FrameData[7] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit7.Q VPWR VGND
+ sg13g2_dlhq_1
X_435_ Inst_N_IO4_switch_matrix.S4BEG1 S4BEG[1] VPWR VGND sg13g2_buf_1
X_366_ FrameData[4] FrameData_O[4] VPWR VGND sg13g2_buf_1
XFILLER_10_155 VPWR VGND sg13g2_fill_1
X_151_ _052_ _002_ _047_ C_I_top VPWR VGND sg13g2_a21o_1
X_220_ Inst_N_IO4_ConfigMem.Inst_frame3_bit18.Q N2MID[0] N4END[0] NN4END[0] NN4END[8]
+ Inst_N_IO4_ConfigMem.Inst_frame3_bit19.Q Inst_N_IO4_switch_matrix.S2BEG7 VPWR VGND
+ sg13g2_mux4_1
X_349_ FrameData[27] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_418_ Inst_N_IO4_switch_matrix.S2BEG0 S2BEG[0] VPWR VGND sg13g2_buf_1
X_134_ _035_ _036_ Inst_N_IO4_ConfigMem.Inst_frame0_bit27.Q _037_ VPWR VGND sg13g2_mux2_1
X_203_ Inst_N_IO4_ConfigMem.Inst_frame2_bit21.Q N4END[13] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ NN4END[13] Inst_C_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame2_bit20.Q
+ Inst_N_IO4_switch_matrix.S4BEG8 VPWR VGND sg13g2_mux4_1
Xclkbuf_0_UserCLK UserCLK clknet_0_UserCLK VPWR VGND sg13g2_buf_8
X_117_ Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q VPWR _021_ VGND N2END[6] Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_o21ai_1
XFILLER_1_238 VPWR VGND sg13g2_fill_1
X_382_ FrameData[20] FrameData_O[20] VPWR VGND sg13g2_buf_1
X_451_ Inst_N_IO4_switch_matrix.SS4BEG1 SS4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_10_315 VPWR VGND sg13g2_fill_1
X_296_ FrameData[6] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit6.Q VPWR VGND
+ sg13g2_dlhq_1
X_434_ Inst_N_IO4_switch_matrix.S4BEG0 S4BEG[0] VPWR VGND sg13g2_buf_1
X_365_ FrameData[3] FrameData_O[3] VPWR VGND sg13g2_buf_1
XFILLER_5_330 VPWR VGND sg13g2_fill_2
X_150_ Inst_N_IO4_ConfigMem.Inst_frame0_bit20.Q _049_ _051_ _048_ _050_ Inst_N_IO4_ConfigMem.Inst_frame0_bit19.Q
+ _052_ VPWR VGND sg13g2_mux4_1
X_348_ FrameData[26] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_279_ FrameData[21] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_417_ Inst_N_IO4_switch_matrix.S1BEG3 S1BEG[3] VPWR VGND sg13g2_buf_1
XFILLER_11_421 VPWR VGND sg13g2_fill_2
XFILLER_2_185 VPWR VGND sg13g2_decap_8
X_202_ Inst_N_IO4_ConfigMem.Inst_frame2_bit23.Q N4END[12] Inst_B_IO_1_bidirectional_frame_config_pass.Q
+ NN4END[12] Inst_D_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame2_bit22.Q
+ Inst_N_IO4_switch_matrix.S4BEG9 VPWR VGND sg13g2_mux4_1
X_133_ Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q N2MID[4] N2MID[5] N2MID[6] N2MID[7]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q _036_ VPWR VGND sg13g2_mux4_1
X_116_ Inst_N_IO4_ConfigMem.Inst_frame0_bit29.Q N2MID[6] N2MID[7] N2END[0] N2END[4]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q _020_ VPWR VGND sg13g2_mux4_1
XFILLER_7_200 VPWR VGND sg13g2_decap_8
X_381_ FrameData[19] FrameData_O[19] VPWR VGND sg13g2_buf_1
X_450_ Inst_N_IO4_switch_matrix.SS4BEG0 SS4BEG[0] VPWR VGND sg13g2_buf_1
X_433_ Inst_N_IO4_switch_matrix.S2BEGb7 S2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_9_158 VPWR VGND sg13g2_fill_1
X_295_ FrameData[5] FrameStrobe[1] Inst_N_IO4_ConfigMem.Inst_frame1_bit5.Q VPWR VGND
+ sg13g2_dlhq_1
X_364_ FrameData[2] FrameData_O[2] VPWR VGND sg13g2_buf_1
X_347_ FrameData[25] FrameStrobe[0] Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_278_ FrameData[20] FrameStrobe[2] Inst_N_IO4_ConfigMem.Inst_frame2_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_416_ Inst_N_IO4_switch_matrix.S1BEG2 S1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_6_139 VPWR VGND sg13g2_decap_8
XFILLER_5_194 VPWR VGND sg13g2_decap_4
X_201_ Inst_N_IO4_ConfigMem.Inst_frame2_bit24.Q N4END[9] NN4END[9] Inst_A_IO_1_bidirectional_frame_config_pass.Q
+ Inst_C_IO_1_bidirectional_frame_config_pass.Q Inst_N_IO4_ConfigMem.Inst_frame2_bit25.Q
+ Inst_N_IO4_switch_matrix.S4BEG10 VPWR VGND sg13g2_mux4_1
X_132_ Inst_N_IO4_ConfigMem.Inst_frame0_bit25.Q N2MID[0] N2MID[1] N2MID[2] N2MID[3]
+ Inst_N_IO4_ConfigMem.Inst_frame0_bit26.Q _035_ VPWR VGND sg13g2_mux4_1
XFILLER_2_164 VPWR VGND sg13g2_decap_8
XFILLER_9_65 VPWR VGND sg13g2_fill_2
XFILLER_0_23 VPWR VGND sg13g2_fill_1
X_115_ _019_ N2END[5] Inst_N_IO4_ConfigMem.Inst_frame0_bit30.Q VPWR VGND sg13g2_nand2b_1
XFILLER_7_245 VPWR VGND sg13g2_fill_2
XFILLER_0_421 VPWR VGND sg13g2_fill_2
X_380_ FrameData[18] FrameData_O[18] VPWR VGND sg13g2_buf_1
.ends

