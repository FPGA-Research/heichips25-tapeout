* NGSPICE file created from LUT4AB.ext - technology: ihp-sg13g2

* Black-box entry subcircuit for sg13g2_nand2_1 abstract view
.subckt sg13g2_nand2_1 Y A B VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_o21ai_1 abstract view
.subckt sg13g2_o21ai_1 B1 VDD Y VSS A1 A2
.ends

* Black-box entry subcircuit for sg13g2_buf_1 abstract view
.subckt sg13g2_buf_1 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dlhq_1 abstract view
.subckt sg13g2_dlhq_1 D GATE Q VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_2 abstract view
.subckt sg13g2_fill_2 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_fill_1 abstract view
.subckt sg13g2_fill_1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux4_1 abstract view
.subckt sg13g2_mux4_1 S0 A0 A1 A2 A3 S1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_mux2_1 abstract view
.subckt sg13g2_mux2_1 A0 A1 S X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand2b_1 abstract view
.subckt sg13g2_nand2b_1 Y B A_N VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a21oi_1 abstract view
.subckt sg13g2_a21oi_1 VSS VDD A1 A2 Y B1
.ends

* Black-box entry subcircuit for sg13g2_nor2_1 abstract view
.subckt sg13g2_nor2_1 A B Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_inv_1 abstract view
.subckt sg13g2_inv_1 VDD Y A VSS
.ends

* Black-box entry subcircuit for sg13g2_or2_1 abstract view
.subckt sg13g2_or2_1 VSS VDD X B A
.ends

* Black-box entry subcircuit for sg13g2_nor2b_1 abstract view
.subckt sg13g2_nor2b_1 A B_N Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_antennanp abstract view
.subckt sg13g2_antennanp VDD VSS A
.ends

* Black-box entry subcircuit for sg13g2_a21o_1 abstract view
.subckt sg13g2_a21o_1 A2 A1 B1 X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a22oi_1 abstract view
.subckt sg13g2_a22oi_1 Y B1 B2 A2 A1 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_a221oi_1 abstract view
.subckt sg13g2_a221oi_1 VDD VSS B2 C1 B1 A1 Y A2
.ends

* Black-box entry subcircuit for sg13g2_nand3_1 abstract view
.subckt sg13g2_nand3_1 B C A Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or3_1 abstract view
.subckt sg13g2_or3_1 A B C X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_tiehi abstract view
.subckt sg13g2_tiehi VDD VSS L_HI
.ends

* Black-box entry subcircuit for sg13g2_and2_1 abstract view
.subckt sg13g2_and2_1 A B X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_dfrbpq_1 abstract view
.subckt sg13g2_dfrbpq_1 RESET_B VSS VDD D Q CLK
.ends

* Black-box entry subcircuit for sg13g2_nor3_1 abstract view
.subckt sg13g2_nor3_1 A B C Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_or4_1 abstract view
.subckt sg13g2_or4_1 A B C D X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_buf_8 abstract view
.subckt sg13g2_buf_8 A X VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_4 abstract view
.subckt sg13g2_decap_4 VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nand3b_1 abstract view
.subckt sg13g2_nand3b_1 B C Y VDD VSS A_N
.ends

* Black-box entry subcircuit for sg13g2_and3_1 abstract view
.subckt sg13g2_and3_1 X A B C VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_nor4_1 abstract view
.subckt sg13g2_nor4_1 A B C D Y VDD VSS
.ends

* Black-box entry subcircuit for sg13g2_decap_8 abstract view
.subckt sg13g2_decap_8 VDD VSS
.ends

.subckt LUT4AB Ci Co E1BEG[0] E1BEG[1] E1BEG[2] E1BEG[3] E1END[0] E1END[1] E1END[2]
+ E1END[3] E2BEG[0] E2BEG[1] E2BEG[2] E2BEG[3] E2BEG[4] E2BEG[5] E2BEG[6] E2BEG[7]
+ E2BEGb[0] E2BEGb[1] E2BEGb[2] E2BEGb[3] E2BEGb[4] E2BEGb[5] E2BEGb[6] E2BEGb[7]
+ E2END[0] E2END[1] E2END[2] E2END[3] E2END[4] E2END[5] E2END[6] E2END[7] E2MID[0]
+ E2MID[1] E2MID[2] E2MID[3] E2MID[4] E2MID[5] E2MID[6] E2MID[7] E6BEG[0] E6BEG[10]
+ E6BEG[11] E6BEG[1] E6BEG[2] E6BEG[3] E6BEG[4] E6BEG[5] E6BEG[6] E6BEG[7] E6BEG[8]
+ E6BEG[9] E6END[0] E6END[10] E6END[11] E6END[1] E6END[2] E6END[3] E6END[4] E6END[5]
+ E6END[6] E6END[7] E6END[8] E6END[9] EE4BEG[0] EE4BEG[10] EE4BEG[11] EE4BEG[12] EE4BEG[13]
+ EE4BEG[14] EE4BEG[15] EE4BEG[1] EE4BEG[2] EE4BEG[3] EE4BEG[4] EE4BEG[5] EE4BEG[6]
+ EE4BEG[7] EE4BEG[8] EE4BEG[9] EE4END[0] EE4END[10] EE4END[11] EE4END[12] EE4END[13]
+ EE4END[14] EE4END[15] EE4END[1] EE4END[2] EE4END[3] EE4END[4] EE4END[5] EE4END[6]
+ EE4END[7] EE4END[8] EE4END[9] FrameData[0] FrameData[10] FrameData[11] FrameData[12]
+ FrameData[13] FrameData[14] FrameData[15] FrameData[16] FrameData[17] FrameData[18]
+ FrameData[19] FrameData[1] FrameData[20] FrameData[21] FrameData[22] FrameData[23]
+ FrameData[24] FrameData[25] FrameData[26] FrameData[27] FrameData[28] FrameData[29]
+ FrameData[2] FrameData[30] FrameData[31] FrameData[3] FrameData[4] FrameData[5]
+ FrameData[6] FrameData[7] FrameData[8] FrameData[9] FrameData_O[0] FrameData_O[10]
+ FrameData_O[11] FrameData_O[12] FrameData_O[13] FrameData_O[14] FrameData_O[15]
+ FrameData_O[16] FrameData_O[17] FrameData_O[18] FrameData_O[19] FrameData_O[1] FrameData_O[20]
+ FrameData_O[21] FrameData_O[22] FrameData_O[23] FrameData_O[24] FrameData_O[25]
+ FrameData_O[26] FrameData_O[27] FrameData_O[28] FrameData_O[29] FrameData_O[2] FrameData_O[30]
+ FrameData_O[31] FrameData_O[3] FrameData_O[4] FrameData_O[5] FrameData_O[6] FrameData_O[7]
+ FrameData_O[8] FrameData_O[9] FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N1END[0] N1END[1] N1END[2] N1END[3] N2BEG[0] N2BEG[1] N2BEG[2]
+ N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6] N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3]
+ N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7] N2END[0] N2END[1] N2END[2] N2END[3] N2END[4]
+ N2END[5] N2END[6] N2END[7] N2MID[0] N2MID[1] N2MID[2] N2MID[3] N2MID[4] N2MID[5]
+ N2MID[6] N2MID[7] N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15]
+ N4BEG[1] N4BEG[2] N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9]
+ N4END[0] N4END[10] N4END[11] N4END[12] N4END[13] N4END[14] N4END[15] N4END[1] N4END[2]
+ N4END[3] N4END[4] N4END[5] N4END[6] N4END[7] N4END[8] N4END[9] NN4BEG[0] NN4BEG[10]
+ NN4BEG[11] NN4BEG[12] NN4BEG[13] NN4BEG[14] NN4BEG[15] NN4BEG[1] NN4BEG[2] NN4BEG[3]
+ NN4BEG[4] NN4BEG[5] NN4BEG[6] NN4BEG[7] NN4BEG[8] NN4BEG[9] NN4END[0] NN4END[10]
+ NN4END[11] NN4END[12] NN4END[13] NN4END[14] NN4END[15] NN4END[1] NN4END[2] NN4END[3]
+ NN4END[4] NN4END[5] NN4END[6] NN4END[7] NN4END[8] NN4END[9] S1BEG[0] S1BEG[1] S1BEG[2]
+ S1BEG[3] S1END[0] S1END[1] S1END[2] S1END[3] S2BEG[0] S2BEG[1] S2BEG[2] S2BEG[3]
+ S2BEG[4] S2BEG[5] S2BEG[6] S2BEG[7] S2BEGb[0] S2BEGb[1] S2BEGb[2] S2BEGb[3] S2BEGb[4]
+ S2BEGb[5] S2BEGb[6] S2BEGb[7] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5]
+ S2END[6] S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6]
+ S2MID[7] S4BEG[0] S4BEG[10] S4BEG[11] S4BEG[12] S4BEG[13] S4BEG[14] S4BEG[15] S4BEG[1]
+ S4BEG[2] S4BEG[3] S4BEG[4] S4BEG[5] S4BEG[6] S4BEG[7] S4BEG[8] S4BEG[9] S4END[0]
+ S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2] S4END[3]
+ S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] SS4BEG[0] SS4BEG[10] SS4BEG[11]
+ SS4BEG[12] SS4BEG[13] SS4BEG[14] SS4BEG[15] SS4BEG[1] SS4BEG[2] SS4BEG[3] SS4BEG[4]
+ SS4BEG[5] SS4BEG[6] SS4BEG[7] SS4BEG[8] SS4BEG[9] SS4END[0] SS4END[10] SS4END[11]
+ SS4END[12] SS4END[13] SS4END[14] SS4END[15] SS4END[1] SS4END[2] SS4END[3] SS4END[4]
+ SS4END[5] SS4END[6] SS4END[7] SS4END[8] SS4END[9] UserCLK UserCLKo VGND VPWR W1BEG[0]
+ W1BEG[1] W1BEG[2] W1BEG[3] W1END[0] W1END[1] W1END[2] W1END[3] W2BEG[0] W2BEG[1]
+ W2BEG[2] W2BEG[3] W2BEG[4] W2BEG[5] W2BEG[6] W2BEG[7] W2BEGb[0] W2BEGb[1] W2BEGb[2]
+ W2BEGb[3] W2BEGb[4] W2BEGb[5] W2BEGb[6] W2BEGb[7] W2END[0] W2END[1] W2END[2] W2END[3]
+ W2END[4] W2END[5] W2END[6] W2END[7] W2MID[0] W2MID[1] W2MID[2] W2MID[3] W2MID[4]
+ W2MID[5] W2MID[6] W2MID[7] W6BEG[0] W6BEG[10] W6BEG[11] W6BEG[1] W6BEG[2] W6BEG[3]
+ W6BEG[4] W6BEG[5] W6BEG[6] W6BEG[7] W6BEG[8] W6BEG[9] W6END[0] W6END[10] W6END[11]
+ W6END[1] W6END[2] W6END[3] W6END[4] W6END[5] W6END[6] W6END[7] W6END[8] W6END[9]
+ WW4BEG[0] WW4BEG[10] WW4BEG[11] WW4BEG[12] WW4BEG[13] WW4BEG[14] WW4BEG[15] WW4BEG[1]
+ WW4BEG[2] WW4BEG[3] WW4BEG[4] WW4BEG[5] WW4BEG[6] WW4BEG[7] WW4BEG[8] WW4BEG[9]
+ WW4END[0] WW4END[10] WW4END[11] WW4END[12] WW4END[13] WW4END[14] WW4END[15] WW4END[1]
+ WW4END[2] WW4END[3] WW4END[4] WW4END[5] WW4END[6] WW4END[7] WW4END[8] WW4END[9]
X_2106_ _0754_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0670_ VPWR VGND sg13g2_nand2_1
X_2037_ _0689_ VPWR _0690_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q _0230_ sg13g2_o21ai_1
X_3086_ Inst_LUT4AB_switch_matrix.E6BEG1 E6BEG[11] VPWR VGND sg13g2_buf_1
X_3155_ Inst_LUT4AB_switch_matrix.N1BEG0 N1BEG[0] VPWR VGND sg13g2_buf_1
X_2939_ FrameData[28] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_321 VPWR VGND sg13g2_fill_2
XFILLER_13_144 VPWR VGND sg13g2_fill_1
X_1270_ _1107_ VPWR _1108_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _1106_ sg13g2_o21ai_1
X_2655_ FrameData[0] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_2724_ FrameData[5] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1606_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q _1021_ _1026_ _1034_ _0275_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q
+ _0276_ VPWR VGND sg13g2_mux4_1
X_1468_ S1END[1] S1END[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q _0143_ VPWR VGND
+ sg13g2_mux2_1
X_3207_ Inst_LUT4AB_switch_matrix.S1BEG0 S1BEG[0] VPWR VGND sg13g2_buf_1
X_2586_ FrameData[27] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_1399_ _0076_ _0075_ _0074_ VPWR VGND sg13g2_nand2b_1
X_1537_ _0201_ VPWR _0209_ VGND _0200_ _0208_ sg13g2_o21ai_1
X_3138_ FrameStrobe[3] FrameStrobe_O[3] VPWR VGND sg13g2_buf_1
X_3069_ E2MID[2] E2BEGb[2] VPWR VGND sg13g2_buf_1
XFILLER_37_62 VPWR VGND sg13g2_fill_1
X_2440_ FrameData[9] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_dlhq_1
X_1253_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q _1090_ _1092_ _1091_ sg13g2_a21oi_1
X_2371_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0453_ _0968_ VPWR VGND sg13g2_nor2_1
X_1322_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q N2MID[4] E2MID[4] W2MID[4] Inst_LUT4AB_switch_matrix.JS2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q _1157_ VPWR VGND sg13g2_mux4_1
X_1184_ VPWR _1025_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VGND sg13g2_inv_1
XFILLER_20_423 VPWR VGND sg13g2_fill_1
X_2569_ FrameData[10] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_2638_ FrameData[15] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_2707_ FrameData[20] FrameStrobe[10] Inst_LUT4AB_switch_matrix.DEBUG_select_LB_SR[0]
+ VPWR VGND sg13g2_dlhq_1
XFILLER_15_217 VPWR VGND sg13g2_fill_1
XFILLER_48_83 VPWR VGND sg13g2_fill_1
X_1940_ VGND VPWR _0598_ _0597_ _0595_ sg13g2_or2_1
X_1871_ VGND VPWR _0479_ _0490_ _0531_ _0488_ sg13g2_a21oi_1
XFILLER_14_250 VPWR VGND sg13g2_fill_2
X_2423_ FrameData[24] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VPWR VGND sg13g2_dlhq_1
X_2285_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q _0912_ _0913_ _0914_ _0915_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q
+ Inst_LUT4AB_switch_matrix.E6BEG0 VPWR VGND sg13g2_mux4_1
X_1236_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q N1END[2] N2END[4] N4END[0] E2END[4]
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _1076_ VPWR VGND sg13g2_mux4_1
X_2354_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q F _0237_ Inst_LUT4AB_switch_matrix.E2BEG0
+ _0248_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q Inst_LUT4AB_switch_matrix.S1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1305_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q N2END[4] S2END[4] EE4END[0] W2END[4]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q _1141_ VPWR VGND sg13g2_mux4_1
XFILLER_4_419 VPWR VGND sg13g2_fill_1
XFILLER_28_397 VPWR VGND sg13g2_fill_1
X_2070_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VPWR _0721_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ _0718_ sg13g2_o21ai_1
XFILLER_34_334 VPWR VGND sg13g2_fill_1
X_2972_ FrameData[29] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1923_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VPWR _0582_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ _0581_ sg13g2_o21ai_1
X_1854_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q _0514_ _0515_ VPWR VGND sg13g2_nor2_1
X_1785_ Inst_LUT4AB_switch_matrix.JW2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q
+ _0448_ VPWR VGND sg13g2_nor2b_1
X_2406_ _0999_ Inst_LUT4AB_switch_matrix.DEBUG_select_LD_SR[0] _0985_ VPWR VGND sg13g2_nand2_1
X_2337_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q G _0960_ VPWR VGND sg13g2_nor2b_1
X_2268_ _0898_ _0900_ Inst_LUT4AB_switch_matrix.SS4BEG0 VPWR VGND sg13g2_nor2_1
X_1219_ _1060_ _1059_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q VPWR VGND sg13g2_nand2b_1
XFILLER_25_301 VPWR VGND sg13g2_fill_2
X_2199_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0838_ _0841_ _0840_ sg13g2_a21oi_1
XFILLER_52_164 VPWR VGND sg13g2_fill_1
X_1570_ _0241_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q _0237_ VPWR VGND sg13g2_nand2_1
XANTENNA_5 VPWR VGND EE4END[5] sg13g2_antennanp
X_3240_ Inst_LUT4AB_switch_matrix.S4BEG1 S4BEG[13] VPWR VGND sg13g2_buf_1
X_3171_ N2MID[4] N2BEGb[4] VPWR VGND sg13g2_buf_1
X_2122_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VPWR _0768_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ _0765_ sg13g2_o21ai_1
X_2053_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q N1END[0] N2END[0] E1END[0] E2END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q _0705_ VPWR VGND sg13g2_mux4_1
X_2955_ FrameData[12] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1837_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q Inst_LUT4AB_switch_matrix.M_AH
+ _0498_ _0497_ sg13g2_a21oi_1
X_1906_ _0564_ VPWR _0565_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q _0562_ sg13g2_o21ai_1
X_1768_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q _0425_ _0432_ _0431_
+ sg13g2_a21oi_1
X_2886_ FrameData[7] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1699_ VGND VPWR _0365_ _0364_ _0362_ sg13g2_or2_1
XFILLER_48_234 VPWR VGND sg13g2_fill_2
XFILLER_16_120 VPWR VGND sg13g2_fill_1
X_1622_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q E G H Inst_LUT4AB_switch_matrix.M_AB
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q _0292_ VPWR VGND sg13g2_mux4_1
X_2740_ FrameData[21] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_2671_ FrameData[16] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_1553_ _0224_ VPWR _0225_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q W1END[0]
+ sg13g2_o21ai_1
X_3223_ S2MID[4] S2BEGb[4] VPWR VGND sg13g2_buf_1
X_1484_ _0157_ VPWR _0158_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q H sg13g2_o21ai_1
X_2105_ _0752_ _0693_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0753_ VPWR VGND
+ sg13g2_mux2_1
X_3085_ Inst_LUT4AB_switch_matrix.E6BEG0 E6BEG[10] VPWR VGND sg13g2_buf_1
X_2036_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q Inst_LUT4AB_switch_matrix.E2BEG5
+ _0689_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q sg13g2_a21oi_1
X_3154_ FrameStrobe[19] FrameStrobe_O[19] VPWR VGND sg13g2_buf_1
X_2938_ FrameData[27] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_2869_ FrameData[22] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_7_8 VPWR VGND sg13g2_fill_2
XFILLER_5_399 VPWR VGND sg13g2_fill_2
X_2723_ FrameData[4] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_2654_ FrameData[31] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1605_ VPWR Inst_LUT4AB_switch_matrix.JS2BEG5 _0275_ VGND sg13g2_inv_1
X_2585_ FrameData[26] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_1536_ VGND VPWR _0204_ _0207_ _0208_ _0206_ sg13g2_a21oi_1
X_3206_ Inst_LUT4AB_switch_matrix.NN4BEG3 NN4BEG[15] VPWR VGND sg13g2_buf_1
X_1467_ _0141_ VPWR _0142_ VGND S2END[5] Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q
+ sg13g2_o21ai_1
X_3137_ FrameStrobe[2] FrameStrobe_O[2] VPWR VGND sg13g2_buf_1
X_1398_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q _1157_ _1159_ _1141_ _1140_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q
+ _0075_ VPWR VGND sg13g2_mux4_1
X_2019_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q _0391_ _0673_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q
+ sg13g2_a21oi_1
X_3068_ E2MID[1] E2BEGb[1] VPWR VGND sg13g2_buf_1
X_2370_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0048_ _0967_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q
+ sg13g2_a21oi_1
X_1321_ _1156_ _1153_ _1148_ Inst_LUT4AB_switch_matrix.JS2BEG3 VPWR VGND sg13g2_a21o_1
XFILLER_1_380 VPWR VGND sg13g2_fill_1
X_1252_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VPWR _1091_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ _1088_ sg13g2_o21ai_1
X_1183_ VPWR _1024_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q VGND sg13g2_inv_1
X_2706_ FrameData[19] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_2568_ FrameData[9] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_1519_ Inst_LUT4AB_switch_matrix.JS2BEG4 _0191_ _1035_ _0182_ _0176_ VPWR VGND sg13g2_a22oi_1
X_2499_ FrameData[4] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VPWR VGND sg13g2_dlhq_1
X_2637_ FrameData[14] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_1870_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q _0520_ _0525_ _0529_ _0527_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q
+ _0530_ VPWR VGND sg13g2_mux4_1
X_2422_ _1008_ VPWR _0007_ VGND _1010_ _1011_ sg13g2_o21ai_1
XFILLER_36_2 VPWR VGND sg13g2_fill_1
X_2353_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit15.Q G Inst_LUT4AB_switch_matrix.E2BEG1
+ _0586_ _0623_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit14.Q Inst_LUT4AB_switch_matrix.S1BEG2
+ VPWR VGND sg13g2_mux4_1
X_2284_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q _1084_ _0148_ _0308_ _0586_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0915_ VPWR VGND sg13g2_mux4_1
X_1235_ VPWR VGND _1074_ _1019_ _1072_ _1068_ _1075_ _1070_ sg13g2_a221oi_1
X_1304_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q N4END[1] E6END[1] W6END[1] Inst_LUT4AB_switch_matrix.JS2BEG1
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q _1140_ VPWR VGND sg13g2_mux4_1
XFILLER_37_387 VPWR VGND sg13g2_fill_2
XFILLER_20_210 VPWR VGND sg13g2_fill_1
X_1999_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q _0617_ _0622_ _0626_ _0624_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q
+ _0655_ VPWR VGND sg13g2_mux4_1
XFILLER_47_107 VPWR VGND sg13g2_fill_2
X_1922_ S1END[1] S1END[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q _0581_ VPWR VGND
+ sg13g2_mux2_1
X_2971_ FrameData[28] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_1853_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q _0511_ _0514_ _0513_ sg13g2_a21oi_1
X_1784_ _0440_ _0447_ Inst_LUT4AB_switch_matrix.JW2BEG4 VPWR VGND sg13g2_nor2_1
XFILLER_41_0 VPWR VGND sg13g2_fill_1
X_2336_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q _0589_ _0959_ _0958_ sg13g2_a21oi_1
X_2405_ _0998_ Inst_LUT4AB_switch_matrix.DEBUG_select_LD_EN[0] _0973_ VPWR VGND sg13g2_nand2b_1
X_1218_ E6END[0] S2END[2] Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q _1059_ VPWR VGND
+ sg13g2_mux2_1
X_2267_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q _0899_ _0900_ VPWR VGND sg13g2_nor2_1
X_2198_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q VPWR _0840_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q
+ _0839_ sg13g2_o21ai_1
XANTENNA_6 VPWR VGND EE4END[6] sg13g2_antennanp
X_3170_ N2MID[3] N2BEGb[3] VPWR VGND sg13g2_buf_1
X_2121_ _0766_ VPWR _0767_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q _1052_ sg13g2_o21ai_1
X_2052_ VGND VPWR _1045_ _0702_ _0704_ _0703_ sg13g2_a21oi_1
X_2954_ FrameData[11] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1905_ _0537_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q _0563_ _0564_ VPWR VGND sg13g2_a21o_1
X_2885_ FrameData[6] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_30_360 VPWR VGND sg13g2_fill_1
X_1836_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q VPWR _0497_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q
+ _1052_ sg13g2_o21ai_1
X_1767_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q VPWR _0431_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q
+ _0430_ sg13g2_o21ai_1
X_1698_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q Inst_LUT4AB_switch_matrix.JN2BEG2
+ _0364_ _0363_ sg13g2_a21oi_1
X_2319_ _0944_ VPWR _0945_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _0556_
+ sg13g2_o21ai_1
X_3299_ WW4END[11] WW4BEG[7] VPWR VGND sg13g2_buf_1
X_1621_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ _0291_ VPWR VGND sg13g2_mux4_1
X_1552_ _0224_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q W1END[2] VPWR VGND sg13g2_nand2b_1
X_2670_ FrameData[15] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_3222_ S2MID[3] S2BEGb[3] VPWR VGND sg13g2_buf_1
X_1483_ _0157_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q Inst_LUT4AB_switch_matrix.M_AB
+ VPWR VGND sg13g2_nand2b_1
X_2104_ _0751_ VPWR _0752_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q _0748_ sg13g2_o21ai_1
X_3153_ FrameStrobe[18] FrameStrobe_O[18] VPWR VGND sg13g2_buf_1
X_2035_ _0688_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop Inst_LD_LUT4c_frame_config_dffesr.c_out_mux
+ D VPWR VGND sg13g2_mux2_1
X_3084_ E6END[11] E6BEG[9] VPWR VGND sg13g2_buf_1
X_2868_ FrameData[21] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_2937_ FrameData[26] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_1819_ _0481_ _0480_ _0476_ _0479_ Inst_LF_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_a22oi_1
X_2799_ FrameData[16] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_345 VPWR VGND sg13g2_fill_2
XFILLER_32_422 VPWR VGND sg13g2_fill_2
X_2722_ FrameData[3] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1604_ _0274_ VPWR _0275_ VGND _0257_ _0263_ sg13g2_o21ai_1
X_2653_ FrameData[30] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1535_ _0089_ _0083_ _0080_ _0207_ VPWR VGND sg13g2_a21o_1
X_2584_ FrameData[25] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_3205_ Inst_LUT4AB_switch_matrix.NN4BEG2 NN4BEG[14] VPWR VGND sg13g2_buf_1
X_1466_ _0141_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q W1END[1] VPWR VGND sg13g2_nand2b_1
X_3136_ FrameStrobe[1] FrameStrobe_O[1] VPWR VGND sg13g2_buf_1
X_1397_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q _1083_ _1084_ _1066_ _1065_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q
+ _0074_ VPWR VGND sg13g2_mux4_1
X_3067_ E2MID[0] E2BEGb[0] VPWR VGND sg13g2_buf_1
X_2018_ _0365_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q _0671_ _0672_ VPWR VGND sg13g2_a21o_1
XFILLER_37_20 VPWR VGND sg13g2_fill_1
X_1320_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q _1155_ _1156_ VPWR VGND sg13g2_nor2_1
XFILLER_49_330 VPWR VGND sg13g2_fill_2
X_1182_ VPWR _1023_ WW4END[2] VGND sg13g2_inv_1
X_1251_ _1089_ VPWR _1090_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q H sg13g2_o21ai_1
X_2705_ FrameData[18] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_2636_ FrameData[13] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_2567_ FrameData[8] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_1518_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0190_ _0188_ _0184_ _0186_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q
+ _0191_ VPWR VGND sg13g2_mux4_1
X_2498_ FrameData[3] FrameStrobe[16] Inst_LD_LUT4c_frame_config_dffesr.c_reset_value
+ VPWR VGND sg13g2_dlhq_1
X_1449_ E6END[1] S2END[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q _0125_ VPWR VGND
+ sg13g2_mux2_1
X_3119_ FrameData[16] FrameData_O[16] VPWR VGND sg13g2_buf_1
XFILLER_23_241 VPWR VGND sg13g2_fill_2
XFILLER_23_285 VPWR VGND sg13g2_fill_1
XFILLER_14_252 VPWR VGND sg13g2_fill_1
X_2421_ _1007_ VPWR _1011_ VGND Inst_LG_LUT4c_frame_config_dffesr.c_reset_value _1009_
+ sg13g2_o21ai_1
X_2283_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q G H Inst_LUT4AB_switch_matrix.M_AB
+ Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q _0914_
+ VPWR VGND sg13g2_mux4_1
X_2352_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q H _1159_ Inst_LUT4AB_switch_matrix.E2BEG2
+ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q Inst_LUT4AB_switch_matrix.S1BEG3
+ VPWR VGND sg13g2_mux4_1
X_1303_ _1132_ _1129_ _1139_ Inst_LUT4AB_switch_matrix.JS2BEG1 VPWR VGND sg13g2_a21o_1
XFILLER_49_182 VPWR VGND sg13g2_fill_1
X_1234_ VGND VPWR _1017_ _1073_ _1074_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q sg13g2_a21oi_1
X_1998_ _0645_ _0640_ _0653_ _0654_ VPWR VGND sg13g2_a21o_1
X_2619_ FrameData[28] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_7_226 VPWR VGND sg13g2_fill_1
XFILLER_11_211 VPWR VGND sg13g2_fill_1
XFILLER_11_255 VPWR VGND sg13g2_fill_2
X_1921_ _0579_ VPWR _0580_ VGND S2END[7] Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
+ sg13g2_o21ai_1
X_1852_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VPWR _0513_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ _0512_ sg13g2_o21ai_1
X_2970_ FrameData[27] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_1783_ VPWR VGND _0446_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q _0445_ _1039_ _0447_
+ _0441_ sg13g2_a221oi_1
X_2335_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q VPWR _0958_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ _0148_ sg13g2_o21ai_1
XFILLER_34_0 VPWR VGND sg13g2_fill_2
X_2266_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q N1END[2] W1END[2] E1END[2] F Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q
+ _0899_ VPWR VGND sg13g2_mux4_1
X_2404_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop _0997_ _0995_ _0003_ VPWR VGND
+ sg13g2_mux2_1
X_1217_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q _1057_ _1058_ VPWR VGND sg13g2_nor2_1
X_2197_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q G H Inst_LUT4AB_switch_matrix.M_AD
+ Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q _0839_
+ VPWR VGND sg13g2_mux4_1
XFILLER_45_20 VPWR VGND sg13g2_fill_2
XFILLER_31_339 VPWR VGND sg13g2_fill_1
XANTENNA_7 VPWR VGND EE4END[7] sg13g2_antennanp
X_2120_ _0766_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q Inst_LUT4AB_switch_matrix.M_AD
+ VPWR VGND sg13g2_nand2_1
X_2051_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VPWR _0703_ VGND _0699_ _0701_ sg13g2_o21ai_1
XFILLER_19_141 VPWR VGND sg13g2_fill_1
X_1835_ _0496_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop Inst_LF_LUT4c_frame_config_dffesr.c_out_mux
+ F VPWR VGND sg13g2_mux2_1
X_2953_ FrameData[10] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1904_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q VPWR _0563_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q
+ _0538_ sg13g2_o21ai_1
X_2884_ FrameData[5] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1766_ _0429_ VPWR _0430_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q _0426_ sg13g2_o21ai_1
X_1697_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q VPWR _0363_ VGND _1023_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q
+ sg13g2_o21ai_1
X_2318_ _0944_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _1066_ VPWR VGND sg13g2_nand2_1
X_2249_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q N1END[0] W1END[0] E1END[0] B Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ _0884_ VPWR VGND sg13g2_mux4_1
X_3298_ WW4END[10] WW4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_25_155 VPWR VGND sg13g2_fill_2
XFILLER_31_22 VPWR VGND sg13g2_fill_1
XFILLER_48_236 VPWR VGND sg13g2_fill_1
X_1551_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q _0222_ _0223_ VPWR VGND sg13g2_nor2b_1
X_1620_ VGND VPWR _1041_ _0289_ _0290_ _0288_ sg13g2_a21oi_1
X_1482_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q _1051_ _0156_ _0155_ sg13g2_a21oi_1
X_3152_ FrameStrobe[17] FrameStrobe_O[17] VPWR VGND sg13g2_buf_1
X_3221_ S2MID[2] S2BEGb[2] VPWR VGND sg13g2_buf_1
X_2103_ _0749_ _0750_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q _0751_ VPWR VGND sg13g2_nand3_1
X_3083_ E6END[10] E6BEG[8] VPWR VGND sg13g2_buf_1
X_2034_ _0687_ _0684_ _0682_ _0688_ VPWR VGND sg13g2_a21o_1
X_1818_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q _0478_ _0480_ Inst_LF_LUT4c_frame_config_dffesr.c_I0mux
+ sg13g2_a21oi_1
X_2867_ FrameData[20] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_2936_ FrameData[25] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_2798_ FrameData[15] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_1749_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR _0414_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ _0411_ sg13g2_o21ai_1
XFILLER_45_206 VPWR VGND sg13g2_fill_2
XFILLER_32_412 VPWR VGND sg13g2_fill_2
X_2652_ FrameData[29] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_2721_ FrameData[2] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_3204_ Inst_LUT4AB_switch_matrix.NN4BEG1 NN4BEG[13] VPWR VGND sg13g2_buf_1
X_1465_ _0140_ _0139_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR VGND sg13g2_nand2b_1
X_1603_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q _0268_ _0273_ _0274_ VPWR VGND sg13g2_or3_1
X_2583_ FrameData[24] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1534_ VPWR _0206_ _0205_ VGND sg13g2_inv_1
X_3135_ FrameStrobe[0] FrameStrobe_O[0] VPWR VGND sg13g2_buf_1
X_1396_ _0071_ VPWR _0073_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q _0072_
+ sg13g2_o21ai_1
X_3066_ Inst_LUT4AB_switch_matrix.E2BEG7 E2BEG[7] VPWR VGND sg13g2_buf_1
X_2017_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q VPWR _0671_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q
+ _0366_ sg13g2_o21ai_1
XFILLER_35_261 VPWR VGND sg13g2_fill_1
X_2919_ FrameData[8] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_23_423 VPWR VGND sg13g2_fill_1
X_1181_ VPWR _1022_ S4END[0] VGND sg13g2_inv_1
X_1250_ _1089_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q Inst_LUT4AB_switch_matrix.M_EF
+ VPWR VGND sg13g2_nand2b_1
X_2635_ FrameData[12] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_2704_ FrameData[17] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_2566_ FrameData[7] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_1517_ _0189_ VPWR _0190_ VGND N1END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ sg13g2_o21ai_1
X_2497_ FrameData[2] FrameStrobe[16] Inst_LD_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_dlhq_1
X_1448_ _0123_ VPWR _0124_ VGND W2END[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q
+ sg13g2_o21ai_1
X_3118_ FrameData[15] FrameData_O[15] VPWR VGND sg13g2_buf_1
X_1379_ VPWR VGND _1160_ _0053_ _0056_ _1124_ _0057_ _0008_ sg13g2_a221oi_1
X_3049_ VPWR VGND _1165_ sg13g2_tiehi
XFILLER_23_89 VPWR VGND sg13g2_fill_2
X_2420_ VPWR VGND Inst_LUT4AB_switch_matrix.DEBUG_select_LG_SR[0] _0630_ _0985_ _0632_
+ _1010_ _0635_ sg13g2_a221oi_1
X_2282_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q C D E F Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0913_ VPWR VGND sg13g2_mux4_1
X_2351_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q E6END[1] S4END[1] S2END[2] A Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q
+ Inst_LUT4AB_switch_matrix.S4BEG0 VPWR VGND sg13g2_mux4_1
X_1233_ A B Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1073_ VPWR VGND sg13g2_mux2_1
X_1302_ VPWR VGND _1138_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q _1136_ _1027_ _1139_
+ _1134_ sg13g2_a221oi_1
X_1997_ _0650_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0649_ _0653_ VPWR VGND sg13g2_mux4_1
X_2549_ FrameData[22] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_2618_ FrameData[27] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_43_337 VPWR VGND sg13g2_fill_2
XFILLER_34_55 VPWR VGND sg13g2_fill_2
XFILLER_18_89 VPWR VGND sg13g2_fill_1
X_1920_ _0579_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q W1END[3] VPWR VGND sg13g2_nand2b_1
X_1851_ S1END[3] S2END[7] Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q _0512_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_42_392 VPWR VGND sg13g2_fill_1
X_1782_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q _0443_ _0446_ _1039_ sg13g2_a21oi_1
X_2403_ Inst_LC_LUT4c_frame_config_dffesr.c_reset_value _0467_ _0996_ _0997_ VPWR
+ VGND sg13g2_mux2_1
X_2334_ _0957_ VPWR Inst_LUT4AB_switch_matrix.NN4BEG1 VGND _1050_ _0955_ sg13g2_o21ai_1
X_2196_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q _1158_ _0196_ _0276_ _0556_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0838_ VPWR VGND sg13g2_mux4_1
X_2265_ _0894_ _0897_ _0898_ VPWR VGND sg13g2_nor2_1
X_1216_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q N1END[0] N2END[2] N4END[2] E2END[2]
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q _1057_ VPWR VGND sg13g2_mux4_1
XFILLER_27_0 VPWR VGND sg13g2_fill_2
XFILLER_52_156 VPWR VGND sg13g2_fill_1
XFILLER_33_370 VPWR VGND sg13g2_fill_1
XFILLER_28_197 VPWR VGND sg13g2_fill_1
XFILLER_45_76 VPWR VGND sg13g2_fill_1
XANTENNA_8 VPWR VGND EE4END[8] sg13g2_antennanp
X_2050_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ _0702_ VPWR VGND sg13g2_mux4_1
X_2952_ FrameData[9] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1834_ _0492_ _0495_ _0473_ _0496_ VPWR VGND sg13g2_mux2_1
X_1903_ _0556_ _0561_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q _0562_ VPWR VGND sg13g2_mux2_1
X_2883_ FrameData[4] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_1765_ _0427_ _0428_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q _0429_ VPWR VGND sg13g2_nand3_1
X_1696_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q _0361_ _0362_ VPWR VGND sg13g2_nor2_1
X_2317_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _0276_ _0943_ _0942_
+ sg13g2_a21oi_1
X_2248_ _0879_ _0882_ _0883_ VPWR VGND sg13g2_nor2_1
X_2179_ _0821_ VPWR _0822_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q _1052_ sg13g2_o21ai_1
X_3297_ WW4END[9] WW4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_0_277 VPWR VGND sg13g2_fill_2
XFILLER_16_112 VPWR VGND sg13g2_fill_2
X_1550_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q N1END[2] N2END[6] E1END[2] E2END[6]
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0222_ VPWR VGND sg13g2_mux4_1
X_3220_ S2MID[1] S2BEGb[1] VPWR VGND sg13g2_buf_1
X_1481_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q F _0155_ VPWR VGND sg13g2_nor2_1
X_3151_ FrameStrobe[16] FrameStrobe_O[16] VPWR VGND sg13g2_buf_1
X_2102_ _0750_ Inst_LUT4AB_switch_matrix.JS2BEG7 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ VPWR VGND sg13g2_nand2b_1
X_3082_ E6END[9] E6BEG[7] VPWR VGND sg13g2_buf_1
X_2033_ _0679_ _0686_ _0687_ VPWR VGND sg13g2_and2_1
X_2935_ FrameData[24] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_2866_ FrameData[19] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1817_ _0311_ _0209_ _0312_ _0479_ VPWR VGND sg13g2_a21o_1
X_1748_ _0412_ VPWR _0413_ VGND W2END[3] Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q
+ sg13g2_o21ai_1
X_2797_ FrameData[14] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_1679_ _0344_ _0346_ _0339_ _0347_ VPWR VGND sg13g2_nand3_1
XFILLER_21_170 VPWR VGND sg13g2_fill_2
X_1602_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q _0270_ _0273_ _0272_ sg13g2_a21oi_1
X_2651_ FrameData[28] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_2582_ FrameData[23] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_2720_ FrameData[1] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_3203_ Inst_LUT4AB_switch_matrix.NN4BEG0 NN4BEG[12] VPWR VGND sg13g2_buf_1
X_1464_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q N1END[1] N2END[5] E1END[1] E2END[5]
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q _0139_ VPWR VGND sg13g2_mux4_1
X_1395_ _0043_ _0048_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q _0072_ VPWR VGND
+ sg13g2_mux2_1
X_1533_ _0205_ _0202_ _0203_ VPWR VGND sg13g2_nand2_1
X_2016_ E F _0670_ Inst_LUT4AB_switch_matrix.M_EF VPWR VGND sg13g2_mux2_1
X_3134_ FrameData[31] FrameData_O[31] VPWR VGND sg13g2_buf_1
X_3065_ Inst_LUT4AB_switch_matrix.E2BEG6 E2BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_27_207 VPWR VGND sg13g2_fill_2
X_2918_ FrameData[7] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_2849_ FrameData[2] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_49_332 VPWR VGND sg13g2_fill_1
X_1180_ VPWR _1021_ N2MID[4] VGND sg13g2_inv_1
X_1516_ _0189_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q N2END[5] VPWR VGND sg13g2_nand2b_1
X_2565_ FrameData[6] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VPWR VGND sg13g2_dlhq_1
X_2634_ FrameData[11] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_2703_ FrameData[16] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_3117_ FrameData[14] FrameData_O[14] VPWR VGND sg13g2_buf_1
X_2496_ FrameData[1] FrameStrobe[16] Inst_LD_LUT4c_frame_config_dffesr.c_out_mux VPWR
+ VGND sg13g2_dlhq_1
X_1447_ _0123_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q W6END[1] VPWR VGND sg13g2_nand2b_1
X_1378_ _0055_ _0054_ _1085_ _0056_ VPWR VGND sg13g2_mux2_1
X_3048_ VPWR VGND _1164_ sg13g2_tiehi
XFILLER_2_136 VPWR VGND sg13g2_fill_2
XFILLER_14_298 VPWR VGND sg13g2_fill_1
X_2281_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q E1END[3] W1END[3] A B Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q
+ _0912_ VPWR VGND sg13g2_mux4_1
X_1232_ _1072_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _1071_ VPWR VGND sg13g2_nand2_1
X_1301_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q _1137_ _1138_ _1027_ sg13g2_a21oi_1
X_2350_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q E6END[0] S4END[2] S2END[3] B Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q
+ Inst_LUT4AB_switch_matrix.S4BEG1 VPWR VGND sg13g2_mux4_1
X_1996_ _0649_ _0650_ _0652_ VPWR VGND sg13g2_nor2_1
X_2548_ FrameData[21] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_2617_ FrameData[26] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_2479_ FrameData[16] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.c_reset_value
+ VPWR VGND sg13g2_dlhq_1
XFILLER_28_379 VPWR VGND sg13g2_fill_1
X_1850_ _0510_ VPWR _0511_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q W1END[1]
+ sg13g2_o21ai_1
X_1781_ VGND VPWR _0445_ _0444_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q sg13g2_or2_1
X_2333_ _0957_ _1050_ _0956_ VPWR VGND sg13g2_nand2_1
X_2402_ _0996_ Inst_LUT4AB_switch_matrix.DEBUG_select_LC_SR[0] _0985_ VPWR VGND sg13g2_nand2_1
X_1215_ _1056_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q _1055_ VPWR VGND sg13g2_nand2_1
X_2264_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit28.Q VPWR _0897_ VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q
+ _0896_ sg13g2_o21ai_1
X_2195_ _0826_ VPWR Inst_LUT4AB_switch_matrix.JN2BEG0 VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q
+ _0837_ sg13g2_o21ai_1
X_1979_ VGND VPWR _0632_ _0635_ _0636_ _0630_ sg13g2_a21oi_1
XANTENNA_9 VPWR VGND N4END[12] sg13g2_antennanp
X_1902_ _0560_ VPWR _0561_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q _0557_ sg13g2_o21ai_1
X_2951_ FrameData[8] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1833_ _0493_ _0494_ _0486_ _0495_ VPWR VGND sg13g2_mux2_1
X_2882_ FrameData[3] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1764_ _0428_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q W2END[0] VPWR VGND sg13g2_nand2_1
X_2316_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q E _0942_ VPWR VGND sg13g2_nor2_1
X_3296_ WW4END[8] WW4BEG[4] VPWR VGND sg13g2_buf_1
X_1695_ E2END[3] SS4END[3] Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q _0361_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_53_422 VPWR VGND sg13g2_fill_2
X_2247_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q VPWR _0882_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q
+ _0881_ sg13g2_o21ai_1
X_2178_ _0821_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q Inst_LUT4AB_switch_matrix.M_AB
+ VPWR VGND sg13g2_nand2_1
XFILLER_31_68 VPWR VGND sg13g2_fill_1
XFILLER_0_289 VPWR VGND sg13g2_fill_1
X_3150_ FrameStrobe[15] FrameStrobe_O[15] VPWR VGND sg13g2_buf_1
X_1480_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0151_ _0154_ _0153_ sg13g2_a21oi_1
X_2101_ _0749_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q Inst_LUT4AB_switch_matrix.JW2BEG7
+ VPWR VGND sg13g2_nand2_1
X_2032_ _0686_ _0676_ _0685_ VPWR VGND sg13g2_nand2b_1
X_3081_ E6END[8] E6BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_50_414 VPWR VGND sg13g2_fill_1
X_2865_ FrameData[18] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_2934_ FrameData[23] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_30_171 VPWR VGND sg13g2_fill_1
X_1678_ _0346_ _0247_ _0345_ VPWR VGND sg13g2_nand2b_1
X_1816_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q _0238_ _0478_ _0477_ sg13g2_a21oi_1
X_2796_ FrameData[13] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_1747_ _0412_ _1028_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q VPWR VGND sg13g2_nand2_1
X_3279_ W2MID[7] W2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_17_422 VPWR VGND sg13g2_fill_2
XFILLER_16_90 VPWR VGND sg13g2_fill_1
X_1601_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VPWR _0272_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ _0271_ sg13g2_o21ai_1
X_2650_ FrameData[27] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_2581_ FrameData[22] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1532_ VGND VPWR _0204_ _0203_ _0202_ sg13g2_or2_1
X_3202_ NN4END[15] NN4BEG[11] VPWR VGND sg13g2_buf_1
X_1463_ _0137_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q _0138_ VPWR VGND sg13g2_nor2b_1
X_3133_ FrameData[30] FrameData_O[30] VPWR VGND sg13g2_buf_1
X_1394_ _0022_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q _0070_ _0071_ VPWR VGND
+ sg13g2_a21o_1
X_2015_ _0668_ _0669_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0670_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_35_285 VPWR VGND sg13g2_fill_1
X_3064_ Inst_LUT4AB_switch_matrix.E2BEG5 E2BEG[5] VPWR VGND sg13g2_buf_1
X_2917_ FrameData[6] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_2848_ FrameData[1] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_2779_ FrameData[28] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_18_208 VPWR VGND sg13g2_fill_1
XFILLER_26_296 VPWR VGND sg13g2_fill_2
XFILLER_49_322 VPWR VGND sg13g2_fill_2
X_2702_ FrameData[15] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_2564_ FrameData[5] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VPWR VGND sg13g2_dlhq_1
X_1515_ _0187_ VPWR _0188_ VGND E1END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ sg13g2_o21ai_1
X_2633_ FrameData[10] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_2495_ FrameData[0] FrameStrobe[16] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_3116_ FrameData[13] FrameData_O[13] VPWR VGND sg13g2_buf_1
X_1377_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _1121_ _0055_ VPWR VGND sg13g2_mux2_1
X_1446_ _0122_ _1032_ _0121_ VPWR VGND sg13g2_nand2_1
X_3047_ VPWR VGND _1163_ sg13g2_tiehi
X_2280_ _0907_ _0911_ Inst_LUT4AB_switch_matrix.E6BEG1 VPWR VGND sg13g2_nor2_1
X_1231_ C E Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1071_ VPWR VGND sg13g2_mux2_1
X_1300_ W2END[2] W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q _1137_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_45_380 VPWR VGND sg13g2_fill_1
X_1995_ _0651_ _0649_ _0650_ VPWR VGND sg13g2_nand2_1
X_2616_ FrameData[25] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_2547_ FrameData[20] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_1429_ _0105_ VPWR _0106_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0083_ sg13g2_o21ai_1
X_2478_ FrameData[15] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_dlhq_1
XFILLER_34_57 VPWR VGND sg13g2_fill_1
XFILLER_50_56 VPWR VGND sg13g2_fill_1
X_1780_ S1END[1] S1END[3] Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q _0444_ VPWR VGND
+ sg13g2_mux2_1
X_2332_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q N1END[3] E1END[3] W1END[3] A Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ _0956_ VPWR VGND sg13g2_mux4_1
XFILLER_6_273 VPWR VGND sg13g2_fill_2
X_2401_ _0995_ Inst_LUT4AB_switch_matrix.DEBUG_select_LC_EN[0] _0973_ VPWR VGND sg13g2_nand2b_1
XFILLER_27_2 VPWR VGND sg13g2_fill_1
X_1214_ _1053_ _1054_ _1020_ _1055_ VPWR VGND sg13g2_mux2_1
X_2263_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q _1084_ _0896_ _0895_
+ sg13g2_a21oi_1
X_2194_ _0831_ VPWR _0837_ VGND _0833_ _0836_ sg13g2_o21ai_1
X_1978_ _0627_ _0634_ _0635_ VPWR VGND sg13g2_nor2_1
XFILLER_43_136 VPWR VGND sg13g2_fill_2
XFILLER_28_155 VPWR VGND sg13g2_fill_1
X_1832_ _0481_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ _0487_ _0494_ VPWR VGND sg13g2_mux4_1
X_2881_ FrameData[2] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_1901_ _0558_ _0559_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q _0560_ VPWR VGND sg13g2_nand3_1
X_2950_ FrameData[7] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1694_ Inst_LUT4AB_switch_matrix.JN2BEG2 _0354_ _0360_ _0352_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q
+ VPWR VGND sg13g2_a22oi_1
X_1763_ _0427_ S2END[0] Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q VPWR VGND sg13g2_nand2b_1
X_2315_ W1END[1] D Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _0941_ VPWR VGND sg13g2_mux2_1
XFILLER_32_0 VPWR VGND sg13g2_fill_1
X_2246_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q _0308_ _0881_ _0880_ sg13g2_a21oi_1
X_3295_ WW4END[7] WW4BEG[3] VPWR VGND sg13g2_buf_1
X_2177_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q G _0820_ _0819_ sg13g2_a21oi_1
XFILLER_0_279 VPWR VGND sg13g2_fill_1
XFILLER_16_114 VPWR VGND sg13g2_fill_1
XFILLER_24_191 VPWR VGND sg13g2_fill_2
XFILLER_8_346 VPWR VGND sg13g2_fill_2
XFILLER_39_206 VPWR VGND sg13g2_fill_1
X_3080_ E6END[7] E6BEG[5] VPWR VGND sg13g2_buf_1
X_2100_ Inst_LUT4AB_switch_matrix.JN2BEG7 Inst_LUT4AB_switch_matrix.E2BEG7 Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q
+ _0748_ VPWR VGND sg13g2_mux2_1
X_2031_ _0149_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0199_ _0685_ VPWR VGND sg13g2_mux4_1
X_2795_ FrameData[12] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1815_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q _0239_ _0477_ VPWR VGND sg13g2_nor2b_1
X_2864_ FrameData[17] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_2933_ FrameData[22] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1677_ _0280_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0310_ _0345_ VPWR VGND sg13g2_mux4_1
X_1746_ S4END[3] SS4END[3] Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q _0411_ VPWR VGND
+ sg13g2_mux2_1
X_2229_ _0867_ _1048_ _0866_ VPWR VGND sg13g2_nand2_1
X_3278_ W2MID[6] W2BEGb[6] VPWR VGND sg13g2_buf_1
XFILLER_29_294 VPWR VGND sg13g2_fill_2
X_1462_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q _0135_ _0137_ _0136_ sg13g2_a21oi_1
X_1600_ S1END[2] S2END[6] Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q _0271_ VPWR VGND
+ sg13g2_mux2_1
X_2580_ FrameData[21] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_1531_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q _0197_ _0198_ _0170_ _0169_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q
+ _0203_ VPWR VGND sg13g2_mux4_1
X_3201_ NN4END[14] NN4BEG[10] VPWR VGND sg13g2_buf_1
X_3132_ FrameData[29] FrameData_O[29] VPWR VGND sg13g2_buf_1
X_1393_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit19.Q VPWR _0070_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit18.Q
+ _0023_ sg13g2_o21ai_1
X_3063_ Inst_LUT4AB_switch_matrix.E2BEG4 E2BEG[4] VPWR VGND sg13g2_buf_1
X_2014_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_switch_matrix.E2BEG4 Inst_LUT4AB_switch_matrix.JW2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q _0669_ VPWR VGND sg13g2_mux4_1
X_2778_ FrameData[27] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_2847_ FrameData[0] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_2916_ FrameData[5] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1729_ _0394_ _0393_ _0368_ VPWR VGND sg13g2_nand2b_1
X_2632_ FrameData[9] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_2701_ FrameData[14] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_2563_ FrameData[4] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VPWR VGND sg13g2_dlhq_1
X_1514_ _0187_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q E2END[5] VPWR VGND sg13g2_nand2b_1
X_1445_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q N1END[1] N4END[3] N2END[3] E2END[3]
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q _0121_ VPWR VGND sg13g2_mux4_1
X_2494_ FrameData[31] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_3046_ _1169_ VGND VPWR _0007_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop clknet_1_1__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_3115_ FrameData[12] FrameData_O[12] VPWR VGND sg13g2_buf_1
X_1376_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _1121_ _0054_ VPWR VGND sg13g2_mux2_1
XFILLER_48_67 VPWR VGND sg13g2_fill_1
XFILLER_49_142 VPWR VGND sg13g2_fill_2
XFILLER_49_131 VPWR VGND sg13g2_fill_1
X_1230_ VGND VPWR _1017_ _1069_ _1070_ _1018_ sg13g2_a21oi_1
X_1994_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q _0585_ _0586_ _0588_ _0587_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q
+ _0650_ VPWR VGND sg13g2_mux4_1
X_2615_ FrameData[24] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_2546_ FrameData[19] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VPWR VGND sg13g2_dlhq_1
X_2477_ FrameData[14] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_dlhq_1
X_1428_ _0105_ _0078_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 VPWR
+ VGND sg13g2_nand2b_1
X_3029_ FrameData[22] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1359_ VPWR Inst_LUT4AB_switch_matrix.JW2BEG3 _0037_ VGND sg13g2_inv_1
XFILLER_28_326 VPWR VGND sg13g2_fill_2
X_2400_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop _0994_ _0992_ _0002_ VPWR VGND
+ sg13g2_mux2_1
X_2331_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q _1052_ _1158_ _0196_ _0290_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q
+ _0955_ VPWR VGND sg13g2_mux4_1
X_1213_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q A D C E Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q
+ _1054_ VPWR VGND sg13g2_mux4_1
X_2262_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q G _0895_ VPWR VGND sg13g2_nor2b_1
XFILLER_52_137 VPWR VGND sg13g2_fill_1
X_2193_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VPWR _0836_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ _0835_ sg13g2_o21ai_1
X_1977_ _0532_ _0633_ _0634_ VPWR VGND sg13g2_nor2_1
X_2529_ FrameData[2] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
XFILLER_20_38 VPWR VGND sg13g2_fill_1
XFILLER_16_318 VPWR VGND sg13g2_fill_2
X_1831_ _0481_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ _0487_ _0493_ VPWR VGND sg13g2_mux4_1
XFILLER_42_170 VPWR VGND sg13g2_fill_2
X_1900_ _0559_ W2MID[5] Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q VPWR VGND sg13g2_nand2_1
X_2880_ FrameData[1] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_15_351 VPWR VGND sg13g2_fill_1
X_1693_ VGND VPWR _0356_ _0359_ _0360_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit5.Q sg13g2_a21oi_1
X_1762_ N2END[0] EE4END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q _0426_ VPWR VGND
+ sg13g2_mux2_1
X_2314_ N1END[1] E1END[1] Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q _0940_ VPWR VGND
+ sg13g2_mux2_1
X_2245_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q C _0880_ VPWR VGND sg13g2_nor2b_1
X_2176_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q F _0819_ VPWR VGND sg13g2_nor2b_1
X_3294_ WW4END[6] WW4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_25_0 VPWR VGND sg13g2_fill_2
XFILLER_21_321 VPWR VGND sg13g2_fill_1
XFILLER_21_343 VPWR VGND sg13g2_fill_2
XFILLER_16_159 VPWR VGND sg13g2_fill_2
XFILLER_12_398 VPWR VGND sg13g2_fill_2
X_2030_ VGND VPWR _0684_ _0683_ _0676_ sg13g2_or2_1
X_2932_ FrameData[21] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_1814_ VGND VPWR _0476_ _0475_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit21.Q sg13g2_or2_1
X_2794_ FrameData[11] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_2863_ FrameData[16] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_1745_ _0409_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q _0410_ VPWR VGND sg13g2_nor2b_1
X_1676_ VGND VPWR _0344_ _0343_ _0247_ sg13g2_or2_1
XFILLER_7_391 VPWR VGND sg13g2_fill_2
XFILLER_38_251 VPWR VGND sg13g2_fill_1
X_2228_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q N1END[3] S1END[3] W1END[3] A Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ _0866_ VPWR VGND sg13g2_mux4_1
X_3277_ W2MID[5] W2BEGb[5] VPWR VGND sg13g2_buf_1
X_2159_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q C _0803_ _0802_ sg13g2_a21oi_1
XFILLER_26_48 VPWR VGND sg13g2_fill_1
XFILLER_29_273 VPWR VGND sg13g2_fill_2
X_3200_ NN4END[13] NN4BEG[9] VPWR VGND sg13g2_buf_1
X_1461_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR _0136_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ _0133_ sg13g2_o21ai_1
X_1392_ _0069_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop Inst_LA_LUT4c_frame_config_dffesr.c_out_mux
+ A VPWR VGND sg13g2_mux2_1
XFILLER_8_199 VPWR VGND sg13g2_fill_1
X_1530_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q _0147_ _0148_ _0130_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q
+ _0202_ VPWR VGND sg13g2_mux4_1
X_2013_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q Inst_LUT4AB_switch_matrix.JN2BEG6
+ Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_switch_matrix.E2BEG6 Inst_LUT4AB_switch_matrix.JW2BEG6
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q _0668_ VPWR VGND sg13g2_mux4_1
X_3131_ FrameData[28] FrameData_O[28] VPWR VGND sg13g2_buf_1
X_3062_ Inst_LUT4AB_switch_matrix.E2BEG3 E2BEG[3] VPWR VGND sg13g2_buf_1
X_2915_ FrameData[4] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_2777_ FrameData[26] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_2846_ FrameData[31] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1728_ _0392_ VPWR _0393_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q _0389_
+ sg13g2_o21ai_1
X_1659_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q _0327_ _0328_ VPWR VGND sg13g2_nor2_1
XFILLER_49_324 VPWR VGND sg13g2_fill_1
XFILLER_32_257 VPWR VGND sg13g2_fill_1
XFILLER_17_276 VPWR VGND sg13g2_fill_1
XFILLER_17_298 VPWR VGND sg13g2_fill_1
X_2631_ FrameData[8] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_2562_ FrameData[3] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VPWR VGND sg13g2_dlhq_1
X_2700_ FrameData[13] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_1513_ _0185_ VPWR _0186_ VGND W1END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ sg13g2_o21ai_1
X_1375_ VGND VPWR _0049_ _0050_ _0053_ _0052_ sg13g2_a21oi_1
X_2493_ FrameData[30] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_1444_ _1033_ _0114_ _0119_ _0120_ VPWR VGND sg13g2_nor3_1
X_3045_ _1170_ VGND VPWR _0006_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop clknet_1_1__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_3114_ FrameData[11] FrameData_O[11] VPWR VGND sg13g2_buf_1
X_2829_ FrameData[14] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_49_110 VPWR VGND sg13g2_fill_1
XFILLER_49_165 VPWR VGND sg13g2_fill_2
XFILLER_45_371 VPWR VGND sg13g2_fill_1
X_1993_ _0648_ VPWR _0649_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q _0646_ sg13g2_o21ai_1
X_2545_ FrameData[18] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VPWR VGND sg13g2_dlhq_1
X_2614_ FrameData[23] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1358_ _0027_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q _0036_ _0037_ VPWR VGND sg13g2_a21o_1
X_1427_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0081_ _0104_ VPWR
+ VGND sg13g2_nor2_1
X_2476_ FrameData[13] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_3028_ FrameData[21] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_1289_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q G _1126_ _1125_ sg13g2_a21oi_1
XFILLER_1_5 VPWR VGND sg13g2_fill_2
XFILLER_6_264 VPWR VGND sg13g2_fill_1
X_2192_ VGND VPWR SS4END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q _0835_ _0834_
+ sg13g2_a21oi_1
X_1212_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q F G H Inst_LUT4AB_switch_matrix.M_AB
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q _1053_ VPWR VGND sg13g2_mux4_1
X_2261_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q _0626_ _0894_ _0893_
+ sg13g2_a21oi_1
X_2330_ VGND VPWR _0948_ _0952_ Inst_LUT4AB_switch_matrix.NN4BEG2 _0954_ sg13g2_a21oi_1
XFILLER_33_341 VPWR VGND sg13g2_fill_1
X_1976_ _0590_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0565_ _0633_ VPWR VGND sg13g2_mux4_1
X_2528_ FrameData[1] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_2459_ FrameData[28] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_dlhq_1
XFILLER_43_138 VPWR VGND sg13g2_fill_1
XFILLER_6_19 VPWR VGND sg13g2_fill_2
XFILLER_3_234 VPWR VGND sg13g2_fill_2
XFILLER_47_422 VPWR VGND sg13g2_fill_2
X_1830_ _0489_ _0491_ _0486_ _0492_ VPWR VGND sg13g2_mux2_1
X_1761_ VPWR _0425_ _0424_ VGND sg13g2_inv_1
XFILLER_15_374 VPWR VGND sg13g2_fill_1
X_2313_ _0937_ _0939_ Inst_LUT4AB_switch_matrix.EE4BEG0 VPWR VGND sg13g2_nor2_1
X_1692_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q _0358_ _0359_ _1031_ sg13g2_a21oi_1
X_2244_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q _0430_ _0879_ _0878_ sg13g2_a21oi_1
X_2175_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q B D C E Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ _0818_ VPWR VGND sg13g2_mux4_1
X_3293_ WW4END[5] WW4BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_18_0 VPWR VGND sg13g2_fill_2
XFILLER_40_108 VPWR VGND sg13g2_fill_2
X_1959_ N2MID[0] E2MID[0] Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q _0616_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_31_49 VPWR VGND sg13g2_fill_2
XFILLER_24_160 VPWR VGND sg13g2_fill_2
XFILLER_47_230 VPWR VGND sg13g2_fill_1
X_2931_ FrameData[20] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_1813_ _0474_ VPWR _0475_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q _0236_ sg13g2_o21ai_1
X_2862_ FrameData[15] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_2793_ FrameData[10] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1744_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q _0407_ _0409_ _0408_ sg13g2_a21oi_1
XFILLER_30_152 VPWR VGND sg13g2_fill_2
X_1675_ _0280_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0310_ _0343_ VPWR VGND sg13g2_mux4_1
X_3276_ W2MID[4] W2BEGb[4] VPWR VGND sg13g2_buf_1
X_2227_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q _1052_ _1158_ _0196_ _0253_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q
+ _0865_ VPWR VGND sg13g2_mux4_1
X_2158_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q B _0802_ VPWR VGND sg13g2_nor2b_1
X_2089_ _0738_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0737_ VPWR VGND sg13g2_nand2b_1
XFILLER_12_163 VPWR VGND sg13g2_fill_1
XFILLER_12_185 VPWR VGND sg13g2_fill_1
X_1460_ _0134_ VPWR _0135_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q H sg13g2_o21ai_1
X_3130_ FrameData[27] FrameData_O[27] VPWR VGND sg13g2_buf_1
X_1391_ VGND VPWR _0061_ _0068_ _0069_ _0057_ sg13g2_a21oi_1
X_2012_ _0667_ VPWR H VGND Inst_LH_LUT4c_frame_config_dffesr.c_out_mux _0666_ sg13g2_o21ai_1
X_3061_ Inst_LUT4AB_switch_matrix.E2BEG2 E2BEG[2] VPWR VGND sg13g2_buf_1
X_2845_ FrameData[30] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_2914_ FrameData[3] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1658_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q _0324_ _0327_ _0326_ sg13g2_a21oi_1
X_2776_ FrameData[25] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1727_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q _0391_ _0392_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q
+ sg13g2_a21oi_1
X_1589_ H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ _0260_ VPWR VGND sg13g2_mux2_1
X_3259_ clknet_1_0__leaf_UserCLK UserCLKo VPWR VGND sg13g2_buf_1
XFILLER_53_36 VPWR VGND sg13g2_fill_1
XFILLER_26_277 VPWR VGND sg13g2_fill_2
XFILLER_49_303 VPWR VGND sg13g2_fill_2
X_1512_ _0185_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q W1END[3] VPWR VGND sg13g2_nand2b_1
X_2630_ FrameData[7] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_2561_ FrameData[2] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VPWR VGND sg13g2_dlhq_1
X_2492_ FrameData[29] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_3113_ FrameData[10] FrameData_O[10] VPWR VGND sg13g2_buf_1
X_1374_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q _0022_ _0052_ _0051_ sg13g2_a21oi_1
X_1443_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0116_ _0119_ _0118_ sg13g2_a21oi_1
X_3044_ _1163_ VGND VPWR _0005_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop clknet_1_1__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_2828_ FrameData[13] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_2759_ FrameData[8] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1992_ _0537_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q _0647_ _0648_ VPWR VGND sg13g2_a21o_1
XFILLER_9_251 VPWR VGND sg13g2_fill_1
X_2544_ FrameData[17] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VPWR VGND sg13g2_dlhq_1
X_2613_ FrameData[22] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_2475_ FrameData[12] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_1357_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q _0029_ _0035_ _0036_ VPWR VGND sg13g2_nor3_1
X_1426_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0076_ _0103_ VPWR
+ VGND sg13g2_nor2_1
X_1288_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q F _1125_ VPWR VGND sg13g2_nor2b_1
X_3027_ FrameData[20] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_1211_ VPWR _1052_ H VGND sg13g2_inv_1
X_2260_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit27.Q VPWR _0893_ VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q
+ _0148_ sg13g2_o21ai_1
X_2191_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q E6END[1] _0834_ VPWR VGND sg13g2_nor2b_1
X_1975_ _0632_ _0532_ _0631_ VPWR VGND sg13g2_nand2b_1
X_2527_ FrameData[0] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VPWR VGND sg13g2_dlhq_1
X_1409_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q _1102_ _1103_ _1119_ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit13.Q
+ _0086_ VPWR VGND sg13g2_mux4_1
X_2458_ FrameData[27] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_dlhq_1
XFILLER_29_38 VPWR VGND sg13g2_fill_2
X_2389_ _0986_ Inst_LUT4AB_switch_matrix.DEBUG_select_LH_SR[0] _0985_ VPWR VGND sg13g2_nand2_1
XFILLER_35_92 VPWR VGND sg13g2_fill_2
X_1691_ _0357_ VPWR _0358_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q W2END[3]
+ sg13g2_o21ai_1
X_1760_ _0423_ VPWR _0424_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q _0420_ sg13g2_o21ai_1
X_2312_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q _0938_ _0939_ VPWR VGND sg13g2_nor2_1
X_3292_ WW4END[4] WW4BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_38_423 VPWR VGND sg13g2_fill_1
X_2243_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q VPWR _0878_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit0.Q
+ _0586_ sg13g2_o21ai_1
X_2174_ _0806_ VPWR Inst_LUT4AB_switch_matrix.E2BEG0 VGND _0816_ _0817_ sg13g2_o21ai_1
X_1889_ S1END[3] S2END[7] Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q _0549_ VPWR VGND
+ sg13g2_mux2_1
X_1958_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q VPWR _0615_ VGND _0613_ _0614_ sg13g2_o21ai_1
XFILLER_0_227 VPWR VGND sg13g2_fill_2
X_2930_ FrameData[19] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_2861_ FrameData[14] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_1674_ _0314_ _0339_ _0341_ _0342_ VPWR VGND sg13g2_nor3_1
X_1812_ _0474_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q _0237_ VPWR VGND sg13g2_nand2_1
X_2792_ FrameData[9] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_7_393 VPWR VGND sg13g2_fill_1
X_1743_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR _0408_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ _0405_ sg13g2_o21ai_1
XFILLER_30_197 VPWR VGND sg13g2_fill_2
X_3275_ W2MID[3] W2BEGb[3] VPWR VGND sg13g2_buf_1
X_2226_ _0862_ _0864_ Inst_LUT4AB_switch_matrix.WW4BEG2 VPWR VGND sg13g2_nor2_1
XFILLER_30_0 VPWR VGND sg13g2_fill_2
XFILLER_53_234 VPWR VGND sg13g2_fill_1
XFILLER_53_212 VPWR VGND sg13g2_fill_2
X_2157_ D E Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q _0801_ VPWR VGND sg13g2_mux2_1
X_2088_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q E G F Inst_LUT4AB_switch_matrix.M_AH
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q _0737_ VPWR VGND sg13g2_mux4_1
X_1390_ VPWR VGND _1160_ _0052_ _0067_ _0049_ _0068_ _0050_ sg13g2_a221oi_1
X_3060_ Inst_LUT4AB_switch_matrix.E2BEG1 E2BEG[1] VPWR VGND sg13g2_buf_1
X_2011_ _0667_ Inst_LH_LUT4c_frame_config_dffesr.LUT_flop Inst_LH_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_nand2_1
XFILLER_35_267 VPWR VGND sg13g2_fill_2
X_2844_ FrameData[29] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_2913_ FrameData[2] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_1588_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q _1051_ _0259_ _0258_ sg13g2_a21oi_1
X_1657_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VPWR _0326_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ _0325_ sg13g2_o21ai_1
X_2775_ FrameData[24] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1726_ VPWR _0391_ _0390_ VGND sg13g2_inv_1
X_3189_ Inst_LUT4AB_switch_matrix.N4BEG2 N4BEG[14] VPWR VGND sg13g2_buf_1
X_3258_ Inst_LUT4AB_switch_matrix.SS4BEG3 SS4BEG[15] VPWR VGND sg13g2_buf_1
X_2209_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q _1084_ _0148_ _0308_ _0586_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0850_ VPWR VGND sg13g2_mux4_1
X_1511_ _0183_ VPWR _0184_ VGND S1END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q
+ sg13g2_o21ai_1
X_2560_ FrameData[1] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VPWR VGND sg13g2_dlhq_1
X_2491_ FrameData[28] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_1442_ _1032_ VPWR _0118_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0117_ sg13g2_o21ai_1
X_3043_ _1164_ VGND VPWR _0004_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop clknet_1_0__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_1373_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q VPWR _0051_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q
+ _0023_ sg13g2_o21ai_1
XFILLER_4_97 VPWR VGND sg13g2_fill_2
X_3112_ FrameData[9] FrameData_O[9] VPWR VGND sg13g2_buf_1
XFILLER_23_18 VPWR VGND sg13g2_fill_1
X_2758_ FrameData[7] FrameStrobe[8] Inst_LUT4AB_switch_matrix.DEBUG_select_LG_EN[0]
+ VPWR VGND sg13g2_dlhq_1
X_2827_ FrameData[12] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1709_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VPWR _0375_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ _0372_ sg13g2_o21ai_1
X_2689_ FrameData[2] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_14_215 VPWR VGND sg13g2_fill_2
XFILLER_8_0 VPWR VGND sg13g2_fill_1
X_1991_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q VPWR _0647_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q
+ _0538_ sg13g2_o21ai_1
X_2612_ FrameData[21] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_2543_ FrameData[16] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VPWR VGND sg13g2_dlhq_1
X_1425_ _0098_ _0099_ _0101_ _0102_ VPWR VGND sg13g2_nor3_1
X_2474_ FrameData[11] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_3026_ FrameData[19] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1356_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q _0033_ _0035_ _0034_ sg13g2_a21oi_1
X_1287_ _1122_ _1123_ _1085_ _1124_ VPWR VGND sg13g2_nand3_1
XFILLER_1_87 VPWR VGND sg13g2_fill_1
X_1210_ VPWR _1051_ G VGND sg13g2_inv_1
X_2190_ VGND VPWR _1028_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q _0833_ _0832_ sg13g2_a21oi_1
X_1974_ _0590_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0565_ _0631_ VPWR VGND sg13g2_mux4_1
XFILLER_33_376 VPWR VGND sg13g2_fill_2
X_2526_ FrameData[31] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_409 VPWR VGND sg13g2_fill_1
X_1408_ _0077_ _0079_ _0082_ _0084_ _0085_ VPWR VGND sg13g2_or4_1
X_2457_ FrameData[26] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_2388_ VGND VPWR _0983_ _0984_ _0985_ _0979_ sg13g2_a21oi_1
X_1339_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q _0017_ _0019_ _0018_ sg13g2_a21oi_1
XFILLER_24_343 VPWR VGND sg13g2_fill_2
X_3009_ FrameData[2] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_1690_ _0357_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q _1030_ VPWR VGND sg13g2_nand2_1
X_2311_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q N1END[2] S1END[2] E1END[2] F Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
+ _0938_ VPWR VGND sg13g2_mux4_1
X_3291_ Inst_LUT4AB_switch_matrix.W6BEG1 W6BEG[11] VPWR VGND sg13g2_buf_1
X_2242_ _0871_ _0877_ Inst_LUT4AB_switch_matrix.SS4BEG3 VPWR VGND sg13g2_nor2_1
X_2173_ _0817_ _0811_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q VPWR VGND sg13g2_nand2b_1
X_1957_ W2MID[0] Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q _0614_ VPWR VGND sg13g2_nor2_1
XFILLER_21_302 VPWR VGND sg13g2_fill_2
X_1888_ _0547_ VPWR _0548_ VGND W1END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ sg13g2_o21ai_1
X_2509_ FrameData[14] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
XFILLER_50_419 VPWR VGND sg13g2_fill_1
X_2860_ FrameData[13] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_1811_ _0473_ _0470_ _0472_ _0469_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q VPWR
+ VGND sg13g2_a22oi_1
X_2791_ FrameData[8] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1673_ _0247_ _0340_ _0341_ VPWR VGND sg13g2_nor2_1
X_1742_ _0406_ VPWR _0407_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q H sg13g2_o21ai_1
X_2225_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q _0863_ _0864_ VPWR VGND sg13g2_nor2_1
X_3274_ W2MID[2] W2BEGb[2] VPWR VGND sg13g2_buf_1
XFILLER_23_0 VPWR VGND sg13g2_fill_1
X_2156_ _0798_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0799_ _0800_ VPWR VGND sg13g2_a21o_1
X_2087_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ _0736_ VPWR VGND sg13g2_mux4_1
X_2989_ FrameData[14] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_32_408 VPWR VGND sg13g2_fill_1
XFILLER_32_72 VPWR VGND sg13g2_fill_2
XFILLER_32_50 VPWR VGND sg13g2_fill_1
X_2010_ VGND VPWR _0661_ _0665_ _0666_ _0659_ sg13g2_a21oi_1
XFILLER_35_202 VPWR VGND sg13g2_fill_2
X_2912_ FrameData[1] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_2774_ FrameData[23] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_2843_ FrameData[28] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_1725_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q N2MID[7] E2MID[7] S2MID[7] W2MID[7]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q _0390_ VPWR VGND sg13g2_mux4_1
X_1587_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q E _0258_ VPWR VGND sg13g2_nor2_1
X_1656_ S1END[0] S1END[2] Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q _0325_ VPWR VGND
+ sg13g2_mux2_1
X_3188_ Inst_LUT4AB_switch_matrix.N4BEG1 N4BEG[13] VPWR VGND sg13g2_buf_1
X_2139_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q VPWR _0784_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ _0783_ sg13g2_o21ai_1
X_2208_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q G H Inst_LUT4AB_switch_matrix.M_AB
+ Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q _0849_
+ VPWR VGND sg13g2_mux4_1
X_3257_ Inst_LUT4AB_switch_matrix.SS4BEG2 SS4BEG[14] VPWR VGND sg13g2_buf_1
XFILLER_1_378 VPWR VGND sg13g2_fill_2
X_1510_ _0183_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q S2END[5] VPWR VGND sg13g2_nand2b_1
X_2490_ FrameData[27] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_1441_ A B Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q _0117_ VPWR VGND sg13g2_mux2_1
X_1372_ VGND VPWR _1029_ _0043_ _0050_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q sg13g2_a21oi_1
X_3042_ _1165_ VGND VPWR _0003_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop clknet_1_0__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_3111_ FrameData[8] FrameData_O[8] VPWR VGND sg13g2_buf_1
X_1708_ _0373_ VPWR _0374_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q H sg13g2_o21ai_1
X_2757_ FrameData[6] FrameStrobe[8] Inst_LUT4AB_switch_matrix.DEBUG_select_LG_SR[0]
+ VPWR VGND sg13g2_dlhq_1
X_2826_ FrameData[11] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_2688_ FrameData[1] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_48_49 VPWR VGND sg13g2_fill_1
X_1639_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit12.Q N2MID[3] E2MID[3] S2MID[3] W2MID[3]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit13.Q _0308_ VPWR VGND sg13g2_mux4_1
XFILLER_46_308 VPWR VGND sg13g2_fill_1
XFILLER_14_227 VPWR VGND sg13g2_fill_2
X_1990_ _0556_ _0561_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q _0646_ VPWR VGND sg13g2_mux2_1
X_2542_ FrameData[15] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VPWR VGND sg13g2_dlhq_1
X_2611_ FrameData[20] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_1355_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q VPWR _0034_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ _0031_ sg13g2_o21ai_1
X_1424_ _0100_ VPWR _0101_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ _0076_ sg13g2_o21ai_1
X_2473_ FrameData[10] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_3025_ FrameData[18] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_1286_ _1123_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 _1121_ VPWR
+ VGND sg13g2_nand2_1
XFILLER_18_19 VPWR VGND sg13g2_fill_2
X_2809_ FrameData[26] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_46_105 VPWR VGND sg13g2_fill_2
XFILLER_6_289 VPWR VGND sg13g2_fill_1
X_1973_ VGND VPWR _0532_ _0593_ _0630_ _0629_ sg13g2_a21oi_1
XFILLER_53_0 VPWR VGND sg13g2_fill_2
X_2525_ FrameData[30] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VPWR VGND sg13g2_dlhq_1
X_2456_ FrameData[25] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_2387_ _0981_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q _0984_ VPWR VGND sg13g2_nor2b_1
X_1338_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q VPWR _0018_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q
+ _0015_ sg13g2_o21ai_1
X_1407_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 _0083_ _0084_ VPWR
+ VGND sg13g2_nor2_1
X_3008_ FrameData[1] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1269_ _1107_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q _1105_ VPWR VGND sg13g2_nand2b_1
XFILLER_30_336 VPWR VGND sg13g2_fill_2
X_2310_ _0933_ _0936_ _0937_ VPWR VGND sg13g2_nor2_1
X_2172_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0814_ _0816_ _0815_ sg13g2_a21oi_1
X_3290_ Inst_LUT4AB_switch_matrix.W6BEG0 W6BEG[10] VPWR VGND sg13g2_buf_1
X_2241_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q _0875_ _0877_ _0876_ sg13g2_a21oi_1
X_1887_ _0547_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q W1END[3] VPWR VGND sg13g2_nand2b_1
X_1956_ Inst_LUT4AB_switch_matrix.JW2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q
+ _0613_ VPWR VGND sg13g2_nor2b_1
X_2508_ FrameData[13] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_229 VPWR VGND sg13g2_fill_1
X_2439_ FrameData[8] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.c_out_mux VPWR
+ VGND sg13g2_dlhq_1
XFILLER_8_318 VPWR VGND sg13g2_fill_1
XFILLER_12_325 VPWR VGND sg13g2_fill_1
XFILLER_46_93 VPWR VGND sg13g2_fill_2
X_2790_ FrameData[7] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1810_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q _0471_ _0472_ VPWR VGND sg13g2_nor2_1
X_1741_ _0406_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q Inst_LUT4AB_switch_matrix.M_EF
+ VPWR VGND sg13g2_nand2b_1
X_1672_ _0280_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ _0310_ _0340_ VPWR VGND sg13g2_mux4_1
XFILLER_30_2 VPWR VGND sg13g2_fill_1
X_3273_ W2MID[1] W2BEGb[1] VPWR VGND sg13g2_buf_1
X_2155_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VPWR _0799_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ _0796_ sg13g2_o21ai_1
X_2224_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q N1END[0] W1END[0] S1END[0] B Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ _0863_ VPWR VGND sg13g2_mux4_1
Xclkbuf_1_0__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_0__leaf_UserCLK_regs VPWR
+ VGND sg13g2_buf_8
X_2086_ Inst_LUT4AB_switch_matrix.JN2BEG7 _0734_ _0735_ _0727_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q
+ VPWR VGND sg13g2_a22oi_1
X_1939_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VPWR _0597_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ _0596_ sg13g2_o21ai_1
X_2988_ FrameData[13] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_44_236 VPWR VGND sg13g2_fill_2
XFILLER_52_291 VPWR VGND sg13g2_fill_2
XFILLER_52_280 VPWR VGND sg13g2_fill_1
XFILLER_35_269 VPWR VGND sg13g2_fill_1
X_2911_ FrameData[0] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_2773_ FrameData[22] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1724_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q E2MID[6] W2MID[6] S2MID[6] Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q _0389_ VPWR VGND sg13g2_mux4_1
X_2842_ FrameData[27] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_1586_ _1042_ _0256_ _0257_ VPWR VGND sg13g2_and2_1
X_1655_ _0323_ VPWR _0324_ VGND S2END[6] Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q
+ sg13g2_o21ai_1
X_3256_ Inst_LUT4AB_switch_matrix.SS4BEG1 SS4BEG[13] VPWR VGND sg13g2_buf_1
X_3187_ Inst_LUT4AB_switch_matrix.N4BEG0 N4BEG[12] VPWR VGND sg13g2_buf_1
X_2138_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q G _0783_ _0782_ sg13g2_a21oi_1
X_2207_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q C D E F Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0848_ VPWR VGND sg13g2_mux4_1
X_2069_ _0719_ VPWR _0720_ VGND S2END[0] Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q
+ sg13g2_o21ai_1
XFILLER_5_129 VPWR VGND sg13g2_fill_2
XFILLER_17_269 VPWR VGND sg13g2_fill_2
XFILLER_27_95 VPWR VGND sg13g2_fill_2
XFILLER_40_250 VPWR VGND sg13g2_fill_2
X_1371_ _0049_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q _0048_ VPWR VGND sg13g2_nand2_1
X_3110_ FrameData[7] FrameData_O[7] VPWR VGND sg13g2_buf_1
X_1440_ _0115_ VPWR _0116_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q D sg13g2_o21ai_1
XFILLER_48_350 VPWR VGND sg13g2_fill_1
X_3041_ _1166_ VGND VPWR _0002_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop clknet_1_0__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
XFILLER_23_217 VPWR VGND sg13g2_fill_2
X_2825_ FrameData[10] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1707_ _0373_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q Inst_LUT4AB_switch_matrix.M_AB
+ VPWR VGND sg13g2_nand2b_1
X_1638_ _0306_ VPWR _0307_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q _0303_ sg13g2_o21ai_1
X_2756_ FrameData[5] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_2687_ FrameData[0] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1569_ _0240_ Inst_LE_LUT4c_frame_config_dffesr.c_I0mux _0209_ VPWR VGND sg13g2_nand2_1
X_3239_ Inst_LUT4AB_switch_matrix.S4BEG0 S4BEG[12] VPWR VGND sg13g2_buf_1
XFILLER_1_143 VPWR VGND sg13g2_fill_2
X_2541_ FrameData[14] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VPWR VGND sg13g2_dlhq_1
X_2610_ FrameData[19] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_2472_ FrameData[9] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_1354_ _0032_ VPWR _0033_ VGND W2END[4] Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q
+ sg13g2_o21ai_1
X_1285_ _1122_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _1121_ VPWR
+ VGND sg13g2_nand2b_1
X_1423_ _0100_ _0078_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 VPWR
+ VGND sg13g2_nand2b_1
XFILLER_48_180 VPWR VGND sg13g2_fill_2
X_3024_ FrameData[17] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_50_18 VPWR VGND sg13g2_fill_2
X_2808_ FrameData[25] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_2739_ FrameData[20] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_3_419 VPWR VGND sg13g2_fill_1
XFILLER_27_320 VPWR VGND sg13g2_fill_2
XFILLER_42_312 VPWR VGND sg13g2_fill_2
XFILLER_27_386 VPWR VGND sg13g2_fill_1
XFILLER_18_386 VPWR VGND sg13g2_fill_2
X_1972_ _0627_ VPWR _0629_ VGND _0532_ _0628_ sg13g2_o21ai_1
X_2524_ FrameData[29] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VPWR VGND sg13g2_dlhq_1
XFILLER_46_0 VPWR VGND sg13g2_fill_2
X_2455_ FrameData[24] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_1268_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q A D C E Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q
+ _1106_ VPWR VGND sg13g2_mux4_1
X_1406_ VGND VPWR _0083_ _0075_ _0074_ sg13g2_or2_1
X_1337_ _0016_ VPWR _0017_ VGND W2END[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ sg13g2_o21ai_1
X_2386_ _0982_ VPWR _0983_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q Inst_LUT4AB_switch_matrix.JN2BEG1
+ sg13g2_o21ai_1
XFILLER_28_128 VPWR VGND sg13g2_fill_2
X_3007_ FrameData[0] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1199_ VPWR _1040_ EE4END[3] VGND sg13g2_inv_1
XFILLER_15_323 VPWR VGND sg13g2_fill_1
XFILLER_51_72 VPWR VGND sg13g2_fill_1
X_2171_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VPWR _0815_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q
+ _0813_ sg13g2_o21ai_1
X_2240_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q VPWR _0876_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ _0873_ sg13g2_o21ai_1
XFILLER_33_153 VPWR VGND sg13g2_fill_2
X_1955_ Inst_LUT4AB_switch_matrix.JW2BEG6 _0611_ _0612_ _0604_ _0598_ VPWR VGND sg13g2_a22oi_1
X_1886_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q N1END[3] N2END[7] E1END[3] E2END[7]
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q _0546_ VPWR VGND sg13g2_mux4_1
X_2507_ FrameData[12] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VPWR VGND sg13g2_dlhq_1
X_2438_ FrameData[7] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_2369_ _0966_ _0617_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VPWR VGND sg13g2_nand2b_1
XFILLER_47_289 VPWR VGND sg13g2_fill_1
XFILLER_46_50 VPWR VGND sg13g2_fill_2
XFILLER_7_88 VPWR VGND sg13g2_fill_2
X_1671_ _0336_ VPWR _0339_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q _0338_ sg13g2_o21ai_1
X_1740_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q _1051_ _0405_ _0404_ sg13g2_a21oi_1
XFILLER_30_134 VPWR VGND sg13g2_fill_1
X_3272_ W2MID[0] W2BEGb[0] VPWR VGND sg13g2_buf_1
X_2154_ _0797_ VPWR _0798_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q _1052_ sg13g2_o21ai_1
X_2223_ _0858_ _0861_ _0862_ VPWR VGND sg13g2_nor2_1
X_2085_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q _0732_ _0735_ VPWR VGND sg13g2_nor2_1
X_2987_ FrameData[12] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1938_ E F Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q _0596_ VPWR VGND sg13g2_mux2_1
X_1869_ VPWR _0529_ _0528_ VGND sg13g2_inv_1
XFILLER_29_201 VPWR VGND sg13g2_fill_2
XFILLER_12_112 VPWR VGND sg13g2_fill_1
XFILLER_4_399 VPWR VGND sg13g2_fill_2
XFILLER_35_259 VPWR VGND sg13g2_fill_2
XFILLER_35_248 VPWR VGND sg13g2_fill_1
X_2910_ FrameData[31] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_2841_ FrameData[26] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_1723_ Inst_LUT4AB_switch_matrix.JN2BEG4 _0382_ _0388_ _0377_ _0370_ VPWR VGND sg13g2_a22oi_1
X_2772_ FrameData[21] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_1654_ _0323_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q W1END[2] VPWR VGND sg13g2_nand2b_1
X_1585_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ _0256_ VPWR VGND sg13g2_mux4_1
X_2206_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q E1END[3] W1END[3] A B Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q
+ _0847_ VPWR VGND sg13g2_mux4_1
X_3255_ Inst_LUT4AB_switch_matrix.SS4BEG0 SS4BEG[12] VPWR VGND sg13g2_buf_1
X_3186_ N4END[15] N4BEG[11] VPWR VGND sg13g2_buf_1
X_2137_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q F _0782_ VPWR VGND sg13g2_nor2b_1
X_2068_ _0719_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q W1END[0] VPWR VGND sg13g2_nand2b_1
X_1370_ _0047_ VPWR _0048_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q _0044_ sg13g2_o21ai_1
X_3040_ _1167_ VGND VPWR _0001_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop clknet_1_0__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_2824_ FrameData[9] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1706_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q _1051_ _0372_ _0371_ sg13g2_a21oi_1
X_1637_ _0304_ _0305_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit13.Q _0306_ VPWR VGND sg13g2_nand3_1
X_2755_ FrameData[4] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_2686_ FrameData[31] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_3238_ S4END[15] S4BEG[11] VPWR VGND sg13g2_buf_1
X_1499_ _0172_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q D VPWR VGND sg13g2_nand2b_1
X_1568_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q N2END[7] S2END[7] EE4END[2] W2END[7]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q _0239_ VPWR VGND sg13g2_mux4_1
X_3307_ Inst_LUT4AB_switch_matrix.WW4BEG3 WW4BEG[15] VPWR VGND sg13g2_buf_1
X_3169_ N2MID[2] N2BEGb[2] VPWR VGND sg13g2_buf_1
X_2540_ FrameData[13] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VPWR VGND sg13g2_dlhq_1
X_1422_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 _0083_ _0099_ VPWR
+ VGND sg13g2_nor2_1
X_2471_ FrameData[8] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_3023_ FrameData[16] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_1353_ _0032_ _1023_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q VPWR VGND sg13g2_nand2_1
X_1284_ _1120_ Ci Inst_LA_LUT4c_frame_config_dffesr.c_I0mux _1121_ VPWR VGND sg13g2_mux2_1
X_2738_ FrameData[19] FrameStrobe[9] Inst_LUT4AB_switch_matrix.DEBUG_select_LE_EN[0]
+ VPWR VGND sg13g2_dlhq_1
X_2807_ FrameData[24] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_2669_ FrameData[14] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_27_343 VPWR VGND sg13g2_fill_2
XFILLER_6_0 VPWR VGND sg13g2_fill_2
X_1971_ _0590_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0565_ _0628_ VPWR VGND sg13g2_mux4_1
X_2523_ FrameData[28] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VPWR VGND sg13g2_dlhq_1
XFILLER_39_0 VPWR VGND sg13g2_fill_1
X_2454_ FrameData[23] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_2385_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _1064_ _0982_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ sg13g2_a21oi_1
X_1405_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14 _0081_ _0082_ VPWR
+ VGND sg13g2_nor2_1
X_1198_ VPWR _1039_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VGND sg13g2_inv_1
X_1267_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q F G H Inst_LUT4AB_switch_matrix.M_AD
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q _1105_ VPWR VGND sg13g2_mux4_1
X_3006_ FrameData[31] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1336_ _0016_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q W6END[0] VPWR VGND sg13g2_nand2b_1
XFILLER_51_84 VPWR VGND sg13g2_fill_1
X_2170_ W2END[1] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q _0814_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_33_121 VPWR VGND sg13g2_fill_2
X_1954_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q _0609_ _0612_ VPWR VGND sg13g2_nor2_1
X_1885_ VGND VPWR _1044_ _0539_ _0545_ _0544_ sg13g2_a21oi_1
X_2368_ _0651_ VPWR Co VGND _0639_ _0652_ sg13g2_o21ai_1
X_2506_ FrameData[11] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VPWR VGND sg13g2_dlhq_1
X_2437_ FrameData[6] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_1319_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit8.Q _1154_ _1155_ VPWR VGND sg13g2_nor2_1
X_2299_ S1END[0] B Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q _0928_ VPWR VGND sg13g2_mux2_1
XFILLER_24_187 VPWR VGND sg13g2_decap_4
Xclkbuf_1_0__f_UserCLK clknet_0_UserCLK clknet_1_0__leaf_UserCLK VPWR VGND sg13g2_buf_8
X_1670_ _0337_ VPWR _0338_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q _0329_ sg13g2_o21ai_1
XFILLER_38_202 VPWR VGND sg13g2_fill_2
X_3271_ Inst_LUT4AB_switch_matrix.JW2BEG7 W2BEG[7] VPWR VGND sg13g2_buf_1
X_2222_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q VPWR _0861_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q
+ _0860_ sg13g2_o21ai_1
X_2153_ _0797_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q Inst_LUT4AB_switch_matrix.M_EF
+ VPWR VGND sg13g2_nand2_1
X_2084_ _0734_ _0733_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VPWR VGND sg13g2_nand2b_1
X_1937_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q Inst_LUT4AB_switch_matrix.M_EF
+ _0595_ _0594_ sg13g2_a21oi_1
X_2986_ FrameData[11] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1868_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit18.Q N2END[7] E2END[7] S2END[7] WW4END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit19.Q _0528_ VPWR VGND sg13g2_mux4_1
X_1799_ _0398_ VPWR _0462_ VGND _0204_ _0461_ sg13g2_o21ai_1
XFILLER_52_293 VPWR VGND sg13g2_fill_1
XFILLER_44_238 VPWR VGND sg13g2_fill_1
XFILLER_16_21 VPWR VGND sg13g2_fill_1
XFILLER_16_32 VPWR VGND sg13g2_fill_2
XFILLER_43_271 VPWR VGND sg13g2_fill_2
X_2771_ FrameData[20] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_422 VPWR VGND sg13g2_fill_2
X_2840_ FrameData[25] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1653_ _0322_ _0321_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VPWR VGND sg13g2_nand2b_1
X_1584_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q _0248_ _0255_ _0254_ sg13g2_a21oi_1
X_1722_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q _0387_ _0388_ VPWR VGND sg13g2_nor2_1
X_3185_ N4END[14] N4BEG[10] VPWR VGND sg13g2_buf_1
X_3254_ SS4END[15] SS4BEG[11] VPWR VGND sg13g2_buf_1
X_2205_ Inst_LUT4AB_switch_matrix.W6BEG1 _0846_ _0841_ VPWR VGND sg13g2_nand2b_1
XFILLER_41_219 VPWR VGND sg13g2_fill_2
X_2136_ _0780_ VPWR _0781_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q _1052_ sg13g2_o21ai_1
XFILLER_22_422 VPWR VGND sg13g2_fill_2
X_2067_ S1END[0] S1END[2] Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q _0718_ VPWR VGND
+ sg13g2_mux2_1
X_2969_ FrameData[26] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_1_304 VPWR VGND sg13g2_fill_2
XFILLER_27_20 VPWR VGND sg13g2_fill_2
XFILLER_40_252 VPWR VGND sg13g2_fill_1
XFILLER_23_219 VPWR VGND sg13g2_fill_1
X_2754_ FrameData[3] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_296 VPWR VGND sg13g2_fill_2
X_2823_ FrameData[8] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1705_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q F _0371_ VPWR VGND sg13g2_nor2_1
X_1636_ _0305_ S2MID[2] Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q VPWR VGND sg13g2_nand2b_1
X_1567_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q N4END[3] W2END[3] E2END[3] Inst_LUT4AB_switch_matrix.JN2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q _0238_ VPWR VGND sg13g2_mux4_1
X_3306_ Inst_LUT4AB_switch_matrix.WW4BEG2 WW4BEG[14] VPWR VGND sg13g2_buf_1
X_2685_ FrameData[30] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_3237_ S4END[14] S4BEG[10] VPWR VGND sg13g2_buf_1
X_3168_ N2MID[1] N2BEGb[1] VPWR VGND sg13g2_buf_1
XFILLER_39_385 VPWR VGND sg13g2_fill_1
X_2119_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q G _0765_ _0764_ sg13g2_a21oi_1
X_1498_ VPWR _0171_ _0170_ VGND sg13g2_inv_1
X_3099_ Inst_LUT4AB_switch_matrix.EE4BEG0 EE4BEG[12] VPWR VGND sg13g2_buf_1
X_1421_ _0073_ VPWR _0098_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0081_ sg13g2_o21ai_1
X_2470_ FrameData[7] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VPWR VGND sg13g2_dlhq_1
X_1352_ VGND VPWR _1022_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q _0031_ _0030_ sg13g2_a21oi_1
X_3022_ FrameData[15] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_1283_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit2.Q _1102_ _1103_ _1119_ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q
+ _1120_ VPWR VGND sg13g2_mux4_1
X_2737_ FrameData[18] FrameStrobe[9] Inst_LUT4AB_switch_matrix.DEBUG_select_LE_SR[0]
+ VPWR VGND sg13g2_dlhq_1
X_2668_ FrameData[13] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_2806_ FrameData[23] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1619_ N2END[3] E2END[3] Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q _0289_ VPWR VGND
+ sg13g2_mux2_1
X_2599_ FrameData[8] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_42_314 VPWR VGND sg13g2_fill_1
X_1970_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit4.Q _0617_ _0622_ _0626_ _0624_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit5.Q
+ _0627_ VPWR VGND sg13g2_mux4_1
XFILLER_18_388 VPWR VGND sg13g2_fill_1
X_2522_ FrameData[27] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VPWR VGND sg13g2_dlhq_1
X_1404_ _0081_ _0074_ _0075_ VPWR VGND sg13g2_nand2_1
X_1335_ S2END[2] S4END[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q _0015_ VPWR VGND
+ sg13g2_mux2_1
X_2453_ FrameData[22] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_2384_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0021_ _0981_ _0980_ sg13g2_a21oi_1
X_3005_ FrameData[30] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1266_ VPWR _1104_ _1103_ VGND sg13g2_inv_1
X_1197_ VPWR _1038_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q VGND sg13g2_inv_1
XFILLER_51_177 VPWR VGND sg13g2_fill_1
XFILLER_19_21 VPWR VGND sg13g2_fill_2
XFILLER_35_42 VPWR VGND sg13g2_fill_2
XFILLER_35_20 VPWR VGND sg13g2_fill_1
X_1953_ _0611_ _0610_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VPWR VGND sg13g2_nand2b_1
X_1884_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q VPWR _0544_ VGND _0542_ _0543_ sg13g2_o21ai_1
XFILLER_51_0 VPWR VGND sg13g2_fill_1
X_2505_ FrameData[10] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VPWR VGND sg13g2_dlhq_1
X_2367_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q C Inst_LUT4AB_switch_matrix.JW2BEG3
+ _0453_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q Inst_LUT4AB_switch_matrix.N1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1318_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q N2END[4] E1END[2] E2END[4] E6END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _1154_ VPWR VGND sg13g2_mux4_1
X_2436_ FrameData[5] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_2298_ _0926_ VPWR _0927_ VGND N1END[0] Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q
+ sg13g2_o21ai_1
X_1249_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _1051_ _1088_ _1087_ sg13g2_a21oi_1
XANTENNA_40 VPWR VGND EE4END[9] sg13g2_antennanp
XFILLER_38_225 VPWR VGND sg13g2_fill_1
X_2152_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q G _0796_ _0795_ sg13g2_a21oi_1
X_2221_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q _0308_ _0860_ _0859_
+ sg13g2_a21oi_1
X_3270_ Inst_LUT4AB_switch_matrix.JW2BEG6 W2BEG[6] VPWR VGND sg13g2_buf_1
X_2083_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q N1END[0] N2END[0] E1END[0] EE4END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q _0733_ VPWR VGND sg13g2_mux4_1
X_1936_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q VPWR _0594_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
+ _1052_ sg13g2_o21ai_1
X_1867_ VPWR _0527_ _0526_ VGND sg13g2_inv_1
X_2985_ FrameData[10] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1798_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _0395_ _0461_ VPWR VGND sg13g2_mux2_1
X_2419_ _1009_ Inst_LUT4AB_switch_matrix.DEBUG_select_LG_SR[0] _0985_ VPWR VGND sg13g2_nand2_1
XFILLER_4_346 VPWR VGND sg13g2_fill_1
X_1721_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0384_ _0387_ _0386_ sg13g2_a21oi_1
X_2770_ FrameData[19] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1652_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q N1END[2] N2END[6] E1END[2] E2END[6]
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q _0321_ VPWR VGND sg13g2_mux4_1
X_1583_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q VPWR _0254_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q
+ _0253_ sg13g2_o21ai_1
X_3184_ N4END[13] N4BEG[9] VPWR VGND sg13g2_buf_1
X_3253_ SS4END[14] SS4BEG[10] VPWR VGND sg13g2_buf_1
X_2135_ _0780_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q Inst_LUT4AB_switch_matrix.M_AH
+ VPWR VGND sg13g2_nand2_1
X_2204_ _0845_ VPWR _0846_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0842_ sg13g2_o21ai_1
X_2066_ _0717_ _0716_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VPWR VGND sg13g2_nand2b_1
X_1919_ _0577_ VPWR _0578_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0576_ sg13g2_o21ai_1
X_2899_ FrameData[20] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_2968_ FrameData[25] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_16_261 VPWR VGND sg13g2_fill_2
X_1704_ _0370_ _0369_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VPWR VGND sg13g2_nand2b_1
X_2753_ FrameData[2] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_2684_ FrameData[29] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_2822_ FrameData[7] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1635_ _0304_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q Inst_LUT4AB_switch_matrix.E2BEG5
+ VPWR VGND sg13g2_nand2_1
X_3305_ Inst_LUT4AB_switch_matrix.WW4BEG1 WW4BEG[13] VPWR VGND sg13g2_buf_1
X_1497_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q N2END[4] E2END[4] SS4END[2] W2END[4]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q _0170_ VPWR VGND sg13g2_mux4_1
X_1566_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit10.Q N2MID[7] E2MID[7] S2MID[7] W2MID[7]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit11.Q _0237_ VPWR VGND sg13g2_mux4_1
X_3236_ S4END[13] S4BEG[9] VPWR VGND sg13g2_buf_1
X_3167_ N2MID[0] N2BEGb[0] VPWR VGND sg13g2_buf_1
X_3098_ EE4END[15] EE4BEG[11] VPWR VGND sg13g2_buf_1
X_2118_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q F _0764_ VPWR VGND sg13g2_nor2b_1
X_2049_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VPWR _0701_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ _0700_ sg13g2_o21ai_1
XFILLER_13_89 VPWR VGND sg13g2_fill_2
XFILLER_13_220 VPWR VGND sg13g2_fill_2
X_1351_ S2END[4] Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q _0030_ VPWR VGND sg13g2_nor2_1
X_1420_ _0091_ _0096_ _0097_ VPWR VGND sg13g2_and2_1
XFILLER_36_356 VPWR VGND sg13g2_fill_2
X_3021_ FrameData[14] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_1282_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit27.Q N2END[6] SS4END[3] E2END[6] W2END[6]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit26.Q _1119_ VPWR VGND sg13g2_mux4_1
XFILLER_51_337 VPWR VGND sg13g2_fill_2
X_2805_ FrameData[22] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1618_ VGND VPWR _1030_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q _0288_ _0287_ sg13g2_a21oi_1
X_2736_ FrameData[17] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_2667_ FrameData[12] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_2598_ FrameData[7] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1549_ _0221_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q _0220_ VPWR VGND sg13g2_nand2_1
X_3219_ S2MID[0] S2BEGb[0] VPWR VGND sg13g2_buf_1
XFILLER_42_337 VPWR VGND sg13g2_fill_1
XFILLER_27_345 VPWR VGND sg13g2_fill_1
Xclkbuf_regs_0_UserCLK UserCLK UserCLK_regs VPWR VGND sg13g2_buf_8
XFILLER_33_359 VPWR VGND sg13g2_fill_1
X_2521_ FrameData[26] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VPWR VGND sg13g2_dlhq_1
X_1334_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0013_ _0014_ VPWR VGND sg13g2_nor2b_1
X_1403_ _0074_ _0075_ _0080_ VPWR VGND sg13g2_and2_1
X_1265_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit26.Q N2MID[7] E2MID[7] S2MID[7] W2MID[7]
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q _1103_ VPWR VGND sg13g2_mux4_1
X_2452_ FrameData[21] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_2383_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q VPWR _0980_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q
+ Inst_LUT4AB_switch_matrix.JS2BEG1 sg13g2_o21ai_1
X_3004_ FrameData[29] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1196_ VPWR _1037_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VGND sg13g2_inv_1
X_2719_ FrameData[0] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_10_68 VPWR VGND sg13g2_fill_1
XFILLER_33_123 VPWR VGND sg13g2_fill_1
XFILLER_18_186 VPWR VGND sg13g2_fill_2
X_1883_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VPWR _0543_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ _0540_ sg13g2_o21ai_1
X_1952_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q N1END[3] N2END[7] E1END[3] E2END[7]
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0610_ VPWR VGND sg13g2_mux4_1
XFILLER_44_0 VPWR VGND sg13g2_fill_2
X_2504_ FrameData[9] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VPWR VGND sg13g2_dlhq_1
X_2435_ FrameData[4] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
X_2366_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q D _0237_ Inst_LUT4AB_switch_matrix.JW2BEG0
+ _0248_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit21.Q Inst_LUT4AB_switch_matrix.N1BEG1
+ VPWR VGND sg13g2_mux4_1
X_1317_ _1152_ VPWR _1153_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _1150_ sg13g2_o21ai_1
X_1248_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q F _1087_ VPWR VGND sg13g2_nor2_1
X_2297_ VGND VPWR _1016_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q _0926_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
+ sg13g2_a21oi_1
X_1179_ VPWR _1020_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit0.Q VGND sg13g2_inv_1
XFILLER_12_307 VPWR VGND sg13g2_fill_1
XANTENNA_30 VPWR VGND S4END[0] sg13g2_antennanp
XFILLER_15_156 VPWR VGND sg13g2_fill_2
X_2151_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q F _0795_ VPWR VGND sg13g2_nor2b_1
X_2220_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q C _0859_ VPWR VGND sg13g2_nor2b_1
X_2082_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q _0729_ _0732_ _0731_ sg13g2_a21oi_1
X_2984_ FrameData[9] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1935_ VPWR _0593_ _0592_ VGND sg13g2_inv_1
X_1866_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit18.Q N4END[3] EE4END[0] S4END[3] Inst_LUT4AB_switch_matrix.JN2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit19.Q _0526_ VPWR VGND sg13g2_mux4_1
X_1797_ VGND VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 _0395_
+ _0460_ _0459_ sg13g2_a21oi_1
X_2418_ Inst_LUT4AB_switch_matrix.DEBUG_select_LG_EN[0] Inst_LG_LUT4c_frame_config_dffesr.LUT_flop
+ _1008_ VPWR VGND _0973_ sg13g2_nand3b_1
X_2349_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q S2END[0] W6END[1] S4END[3] C Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q
+ Inst_LUT4AB_switch_matrix.S4BEG2 VPWR VGND sg13g2_mux4_1
XFILLER_32_22 VPWR VGND sg13g2_fill_1
XFILLER_4_303 VPWR VGND sg13g2_fill_1
X_1720_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VPWR _0386_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ _0385_ sg13g2_o21ai_1
X_1651_ _0319_ VPWR _0320_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0317_ sg13g2_o21ai_1
X_3252_ SS4END[13] SS4BEG[9] VPWR VGND sg13g2_buf_1
X_1582_ _0252_ VPWR _0253_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q _0249_ sg13g2_o21ai_1
X_3183_ N4END[12] N4BEG[8] VPWR VGND sg13g2_buf_1
X_2134_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q B D C E Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ _0779_ VPWR VGND sg13g2_mux4_1
X_2065_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q N1END[0] NN4END[0] E1END[0] E2END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q _0716_ VPWR VGND sg13g2_mux4_1
X_2203_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit0.Q _0844_ _0845_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit1.Q
+ sg13g2_a21oi_1
X_2967_ FrameData[24] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1918_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0575_ _0577_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q
+ sg13g2_a21oi_1
X_2898_ FrameData[19] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1849_ _0510_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q W1END[3] VPWR VGND sg13g2_nand2b_1
XFILLER_27_55 VPWR VGND sg13g2_fill_1
X_2821_ FrameData[6] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1703_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q
+ _0369_ VPWR VGND sg13g2_mux4_1
X_2752_ FrameData[1] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1634_ N2MID[2] E2MID[2] Inst_LUT4AB_ConfigMem.Inst_frame7_bit12.Q _0303_ VPWR VGND
+ sg13g2_mux2_1
X_2683_ FrameData[28] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_3235_ S4END[12] S4BEG[8] VPWR VGND sg13g2_buf_1
X_1565_ _0232_ _0235_ _0236_ VPWR VGND sg13g2_nor2_1
X_3304_ Inst_LUT4AB_switch_matrix.WW4BEG0 WW4BEG[12] VPWR VGND sg13g2_buf_1
X_1496_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q NN4END[1] EE4END[1] S4END[1] Inst_LUT4AB_switch_matrix.JS2BEG2
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q _0169_ VPWR VGND sg13g2_mux4_1
X_3097_ EE4END[14] EE4BEG[10] VPWR VGND sg13g2_buf_1
X_2117_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q B D C E Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q
+ _0763_ VPWR VGND sg13g2_mux4_1
X_2048_ E F Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q _0700_ VPWR VGND sg13g2_mux2_1
X_3166_ Inst_LUT4AB_switch_matrix.JN2BEG7 N2BEG[7] VPWR VGND sg13g2_buf_1
XFILLER_22_276 VPWR VGND sg13g2_fill_1
XFILLER_38_43 VPWR VGND sg13g2_fill_1
X_1350_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0028_ _0029_ VPWR VGND sg13g2_nor2b_1
X_1281_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q NN4END[3] WW4END[0] S4END[3] Inst_LUT4AB_switch_matrix.JN2BEG1
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q _1118_ VPWR VGND sg13g2_mux4_1
X_3020_ FrameData[13] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_2804_ FrameData[21] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_2597_ FrameData[6] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1617_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q VPWR _0287_ VGND S2END[3] Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q
+ sg13g2_o21ai_1
X_2666_ FrameData[11] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_2735_ FrameData[16] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_1548_ _0219_ VPWR _0220_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0218_ sg13g2_o21ai_1
X_3149_ FrameStrobe[14] FrameStrobe_O[14] VPWR VGND sg13g2_buf_1
X_3218_ Inst_LUT4AB_switch_matrix.JS2BEG7 S2BEG[7] VPWR VGND sg13g2_buf_1
X_1479_ _1037_ VPWR _0153_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0152_ sg13g2_o21ai_1
XFILLER_24_89 VPWR VGND sg13g2_fill_2
Xclkbuf_0_UserCLK_regs UserCLK_regs clknet_0_UserCLK_regs VPWR VGND sg13g2_buf_8
XFILLER_2_423 VPWR VGND sg13g2_fill_1
XFILLER_2_401 VPWR VGND sg13g2_fill_1
X_2520_ FrameData[25] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VPWR VGND sg13g2_dlhq_1
X_1402_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10 _0078_ _0079_ VPWR
+ VGND sg13g2_nor2b_1
X_2451_ FrameData[20] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VPWR VGND sg13g2_dlhq_1
X_1333_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q N1END[0] E2END[2] N2END[2] E6END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q _0013_ VPWR VGND sg13g2_mux4_1
X_1264_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit26.Q N2MID[6] S2MID[6] W2MID[6] Inst_LUT4AB_switch_matrix.JN2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit27.Q _1102_ VPWR VGND sg13g2_mux4_1
X_3003_ FrameData[28] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_2382_ VPWR VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q
+ _0978_ _0976_ _0979_ _0977_ sg13g2_a221oi_1
X_1195_ VPWR _1036_ S4END[1] VGND sg13g2_inv_1
X_2718_ FrameData[31] FrameStrobe[10] Inst_LUT4AB_switch_matrix.DEBUG_select_LC_EN[0]
+ VPWR VGND sg13g2_dlhq_1
X_2649_ FrameData[26] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_15_349 VPWR VGND sg13g2_fill_2
XFILLER_4_0 VPWR VGND sg13g2_fill_2
X_1951_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0607_ _0609_ _0608_ sg13g2_a21oi_1
X_1882_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q Inst_LUT4AB_switch_matrix.M_AB
+ _0542_ _0541_ sg13g2_a21oi_1
X_2503_ FrameData[8] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VPWR VGND sg13g2_dlhq_1
XFILLER_37_0 VPWR VGND sg13g2_fill_2
X_2434_ FrameData[3] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_2365_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit23.Q E Inst_LUT4AB_switch_matrix.JW2BEG1
+ _0586_ _0623_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit22.Q Inst_LUT4AB_switch_matrix.N1BEG2
+ VPWR VGND sg13g2_mux4_1
X_1316_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _1151_ _1152_ _1024_ sg13g2_a21oi_1
X_1178_ VPWR _1019_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q VGND sg13g2_inv_1
XFILLER_2_92 VPWR VGND sg13g2_fill_1
X_1247_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q A B C E Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q
+ _1086_ VPWR VGND sg13g2_mux4_1
X_2296_ VPWR _0925_ _0924_ VGND sg13g2_inv_1
XANTENNA_20 VPWR VGND NN4END[7] sg13g2_antennanp
XANTENNA_31 VPWR VGND S4END[0] sg13g2_antennanp
XFILLER_43_422 VPWR VGND sg13g2_fill_2
XFILLER_11_374 VPWR VGND sg13g2_fill_1
X_2150_ _0794_ VPWR Inst_LUT4AB_switch_matrix.JS2BEG0 VGND _0785_ _0786_ sg13g2_o21ai_1
X_2081_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VPWR _0731_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ _0730_ sg13g2_o21ai_1
X_1934_ _0590_ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0565_ _0592_ VPWR VGND sg13g2_mux4_1
XFILLER_34_422 VPWR VGND sg13g2_fill_2
X_2983_ FrameData[8] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1796_ _0458_ _0202_ _0459_ VPWR VGND _0203_ sg13g2_nand3b_1
X_1865_ _0524_ VPWR _0525_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q _0521_ sg13g2_o21ai_1
X_2417_ _1007_ Inst_LUT4AB_switch_matrix.DEBUG_select_LG_EN[0] _0973_ VPWR VGND sg13g2_nand2b_1
X_2348_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q S2END[1] S4END[0] W6END[0] D Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q
+ Inst_LUT4AB_switch_matrix.S4BEG3 VPWR VGND sg13g2_mux4_1
X_2279_ VGND VPWR _1049_ _0909_ _0911_ _0910_ sg13g2_a21oi_1
XFILLER_16_68 VPWR VGND sg13g2_fill_1
XFILLER_25_422 VPWR VGND sg13g2_fill_2
XFILLER_52_285 VPWR VGND sg13g2_fill_1
X_1581_ _0250_ _0251_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit15.Q _0252_ VPWR VGND sg13g2_nand3_1
X_1650_ _0319_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q _0318_ VPWR VGND sg13g2_nand2b_1
X_3182_ N4END[11] N4BEG[7] VPWR VGND sg13g2_buf_1
X_3251_ SS4END[12] SS4BEG[8] VPWR VGND sg13g2_buf_1
X_2202_ VPWR _0844_ _0843_ VGND sg13g2_inv_1
X_2133_ _0771_ VPWR Inst_LUT4AB_switch_matrix.JW2BEG0 VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q
+ _0778_ sg13g2_o21ai_1
X_2064_ _0714_ VPWR _0715_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q _0713_ sg13g2_o21ai_1
X_2897_ FrameData[18] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_1917_ N1END[3] N2END[7] Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q _0576_ VPWR VGND
+ sg13g2_mux2_1
X_2966_ FrameData[23] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1848_ _0509_ _0508_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VPWR VGND sg13g2_nand2b_1
X_1779_ _0442_ VPWR _0443_ VGND S2END[5] Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ sg13g2_o21ai_1
X_2751_ FrameData[0] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_2820_ FrameData[5] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1633_ Inst_LUT4AB_switch_matrix.E2BEG5 _0296_ _0302_ _0294_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q
+ VPWR VGND sg13g2_a22oi_1
X_1564_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q _0233_ _0234_ _0235_ VPWR VGND sg13g2_nor3_1
X_2682_ FrameData[27] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_1702_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q _0365_ _0368_ _0367_
+ sg13g2_a21oi_1
X_3234_ S4END[11] S4BEG[7] VPWR VGND sg13g2_buf_1
X_3165_ Inst_LUT4AB_switch_matrix.JN2BEG6 N2BEG[6] VPWR VGND sg13g2_buf_1
X_1495_ Inst_LUT4AB_switch_matrix.JS2BEG2 _0168_ _1038_ _0161_ _0160_ VPWR VGND sg13g2_a22oi_1
X_3303_ WW4END[15] WW4BEG[11] VPWR VGND sg13g2_buf_1
X_2116_ A B _0669_ Inst_LUT4AB_switch_matrix.M_AB VPWR VGND sg13g2_mux2_1
X_3096_ EE4END[13] EE4BEG[9] VPWR VGND sg13g2_buf_1
X_2047_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q Inst_LUT4AB_switch_matrix.M_AD
+ _0699_ _0698_ sg13g2_a21oi_1
X_2949_ FrameData[6] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_45_369 VPWR VGND sg13g2_fill_2
XFILLER_13_222 VPWR VGND sg13g2_fill_1
X_1280_ Inst_LUT4AB_switch_matrix.JN2BEG1 _1110_ _1117_ _1108_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_51_339 VPWR VGND sg13g2_fill_1
X_2803_ FrameData[20] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_2734_ FrameData[15] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_2596_ FrameData[5] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1547_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0217_ _0219_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q
+ sg13g2_a21oi_1
X_2665_ FrameData[10] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1616_ _0285_ VPWR _0286_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q _0282_ sg13g2_o21ai_1
X_3148_ FrameStrobe[13] FrameStrobe_O[13] VPWR VGND sg13g2_buf_1
X_3217_ Inst_LUT4AB_switch_matrix.JS2BEG6 S2BEG[6] VPWR VGND sg13g2_buf_1
X_1478_ A B Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q _0152_ VPWR VGND sg13g2_mux2_1
X_3079_ E6END[6] E6BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_33_339 VPWR VGND sg13g2_fill_2
XFILLER_41_361 VPWR VGND sg13g2_fill_1
X_2450_ FrameData[19] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VPWR VGND sg13g2_dlhq_1
X_1401_ _0075_ _0074_ _0078_ VPWR VGND sg13g2_nor2b_1
X_2381_ _0390_ _0237_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _0978_ VPWR VGND sg13g2_mux2_1
X_1194_ VPWR _1035_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q VGND sg13g2_inv_1
X_1263_ _1094_ _1101_ Inst_LUT4AB_switch_matrix.JN2BEG3 VPWR VGND sg13g2_nor2_1
X_1332_ _0011_ VPWR _0012_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0010_ sg13g2_o21ai_1
X_3002_ FrameData[27] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_32_361 VPWR VGND sg13g2_fill_1
X_2717_ FrameData[30] FrameStrobe[10] Inst_LUT4AB_switch_matrix.DEBUG_select_LC_SR[0]
+ VPWR VGND sg13g2_dlhq_1
X_2579_ FrameData[20] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_2648_ FrameData[25] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1950_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VPWR _0608_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q
+ _0605_ sg13g2_o21ai_1
X_1881_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q VPWR _0541_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q
+ _1052_ sg13g2_o21ai_1
X_2502_ FrameData[7] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VPWR VGND sg13g2_dlhq_1
X_2433_ FrameData[2] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ VPWR VGND sg13g2_dlhq_1
X_1315_ W2END[4] WW4END[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q _1151_ VPWR VGND
+ sg13g2_mux2_1
X_2364_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit24.Q F _1159_ Inst_LUT4AB_switch_matrix.JW2BEG2
+ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit25.Q Inst_LUT4AB_switch_matrix.N1BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_52_423 VPWR VGND sg13g2_fill_1
XFILLER_52_401 VPWR VGND sg13g2_fill_1
X_1177_ VPWR _1018_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q VGND sg13g2_inv_1
X_1246_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q _1083_ _1084_ _1066_ _1065_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q
+ _1085_ VPWR VGND sg13g2_mux4_1
X_2295_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit28.Q C _0308_ _0586_ _0366_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q
+ _0924_ VPWR VGND sg13g2_mux4_1
XANTENNA_10 VPWR VGND N4END[14] sg13g2_antennanp
XANTENNA_21 VPWR VGND NN4END[8] sg13g2_antennanp
XANTENNA_32 VPWR VGND EE4END[11] sg13g2_antennanp
XFILLER_21_58 VPWR VGND sg13g2_fill_2
XFILLER_11_397 VPWR VGND sg13g2_fill_2
XFILLER_34_412 VPWR VGND sg13g2_fill_2
X_2080_ S1END[0] S2END[0] Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q _0730_ VPWR VGND
+ sg13g2_mux2_1
X_1933_ _0565_ _0590_ _0591_ VPWR VGND sg13g2_nor2_1
X_2982_ FrameData[7] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1795_ _0458_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0395_ VPWR
+ VGND sg13g2_nand2b_1
X_1864_ _0522_ _0523_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q _0524_ VPWR VGND sg13g2_nand3_1
X_2416_ Inst_LF_LUT4c_frame_config_dffesr.LUT_flop _1006_ _1004_ _0006_ VPWR VGND
+ sg13g2_mux2_1
X_2278_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q VPWR _0910_ VGND _1049_ _0908_ sg13g2_o21ai_1
X_2347_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q F Inst_LUT4AB_switch_matrix.JS2BEG3
+ _0453_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q Inst_LUT4AB_switch_matrix.W1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1229_ F G Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1069_ VPWR VGND sg13g2_mux2_1
XFILLER_16_423 VPWR VGND sg13g2_fill_1
X_1580_ _0251_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q W2END[5] VPWR VGND sg13g2_nand2_1
X_3250_ SS4END[11] SS4BEG[7] VPWR VGND sg13g2_buf_1
X_3181_ N4END[10] N4BEG[6] VPWR VGND sg13g2_buf_1
X_2132_ _0777_ VPWR _0778_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0772_ sg13g2_o21ai_1
X_2201_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q C D E F Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0843_ VPWR VGND sg13g2_mux4_1
X_2063_ _0714_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q _0712_ VPWR VGND sg13g2_nand2b_1
X_1916_ _0574_ VPWR _0575_ VGND E1END[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q
+ sg13g2_o21ai_1
X_1847_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q N1END[3] N2END[7] E1END[3] E2END[7]
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q _0508_ VPWR VGND sg13g2_mux4_1
X_2896_ FrameData[17] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_2965_ FrameData[22] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1778_ _0442_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q W1END[1] VPWR VGND sg13g2_nand2b_1
XFILLER_9_408 VPWR VGND sg13g2_fill_1
XFILLER_48_301 VPWR VGND sg13g2_fill_2
X_2750_ FrameData[31] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_2681_ FrameData[26] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_1701_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q VPWR _0367_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q
+ _0366_ sg13g2_o21ai_1
X_1632_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q _0301_ _0302_ VPWR VGND sg13g2_nor2_1
X_1563_ N2MID[6] Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q _0234_ VPWR VGND sg13g2_nor2_1
X_3302_ WW4END[14] WW4BEG[10] VPWR VGND sg13g2_buf_1
X_1494_ VGND VPWR _1037_ _0162_ _0168_ _0167_ sg13g2_a21oi_1
X_3233_ S4END[10] S4BEG[6] VPWR VGND sg13g2_buf_1
X_2115_ _0762_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0761_ Inst_LUT4AB_switch_matrix.M_AH
+ VPWR VGND sg13g2_a21o_1
X_3095_ EE4END[12] EE4BEG[8] VPWR VGND sg13g2_buf_1
X_3164_ Inst_LUT4AB_switch_matrix.JN2BEG5 N2BEG[5] VPWR VGND sg13g2_buf_1
X_2046_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q VPWR _0698_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
+ _1051_ sg13g2_o21ai_1
X_2879_ FrameData[0] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_2948_ FrameData[5] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_9_205 VPWR VGND sg13g2_fill_1
XFILLER_44_381 VPWR VGND sg13g2_fill_2
X_2802_ FrameData[19] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_2733_ FrameData[14] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_2664_ FrameData[9] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_2595_ FrameData[4] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_1546_ A B Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q _0218_ VPWR VGND sg13g2_mux2_1
X_1615_ _0285_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit13.Q _0284_ VPWR VGND sg13g2_nand2_1
X_1477_ _0150_ VPWR _0151_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q D sg13g2_o21ai_1
X_3147_ FrameStrobe[12] FrameStrobe_O[12] VPWR VGND sg13g2_buf_1
X_3078_ E6END[5] E6BEG[3] VPWR VGND sg13g2_buf_1
X_3216_ Inst_LUT4AB_switch_matrix.JS2BEG5 S2BEG[5] VPWR VGND sg13g2_buf_1
X_2029_ _0149_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ _0199_ _0683_ VPWR VGND sg13g2_mux4_1
XFILLER_10_259 VPWR VGND sg13g2_fill_2
XFILLER_41_395 VPWR VGND sg13g2_fill_1
X_1331_ _0011_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q _0009_ VPWR VGND sg13g2_nand2b_1
X_1400_ _0073_ VPWR _0077_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0076_ sg13g2_o21ai_1
X_2380_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q _1104_ _0977_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q
+ sg13g2_a21oi_1
X_1193_ VPWR _1034_ S2MID[4] VGND sg13g2_inv_1
X_1262_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q _1100_ _1101_ VPWR VGND sg13g2_nor2_1
X_3001_ FrameData[26] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_51_159 VPWR VGND sg13g2_fill_1
X_2647_ FrameData[24] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_2716_ FrameData[29] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1529_ _0201_ _0149_ _0199_ VPWR VGND sg13g2_nand2_1
X_2578_ FrameData[19] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_19_69 VPWR VGND sg13g2_fill_1
X_1880_ E F Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q _0540_ VPWR VGND sg13g2_mux2_1
X_2501_ FrameData[6] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VPWR VGND sg13g2_dlhq_1
X_2294_ _0917_ _0923_ Inst_LUT4AB_switch_matrix.EE4BEG3 VPWR VGND sg13g2_nor2_1
XFILLER_37_2 VPWR VGND sg13g2_fill_1
X_1314_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q S4END[0] _1150_ _1149_
+ sg13g2_a21oi_1
X_2432_ FrameData[1] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VPWR VGND sg13g2_dlhq_1
X_2363_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit26.Q N2END[2] N4END[1] E6END[1] E Inst_LUT4AB_ConfigMem.Inst_frame14_bit27.Q
+ Inst_LUT4AB_switch_matrix.N4BEG0 VPWR VGND sg13g2_mux4_1
Xclkbuf_1_1__f_UserCLK_regs clknet_0_UserCLK_regs clknet_1_1__leaf_UserCLK_regs VPWR
+ VGND sg13g2_buf_8
X_1176_ VPWR _1017_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q VGND sg13g2_inv_1
X_1245_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q N2MID[3] E2MID[3] S2MID[3] W2MID[3]
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q _1084_ VPWR VGND sg13g2_mux4_1
XANTENNA_22 VPWR VGND NN4END[9] sg13g2_antennanp
XANTENNA_33 VPWR VGND EE4END[13] sg13g2_antennanp
XANTENNA_11 VPWR VGND N4END[5] sg13g2_antennanp
X_1932_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit0.Q _0585_ _0586_ _0588_ _0587_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit1.Q
+ _0590_ VPWR VGND sg13g2_mux4_1
X_2981_ FrameData[6] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1863_ _0523_ W2MID[7] Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q VPWR VGND sg13g2_nand2_1
X_2415_ Inst_LF_LUT4c_frame_config_dffesr.c_reset_value _0496_ _1005_ _1006_ VPWR
+ VGND sg13g2_mux2_1
X_1794_ _0432_ _0456_ _0457_ VPWR VGND sg13g2_nor2b_1
X_2277_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q G H Inst_LUT4AB_switch_matrix.M_AD
+ Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q _0909_
+ VPWR VGND sg13g2_mux4_1
X_1228_ _1068_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _1067_ VPWR VGND sg13g2_nand2_1
X_2346_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q G _0237_ Inst_LUT4AB_switch_matrix.JS2BEG0
+ _0248_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit9.Q Inst_LUT4AB_switch_matrix.W1BEG1
+ VPWR VGND sg13g2_mux4_1
X_3180_ N4END[9] N4BEG[5] VPWR VGND sg13g2_buf_1
X_2131_ _0773_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q _0776_ _0777_ VPWR VGND sg13g2_a21o_1
X_2062_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q
+ _0713_ VPWR VGND sg13g2_mux4_1
X_2200_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit30.Q E1END[2] W1END[2] A B Inst_LUT4AB_ConfigMem.Inst_frame11_bit31.Q
+ _0842_ VPWR VGND sg13g2_mux4_1
X_2964_ FrameData[21] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_34_210 VPWR VGND sg13g2_fill_1
X_1846_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q _0506_ _0507_ VPWR VGND sg13g2_and2_1
X_1915_ _0574_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q E2END[7] VPWR VGND sg13g2_nand2b_1
X_1777_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q N1END[1] N2END[5] E1END[1] E2END[5]
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q _0441_ VPWR VGND sg13g2_mux4_1
X_2895_ FrameData[16] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_2329_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q _0953_ _0954_ VPWR VGND sg13g2_nor2_1
XFILLER_25_254 VPWR VGND sg13g2_fill_2
X_1631_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q _0299_ _0301_ _0300_ sg13g2_a21oi_1
X_2680_ FrameData[25] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1700_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q NN4END[3] S2END[6] E2END[6] W2END[6]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit2.Q _0366_ VPWR VGND sg13g2_mux4_1
X_3232_ S4END[9] S4BEG[5] VPWR VGND sg13g2_buf_1
X_1562_ E2MID[6] Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q _0233_ VPWR VGND sg13g2_nor2b_1
X_3301_ WW4END[13] WW4BEG[9] VPWR VGND sg13g2_buf_1
X_1493_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0164_ _0167_ _0166_ sg13g2_a21oi_1
X_2114_ _0758_ _0697_ _0752_ _0762_ VPWR VGND sg13g2_mux2_1
X_2045_ _0696_ _0697_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q Inst_LUT4AB_switch_matrix.M_AD
+ VPWR VGND sg13g2_mux2_1
X_3094_ EE4END[11] EE4BEG[7] VPWR VGND sg13g2_buf_1
X_3163_ Inst_LUT4AB_switch_matrix.JN2BEG4 N2BEG[4] VPWR VGND sg13g2_buf_1
X_2947_ FrameData[4] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_1829_ _0481_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ _0487_ _0491_ VPWR VGND sg13g2_mux4_1
X_2878_ FrameData[31] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_38_68 VPWR VGND sg13g2_fill_1
XFILLER_5_401 VPWR VGND sg13g2_fill_1
XFILLER_48_187 VPWR VGND sg13g2_fill_1
XFILLER_36_327 VPWR VGND sg13g2_fill_2
X_2801_ FrameData[18] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_2594_ FrameData[3] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_2732_ FrameData[13] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_2663_ FrameData[8] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1614_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q Inst_LUT4AB_switch_matrix.E2BEG3
+ _0284_ _0283_ sg13g2_a21oi_1
X_1545_ _0216_ VPWR _0217_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q C sg13g2_o21ai_1
X_3215_ Inst_LUT4AB_switch_matrix.JS2BEG4 S2BEG[4] VPWR VGND sg13g2_buf_1
X_1476_ _0150_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q E VPWR VGND sg13g2_nand2b_1
X_3146_ FrameStrobe[11] FrameStrobe_O[11] VPWR VGND sg13g2_buf_1
X_3077_ E6END[4] E6BEG[2] VPWR VGND sg13g2_buf_1
X_2028_ _0678_ _0679_ _0681_ _0682_ VPWR VGND sg13g2_nor3_1
XFILLER_50_352 VPWR VGND sg13g2_fill_2
XFILLER_26_360 VPWR VGND sg13g2_fill_2
XFILLER_5_297 VPWR VGND sg13g2_fill_2
X_1261_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit7.Q _1095_ _1096_ _1099_ _1097_ _1015_
+ _1100_ VPWR VGND sg13g2_mux4_1
X_1330_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q A D C E Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q
+ _0010_ VPWR VGND sg13g2_mux4_1
X_3000_ FrameData[25] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1192_ VPWR _1033_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q VGND sg13g2_inv_1
XFILLER_51_149 VPWR VGND sg13g2_fill_2
X_2577_ FrameData[18] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_2715_ FrameData[28] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_2646_ FrameData[23] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1459_ _0134_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q Inst_LUT4AB_switch_matrix.M_EF
+ VPWR VGND sg13g2_nand2b_1
X_1528_ _0149_ _0199_ _0200_ VPWR VGND sg13g2_nor2_1
X_3129_ FrameData[26] FrameData_O[26] VPWR VGND sg13g2_buf_1
XFILLER_50_193 VPWR VGND sg13g2_fill_2
XFILLER_41_193 VPWR VGND sg13g2_fill_1
X_2500_ FrameData[5] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VPWR VGND sg13g2_dlhq_1
X_2431_ FrameData[0] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VPWR VGND sg13g2_dlhq_1
X_2362_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q N2END[3] N4END[2] E6END[0] F Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q
+ Inst_LUT4AB_switch_matrix.N4BEG1 VPWR VGND sg13g2_mux4_1
X_2293_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q _0919_ _0923_ _0922_ sg13g2_a21oi_1
X_1313_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q S2END[4] _1149_ VPWR VGND sg13g2_nor2b_1
X_1244_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit28.Q E2MID[2] S2MID[2] W2MID[2] Inst_LUT4AB_switch_matrix.E2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q _1083_ VPWR VGND sg13g2_mux4_1
X_1175_ VPWR _1016_ E1END[0] VGND sg13g2_inv_1
XANTENNA_34 VPWR VGND N4END[11] sg13g2_antennanp
XANTENNA_12 VPWR VGND N4END[9] sg13g2_antennanp
XFILLER_32_160 VPWR VGND sg13g2_fill_2
XANTENNA_23 VPWR VGND S2END[1] sg13g2_antennanp
X_2629_ FrameData[6] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_15_105 VPWR VGND sg13g2_fill_1
XFILLER_15_138 VPWR VGND sg13g2_fill_1
XFILLER_19_400 VPWR VGND sg13g2_fill_2
X_2980_ FrameData[5] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1931_ VPWR _0589_ _0588_ VGND sg13g2_inv_1
X_1793_ _0455_ VPWR _0456_ VGND Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q _0452_
+ sg13g2_o21ai_1
X_1862_ _0522_ S2MID[7] Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q VPWR VGND sg13g2_nand2b_1
X_2414_ _1005_ Inst_LUT4AB_switch_matrix.DEBUG_select_LF_SR[0] _0985_ VPWR VGND sg13g2_nand2_1
XFILLER_35_0 VPWR VGND sg13g2_fill_1
X_2276_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q _1158_ _0196_ _0276_ _0556_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ _0908_ VPWR VGND sg13g2_mux4_1
X_1227_ H Inst_LUT4AB_switch_matrix.M_AH Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q
+ _1067_ VPWR VGND sg13g2_mux2_1
X_2345_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit11.Q H Inst_LUT4AB_switch_matrix.JS2BEG1
+ _0586_ _0623_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit10.Q Inst_LUT4AB_switch_matrix.W1BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_32_48 VPWR VGND sg13g2_fill_2
X_2130_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q VPWR _0776_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q
+ _0775_ sg13g2_o21ai_1
X_2061_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q E G F Inst_LUT4AB_switch_matrix.M_AB
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q _0712_ VPWR VGND sg13g2_mux4_1
X_2963_ FrameData[20] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_1914_ _0572_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q _0573_ VPWR VGND sg13g2_nor2b_1
X_1845_ _0505_ VPWR _0506_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q _0504_ sg13g2_o21ai_1
X_1776_ VGND VPWR _1039_ _0433_ _0440_ _0439_ sg13g2_a21oi_1
X_2894_ FrameData[15] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_2328_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q N1END[0] W1END[0] E1END[0] B Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q
+ _0953_ VPWR VGND sg13g2_mux4_1
X_2259_ _0887_ _0892_ Inst_LUT4AB_switch_matrix.SS4BEG1 VPWR VGND sg13g2_nor2_1
XFILLER_43_58 VPWR VGND sg13g2_fill_1
X_1630_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VPWR _0300_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q
+ _0297_ sg13g2_o21ai_1
X_3231_ S4END[8] S4BEG[4] VPWR VGND sg13g2_buf_1
X_3162_ Inst_LUT4AB_switch_matrix.JN2BEG3 N2BEG[3] VPWR VGND sg13g2_buf_1
X_1561_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q _0230_ _0232_ _0231_ sg13g2_a21oi_1
X_3300_ WW4END[12] WW4BEG[8] VPWR VGND sg13g2_buf_1
X_1492_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit4.Q VPWR _0166_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q
+ _0165_ sg13g2_o21ai_1
X_2113_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q _0759_ _0760_ _0761_ VPWR VGND
+ sg13g2_nor3_1
X_2044_ _0696_ Inst_LUT4AB_switch_matrix.M_AB _0693_ _0697_ VPWR VGND sg13g2_mux2_1
X_3093_ EE4END[10] EE4BEG[6] VPWR VGND sg13g2_buf_1
X_2877_ FrameData[30] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_2946_ FrameData[3] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1828_ _0490_ _0486_ _0487_ VPWR VGND sg13g2_nand2_1
X_1759_ _0421_ _0422_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q _0423_ VPWR VGND sg13g2_nand3_1
XFILLER_13_214 VPWR VGND sg13g2_fill_1
X_2731_ FrameData[12] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_2800_ FrameData[17] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_1544_ _0216_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q D VPWR VGND sg13g2_nand2b_1
X_2593_ FrameData[2] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_2662_ FrameData[7] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1613_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q S4END[2] _0283_ VPWR VGND sg13g2_nor2b_1
X_3145_ FrameStrobe[10] FrameStrobe_O[10] VPWR VGND sg13g2_buf_1
X_3214_ Inst_LUT4AB_switch_matrix.JS2BEG3 S2BEG[3] VPWR VGND sg13g2_buf_1
X_1475_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit2.Q _0147_ _0148_ _0130_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit3.Q
+ _0149_ VPWR VGND sg13g2_mux4_1
X_3076_ E6END[3] E6BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_24_49 VPWR VGND sg13g2_fill_2
X_2027_ _0680_ _0676_ _0681_ VPWR VGND sg13g2_nor2b_1
X_2929_ FrameData[18] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_45_103 VPWR VGND sg13g2_fill_2
X_1260_ VGND VPWR _1012_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _1099_ _1098_ sg13g2_a21oi_1
X_1191_ VPWR _1032_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VGND sg13g2_inv_1
X_2714_ FrameData[27] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_2576_ FrameData[17] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_2645_ FrameData[22] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1527_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit4.Q _0197_ _0198_ _0170_ _0169_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit5.Q
+ _0199_ VPWR VGND sg13g2_mux4_1
X_3128_ FrameData[25] FrameData_O[25] VPWR VGND sg13g2_buf_1
X_1458_ F G Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q _0133_ VPWR VGND sg13g2_mux2_1
X_1389_ _0067_ _0064_ _0066_ _0063_ _0062_ VPWR VGND sg13g2_a22oi_1
XFILLER_50_150 VPWR VGND sg13g2_fill_1
X_3059_ Inst_LUT4AB_switch_matrix.E2BEG0 E2BEG[0] VPWR VGND sg13g2_buf_1
X_2361_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q N2END[0] N4END[3] W6END[1] G Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q
+ Inst_LUT4AB_switch_matrix.N4BEG2 VPWR VGND sg13g2_mux4_1
X_2430_ FrameData[31] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VPWR VGND sg13g2_dlhq_1
X_2292_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q VPWR _0922_ VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ _0921_ sg13g2_o21ai_1
X_1312_ VPWR VGND _1147_ _1025_ _1145_ _1024_ _1148_ _1143_ sg13g2_a221oi_1
X_1243_ _1082_ _1019_ _1075_ Inst_LUT4AB_switch_matrix.E2BEG3 VPWR VGND sg13g2_a21o_1
X_1174_ VPWR _1015_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VGND sg13g2_inv_1
XANTENNA_13 VPWR VGND NN4END[11] sg13g2_antennanp
XANTENNA_35 VPWR VGND N4END[13] sg13g2_antennanp
XANTENNA_24 VPWR VGND S2END[1] sg13g2_antennanp
X_2559_ FrameData[0] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VPWR VGND sg13g2_dlhq_1
X_2628_ FrameData[5] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_28_423 VPWR VGND sg13g2_fill_1
XFILLER_19_423 VPWR VGND sg13g2_fill_1
X_1930_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit21.Q N2END[3] SS4END[0] E2END[3] W2END[3]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit20.Q _0588_ VPWR VGND sg13g2_mux4_1
X_1792_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame10_bit28.Q _0453_ _0455_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit29.Q
+ sg13g2_a21oi_1
X_1861_ N2MID[7] E2MID[7] Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q _0521_ VPWR VGND
+ sg13g2_mux2_1
X_2413_ _1004_ Inst_LUT4AB_switch_matrix.DEBUG_select_LF_EN[0] _0973_ VPWR VGND sg13g2_nand2b_1
X_2344_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit12.Q A _1159_ Inst_LUT4AB_switch_matrix.JS2BEG2
+ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit13.Q Inst_LUT4AB_switch_matrix.W1BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_28_0 VPWR VGND sg13g2_fill_1
XFILLER_52_212 VPWR VGND sg13g2_fill_2
X_2275_ VPWR VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q Inst_LUT4AB_ConfigMem.Inst_frame12_bit9.Q
+ _0906_ _0902_ _0907_ _0905_ sg13g2_a221oi_1
X_1226_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit29.Q NN4END[0] S2END[2] E2END[2] W2END[2]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit28.Q _1066_ VPWR VGND sg13g2_mux4_1
XFILLER_52_278 VPWR VGND sg13g2_fill_2
XFILLER_7_168 VPWR VGND sg13g2_fill_1
X_2060_ VGND VPWR _1046_ _0711_ Inst_LUT4AB_switch_matrix.JS2BEG7 _0704_ sg13g2_a21oi_1
X_1913_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0570_ _0572_ _0571_ sg13g2_a21oi_1
X_2962_ FrameData[19] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_2893_ FrameData[14] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_1844_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q _0503_ _0505_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q
+ sg13g2_a21oi_1
X_1775_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit13.Q VPWR _0439_ VGND _0437_ _0438_ sg13g2_o21ai_1
X_2258_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q _0888_ _0892_ _0891_
+ sg13g2_a21oi_1
X_2327_ VPWR _0952_ _0951_ VGND sg13g2_inv_1
X_1209_ VPWR _1050_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit7.Q VGND sg13g2_inv_1
X_2189_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q VPWR _0832_ VGND W2END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q
+ sg13g2_o21ai_1
X_1560_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit11.Q VPWR _0231_ VGND W2MID[6] Inst_LUT4AB_ConfigMem.Inst_frame7_bit10.Q
+ sg13g2_o21ai_1
X_3230_ S4END[7] S4BEG[3] VPWR VGND sg13g2_buf_1
X_2112_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0757_ _0760_ VPWR VGND sg13g2_nor2_1
X_3161_ Inst_LUT4AB_switch_matrix.JN2BEG2 N2BEG[2] VPWR VGND sg13g2_buf_1
X_1491_ S2END[3] S4END[3] Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q _0165_ VPWR VGND
+ sg13g2_mux2_1
X_2043_ C D _0695_ _0696_ VPWR VGND sg13g2_mux2_1
X_3092_ EE4END[9] EE4BEG[5] VPWR VGND sg13g2_buf_1
X_1827_ _0481_ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ _0487_ _0489_ VPWR VGND sg13g2_mux4_1
X_2876_ FrameData[29] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_2945_ FrameData[2] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_1689_ VGND VPWR _0356_ _0355_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q sg13g2_or2_1
X_1758_ _0422_ W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VPWR VGND sg13g2_nand2b_1
XFILLER_38_37 VPWR VGND sg13g2_fill_1
XFILLER_36_307 VPWR VGND sg13g2_fill_2
X_2730_ FrameData[11] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_2661_ FrameData[6] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1543_ _0211_ _0214_ _0215_ VPWR VGND sg13g2_nor2_1
X_2592_ FrameData[1] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1612_ NN4END[2] E2END[2] Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q _0282_ VPWR VGND
+ sg13g2_mux2_1
X_1474_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q N2MID[3] E2MID[3] S2MID[3] W2MID[3]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit5.Q _0148_ VPWR VGND sg13g2_mux4_1
X_3144_ FrameStrobe[9] FrameStrobe_O[9] VPWR VGND sg13g2_buf_1
X_3075_ E6END[2] E6BEG[0] VPWR VGND sg13g2_buf_1
X_3213_ Inst_LUT4AB_switch_matrix.JS2BEG2 S2BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_10_0 VPWR VGND sg13g2_fill_1
XFILLER_50_354 VPWR VGND sg13g2_fill_1
X_2026_ _0149_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0199_ _0680_ VPWR VGND sg13g2_mux4_1
X_2928_ FrameData[17] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_40_27 VPWR VGND sg13g2_fill_1
X_2859_ FrameData[12] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_5_222 VPWR VGND sg13g2_fill_2
XFILLER_30_82 VPWR VGND sg13g2_fill_2
X_1190_ VPWR _1031_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit4.Q VGND sg13g2_inv_1
XFILLER_36_115 VPWR VGND sg13g2_fill_2
X_2644_ FrameData[21] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_2713_ FrameData[26] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_2575_ FrameData[16] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_1457_ _0132_ _0131_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR VGND sg13g2_nand2b_1
X_1526_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit6.Q N2MID[5] E2MID[5] S2MID[5] W2MID[5]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit7.Q _0198_ VPWR VGND sg13g2_mux4_1
X_3127_ FrameData[24] FrameData_O[24] VPWR VGND sg13g2_buf_1
X_1388_ _1085_ _0065_ _0066_ VPWR VGND sg13g2_and2_1
X_3058_ Inst_LUT4AB_switch_matrix.E1BEG3 E1BEG[3] VPWR VGND sg13g2_buf_1
X_2009_ _0655_ _0664_ _0665_ VPWR VGND sg13g2_nor2b_1
X_2291_ _0920_ VPWR _0921_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q E sg13g2_o21ai_1
X_2360_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit1.Q N2END[1] W6END[0] N4END[0] H Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q
+ Inst_LUT4AB_switch_matrix.N4BEG3 VPWR VGND sg13g2_mux4_1
X_1311_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q _1146_ _1147_ _1024_ sg13g2_a21oi_1
X_1173_ VPWR _1014_ E6END[0] VGND sg13g2_inv_1
X_1242_ VGND VPWR _1080_ _1081_ _1082_ _1077_ sg13g2_a21oi_1
XANTENNA_36 VPWR VGND N4END[13] sg13g2_antennanp
XANTENNA_14 VPWR VGND NN4END[12] sg13g2_antennanp
XANTENNA_25 VPWR VGND S2END[1] sg13g2_antennanp
X_2627_ FrameData[4] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_2558_ FrameData[31] FrameStrobe[15] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VPWR VGND sg13g2_dlhq_1
X_1509_ _1035_ _0181_ _0182_ VPWR VGND sg13g2_nor2_1
X_2489_ FrameData[26] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ VPWR VGND sg13g2_dlhq_1
XFILLER_23_173 VPWR VGND sg13g2_fill_1
X_1860_ _0518_ VPWR _0520_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q _0519_ sg13g2_o21ai_1
X_1791_ VPWR _0454_ _0453_ VGND sg13g2_inv_1
X_2343_ _0963_ _0965_ Inst_LUT4AB_switch_matrix.NN4BEG0 VPWR VGND sg13g2_nor2_1
X_2274_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q C D E F Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ _0906_ VPWR VGND sg13g2_mux4_1
X_2412_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop _1003_ _1001_ _0005_ VPWR VGND
+ sg13g2_mux2_1
X_1225_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit28.Q EE4END[2] S4END[2] W2END[7] Inst_LUT4AB_switch_matrix.E2BEG1
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit29.Q _1065_ VPWR VGND sg13g2_mux4_1
X_1989_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux _0642_ _0644_ _0645_ VPWR VGND sg13g2_or3_1
XFILLER_43_235 VPWR VGND sg13g2_fill_2
X_1912_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VPWR _0571_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ _0568_ sg13g2_o21ai_1
X_2961_ FrameData[18] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_1843_ A B Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q _0504_ VPWR VGND sg13g2_mux2_1
X_2892_ FrameData[13] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_42_290 VPWR VGND sg13g2_fill_1
XFILLER_34_279 VPWR VGND sg13g2_fill_1
X_1774_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit12.Q VPWR _0438_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ _0435_ sg13g2_o21ai_1
X_1208_ VPWR _1049_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q VGND sg13g2_inv_1
X_2257_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q VPWR _0891_ VGND Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ _0890_ sg13g2_o21ai_1
X_2326_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q VPWR _0951_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q
+ _0950_ sg13g2_o21ai_1
X_2188_ _0830_ VPWR _0831_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q _0829_ sg13g2_o21ai_1
X_1490_ _0163_ VPWR _0164_ VGND W2END[3] Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q
+ sg13g2_o21ai_1
X_2111_ _0758_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0759_ VPWR VGND sg13g2_nor2b_1
X_2042_ _0694_ VPWR _0695_ VGND Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0693_
+ sg13g2_o21ai_1
X_3091_ EE4END[8] EE4BEG[4] VPWR VGND sg13g2_buf_1
X_3160_ Inst_LUT4AB_switch_matrix.JN2BEG1 N2BEG[1] VPWR VGND sg13g2_buf_1
X_1826_ _0486_ _0487_ _0488_ VPWR VGND sg13g2_nor2_1
X_2875_ FrameData[28] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_2944_ FrameData[1] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1688_ E6END[1] S2END[3] Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q _0355_ VPWR VGND
+ sg13g2_mux2_1
X_1757_ _0421_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q Inst_LUT4AB_switch_matrix.JW2BEG2
+ VPWR VGND sg13g2_nand2_1
X_2309_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit24.Q VPWR _0936_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q
+ _0935_ sg13g2_o21ai_1
XFILLER_38_49 VPWR VGND sg13g2_fill_2
X_3289_ W6END[11] W6BEG[9] VPWR VGND sg13g2_buf_1
XFILLER_28_60 VPWR VGND sg13g2_fill_1
X_1611_ VPWR _0281_ _0280_ VGND sg13g2_inv_1
X_2660_ FrameData[5] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1542_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VPWR _0214_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ _0213_ sg13g2_o21ai_1
X_2591_ FrameData[0] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_3212_ Inst_LUT4AB_switch_matrix.JS2BEG1 S2BEG[1] VPWR VGND sg13g2_buf_1
X_1473_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q N2MID[2] W2MID[2] E2MID[2] Inst_LUT4AB_switch_matrix.E2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q _0147_ VPWR VGND sg13g2_mux4_1
XFILLER_39_168 VPWR VGND sg13g2_fill_1
X_3143_ FrameStrobe[8] FrameStrobe_O[8] VPWR VGND sg13g2_buf_1
X_2025_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q _0452_ _0454_ _0430_ _0424_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q
+ _0679_ VPWR VGND sg13g2_mux4_1
X_3074_ E2MID[7] E2BEGb[7] VPWR VGND sg13g2_buf_1
XFILLER_50_377 VPWR VGND sg13g2_fill_2
X_2927_ FrameData[16] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_2858_ FrameData[11] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_2789_ FrameData[6] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1809_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q _0329_ _0471_ VPWR VGND sg13g2_nor2_1
XFILLER_45_105 VPWR VGND sg13g2_fill_1
XFILLER_41_377 VPWR VGND sg13g2_fill_1
X_2574_ FrameData[15] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.c_reset_value
+ VPWR VGND sg13g2_dlhq_1
X_2643_ FrameData[20] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_2712_ FrameData[25] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1456_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ _0131_ VPWR VGND sg13g2_mux4_1
X_1525_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q N2MID[4] E2MID[4] S2MID[4] Inst_LUT4AB_switch_matrix.JS2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q _0197_ VPWR VGND sg13g2_mux4_1
X_1387_ _0065_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _1121_ VPWR
+ VGND sg13g2_nand2b_1
X_2008_ _0645_ _0663_ _0640_ _0664_ VPWR VGND sg13g2_nand3_1
X_3126_ FrameData[23] FrameData_O[23] VPWR VGND sg13g2_buf_1
X_3057_ Inst_LUT4AB_switch_matrix.E1BEG2 E1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_27_116 VPWR VGND sg13g2_fill_2
XFILLER_23_399 VPWR VGND sg13g2_fill_2
XFILLER_41_141 VPWR VGND sg13g2_fill_1
X_2290_ _0920_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q _0276_ VPWR VGND sg13g2_nand2_1
X_1310_ H Inst_LUT4AB_switch_matrix.M_AD Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q
+ _1146_ VPWR VGND sg13g2_mux2_1
X_1241_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit7.Q _1078_ _1081_ _1018_ sg13g2_a21oi_1
X_1172_ VPWR _1013_ E1END[2] VGND sg13g2_inv_1
XANTENNA_15 VPWR VGND NN4END[14] sg13g2_antennanp
XANTENNA_37 VPWR VGND N4END[7] sg13g2_antennanp
XANTENNA_26 VPWR VGND S2END[1] sg13g2_antennanp
X_2557_ FrameData[30] FrameStrobe[15] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VPWR VGND sg13g2_dlhq_1
X_2626_ FrameData[3] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1508_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0179_ _0181_ _0180_ sg13g2_a21oi_1
X_1439_ _0115_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q E VPWR VGND sg13g2_nand2b_1
X_2488_ FrameData[25] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VPWR VGND sg13g2_dlhq_1
XFILLER_43_417 VPWR VGND sg13g2_fill_1
X_3109_ FrameData[6] FrameData_O[6] VPWR VGND sg13g2_buf_1
X_1790_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit8.Q N2MID[1] E2MID[1] S2MID[1] W2MID[1]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit9.Q _0453_ VPWR VGND sg13g2_mux4_1
X_2411_ Inst_LE_LUT4c_frame_config_dffesr.c_reset_value _0348_ _1002_ _1003_ VPWR
+ VGND sg13g2_mux2_1
X_2342_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q _0964_ _0965_ VPWR VGND sg13g2_nor2_1
X_2273_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q _0904_ _0905_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit8.Q
+ sg13g2_a21oi_1
X_1224_ VPWR _1064_ Inst_LUT4AB_switch_matrix.E2BEG1 VGND sg13g2_inv_1
XFILLER_52_236 VPWR VGND sg13g2_fill_2
X_1988_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q _0643_ _0644_ VPWR VGND sg13g2_nor2_1
X_2609_ FrameData[18] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_2960_ FrameData[17] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_19_233 VPWR VGND sg13g2_fill_1
X_1842_ _0502_ VPWR _0503_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q C sg13g2_o21ai_1
X_1911_ _0569_ VPWR _0570_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q H sg13g2_o21ai_1
X_2891_ FrameData[12] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_1773_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q Inst_LUT4AB_switch_matrix.M_AD
+ _0437_ _0436_ sg13g2_a21oi_1
X_1207_ VPWR _1048_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q VGND sg13g2_inv_1
X_2256_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q _1157_ _0890_ _0889_
+ sg13g2_a21oi_1
X_2187_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q _0827_ _0830_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q
+ sg13g2_a21oi_1
X_2325_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q _0308_ _0950_ _0949_ sg13g2_a21oi_1
XFILLER_25_236 VPWR VGND sg13g2_fill_1
X_2041_ _0694_ Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0669_ VPWR VGND sg13g2_nand2_1
X_2110_ _0757_ Inst_LUT4AB_switch_matrix.M_EF _0753_ _0758_ VPWR VGND sg13g2_mux2_1
X_3090_ EE4END[7] EE4BEG[3] VPWR VGND sg13g2_buf_1
X_2943_ FrameData[0] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1825_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q _0307_ _0309_ _0290_ _0286_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q
+ _0487_ VPWR VGND sg13g2_mux4_1
X_1756_ _0419_ VPWR _0420_ VGND _1012_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q sg13g2_o21ai_1
X_2874_ FrameData[27] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_30_272 VPWR VGND sg13g2_fill_2
X_2308_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q _1084_ _0935_ _0934_
+ sg13g2_a21oi_1
X_1687_ _0354_ _1031_ _0353_ VPWR VGND sg13g2_nand2_1
X_3288_ W6END[10] W6BEG[8] VPWR VGND sg13g2_buf_1
X_2239_ _0874_ VPWR _0875_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q _0556_ sg13g2_o21ai_1
XFILLER_36_309 VPWR VGND sg13g2_fill_1
XFILLER_29_350 VPWR VGND sg13g2_fill_1
XFILLER_44_342 VPWR VGND sg13g2_fill_1
X_1610_ _0255_ _0279_ _0280_ VPWR VGND sg13g2_nor2b_1
X_2590_ FrameData[31] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1472_ Inst_LUT4AB_switch_matrix.E2BEG4 _0140_ _0146_ _0138_ _0132_ VPWR VGND sg13g2_a22oi_1
X_3142_ FrameStrobe[7] FrameStrobe_O[7] VPWR VGND sg13g2_buf_1
X_1541_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q _1051_ _0213_ _0212_ sg13g2_a21oi_1
X_3211_ Inst_LUT4AB_switch_matrix.JS2BEG0 S2BEG[0] VPWR VGND sg13g2_buf_1
X_2024_ _0676_ _0677_ _0678_ VPWR VGND sg13g2_nor2_1
X_3073_ E2MID[6] E2BEGb[6] VPWR VGND sg13g2_buf_1
X_2926_ FrameData[15] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_2857_ FrameData[10] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1808_ _0470_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q _0334_ VPWR VGND sg13g2_nand2_1
X_1739_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q F _0404_ VPWR VGND sg13g2_nor2_1
X_2788_ FrameData[5] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_30_84 VPWR VGND sg13g2_fill_1
XFILLER_36_117 VPWR VGND sg13g2_fill_1
X_2711_ FrameData[24] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_2573_ FrameData[14] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_dlhq_1
X_1524_ _0193_ VPWR _0196_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q _0195_ sg13g2_o21ai_1
X_2642_ FrameData[19] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_3125_ FrameData[22] FrameData_O[22] VPWR VGND sg13g2_buf_1
X_1386_ _0064_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _1121_ VPWR
+ VGND sg13g2_nand2_1
X_1455_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q N2END[2] E2END[2] S2END[2] WW4END[2]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q _0130_ VPWR VGND sg13g2_mux4_1
X_2007_ VPWR _0663_ _0662_ VGND sg13g2_inv_1
XFILLER_35_18 VPWR VGND sg13g2_fill_2
X_3056_ Inst_LUT4AB_switch_matrix.E1BEG1 E1BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_50_186 VPWR VGND sg13g2_fill_2
X_2909_ FrameData[30] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_2_238 VPWR VGND sg13g2_fill_1
X_1240_ _1080_ _1017_ _1079_ VPWR VGND sg13g2_nand2_1
X_1171_ VPWR _1012_ N4END[0] VGND sg13g2_inv_1
XANTENNA_16 VPWR VGND NN4END[14] sg13g2_antennanp
XANTENNA_38 VPWR VGND NN4END[15] sg13g2_antennanp
XANTENNA_27 VPWR VGND S2END[1] sg13g2_antennanp
X_1507_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q VPWR _0180_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q
+ _0177_ sg13g2_o21ai_1
X_2556_ FrameData[29] FrameStrobe[15] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VPWR VGND sg13g2_dlhq_1
X_2625_ FrameData[2] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_2487_ FrameData[24] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VPWR VGND sg13g2_dlhq_1
X_1369_ _0045_ _0046_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q _0047_ VPWR VGND sg13g2_nand3_1
X_3108_ FrameData[5] FrameData_O[5] VPWR VGND sg13g2_buf_1
X_1438_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0111_ _0114_ _0113_ sg13g2_a21oi_1
X_3039_ _1168_ VGND VPWR _0000_ Inst_LH_LUT4c_frame_config_dffesr.LUT_flop clknet_1_1__leaf_UserCLK_regs
+ sg13g2_dfrbpq_1
X_2410_ _1002_ Inst_LUT4AB_switch_matrix.DEBUG_select_LE_SR[0] _0985_ VPWR VGND sg13g2_nand2_1
X_2341_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q N1END[2] W1END[2] E1END[2] F Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q
+ _0964_ VPWR VGND sg13g2_mux4_1
X_2272_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q B _0904_ _0903_ sg13g2_a21oi_1
X_1223_ _1056_ VPWR Inst_LUT4AB_switch_matrix.E2BEG1 VGND _1058_ _1063_ sg13g2_o21ai_1
X_1987_ _0520_ _0525_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0643_ VPWR VGND sg13g2_mux2_1
X_2539_ FrameData[12] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VPWR VGND sg13g2_dlhq_1
X_2608_ FrameData[17] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_11_167 VPWR VGND sg13g2_fill_1
X_2890_ FrameData[11] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1910_ _0569_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q Inst_LUT4AB_switch_matrix.M_AD
+ VPWR VGND sg13g2_nand2b_1
X_1841_ _0502_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q D VPWR VGND sg13g2_nand2b_1
X_1772_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q VPWR _0436_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q
+ _1052_ sg13g2_o21ai_1
X_2324_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q C _0949_ VPWR VGND sg13g2_nor2b_1
X_1206_ VPWR _1047_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit21.Q VGND sg13g2_inv_1
X_2255_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q _1052_ _0889_ VPWR VGND sg13g2_nor2_1
X_2186_ VGND VPWR N4END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q _0829_ _0828_
+ sg13g2_a21oi_1
XFILLER_4_119 VPWR VGND sg13g2_fill_1
X_2040_ _0693_ _0690_ _0692_ VPWR VGND sg13g2_nand2_1
X_2873_ FrameData[26] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_2942_ FrameData[31] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1686_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q N2END[3] N4END[3] E1END[1] E2END[3]
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q _0353_ VPWR VGND sg13g2_mux4_1
X_1824_ _0486_ _0485_ _0483_ VPWR VGND sg13g2_nand2b_1
X_1755_ _0419_ SS4END[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VPWR VGND sg13g2_nand2_1
X_2307_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q G _0934_ VPWR VGND sg13g2_nor2b_1
X_3287_ W6END[9] W6BEG[7] VPWR VGND sg13g2_buf_1
X_2238_ _0874_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q _0023_ VPWR VGND sg13g2_nand2_1
X_2169_ VGND VPWR S2END[1] Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q _0813_ _0812_
+ sg13g2_a21oi_1
XFILLER_44_72 VPWR VGND sg13g2_fill_2
XFILLER_12_262 VPWR VGND sg13g2_fill_2
X_1540_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q E _0212_ VPWR VGND sg13g2_nor2_1
X_1471_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q _0145_ _0146_ VPWR VGND sg13g2_nor2_1
X_3141_ FrameStrobe[6] FrameStrobe_O[6] VPWR VGND sg13g2_buf_1
X_3210_ Inst_LUT4AB_switch_matrix.S1BEG3 S1BEG[3] VPWR VGND sg13g2_buf_1
X_3072_ E2MID[5] E2BEGb[5] VPWR VGND sg13g2_buf_1
X_2023_ _0149_ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0199_ _0677_ VPWR VGND sg13g2_mux4_1
XFILLER_50_379 VPWR VGND sg13g2_fill_1
X_2925_ FrameData[14] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_1807_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q _0315_ _0469_ _0468_ sg13g2_a21oi_1
X_2856_ FrameData[9] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1669_ _0337_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q _0334_ VPWR VGND sg13g2_nand2_1
X_1738_ _0403_ _0402_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR VGND sg13g2_nand2b_1
X_2787_ FrameData[4] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_26_321 VPWR VGND sg13g2_fill_1
X_2710_ FrameData[23] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_2572_ FrameData[13] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_dlhq_1
X_2641_ FrameData[18] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_1454_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q N4END[2] E2END[2] W2END[7] Inst_LUT4AB_switch_matrix.E2BEG2
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q _0129_ VPWR VGND sg13g2_mux4_1
X_1523_ _0194_ VPWR _0195_ VGND _1021_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q sg13g2_o21ai_1
X_3124_ FrameData[21] FrameData_O[21] VPWR VGND sg13g2_buf_1
X_1385_ VGND VPWR Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _1121_
+ _0063_ _1085_ sg13g2_a21oi_1
X_3055_ Inst_LUT4AB_switch_matrix.E1BEG0 E1BEG[0] VPWR VGND sg13g2_buf_1
X_2006_ _0650_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0649_ _0662_ VPWR VGND sg13g2_mux4_1
X_2839_ FrameData[24] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_2908_ FrameData[29] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_18_107 VPWR VGND sg13g2_fill_1
XFILLER_22_390 VPWR VGND sg13g2_fill_1
XANTENNA_17 VPWR VGND NN4END[4] sg13g2_antennanp
X_2624_ FrameData[1] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
XANTENNA_39 VPWR VGND EE4END[12] sg13g2_antennanp
XANTENNA_28 VPWR VGND S2END[1] sg13g2_antennanp
X_2555_ FrameData[28] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.c_reset_value
+ VPWR VGND sg13g2_dlhq_1
X_1506_ _0178_ VPWR _0179_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q H sg13g2_o21ai_1
X_2486_ FrameData[23] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VPWR VGND sg13g2_dlhq_1
X_1437_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VPWR _0113_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ _0112_ sg13g2_o21ai_1
X_3107_ FrameData[4] FrameData_O[4] VPWR VGND sg13g2_buf_1
X_3038_ FrameData[31] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1299_ _1136_ _1135_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q VPWR VGND sg13g2_nand2b_1
X_1368_ _0046_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q W2MID[1] VPWR VGND sg13g2_nand2_1
X_2340_ _0959_ _0962_ _0963_ VPWR VGND sg13g2_nor2_1
X_2271_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q A _0903_ VPWR VGND sg13g2_nor2b_1
X_1222_ _1062_ _1060_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit1.Q _1063_ VPWR VGND sg13g2_a21o_1
XFILLER_52_238 VPWR VGND sg13g2_fill_1
X_1986_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q _0527_ _0642_ _0641_ sg13g2_a21oi_1
X_2607_ FrameData[16] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_2538_ FrameData[11] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VPWR VGND sg13g2_dlhq_1
X_2469_ FrameData[6] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8
+ VPWR VGND sg13g2_dlhq_1
XFILLER_47_72 VPWR VGND sg13g2_fill_1
XFILLER_19_268 VPWR VGND sg13g2_fill_2
X_1840_ VGND VPWR _0501_ _0500_ _0498_ sg13g2_or2_1
XFILLER_30_400 VPWR VGND sg13g2_fill_1
XFILLER_30_422 VPWR VGND sg13g2_fill_2
X_1771_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q _1051_ _0435_ _0434_ sg13g2_a21oi_1
X_2254_ _0197_ _0316_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q _0888_ VPWR VGND
+ sg13g2_mux2_1
X_2323_ _0946_ _0947_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q _0948_ VPWR VGND sg13g2_nand3_1
X_2185_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q N2END[1] _0828_ VPWR VGND sg13g2_nor2b_1
X_1205_ VPWR _1046_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit25.Q VGND sg13g2_inv_1
X_1969_ VPWR _0626_ _0625_ VGND sg13g2_inv_1
XFILLER_33_74 VPWR VGND sg13g2_fill_1
X_1823_ _0484_ VPWR _0485_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q _0276_ sg13g2_o21ai_1
X_2872_ FrameData[25] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_2941_ FrameData[30] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1685_ _0351_ VPWR _0352_ VGND _1031_ _0350_ sg13g2_o21ai_1
X_1754_ Inst_LUT4AB_switch_matrix.JW2BEG2 _0417_ _0418_ _0410_ _0403_ VPWR VGND sg13g2_a22oi_1
XFILLER_38_352 VPWR VGND sg13g2_fill_1
X_2306_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q _0529_ _0933_ _0932_
+ sg13g2_a21oi_1
X_3286_ W6END[8] W6BEG[6] VPWR VGND sg13g2_buf_1
X_2237_ _0872_ VPWR _0873_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q E sg13g2_o21ai_1
X_2168_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q E6END[1] _0812_ VPWR VGND sg13g2_nor2b_1
X_2099_ Inst_LUT4AB_switch_matrix.E2BEG7 _0741_ _0747_ _0739_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q
+ VPWR VGND sg13g2_a22oi_1
XFILLER_0_145 VPWR VGND sg13g2_fill_2
XFILLER_8_234 VPWR VGND sg13g2_fill_2
X_1470_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q _0142_ _0145_ _0144_ sg13g2_a21oi_1
X_3140_ FrameStrobe[5] FrameStrobe_O[5] VPWR VGND sg13g2_buf_1
X_3071_ E2MID[4] E2BEGb[4] VPWR VGND sg13g2_buf_1
X_2022_ _0676_ _0672_ _0675_ _0208_ Inst_LD_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_a22oi_1
X_2924_ FrameData[13] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_2786_ FrameData[3] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_2855_ FrameData[8] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1806_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q _0316_ _0468_ VPWR VGND sg13g2_nor2_1
X_1599_ _0269_ VPWR _0270_ VGND W1END[0] Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ sg13g2_o21ai_1
X_1668_ _0335_ VPWR _0336_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q _0316_ sg13g2_o21ai_1
X_1737_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q A B D E Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q
+ _0402_ VPWR VGND sg13g2_mux4_1
X_3269_ Inst_LUT4AB_switch_matrix.JW2BEG5 W2BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_5_204 VPWR VGND sg13g2_fill_1
XFILLER_39_95 VPWR VGND sg13g2_fill_2
XFILLER_39_62 VPWR VGND sg13g2_fill_1
XFILLER_36_108 VPWR VGND sg13g2_fill_2
X_2640_ FrameData[17] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_2571_ FrameData[12] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_1453_ VGND VPWR _0122_ _0128_ Inst_LUT4AB_switch_matrix.E2BEG2 _0120_ sg13g2_a21oi_1
X_1522_ _0194_ E2MID[4] Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q VPWR VGND sg13g2_nand2_1
X_2005_ _0645_ _0640_ _0660_ _0661_ VPWR VGND sg13g2_a21o_1
X_3123_ FrameData[20] FrameData_O[20] VPWR VGND sg13g2_buf_1
X_3054_ VPWR VGND _1170_ sg13g2_tiehi
X_1384_ _0062_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _1121_ VPWR
+ VGND sg13g2_nand2b_1
XFILLER_50_111 VPWR VGND sg13g2_fill_1
XFILLER_35_141 VPWR VGND sg13g2_fill_2
X_2907_ FrameData[28] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_2769_ FrameData[18] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_2838_ FrameData[23] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_18_119 VPWR VGND sg13g2_fill_2
XFILLER_26_141 VPWR VGND sg13g2_fill_2
XFILLER_26_174 VPWR VGND sg13g2_fill_2
XFILLER_25_86 VPWR VGND sg13g2_fill_2
XFILLER_2_57 VPWR VGND sg13g2_fill_1
XANTENNA_18 VPWR VGND NN4END[5] sg13g2_antennanp
XFILLER_32_100 VPWR VGND sg13g2_fill_2
XANTENNA_29 VPWR VGND S4END[0] sg13g2_antennanp
X_2554_ FrameData[27] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_dlhq_1
X_2623_ FrameData[0] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_49_0 VPWR VGND sg13g2_fill_1
X_1505_ _0178_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q Inst_LUT4AB_switch_matrix.M_AH
+ VPWR VGND sg13g2_nand2b_1
X_1367_ _0045_ S2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q VPWR VGND sg13g2_nand2b_1
X_2485_ FrameData[22] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VPWR VGND sg13g2_dlhq_1
X_1436_ F G Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q _0112_ VPWR VGND sg13g2_mux2_1
X_3106_ FrameData[3] FrameData_O[3] VPWR VGND sg13g2_buf_1
X_3037_ FrameData[30] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1298_ S4END[2] SS4END[2] Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q _1135_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_14_188 VPWR VGND sg13g2_fill_1
X_2270_ _0901_ VPWR _0902_ VGND _1013_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q sg13g2_o21ai_1
X_1221_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit31.Q _1061_ _1062_ _1020_ sg13g2_a21oi_1
X_1985_ Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q VPWR _0641_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit8.Q
+ _0528_ sg13g2_o21ai_1
X_2537_ FrameData[10] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VPWR VGND sg13g2_dlhq_1
X_2606_ FrameData[15] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_1419_ _0073_ _0092_ _0093_ _0095_ _0096_ VPWR VGND sg13g2_or4_1
X_2399_ Inst_LB_LUT4c_frame_config_dffesr.c_reset_value _0109_ _0993_ _0994_ VPWR
+ VGND sg13g2_mux2_1
X_2468_ FrameData[5] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_283 VPWR VGND sg13g2_fill_1
X_1770_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q F _0434_ VPWR VGND sg13g2_nor2_1
XFILLER_6_195 VPWR VGND sg13g2_fill_1
X_2253_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit31.Q _0886_ _0887_ VPWR VGND sg13g2_nor2_1
X_2184_ E1END[3] E2END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit26.Q _0827_ VPWR VGND
+ sg13g2_mux2_1
X_1204_ VPWR _1045_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VGND sg13g2_inv_1
X_2322_ _0947_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q _0130_ VPWR VGND sg13g2_nand2b_1
X_1899_ _0558_ S2MID[5] Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q VPWR VGND sg13g2_nand2b_1
X_1968_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit25.Q N2END[1] S2END[1] EE4END[3] W2END[1]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q _0625_ VPWR VGND sg13g2_mux4_1
X_2940_ FrameData[29] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1822_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q _0277_ _0484_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q
+ sg13g2_a21oi_1
X_2871_ FrameData[24] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1753_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit5.Q _0415_ _0418_ VPWR VGND sg13g2_nor2_1
XFILLER_30_220 VPWR VGND sg13g2_fill_2
X_1684_ _0351_ _1031_ _0349_ VPWR VGND sg13g2_nand2b_1
XFILLER_31_0 VPWR VGND sg13g2_fill_1
X_2305_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit23.Q VPWR _0932_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit22.Q
+ _0148_ sg13g2_o21ai_1
X_3285_ W6END[7] W6BEG[5] VPWR VGND sg13g2_buf_1
X_2167_ _0810_ VPWR _0811_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0809_ sg13g2_o21ai_1
X_2236_ _0872_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q _0276_ VPWR VGND sg13g2_nand2_1
XFILLER_21_220 VPWR VGND sg13g2_fill_1
X_2098_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit25.Q _0746_ _0747_ VPWR VGND sg13g2_nor2_1
X_3070_ E2MID[3] E2BEGb[3] VPWR VGND sg13g2_buf_1
X_2021_ Inst_LD_LUT4c_frame_config_dffesr.c_I0mux _0674_ _0675_ VPWR VGND sg13g2_nor2b_1
X_2923_ FrameData[12] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_2785_ FrameData[2] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_1805_ _0467_ Inst_LC_LUT4c_frame_config_dffesr.LUT_flop Inst_LC_LUT4c_frame_config_dffesr.c_out_mux
+ C VPWR VGND sg13g2_mux2_1
X_2854_ FrameData[7] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1736_ VGND VPWR Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 _0395_
+ _0401_ _0400_ sg13g2_a21oi_1
X_1598_ _0269_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q W1END[2] VPWR VGND sg13g2_nand2b_1
X_1667_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit16.Q _0315_ _0335_ _1043_ sg13g2_a21oi_1
X_3199_ NN4END[12] NN4BEG[8] VPWR VGND sg13g2_buf_1
XFILLER_38_183 VPWR VGND sg13g2_fill_2
X_2219_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q _0171_ _0858_ _0857_
+ sg13g2_a21oi_1
X_3268_ Inst_LUT4AB_switch_matrix.JW2BEG4 W2BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_26_389 VPWR VGND sg13g2_fill_1
XFILLER_53_186 VPWR VGND sg13g2_fill_1
XFILLER_41_337 VPWR VGND sg13g2_fill_2
X_2570_ FrameData[11] FrameStrobe[14] Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_3122_ FrameData[19] FrameData_O[19] VPWR VGND sg13g2_buf_1
X_1383_ _0061_ _0060_ _1160_ VPWR VGND sg13g2_nand2b_1
X_1452_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit5.Q _0127_ _0128_ VPWR VGND sg13g2_nor2_1
X_1521_ Inst_LUT4AB_switch_matrix.JS2BEG4 Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q
+ _0192_ _0193_ VPWR VGND sg13g2_a21o_1
X_2004_ _0650_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ _0649_ _0660_ VPWR VGND sg13g2_mux4_1
X_3053_ VPWR VGND _1169_ sg13g2_tiehi
X_2906_ FrameData[27] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_23_315 VPWR VGND sg13g2_fill_1
X_2768_ FrameData[17] FrameStrobe[8] Inst_LUT4AB_switch_matrix.DEBUG_select_LH_EN[0]
+ VPWR VGND sg13g2_dlhq_1
X_1719_ S1END[1] S2END[5] Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q _0385_ VPWR VGND
+ sg13g2_mux2_1
X_2837_ FrameData[22] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_2699_ FrameData[12] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_14_337 VPWR VGND sg13g2_fill_2
XFILLER_41_97 VPWR VGND sg13g2_fill_1
XFILLER_41_75 VPWR VGND sg13g2_fill_2
XFILLER_1_285 VPWR VGND sg13g2_fill_2
XFILLER_9_0 VPWR VGND sg13g2_fill_1
XFILLER_17_131 VPWR VGND sg13g2_fill_1
XANTENNA_19 VPWR VGND NN4END[6] sg13g2_antennanp
X_2553_ FrameData[26] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_dlhq_1
X_1504_ F G Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q _0177_ VPWR VGND sg13g2_mux2_1
X_2622_ FrameData[31] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_3105_ FrameData[2] FrameData_O[2] VPWR VGND sg13g2_buf_1
X_1366_ N2MID[1] E2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q _0044_ VPWR VGND
+ sg13g2_mux2_1
X_1435_ _0110_ VPWR _0111_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q H sg13g2_o21ai_1
X_2484_ FrameData[21] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VPWR VGND sg13g2_dlhq_1
X_3036_ FrameData[29] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1297_ VPWR _1134_ _1133_ VGND sg13g2_inv_1
XFILLER_6_344 VPWR VGND sg13g2_fill_1
X_1220_ W2END[2] WW4END[3] Inst_LUT4AB_ConfigMem.Inst_frame4_bit30.Q _1061_ VPWR VGND
+ sg13g2_mux2_1
X_1984_ Inst_LH_LUT4c_frame_config_dffesr.c_I0mux VPWR _0640_ VGND _0591_ _0638_ sg13g2_o21ai_1
X_2536_ FrameData[9] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.c_reset_value
+ VPWR VGND sg13g2_dlhq_1
X_2605_ FrameData[14] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_2467_ FrameData[4] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VPWR VGND sg13g2_dlhq_1
X_1349_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q N1END[2] E2END[4] N2END[4] E6END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q _0028_ VPWR VGND sg13g2_mux4_1
X_1418_ _0094_ VPWR _0095_ VGND Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ _0083_ sg13g2_o21ai_1
X_2398_ _0993_ Inst_LUT4AB_switch_matrix.DEBUG_select_LB_SR[0] _0985_ VPWR VGND sg13g2_nand2_1
XFILLER_28_215 VPWR VGND sg13g2_fill_2
X_3019_ FrameData[12] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_3_325 VPWR VGND sg13g2_fill_1
X_2321_ VGND VPWR _0946_ _0586_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit8.Q sg13g2_or2_1
X_1203_ VPWR _1044_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit20.Q VGND sg13g2_inv_1
X_2252_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit29.Q N1END[3] E1END[3] W1END[3] A Inst_LUT4AB_ConfigMem.Inst_frame12_bit30.Q
+ _0886_ VPWR VGND sg13g2_mux4_1
X_2183_ _0825_ VPWR _0826_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q _0818_ sg13g2_o21ai_1
X_1898_ N2MID[5] E2MID[5] Inst_LUT4AB_ConfigMem.Inst_frame6_bit22.Q _0557_ VPWR VGND
+ sg13g2_mux2_1
X_1967_ VPWR _0624_ _0623_ VGND sg13g2_inv_1
X_2519_ FrameData[24] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VPWR VGND sg13g2_dlhq_1
X_2870_ FrameData[23] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_15_240 VPWR VGND sg13g2_fill_1
X_1821_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q _0248_ _0483_ _0482_ sg13g2_a21oi_1
X_1683_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q F G H Inst_LUT4AB_switch_matrix.M_AH
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q _0350_ VPWR VGND sg13g2_mux4_1
X_1752_ _0417_ _0416_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR VGND sg13g2_nand2b_1
X_2304_ _0931_ _0930_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit27.Q Inst_LUT4AB_switch_matrix.EE4BEG1
+ VPWR VGND sg13g2_mux2_1
X_3284_ W6END[6] W6BEG[4] VPWR VGND sg13g2_buf_1
XFILLER_24_0 VPWR VGND sg13g2_fill_2
XFILLER_38_387 VPWR VGND sg13g2_fill_2
X_2166_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0807_ _0810_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q
+ sg13g2_a21oi_1
X_2235_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit5.Q _0870_ _0871_ VPWR VGND sg13g2_nor2_1
X_2097_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q _0743_ _0746_ _0745_ sg13g2_a21oi_1
X_2999_ FrameData[24] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_29_321 VPWR VGND sg13g2_fill_2
XFILLER_8_258 VPWR VGND sg13g2_fill_2
XFILLER_12_243 VPWR VGND sg13g2_fill_2
XFILLER_5_47 VPWR VGND sg13g2_fill_1
X_2020_ _0673_ VPWR _0674_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit0.Q _0389_ sg13g2_o21ai_1
X_2922_ FrameData[11] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_2853_ FrameData[6] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_2784_ FrameData[1] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1666_ _0333_ VPWR _0334_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q _0330_ sg13g2_o21ai_1
X_1735_ _0203_ _0399_ _0400_ VPWR VGND _0202_ sg13g2_nand3b_1
X_1804_ _0466_ _0457_ _0463_ _0467_ VPWR VGND sg13g2_a21o_1
X_1597_ _0265_ _0267_ _0268_ VPWR VGND sg13g2_nor2_1
X_3267_ Inst_LUT4AB_switch_matrix.JW2BEG3 W2BEG[3] VPWR VGND sg13g2_buf_1
X_3198_ NN4END[11] NN4BEG[7] VPWR VGND sg13g2_buf_1
X_2149_ _0793_ VPWR _0794_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0787_ sg13g2_o21ai_1
X_2218_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q VPWR _0857_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q
+ _0586_ sg13g2_o21ai_1
XFILLER_30_11 VPWR VGND sg13g2_fill_2
XFILLER_1_423 VPWR VGND sg13g2_fill_1
XFILLER_39_97 VPWR VGND sg13g2_fill_1
X_1520_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit7.Q VPWR _0192_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit6.Q
+ _1034_ sg13g2_o21ai_1
X_3121_ FrameData[18] FrameData_O[18] VPWR VGND sg13g2_buf_1
X_1382_ _0059_ _0058_ _1085_ _0060_ VPWR VGND sg13g2_mux2_1
X_1451_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q _0124_ _0127_ _0126_ sg13g2_a21oi_1
X_3052_ VPWR VGND _1168_ sg13g2_tiehi
X_2003_ _0659_ _0654_ _0655_ _0658_ VPWR VGND sg13g2_and3_1
XFILLER_50_146 VPWR VGND sg13g2_fill_1
X_2905_ FrameData[26] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_2836_ FrameData[21] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_2767_ FrameData[16] FrameStrobe[8] Inst_LUT4AB_switch_matrix.DEBUG_select_LH_SR[0]
+ VPWR VGND sg13g2_dlhq_1
X_1718_ _0383_ VPWR _0384_ VGND W1END[1] Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q
+ sg13g2_o21ai_1
X_1649_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q E G H Inst_LUT4AB_switch_matrix.M_AH
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q _0318_ VPWR VGND sg13g2_mux4_1
X_2698_ FrameData[11] FrameStrobe[10] Inst_LUT4AB_switch_matrix.DEBUG_select_LA_EN[0]
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_224 VPWR VGND sg13g2_fill_1
XFILLER_9_375 VPWR VGND sg13g2_fill_1
X_2552_ FrameData[25] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_1503_ _0175_ VPWR _0176_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0174_ sg13g2_o21ai_1
X_2621_ FrameData[30] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_2483_ FrameData[20] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VPWR VGND sg13g2_dlhq_1
X_3104_ FrameData[1] FrameData_O[1] VPWR VGND sg13g2_buf_1
X_1365_ _0039_ _0042_ _0043_ VPWR VGND sg13g2_nor2_1
X_1296_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q NN4END[2] EE4END[2] E1END[0] E6END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q _1133_ VPWR VGND sg13g2_mux4_1
X_3035_ FrameData[28] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_1434_ _0110_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit2.Q Inst_LUT4AB_switch_matrix.M_AD
+ VPWR VGND sg13g2_nand2b_1
X_2819_ FrameData[4] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_33_422 VPWR VGND sg13g2_fill_2
XFILLER_20_105 VPWR VGND sg13g2_fill_2
X_1983_ VGND VPWR _0639_ _0638_ _0591_ sg13g2_or2_1
X_2604_ FrameData[13] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_2535_ FrameData[8] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_dlhq_1
X_1417_ VGND VPWR _0094_ _0076_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ sg13g2_or2_1
X_2466_ FrameData[3] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VPWR VGND sg13g2_dlhq_1
X_3018_ FrameData[11] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_1348_ _0026_ VPWR _0027_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0024_ sg13g2_o21ai_1
X_1279_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit1.Q _1116_ _1117_ VPWR VGND sg13g2_nor2_1
X_2397_ _0992_ Inst_LUT4AB_switch_matrix.DEBUG_select_LB_EN[0] _0973_ VPWR VGND sg13g2_nand2b_1
XFILLER_28_238 VPWR VGND sg13g2_fill_1
XFILLER_22_89 VPWR VGND sg13g2_fill_2
XFILLER_34_208 VPWR VGND sg13g2_fill_2
X_2320_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q _0940_ _0941_ _0943_ _0945_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit13.Q
+ Inst_LUT4AB_switch_matrix.NN4BEG3 VPWR VGND sg13g2_mux4_1
X_2251_ _0883_ _0885_ Inst_LUT4AB_switch_matrix.SS4BEG2 VPWR VGND sg13g2_nor2_1
X_1202_ VPWR _1043_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit17.Q VGND sg13g2_inv_1
X_2182_ _0824_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit29.Q _0825_ VPWR VGND sg13g2_nor2b_1
X_1966_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q NN4END[0] W2END[0] E6END[0] Inst_LUT4AB_switch_matrix.JW2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q _0623_ VPWR VGND sg13g2_mux4_1
X_1897_ _0554_ VPWR _0556_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q _0555_ sg13g2_o21ai_1
X_2518_ FrameData[23] FrameStrobe[16] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VPWR VGND sg13g2_dlhq_1
XFILLER_0_307 VPWR VGND sg13g2_fill_2
X_2449_ FrameData[18] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ VPWR VGND sg13g2_dlhq_1
XFILLER_17_23 VPWR VGND sg13g2_fill_1
X_1820_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q VPWR _0482_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q
+ _0253_ sg13g2_o21ai_1
X_1682_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit2.Q A B D E Inst_LUT4AB_ConfigMem.Inst_frame4_bit3.Q
+ _0349_ VPWR VGND sg13g2_mux4_1
X_1751_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q N1END[1] N2END[3] EE4END[3] E6END[1]
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q _0416_ VPWR VGND sg13g2_mux4_1
XFILLER_38_322 VPWR VGND sg13g2_fill_1
X_2303_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q N1END[3] E1END[3] S1END[3] A Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ _0931_ VPWR VGND sg13g2_mux4_1
X_3283_ W6END[5] W6BEG[3] VPWR VGND sg13g2_buf_1
X_2234_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q N1END[1] E1END[1] W1END[1] D Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q
+ _0870_ VPWR VGND sg13g2_mux4_1
X_2165_ VGND VPWR N2END[1] Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q _0809_ _0808_
+ sg13g2_a21oi_1
XFILLER_17_0 VPWR VGND sg13g2_fill_1
X_2096_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VPWR _0745_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q
+ _0744_ sg13g2_o21ai_1
X_1949_ _0606_ VPWR _0607_ VGND S2END[7] Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q
+ sg13g2_o21ai_1
X_2998_ FrameData[23] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_28_22 VPWR VGND sg13g2_fill_1
X_2921_ FrameData[10] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_2783_ FrameData[0] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_2852_ FrameData[5] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_1803_ _0464_ _0465_ _0203_ _0466_ VPWR VGND sg13g2_mux2_1
X_1596_ _1042_ VPWR _0267_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q _0266_ sg13g2_o21ai_1
X_1665_ _0331_ _0332_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q _0333_ VPWR VGND sg13g2_nand3_1
X_1734_ _0399_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4 _0395_ VPWR
+ VGND sg13g2_nand2b_1
X_3197_ NN4END[10] NN4BEG[6] VPWR VGND sg13g2_buf_1
X_3266_ Inst_LUT4AB_switch_matrix.JW2BEG2 W2BEG[2] VPWR VGND sg13g2_buf_1
X_2217_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q _0851_ _0852_ _0854_ _0856_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit25.Q
+ Inst_LUT4AB_switch_matrix.WW4BEG3 VPWR VGND sg13g2_mux4_1
X_2148_ VGND VPWR _0789_ _0792_ _0793_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q sg13g2_a21oi_1
X_2079_ _0728_ VPWR _0729_ VGND W1END[0] Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q
+ sg13g2_o21ai_1
XFILLER_4_273 VPWR VGND sg13g2_fill_2
X_1450_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit4.Q VPWR _0126_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit3.Q
+ _0125_ sg13g2_o21ai_1
X_3120_ FrameData[17] FrameData_O[17] VPWR VGND sg13g2_buf_1
X_1381_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ _1121_ _0059_ VPWR VGND sg13g2_mux2_1
X_3051_ VPWR VGND _1167_ sg13g2_tiehi
X_2002_ _0645_ _0657_ _0640_ _0658_ VPWR VGND sg13g2_nand3_1
XFILLER_35_111 VPWR VGND sg13g2_fill_1
X_2766_ FrameData[15] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_2835_ FrameData[20] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_2904_ FrameData[25] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_1717_ _0383_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q W1END[3] VPWR VGND sg13g2_nand2b_1
X_1579_ _0250_ SS4END[1] Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q VPWR VGND sg13g2_nand2b_1
X_1648_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit14.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q
+ _0317_ VPWR VGND sg13g2_mux4_1
X_2697_ FrameData[10] FrameStrobe[10] Inst_LUT4AB_switch_matrix.DEBUG_select_LA_SR[0]
+ VPWR VGND sg13g2_dlhq_1
X_3249_ SS4END[10] SS4BEG[6] VPWR VGND sg13g2_buf_1
XFILLER_14_339 VPWR VGND sg13g2_fill_1
X_2620_ FrameData[29] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_2551_ FrameData[24] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_1502_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit11.Q _0173_ _0175_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit12.Q
+ sg13g2_a21oi_1
X_2482_ FrameData[19] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VPWR VGND sg13g2_dlhq_1
X_1433_ _0109_ Inst_LB_LUT4c_frame_config_dffesr.LUT_flop Inst_LB_LUT4c_frame_config_dffesr.c_out_mux
+ B VPWR VGND sg13g2_mux2_1
XFILLER_48_280 VPWR VGND sg13g2_fill_1
X_3103_ FrameData[0] FrameData_O[0] VPWR VGND sg13g2_buf_1
X_1364_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q _0040_ _0041_ _0042_ VPWR VGND sg13g2_nor3_1
X_1295_ _1131_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit1.Q _1132_ VPWR VGND sg13g2_nor2b_1
X_3034_ FrameData[27] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_51_423 VPWR VGND sg13g2_fill_1
X_2749_ FrameData[30] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_180 VPWR VGND sg13g2_fill_2
X_2818_ FrameData[3] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_46_217 VPWR VGND sg13g2_fill_2
X_1982_ VPWR VGND _0590_ _0488_ _0565_ _0479_ _0638_ _0490_ sg13g2_a221oi_1
X_2534_ FrameData[7] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.c_out_mux VPWR
+ VGND sg13g2_dlhq_1
X_2603_ FrameData[12] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_47_0 VPWR VGND sg13g2_fill_1
X_2396_ Inst_LA_LUT4c_frame_config_dffesr.LUT_flop _0991_ _0990_ _0001_ VPWR VGND
+ sg13g2_mux2_1
X_1347_ _0026_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit8.Q _0025_ VPWR VGND sg13g2_nand2b_1
X_1416_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0081_ _0093_ VPWR
+ VGND sg13g2_nor2_1
X_2465_ FrameData[2] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VPWR VGND sg13g2_dlhq_1
X_3017_ FrameData[10] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_1278_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q _1114_ _1116_ _1115_ sg13g2_a21oi_1
XFILLER_24_423 VPWR VGND sg13g2_fill_1
XFILLER_51_275 VPWR VGND sg13g2_fill_2
XFILLER_47_65 VPWR VGND sg13g2_fill_2
XFILLER_15_423 VPWR VGND sg13g2_fill_1
XFILLER_6_121 VPWR VGND sg13g2_fill_2
X_1201_ VPWR _1042_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VGND sg13g2_inv_1
X_2250_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q _0884_ _0885_ VPWR VGND sg13g2_nor2_1
X_2181_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q _0822_ _0824_ _0823_ sg13g2_a21oi_1
X_1965_ _0621_ VPWR _0622_ VGND Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q _0618_ sg13g2_o21ai_1
X_2517_ FrameData[22] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.c_reset_value
+ VPWR VGND sg13g2_dlhq_1
X_1896_ E2MID[4] S2MID[4] Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q _0555_ VPWR VGND
+ sg13g2_mux2_1
X_2448_ FrameData[17] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VPWR VGND sg13g2_dlhq_1
X_2379_ _0976_ _0520_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q VPWR VGND sg13g2_nand2b_1
XFILLER_24_242 VPWR VGND sg13g2_fill_2
X_1750_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q _0413_ _0415_ _0414_ sg13g2_a21oi_1
X_1681_ _0348_ Inst_LE_LUT4c_frame_config_dffesr.LUT_flop Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ E VPWR VGND sg13g2_mux2_1
X_2233_ _0868_ _0869_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit16.Q Inst_LUT4AB_switch_matrix.WW4BEG0
+ VPWR VGND sg13g2_mux2_1
X_2302_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit25.Q H _1157_ _0197_ _0239_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit26.Q
+ _0930_ VPWR VGND sg13g2_mux4_1
X_2164_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q N1END[3] _0808_ VPWR VGND sg13g2_nor2b_1
X_3282_ W6END[4] W6BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_53_315 VPWR VGND sg13g2_fill_2
X_2095_ S1END[0] S1END[2] Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q _0744_ VPWR VGND
+ sg13g2_mux2_1
X_1948_ _0606_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q W1END[3] VPWR VGND sg13g2_nand2b_1
X_1879_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit18.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q
+ _0539_ VPWR VGND sg13g2_mux4_1
XFILLER_21_245 VPWR VGND sg13g2_fill_2
X_2997_ FrameData[22] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_2920_ FrameData[9] FrameStrobe[3] Inst_LUT4AB_ConfigMem.Inst_frame3_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_2851_ FrameData[4] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_2782_ FrameData[31] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1802_ _0202_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ _0395_ _0465_ VPWR VGND sg13g2_mux4_1
X_1733_ _0396_ _0397_ _0206_ _0398_ VPWR VGND sg13g2_nand3_1
X_1595_ N1END[2] N2END[6] Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q _0266_ VPWR VGND
+ sg13g2_mux2_1
X_1664_ _0332_ W2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q VPWR VGND sg13g2_nand2_1
X_3196_ NN4END[9] NN4BEG[5] VPWR VGND sg13g2_buf_1
XFILLER_53_123 VPWR VGND sg13g2_fill_2
X_2147_ _0791_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q _0792_ VPWR VGND sg13g2_nor2b_1
X_3265_ Inst_LUT4AB_switch_matrix.JW2BEG1 W2BEG[1] VPWR VGND sg13g2_buf_1
X_2216_ _0855_ VPWR _0856_ VGND Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _0556_
+ sg13g2_o21ai_1
XFILLER_14_47 VPWR VGND sg13g2_fill_2
X_2078_ _0728_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q W1END[2] VPWR VGND sg13g2_nand2b_1
XFILLER_30_13 VPWR VGND sg13g2_fill_1
XFILLER_29_131 VPWR VGND sg13g2_fill_1
X_1380_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ _1121_ _0058_ VPWR VGND sg13g2_mux2_1
X_2001_ VPWR _0657_ _0656_ VGND sg13g2_inv_1
X_3050_ VPWR VGND _1166_ sg13g2_tiehi
X_2903_ FrameData[24] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1716_ _0381_ VPWR _0382_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0380_ sg13g2_o21ai_1
X_2696_ FrameData[9] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_2765_ FrameData[14] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_2834_ FrameData[19] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1578_ N2END[5] E2END[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit14.Q _0249_ VPWR VGND
+ sg13g2_mux2_1
X_1647_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit16.Q NN4END[2] E2END[1] S2END[1] W2END[1]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit17.Q _0316_ VPWR VGND sg13g2_mux4_1
X_3248_ SS4END[9] SS4BEG[5] VPWR VGND sg13g2_buf_1
X_3179_ N4END[8] N4BEG[4] VPWR VGND sg13g2_buf_1
X_2550_ FrameData[23] FrameStrobe[15] Inst_LG_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
XFILLER_9_322 VPWR VGND sg13g2_fill_1
X_1501_ A B Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q _0174_ VPWR VGND sg13g2_mux2_1
X_1363_ N2MID[0] Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q _0041_ VPWR VGND sg13g2_nor2_1
X_1432_ VGND VPWR _0085_ _0097_ _0109_ _0108_ sg13g2_a21oi_1
X_2481_ FrameData[18] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VPWR VGND sg13g2_dlhq_1
X_3102_ Inst_LUT4AB_switch_matrix.EE4BEG3 EE4BEG[15] VPWR VGND sg13g2_buf_1
X_1294_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q _1130_ _1131_ VPWR VGND sg13g2_nor2_1
X_3033_ FrameData[26] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_2748_ FrameData[29] FrameStrobe[9] Inst_LUT4AB_switch_matrix.DEBUG_select_LF_EN[0]
+ VPWR VGND sg13g2_dlhq_1
X_2679_ FrameData[24] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_2817_ FrameData[2] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_36_12 VPWR VGND sg13g2_fill_2
XFILLER_36_56 VPWR VGND sg13g2_fill_1
XFILLER_27_421 VPWR VGND sg13g2_fill_2
XFILLER_6_369 VPWR VGND sg13g2_fill_2
XFILLER_10_398 VPWR VGND sg13g2_fill_1
X_1981_ _0637_ VPWR G VGND Inst_LG_LUT4c_frame_config_dffesr.c_out_mux _0636_ sg13g2_o21ai_1
XFILLER_20_107 VPWR VGND sg13g2_fill_1
X_2533_ FrameData[6] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_2602_ FrameData[11] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_9_163 VPWR VGND sg13g2_fill_1
X_1346_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q F G H Inst_LUT4AB_switch_matrix.M_AB
+ Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q _0025_ VPWR VGND sg13g2_mux4_1
X_2395_ Inst_LA_LUT4c_frame_config_dffesr.c_reset_value _0069_ _0989_ _0991_ VPWR
+ VGND sg13g2_mux2_1
X_1415_ Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2 _0078_ _0092_ VPWR
+ VGND sg13g2_nor2b_1
X_2464_ FrameData[1] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VPWR VGND sg13g2_dlhq_1
XFILLER_51_254 VPWR VGND sg13g2_fill_1
X_3016_ FrameData[9] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1277_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VPWR _1115_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q
+ _1112_ sg13g2_o21ai_1
X_1200_ VPWR _1041_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit13.Q VGND sg13g2_inv_1
X_2180_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit28.Q VPWR _0823_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit27.Q
+ _0820_ sg13g2_o21ai_1
X_1964_ _0619_ _0620_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit25.Q _0621_ VPWR VGND sg13g2_nand3_1
X_1895_ Inst_LUT4AB_switch_matrix.JS2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q
+ _0553_ _0554_ VPWR VGND sg13g2_a21o_1
X_2516_ FrameData[21] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.c_I0mux VPWR
+ VGND sg13g2_dlhq_1
X_2447_ FrameData[16] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VPWR VGND sg13g2_dlhq_1
X_2378_ Inst_LUT4AB_switch_matrix.DEBUG_select_LH_EN[0] Inst_LH_LUT4c_frame_config_dffesr.LUT_flop
+ _0975_ VPWR VGND _0973_ sg13g2_nand3b_1
X_1329_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q F G H Inst_LUT4AB_switch_matrix.M_AH
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q _0009_ VPWR VGND sg13g2_mux4_1
XFILLER_24_210 VPWR VGND sg13g2_fill_1
XFILLER_47_302 VPWR VGND sg13g2_fill_2
X_1680_ _0348_ _0347_ _0342_ VPWR VGND sg13g2_nand2b_1
X_2301_ Inst_LUT4AB_switch_matrix.EE4BEG2 _0927_ _0929_ _0925_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
+ VPWR VGND sg13g2_a22oi_1
X_3281_ W6END[3] W6BEG[1] VPWR VGND sg13g2_buf_1
X_2163_ N4END[1] EE4END[1] Inst_LUT4AB_ConfigMem.Inst_frame4_bit26.Q _0807_ VPWR VGND
+ sg13g2_mux2_1
X_2232_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q G _1084_ _0148_ _0538_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ _0869_ VPWR VGND sg13g2_mux4_1
X_2094_ _0742_ VPWR _0743_ VGND SS4END[0] Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q
+ sg13g2_o21ai_1
X_1947_ S1END[1] S1END[3] Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q _0605_ VPWR VGND
+ sg13g2_mux2_1
X_2996_ FrameData[21] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_1878_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit23.Q NN4END[1] S2END[5] E2END[5] W2END[5]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit22.Q _0538_ VPWR VGND sg13g2_mux4_1
XFILLER_29_313 VPWR VGND sg13g2_fill_1
XFILLER_4_401 VPWR VGND sg13g2_fill_1
XFILLER_47_198 VPWR VGND sg13g2_fill_2
X_2850_ FrameData[3] FrameStrobe[5] Inst_LUT4AB_ConfigMem.Inst_frame5_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_1663_ _0331_ S2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q VPWR VGND sg13g2_nand2b_1
X_2781_ FrameData[30] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1801_ _0202_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A10
+ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9 Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ _0395_ _0464_ VPWR VGND sg13g2_mux4_1
X_1732_ _0397_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6 _0395_ VPWR
+ VGND sg13g2_nand2b_1
X_1594_ VGND VPWR E2END[6] Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q _0265_ _0264_
+ sg13g2_a21oi_1
XFILLER_22_0 VPWR VGND sg13g2_fill_1
X_3264_ Inst_LUT4AB_switch_matrix.JW2BEG0 W2BEG[0] VPWR VGND sg13g2_buf_1
X_3195_ NN4END[8] NN4BEG[4] VPWR VGND sg13g2_buf_1
X_2146_ VGND VPWR _1028_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q _0791_ _0790_ sg13g2_a21oi_1
X_2215_ _0855_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _1141_ VPWR VGND sg13g2_nand2_1
X_2077_ _0726_ VPWR _0727_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0724_ sg13g2_o21ai_1
X_2979_ FrameData[4] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_4_275 VPWR VGND sg13g2_fill_1
X_2000_ _0650_ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5 Inst_LH_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ _0649_ _0656_ VPWR VGND sg13g2_mux4_1
X_2833_ FrameData[18] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_2902_ FrameData[23] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1715_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0379_ _0381_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit12.Q
+ sg13g2_a21oi_1
X_2764_ FrameData[13] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_1646_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit17.Q _1040_ _1030_ _1022_ _0037_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit16.Q
+ _0315_ VPWR VGND sg13g2_mux4_1
X_2695_ FrameData[8] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_3247_ SS4END[8] SS4BEG[4] VPWR VGND sg13g2_buf_1
X_1577_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit14.Q N4END[1] SS4END[1] W2END[4] Inst_LUT4AB_switch_matrix.JS2BEG3
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit15.Q _0248_ VPWR VGND sg13g2_mux4_1
X_3178_ N4END[7] N4BEG[3] VPWR VGND sg13g2_buf_1
X_2129_ VGND VPWR S4END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q _0775_ _0774_
+ sg13g2_a21oi_1
XFILLER_41_57 VPWR VGND sg13g2_fill_1
X_1500_ _0172_ VPWR _0173_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit10.Q C sg13g2_o21ai_1
XFILLER_9_345 VPWR VGND sg13g2_fill_2
X_2480_ FrameData[17] FrameStrobe[17] Inst_LD_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VPWR VGND sg13g2_dlhq_1
X_3101_ Inst_LUT4AB_switch_matrix.EE4BEG2 EE4BEG[14] VPWR VGND sg13g2_buf_1
X_1362_ E2MID[0] Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q _0040_ VPWR VGND sg13g2_nor2b_1
X_1431_ _0091_ _0102_ _0107_ _0108_ VPWR VGND sg13g2_nor3_1
X_1293_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q A D C E Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ _1130_ VPWR VGND sg13g2_mux4_1
X_3032_ FrameData[25] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_2816_ FrameData[1] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_2747_ FrameData[28] FrameStrobe[9] Inst_LUT4AB_switch_matrix.DEBUG_select_LF_SR[0]
+ VPWR VGND sg13g2_dlhq_1
X_1629_ _0298_ VPWR _0299_ VGND S2END[6] Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q
+ sg13g2_o21ai_1
X_2678_ FrameData[23] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_46_219 VPWR VGND sg13g2_fill_1
XFILLER_36_35 VPWR VGND sg13g2_fill_1
X_1980_ _0637_ Inst_LG_LUT4c_frame_config_dffesr.LUT_flop Inst_LG_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_nand2_1
X_2532_ FrameData[5] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
X_2463_ FrameData[0] FrameStrobe[17] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VPWR VGND sg13g2_dlhq_1
X_2601_ FrameData[10] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
X_3015_ FrameData[8] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1345_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit6.Q A B C E Inst_LUT4AB_ConfigMem.Inst_frame1_bit7.Q
+ _0024_ VPWR VGND sg13g2_mux4_1
X_2394_ _0990_ Inst_LUT4AB_switch_matrix.DEBUG_select_LA_EN[0] _0973_ VPWR VGND sg13g2_nand2b_1
X_1276_ _1113_ VPWR _1114_ VGND Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q W2END[2]
+ sg13g2_o21ai_1
X_1414_ VGND VPWR Inst_LB_LUT4c_frame_config_dffesr.c_I0mux _0089_ _0091_ _0090_ sg13g2_a21oi_1
XFILLER_51_277 VPWR VGND sg13g2_fill_1
XFILLER_47_34 VPWR VGND sg13g2_fill_1
XFILLER_47_23 VPWR VGND sg13g2_fill_1
XFILLER_6_112 VPWR VGND sg13g2_fill_1
X_1963_ _0620_ W2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q VPWR VGND sg13g2_nand2_1
X_1894_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit23.Q VPWR _0553_ VGND _1026_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit22.Q
+ sg13g2_o21ai_1
XFILLER_52_0 VPWR VGND sg13g2_fill_2
X_2515_ FrameData[20] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.c_out_mux
+ VPWR VGND sg13g2_dlhq_1
X_2446_ FrameData[15] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VPWR VGND sg13g2_dlhq_1
X_2377_ _0974_ Inst_LUT4AB_switch_matrix.DEBUG_select_LH_EN[0] _0973_ VPWR VGND sg13g2_nand2b_1
X_1259_ N2END[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _1098_ VPWR VGND sg13g2_nor2_1
X_1328_ _1160_ _1162_ _0008_ VPWR VGND sg13g2_nor2_1
XFILLER_12_417 VPWR VGND sg13g2_fill_2
XFILLER_24_222 VPWR VGND sg13g2_fill_2
XFILLER_24_244 VPWR VGND sg13g2_fill_1
XFILLER_47_358 VPWR VGND sg13g2_fill_2
XFILLER_23_91 VPWR VGND sg13g2_fill_1
X_2231_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit14.Q N1END[2] S1END[2] W1END[2] F Inst_LUT4AB_ConfigMem.Inst_frame11_bit15.Q
+ _0868_ VPWR VGND sg13g2_mux4_1
X_3280_ W6END[2] W6BEG[0] VPWR VGND sg13g2_buf_1
X_2300_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit29.Q _0928_ _0929_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit30.Q
+ sg13g2_a21oi_1
XFILLER_53_317 VPWR VGND sg13g2_fill_1
X_2162_ _0800_ _0805_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit29.Q _0806_ VPWR VGND sg13g2_nand3_1
X_2093_ _0742_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q WW4END[0] VPWR VGND sg13g2_nand2b_1
X_2995_ FrameData[20] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_1946_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit21.Q _0603_ _0604_ VPWR VGND sg13g2_and2_1
X_1877_ _0536_ VPWR _0537_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q _0533_ sg13g2_o21ai_1
X_2429_ FrameData[30] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A6
+ VPWR VGND sg13g2_dlhq_1
XFILLER_8_218 VPWR VGND sg13g2_fill_2
X_1800_ _0401_ _0457_ _0460_ _0462_ _0463_ VPWR VGND sg13g2_nor4_1
X_1662_ N2MID[1] E2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q _0330_ VPWR VGND
+ sg13g2_mux2_1
X_2780_ FrameData[29] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1731_ _0396_ Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7 _0395_ VPWR
+ VGND sg13g2_nand2_1
X_3194_ NN4END[7] NN4BEG[3] VPWR VGND sg13g2_buf_1
X_1593_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q VPWR _0264_ VGND _1013_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q
+ sg13g2_o21ai_1
X_3263_ Inst_LUT4AB_switch_matrix.W1BEG3 W1BEG[3] VPWR VGND sg13g2_buf_1
X_2214_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _0276_ _0854_ _0853_
+ sg13g2_a21oi_1
XFILLER_53_169 VPWR VGND sg13g2_fill_1
X_2145_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q VPWR _0790_ VGND W2END[1] Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ sg13g2_o21ai_1
X_2076_ _0726_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit24.Q _0725_ VPWR VGND sg13g2_nand2b_1
X_1929_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit21.Q N4END[2] W2END[2] SS4END[2] Inst_LUT4AB_switch_matrix.E2BEG4
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit20.Q _0587_ VPWR VGND sg13g2_mux4_1
X_2978_ FrameData[3] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_40_397 VPWR VGND sg13g2_fill_2
XFILLER_4_210 VPWR VGND sg13g2_fill_2
X_2763_ FrameData[12] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit12.Q VPWR
+ VGND sg13g2_dlhq_1
X_2901_ FrameData[22] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_320 VPWR VGND sg13g2_fill_2
X_2832_ FrameData[17] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_1714_ N1END[1] N2END[5] Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q _0380_ VPWR VGND
+ sg13g2_mux2_1
X_1576_ _0247_ _0240_ _0246_ VPWR VGND sg13g2_nand2_1
X_1645_ _0313_ _0247_ _0314_ VPWR VGND sg13g2_nor2b_1
X_2694_ FrameData[7] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_3246_ SS4END[7] SS4BEG[3] VPWR VGND sg13g2_buf_1
X_3177_ N4END[6] N4BEG[2] VPWR VGND sg13g2_buf_1
X_2128_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q S2END[1] _0774_ VPWR VGND sg13g2_nor2b_1
X_2059_ VGND VPWR _1045_ _0705_ _0711_ _0710_ sg13g2_a21oi_1
XFILLER_45_423 VPWR VGND sg13g2_fill_1
XFILLER_17_114 VPWR VGND sg13g2_fill_2
XFILLER_13_353 VPWR VGND sg13g2_fill_2
X_1430_ _0073_ _0103_ _0104_ _0106_ _0107_ VPWR VGND sg13g2_nor4_1
X_3100_ Inst_LUT4AB_switch_matrix.EE4BEG1 EE4BEG[13] VPWR VGND sg13g2_buf_1
XFILLER_36_401 VPWR VGND sg13g2_fill_2
X_1361_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q _0037_ _0039_ _0038_ sg13g2_a21oi_1
X_3031_ FrameData[24] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_1292_ _1128_ VPWR _1129_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q _1126_ sg13g2_o21ai_1
X_2746_ FrameData[27] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_2815_ FrameData[0] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1559_ VPWR Inst_LUT4AB_switch_matrix.JN2BEG5 _0230_ VGND sg13g2_inv_1
X_1628_ _0298_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q W1END[2] VPWR VGND sg13g2_nand2b_1
X_2677_ FrameData[22] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_3229_ S4END[6] S4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_27_423 VPWR VGND sg13g2_fill_1
XFILLER_14_139 VPWR VGND sg13g2_fill_2
XFILLER_18_423 VPWR VGND sg13g2_fill_1
X_2600_ FrameData[9] FrameStrobe[13] Inst_LUT4AB_ConfigMem.Inst_frame13_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_2531_ FrameData[4] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_1413_ Inst_LB_LUT4c_frame_config_dffesr.c_I0mux _0086_ _0090_ VPWR VGND sg13g2_nor2b_1
X_2393_ _0989_ Inst_LUT4AB_switch_matrix.DEBUG_select_LA_SR[0] _0985_ VPWR VGND sg13g2_nand2_1
X_2462_ FrameData[31] FrameStrobe[18] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VPWR VGND sg13g2_dlhq_1
XFILLER_36_242 VPWR VGND sg13g2_fill_2
X_1275_ _1113_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q W6END[0] VPWR VGND sg13g2_nand2b_1
X_3014_ FrameData[7] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1344_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit1.Q N2END[0] S2END[0] E2END[0] WW4END[3]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit0.Q _0023_ VPWR VGND sg13g2_mux4_1
XFILLER_51_289 VPWR VGND sg13g2_fill_1
X_2729_ FrameData[10] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_27_253 VPWR VGND sg13g2_fill_1
XFILLER_27_297 VPWR VGND sg13g2_fill_1
XFILLER_33_289 VPWR VGND sg13g2_fill_2
X_1962_ _0619_ S2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q VPWR VGND sg13g2_nand2b_1
XFILLER_18_253 VPWR VGND sg13g2_fill_2
X_1893_ _0545_ _0552_ Inst_LUT4AB_switch_matrix.JS2BEG6 VPWR VGND sg13g2_nor2_1
X_2514_ FrameData[19] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A15
+ VPWR VGND sg13g2_dlhq_1
X_2376_ _0971_ VPWR _0973_ VGND Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q _0972_ sg13g2_o21ai_1
X_2445_ FrameData[14] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VPWR VGND sg13g2_dlhq_1
X_1258_ E1END[2] E2END[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _1097_ VPWR VGND
+ sg13g2_mux2_1
X_1189_ VPWR _1030_ WW4END[1] VGND sg13g2_inv_1
X_1327_ _1085_ _1161_ _1162_ VPWR VGND sg13g2_nor2_1
XFILLER_47_304 VPWR VGND sg13g2_fill_1
X_2230_ _0867_ VPWR Inst_LUT4AB_switch_matrix.WW4BEG1 VGND _1048_ _0865_ sg13g2_o21ai_1
X_2161_ _0804_ VPWR _0805_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0803_ sg13g2_o21ai_1
X_2092_ _0741_ _0740_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q VPWR VGND sg13g2_nand2b_1
X_2994_ FrameData[19] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_1945_ _0602_ VPWR _0603_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0601_ sg13g2_o21ai_1
X_1876_ _0534_ _0535_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q _0536_ VPWR VGND sg13g2_nand3_1
X_2428_ FrameData[29] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ VPWR VGND sg13g2_dlhq_1
X_2359_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit15.Q D Inst_LUT4AB_switch_matrix.JN2BEG3
+ _0453_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit14.Q Inst_LUT4AB_switch_matrix.E1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1592_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit17.Q VPWR _0263_ VGND _0261_ _0262_ sg13g2_o21ai_1
X_1661_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit16.Q E2MID[0] S2MID[0] W2MID[0] Inst_LUT4AB_switch_matrix.JW2BEG5
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit17.Q _0329_ VPWR VGND sg13g2_mux4_1
X_1730_ _0394_ _0207_ Inst_LC_LUT4c_frame_config_dffesr.c_I0mux _0395_ VPWR VGND sg13g2_mux2_1
X_3193_ NN4END[6] NN4BEG[2] VPWR VGND sg13g2_buf_1
X_2144_ _0788_ VPWR _0789_ VGND S2END[1] Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q
+ sg13g2_o21ai_1
X_3262_ Inst_LUT4AB_switch_matrix.W1BEG2 W1BEG[2] VPWR VGND sg13g2_buf_1
X_2213_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q E _0853_ VPWR VGND sg13g2_nor2_1
X_2075_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q E G F Inst_LUT4AB_switch_matrix.M_EF
+ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q _0725_ VPWR VGND sg13g2_mux4_1
X_1859_ N2MID[6] E2MID[6] Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q _0519_ VPWR VGND
+ sg13g2_mux2_1
X_2977_ FrameData[2] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_1928_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit20.Q N2MID[3] E2MID[3] S2MID[3] W2MID[3]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit21.Q _0586_ VPWR VGND sg13g2_mux4_1
XFILLER_40_343 VPWR VGND sg13g2_fill_2
X_2900_ FrameData[21] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_1713_ _0378_ VPWR _0379_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q E1END[1]
+ sg13g2_o21ai_1
X_2762_ FrameData[11] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit11.Q VPWR
+ VGND sg13g2_dlhq_1
X_2831_ FrameData[16] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_1575_ _0245_ VPWR _0246_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q _0242_ sg13g2_o21ai_1
X_1644_ _0280_ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A7
+ Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1 Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A5
+ _0310_ _0313_ VPWR VGND sg13g2_mux4_1
X_2693_ FrameData[6] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_3245_ SS4END[6] SS4BEG[2] VPWR VGND sg13g2_buf_1
X_3176_ N4END[5] N4BEG[1] VPWR VGND sg13g2_buf_1
X_2127_ W2END[1] W6END[1] Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q _0773_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_41_129 VPWR VGND sg13g2_fill_1
X_2058_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q _0707_ _0710_ _0709_ sg13g2_a21oi_1
XFILLER_9_303 VPWR VGND sg13g2_fill_2
XFILLER_9_347 VPWR VGND sg13g2_fill_1
X_1360_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit1.Q VPWR _0038_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit0.Q
+ S2MID[0] sg13g2_o21ai_1
XFILLER_48_262 VPWR VGND sg13g2_fill_1
X_3030_ FrameData[23] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
X_1291_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit31.Q _1127_ _1128_ _1027_ sg13g2_a21oi_1
XFILLER_51_416 VPWR VGND sg13g2_fill_2
X_2745_ FrameData[26] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit26.Q VPWR
+ VGND sg13g2_dlhq_1
X_2676_ FrameData[21] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit21.Q VPWR
+ VGND sg13g2_dlhq_1
X_2814_ FrameData[31] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1627_ S1END[0] S1END[2] Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q _0297_ VPWR VGND
+ sg13g2_mux2_1
X_1558_ _0229_ VPWR _0230_ VGND _0215_ _0221_ sg13g2_o21ai_1
X_1489_ _0163_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q W6END[1] VPWR VGND sg13g2_nand2b_1
X_3228_ S4END[5] S4BEG[1] VPWR VGND sg13g2_buf_1
X_3159_ Inst_LUT4AB_switch_matrix.JN2BEG0 N2BEG[0] VPWR VGND sg13g2_buf_1
X_2530_ FrameData[3] FrameStrobe[15] Inst_LF_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
XFILLER_13_162 VPWR VGND sg13g2_fill_2
X_2392_ _0975_ VPWR _0000_ VGND _0987_ _0988_ sg13g2_o21ai_1
X_1343_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit0.Q _1012_ _1014_ _1022_ _0021_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit1.Q
+ _0022_ VPWR VGND sg13g2_mux4_1
X_1412_ _0089_ _0087_ _0088_ VPWR VGND sg13g2_nand2_1
X_2461_ FrameData[30] FrameStrobe[18] Inst_LC_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VPWR VGND sg13g2_dlhq_1
X_1274_ _1111_ VPWR _1112_ VGND _1014_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q sg13g2_o21ai_1
X_3013_ FrameData[6] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_2728_ FrameData[9] FrameStrobe[9] Inst_LUT4AB_switch_matrix.DEBUG_select_LD_EN[0]
+ VPWR VGND sg13g2_dlhq_1
X_2659_ FrameData[4] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_10_110 VPWR VGND sg13g2_fill_1
XFILLER_5_0 VPWR VGND sg13g2_fill_1
X_1892_ VPWR VGND _0551_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit21.Q _0550_ _1044_ _0552_
+ _0546_ sg13g2_a221oi_1
X_1961_ N2MID[1] E2MID[1] Inst_LUT4AB_ConfigMem.Inst_frame6_bit24.Q _0618_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_18_287 VPWR VGND sg13g2_fill_2
XFILLER_52_2 VPWR VGND sg13g2_fill_1
X_2513_ FrameData[18] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A14
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_0 VPWR VGND sg13g2_fill_2
X_1326_ Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A8 Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A9
+ _1121_ _1161_ VPWR VGND sg13g2_mux2_1
X_2375_ _0972_ _0969_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q _0967_ _0966_ VPWR
+ VGND sg13g2_a22oi_1
X_2444_ FrameData[13] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VPWR VGND sg13g2_dlhq_1
X_1188_ VPWR _1029_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit8.Q VGND sg13g2_inv_1
X_1257_ W2END[4] W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _1096_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_12_419 VPWR VGND sg13g2_fill_1
XFILLER_24_224 VPWR VGND sg13g2_fill_1
XFILLER_33_38 VPWR VGND sg13g2_fill_2
XFILLER_15_279 VPWR VGND sg13g2_fill_2
X_2160_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit27.Q _0801_ _0804_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit28.Q
+ sg13g2_a21oi_1
X_2091_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit22.Q N1END[0] N2END[0] E1END[0] E2END[0]
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit23.Q _0740_ VPWR VGND sg13g2_mux4_1
X_2993_ FrameData[18] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_1944_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit19.Q _0600_ _0602_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit20.Q
+ sg13g2_a21oi_1
X_1875_ _0535_ WW4END[3] Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q VPWR VGND sg13g2_nand2b_1
XFILLER_9_40 VPWR VGND sg13g2_fill_2
XFILLER_21_238 VPWR VGND sg13g2_decap_8
X_2427_ FrameData[28] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A4
+ VPWR VGND sg13g2_dlhq_1
X_2289_ _0918_ VPWR _0919_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q _0556_
+ sg13g2_o21ai_1
X_1309_ _1145_ _1144_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q VPWR VGND sg13g2_nand2b_1
X_2358_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit16.Q E _0237_ Inst_LUT4AB_switch_matrix.JN2BEG0
+ _0248_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit17.Q Inst_LUT4AB_switch_matrix.E1BEG1
+ VPWR VGND sg13g2_mux4_1
XFILLER_47_124 VPWR VGND sg13g2_fill_2
XFILLER_34_92 VPWR VGND sg13g2_fill_2
X_1591_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VPWR _0262_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q
+ _0259_ sg13g2_o21ai_1
X_1660_ Inst_LUT4AB_switch_matrix.JW2BEG5 _0322_ _0328_ _0320_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q
+ VPWR VGND sg13g2_a22oi_1
X_3192_ NN4END[5] NN4BEG[1] VPWR VGND sg13g2_buf_1
X_2143_ VGND VPWR _1036_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q _0788_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q
+ sg13g2_a21oi_1
X_3261_ Inst_LUT4AB_switch_matrix.W1BEG1 W1BEG[1] VPWR VGND sg13g2_buf_1
XFILLER_26_319 VPWR VGND sg13g2_fill_2
X_2212_ W1END[1] D Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _0852_ VPWR VGND sg13g2_mux2_1
X_2074_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit22.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame4_bit23.Q
+ _0724_ VPWR VGND sg13g2_mux4_1
X_1858_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit19.Q VPWR _0518_ VGND _0516_ _0517_ sg13g2_o21ai_1
X_1927_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit21.Q N2MID[2] W2MID[2] S2MID[2] Inst_LUT4AB_switch_matrix.E2BEG6
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit20.Q _0585_ VPWR VGND sg13g2_mux4_1
X_2976_ FrameData[1] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_1789_ _0450_ VPWR _0452_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q _0451_ sg13g2_o21ai_1
XFILLER_1_418 VPWR VGND sg13g2_fill_1
XFILLER_52_160 VPWR VGND sg13g2_fill_1
XFILLER_48_422 VPWR VGND sg13g2_fill_2
X_2830_ FrameData[15] FrameStrobe[6] Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_344 VPWR VGND sg13g2_fill_2
XFILLER_16_396 VPWR VGND sg13g2_fill_2
X_1712_ _0378_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q E2END[5] VPWR VGND sg13g2_nand2b_1
X_1643_ _0281_ _0310_ _0312_ VPWR VGND sg13g2_nor2_1
X_2761_ FrameData[10] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
XANTENNA_1 VPWR VGND EE4END[10] sg13g2_antennanp
XFILLER_6_41 VPWR VGND sg13g2_fill_2
X_2692_ FrameData[5] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
X_3244_ SS4END[5] SS4BEG[1] VPWR VGND sg13g2_buf_1
X_1574_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit11.Q _0244_ _0245_ Inst_LE_LUT4c_frame_config_dffesr.c_I0mux
+ sg13g2_a21oi_1
X_2126_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q N1END[3] E2END[1] N2END[1] E6END[1]
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit26.Q _0772_ VPWR VGND sg13g2_mux4_1
X_2057_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit24.Q VPWR _0709_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit23.Q
+ _0708_ sg13g2_o21ai_1
X_3175_ N4END[4] N4BEG[0] VPWR VGND sg13g2_buf_1
X_2959_ FrameData[16] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_22_311 VPWR VGND sg13g2_fill_1
XFILLER_17_149 VPWR VGND sg13g2_fill_1
X_1290_ H Inst_LUT4AB_switch_matrix.M_EF Inst_LUT4AB_ConfigMem.Inst_frame3_bit30.Q
+ _1127_ VPWR VGND sg13g2_mux2_1
X_2813_ FrameData[30] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_1626_ _0296_ _0295_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q VPWR VGND sg13g2_nand2b_1
X_2744_ FrameData[25] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit25.Q VPWR
+ VGND sg13g2_dlhq_1
X_2675_ FrameData[20] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit20.Q VPWR
+ VGND sg13g2_dlhq_1
X_3227_ S4END[4] S4BEG[0] VPWR VGND sg13g2_buf_1
X_1557_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit17.Q _0223_ _0228_ _0229_ VPWR VGND sg13g2_or3_1
X_1488_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit2.Q NN4END[3] E1END[1] E2END[3] E6END[1]
+ Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0162_ VPWR VGND sg13g2_mux4_1
X_2109_ VGND VPWR _1052_ _0755_ _0757_ _0756_ sg13g2_a21oi_1
X_3158_ Inst_LUT4AB_switch_matrix.N1BEG3 N1BEG[3] VPWR VGND sg13g2_buf_1
X_3089_ EE4END[6] EE4BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_10_358 VPWR VGND sg13g2_fill_1
XFILLER_10_369 VPWR VGND sg13g2_fill_2
XFILLER_22_141 VPWR VGND sg13g2_fill_1
XFILLER_33_417 VPWR VGND sg13g2_fill_1
X_2460_ FrameData[29] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.c_reset_value
+ VPWR VGND sg13g2_dlhq_1
X_2391_ _0974_ VPWR _0988_ VGND Inst_LH_LUT4c_frame_config_dffesr.c_reset_value _0986_
+ sg13g2_o21ai_1
X_1273_ _1111_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q S2END[2] VPWR VGND sg13g2_nand2_1
X_1411_ _1085_ VPWR _0088_ VGND Ci _1160_ sg13g2_o21ai_1
X_1342_ VPWR Inst_LUT4AB_switch_matrix.JW2BEG1 _0021_ VGND sg13g2_inv_1
XFILLER_51_236 VPWR VGND sg13g2_fill_1
X_3012_ FrameData[5] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit5.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_22_18 VPWR VGND sg13g2_fill_1
XFILLER_22_29 VPWR VGND sg13g2_fill_1
X_1609_ _0278_ VPWR _0279_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q _0276_ sg13g2_o21ai_1
X_2727_ FrameData[8] FrameStrobe[9] Inst_LUT4AB_switch_matrix.DEBUG_select_LD_SR[0]
+ VPWR VGND sg13g2_dlhq_1
X_2589_ FrameData[30] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
X_2658_ FrameData[3] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_42_236 VPWR VGND sg13g2_fill_2
X_1891_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q _0548_ _0551_ _1044_ sg13g2_a21oi_1
X_1960_ _0615_ VPWR _0617_ VGND Inst_LUT4AB_ConfigMem.Inst_frame7_bit25.Q _0616_ sg13g2_o21ai_1
X_2512_ FrameData[17] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A13
+ VPWR VGND sg13g2_dlhq_1
X_2443_ FrameData[12] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VPWR VGND sg13g2_dlhq_1
XFILLER_49_391 VPWR VGND sg13g2_fill_2
X_2374_ _0971_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit31.Q _0970_ VPWR VGND sg13g2_nand2_1
X_1256_ E6END[0] S2END[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit6.Q _1095_ VPWR VGND
+ sg13g2_mux2_1
X_1325_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit6.Q _1157_ _1159_ _1141_ _1140_ Inst_LUT4AB_ConfigMem.Inst_frame10_bit7.Q
+ _1160_ VPWR VGND sg13g2_mux4_1
X_1187_ VPWR _1028_ W6END[1] VGND sg13g2_inv_1
XFILLER_47_339 VPWR VGND sg13g2_fill_2
XFILLER_2_173 VPWR VGND sg13g2_fill_1
X_2090_ _0738_ VPWR _0739_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit24.Q _0736_ sg13g2_o21ai_1
X_2992_ FrameData[17] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_0_65 VPWR VGND sg13g2_fill_1
X_1943_ A B Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q _0601_ VPWR VGND sg13g2_mux2_1
X_1874_ _0534_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q Inst_LUT4AB_switch_matrix.JS2BEG4
+ VPWR VGND sg13g2_nand2_1
Xclkbuf_0_UserCLK UserCLK clknet_0_UserCLK VPWR VGND sg13g2_buf_8
XFILLER_50_0 VPWR VGND sg13g2_fill_1
X_2426_ FrameData[27] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A3
+ VPWR VGND sg13g2_dlhq_1
X_2288_ _0918_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q _1119_ VPWR VGND sg13g2_nand2_1
X_1308_ F G Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q _1144_ VPWR VGND sg13g2_mux2_1
X_1239_ E6END[0] S2END[4] Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1079_ VPWR VGND
+ sg13g2_mux2_1
X_2357_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit19.Q F Inst_LUT4AB_switch_matrix.JN2BEG1
+ _0586_ _0623_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit18.Q Inst_LUT4AB_switch_matrix.E1BEG2
+ VPWR VGND sg13g2_mux4_1
XFILLER_43_364 VPWR VGND sg13g2_fill_2
XFILLER_11_294 VPWR VGND sg13g2_fill_1
XFILLER_50_92 VPWR VGND sg13g2_fill_2
X_1590_ _0260_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q _0261_ VPWR VGND sg13g2_nor2b_1
X_3260_ Inst_LUT4AB_switch_matrix.W1BEG0 W1BEG[0] VPWR VGND sg13g2_buf_1
X_3191_ NN4END[4] NN4BEG[0] VPWR VGND sg13g2_buf_1
XFILLER_38_114 VPWR VGND sg13g2_fill_2
X_2142_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q NN4END[1] E2END[1] E1END[3] E6END[1]
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit26.Q _0787_ VPWR VGND sg13g2_mux4_1
X_2073_ Inst_LUT4AB_switch_matrix.JW2BEG7 _0717_ _0723_ _0715_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q
+ VPWR VGND sg13g2_a22oi_1
X_2211_ N1END[1] S1END[1] Inst_LUT4AB_ConfigMem.Inst_frame11_bit23.Q _0851_ VPWR VGND
+ sg13g2_mux2_1
X_2975_ FrameData[0] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit0.Q VPWR
+ VGND sg13g2_dlhq_1
X_1857_ S2MID[6] Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q _0517_ VPWR VGND sg13g2_nor2_1
X_1926_ Inst_LUT4AB_switch_matrix.E2BEG6 _0578_ _0584_ _0573_ _0567_ VPWR VGND sg13g2_a22oi_1
X_1788_ N2MID[0] S2MID[0] Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q _0451_ VPWR VGND
+ sg13g2_mux2_1
X_2409_ _1001_ Inst_LUT4AB_switch_matrix.DEBUG_select_LE_EN[0] _0973_ VPWR VGND sg13g2_nand2b_1
XFILLER_52_194 VPWR VGND sg13g2_fill_1
XFILLER_31_367 VPWR VGND sg13g2_fill_2
X_2760_ FrameData[9] FrameStrobe[8] Inst_LUT4AB_ConfigMem.Inst_frame8_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
X_1642_ _0311_ _0281_ _0310_ VPWR VGND sg13g2_nand2_1
XANTENNA_2 VPWR VGND EE4END[14] sg13g2_antennanp
X_1711_ _0376_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit13.Q _0377_ VPWR VGND sg13g2_nor2b_1
X_2691_ FrameData[4] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_3243_ SS4END[4] SS4BEG[0] VPWR VGND sg13g2_buf_1
X_1573_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q _0238_ _0244_ _0243_ sg13g2_a21oi_1
X_2125_ _0770_ VPWR _0771_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit28.Q _0763_ sg13g2_o21ai_1
XFILLER_13_0 VPWR VGND sg13g2_fill_2
X_2056_ S1END[0] S2END[0] Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q _0708_ VPWR VGND
+ sg13g2_mux2_1
X_3174_ N2MID[7] N2BEGb[7] VPWR VGND sg13g2_buf_1
X_1909_ E F Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q _0568_ VPWR VGND sg13g2_mux2_1
X_2958_ FrameData[15] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
X_2889_ FrameData[10] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit10.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_51_418 VPWR VGND sg13g2_fill_1
X_2743_ FrameData[24] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit24.Q VPWR
+ VGND sg13g2_dlhq_1
X_2812_ FrameData[29] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1625_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit14.Q N1END[2] N2END[6] E1END[2] E2END[6]
+ Inst_LUT4AB_ConfigMem.Inst_frame3_bit15.Q _0295_ VPWR VGND sg13g2_mux4_1
X_1556_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q _0225_ _0228_ _0227_ sg13g2_a21oi_1
X_2674_ FrameData[19] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit19.Q VPWR
+ VGND sg13g2_dlhq_1
X_3157_ Inst_LUT4AB_switch_matrix.N1BEG2 N1BEG[2] VPWR VGND sg13g2_buf_1
X_3226_ S2MID[7] S2BEGb[7] VPWR VGND sg13g2_buf_1
X_1487_ _1038_ _0154_ _0161_ VPWR VGND sg13g2_nor2_1
XFILLER_42_418 VPWR VGND sg13g2_fill_2
X_2039_ _0691_ VPWR _0692_ VGND Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q _0275_ sg13g2_o21ai_1
X_3088_ EE4END[5] EE4BEG[1] VPWR VGND sg13g2_buf_1
X_2108_ G _0755_ _0756_ VPWR VGND sg13g2_nor2_1
XFILLER_52_49 VPWR VGND sg13g2_fill_2
XFILLER_22_197 VPWR VGND sg13g2_fill_2
XFILLER_13_142 VPWR VGND sg13g2_fill_2
XFILLER_13_164 VPWR VGND sg13g2_fill_1
XFILLER_13_186 VPWR VGND sg13g2_fill_2
X_1410_ _0087_ Ci _1160_ VPWR VGND sg13g2_nand2_1
X_2390_ VPWR VGND Inst_LUT4AB_switch_matrix.DEBUG_select_LH_SR[0] _0659_ _0985_ _0661_
+ _0987_ _0665_ sg13g2_a221oi_1
XFILLER_3_65 VPWR VGND sg13g2_fill_1
X_1272_ _1110_ _1109_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit0.Q VPWR VGND sg13g2_nand2b_1
X_1341_ _0012_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q _0020_ _0021_ VPWR VGND sg13g2_a21o_1
X_3011_ FrameData[4] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit4.Q VPWR
+ VGND sg13g2_dlhq_1
X_2726_ FrameData[7] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit7.Q VPWR
+ VGND sg13g2_dlhq_1
X_1539_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q Inst_LUT4AB_switch_matrix.M_AD
+ _0211_ _0210_ sg13g2_a21oi_1
X_2588_ FrameData[29] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit29.Q VPWR
+ VGND sg13g2_dlhq_1
X_1608_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame9_bit14.Q _0277_ _0278_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit15.Q
+ sg13g2_a21oi_1
X_2657_ FrameData[2] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit2.Q VPWR
+ VGND sg13g2_dlhq_1
X_3209_ Inst_LUT4AB_switch_matrix.S1BEG2 S1BEG[2] VPWR VGND sg13g2_buf_1
XFILLER_27_234 VPWR VGND sg13g2_fill_2
XFILLER_37_60 VPWR VGND sg13g2_fill_2
X_1890_ VGND VPWR _0550_ _0549_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit19.Q sg13g2_or2_1
X_2511_ FrameData[16] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A12
+ VPWR VGND sg13g2_dlhq_1
XFILLER_38_2 VPWR VGND sg13g2_fill_1
X_2373_ Inst_LUT4AB_ConfigMem.Inst_frame0_bit30.Q Inst_LUT4AB_switch_matrix.JN2BEG2
+ Inst_LUT4AB_switch_matrix.JS2BEG2 Inst_LUT4AB_switch_matrix.E2BEG2 Inst_LUT4AB_switch_matrix.JW2BEG2
+ Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0970_ VPWR VGND sg13g2_mux4_1
X_2442_ FrameData[11] FrameStrobe[18] Inst_LB_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A0
+ VPWR VGND sg13g2_dlhq_1
X_1255_ VGND VPWR _1015_ _1086_ _1094_ _1093_ sg13g2_a21oi_1
X_1186_ VPWR _1027_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit0.Q VGND sg13g2_inv_1
X_1324_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit30.Q N2MID[5] E2MID[5] S2MID[5] W2MID[5]
+ Inst_LUT4AB_ConfigMem.Inst_frame7_bit31.Q _1159_ VPWR VGND sg13g2_mux4_1
X_2709_ FrameData[22] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_1942_ _0599_ VPWR _0600_ VGND Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q C sg13g2_o21ai_1
X_2991_ FrameData[16] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_21_218 VPWR VGND sg13g2_fill_2
X_1873_ E6END[1] S4END[1] Inst_LUT4AB_ConfigMem.Inst_frame0_bit22.Q _0533_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_43_0 VPWR VGND sg13g2_fill_1
X_2425_ FrameData[26] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A2
+ VPWR VGND sg13g2_dlhq_1
X_2356_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit20.Q G _1159_ Inst_LUT4AB_switch_matrix.JN2BEG2
+ _1118_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit21.Q Inst_LUT4AB_switch_matrix.E1BEG3
+ VPWR VGND sg13g2_mux4_1
XFILLER_44_39 VPWR VGND sg13g2_fill_2
X_2287_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit1.Q _0916_ _0917_ VPWR VGND sg13g2_nor2_1
X_1307_ VPWR _1143_ _1142_ VGND sg13g2_inv_1
X_1238_ W2END[4] W6END[0] Inst_LUT4AB_ConfigMem.Inst_frame3_bit6.Q _1078_ VPWR VGND
+ sg13g2_mux2_1
X_3190_ Inst_LUT4AB_switch_matrix.N4BEG3 N4BEG[15] VPWR VGND sg13g2_buf_1
X_2210_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit28.Q _0847_ _0848_ _0849_ _0850_ Inst_LUT4AB_ConfigMem.Inst_frame11_bit29.Q
+ Inst_LUT4AB_switch_matrix.W6BEG0 VPWR VGND sg13g2_mux4_1
X_2141_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit29.Q VPWR _0786_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit28.Q
+ _0779_ sg13g2_o21ai_1
X_2072_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit25.Q _0722_ _0723_ VPWR VGND sg13g2_nor2_1
X_1925_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit21.Q _0583_ _0584_ VPWR VGND sg13g2_nor2_1
X_2974_ FrameData[31] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit31.Q VPWR
+ VGND sg13g2_dlhq_1
X_1856_ Inst_LUT4AB_switch_matrix.JN2BEG6 Inst_LUT4AB_ConfigMem.Inst_frame7_bit18.Q
+ _0516_ VPWR VGND sg13g2_nor2b_1
X_1787_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit9.Q VPWR _0450_ VGND _0448_ _0449_ sg13g2_o21ai_1
X_2339_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit4.Q VPWR _0962_ VGND Inst_LUT4AB_ConfigMem.Inst_frame13_bit3.Q
+ _0961_ sg13g2_o21ai_1
X_2408_ Inst_LD_LUT4c_frame_config_dffesr.LUT_flop _1000_ _0998_ _0004_ VPWR VGND
+ sg13g2_mux2_1
XFILLER_52_151 VPWR VGND sg13g2_fill_1
X_1710_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame4_bit11.Q _0374_ _0376_ _0375_ sg13g2_a21oi_1
X_1641_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit12.Q _0307_ _0309_ _0290_ _0286_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit13.Q
+ _0310_ VPWR VGND sg13g2_mux4_1
XANTENNA_3 VPWR VGND EE4END[15] sg13g2_antennanp
X_1572_ Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q _0239_ _0243_ VPWR VGND sg13g2_nor2b_1
X_2690_ FrameData[3] FrameStrobe[10] Inst_LUT4AB_ConfigMem.Inst_frame10_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_3173_ N2MID[6] N2BEGb[6] VPWR VGND sg13g2_buf_1
X_2124_ _0769_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit29.Q _0770_ VPWR VGND sg13g2_nor2b_1
X_3242_ Inst_LUT4AB_switch_matrix.S4BEG3 S4BEG[15] VPWR VGND sg13g2_buf_1
X_2055_ _0706_ VPWR _0707_ VGND W1END[0] Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q
+ sg13g2_o21ai_1
X_1908_ _0567_ _0566_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit20.Q VPWR VGND sg13g2_nand2b_1
X_1839_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit20.Q VPWR _0500_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit19.Q
+ _0499_ sg13g2_o21ai_1
X_2957_ FrameData[14] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit14.Q VPWR
+ VGND sg13g2_dlhq_1
X_2888_ FrameData[9] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_40_110 VPWR VGND sg13g2_fill_1
X_2742_ FrameData[23] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit23.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_31_187 VPWR VGND sg13g2_fill_1
X_2811_ FrameData[28] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_1624_ _0293_ VPWR _0294_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0291_ sg13g2_o21ai_1
X_1555_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit16.Q VPWR _0227_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q
+ _0226_ sg13g2_o21ai_1
X_2673_ FrameData[18] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit18.Q VPWR
+ VGND sg13g2_dlhq_1
X_2107_ _0754_ VPWR _0755_ VGND Inst_LUT4AB_ConfigMem.Inst_frame14_bit16.Q _0753_
+ sg13g2_o21ai_1
X_3087_ EE4END[4] EE4BEG[0] VPWR VGND sg13g2_buf_1
X_3225_ S2MID[6] S2BEGb[6] VPWR VGND sg13g2_buf_1
X_1486_ _0159_ VPWR _0160_ VGND Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0156_ sg13g2_o21ai_1
X_3156_ Inst_LUT4AB_switch_matrix.N1BEG1 N1BEG[1] VPWR VGND sg13g2_buf_1
X_2038_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame8_bit20.Q Inst_LUT4AB_switch_matrix.JW2BEG5
+ _0691_ _1047_ sg13g2_a21oi_1
X_1340_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit1.Q _0014_ _0019_ _0020_ VPWR VGND sg13g2_nor3_1
X_1271_ Inst_LUT4AB_ConfigMem.Inst_frame5_bit31.Q N2END[2] E1END[0] N4END[2] E2END[2]
+ Inst_LUT4AB_ConfigMem.Inst_frame5_bit30.Q _1109_ VPWR VGND sg13g2_mux4_1
X_3010_ FrameData[3] FrameStrobe[0] Inst_LUT4AB_ConfigMem.Inst_frame0_bit3.Q VPWR
+ VGND sg13g2_dlhq_1
X_2656_ FrameData[1] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit1.Q VPWR
+ VGND sg13g2_dlhq_1
X_2725_ FrameData[6] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit6.Q VPWR
+ VGND sg13g2_dlhq_1
X_1469_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit12.Q VPWR _0144_ VGND Inst_LUT4AB_ConfigMem.Inst_frame3_bit11.Q
+ _0143_ sg13g2_o21ai_1
X_2587_ FrameData[28] FrameStrobe[14] Inst_LUT4AB_ConfigMem.Inst_frame14_bit28.Q VPWR
+ VGND sg13g2_dlhq_1
X_1538_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit15.Q VPWR _0210_ VGND Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q
+ _1052_ sg13g2_o21ai_1
X_1607_ Inst_LUT4AB_ConfigMem.Inst_frame6_bit14.Q N2MID[5] E2MID[5] S2MID[5] W2MID[5]
+ Inst_LUT4AB_ConfigMem.Inst_frame6_bit15.Q _0277_ VPWR VGND sg13g2_mux4_1
X_3208_ Inst_LUT4AB_switch_matrix.S1BEG1 S1BEG[1] VPWR VGND sg13g2_buf_1
X_3139_ FrameStrobe[4] FrameStrobe_O[4] VPWR VGND sg13g2_buf_1
XFILLER_50_260 VPWR VGND sg13g2_fill_1
XFILLER_42_238 VPWR VGND sg13g2_fill_1
XFILLER_6_106 VPWR VGND sg13g2_fill_1
XFILLER_2_378 VPWR VGND sg13g2_fill_1
XFILLER_18_235 VPWR VGND sg13g2_fill_1
X_2510_ FrameData[15] FrameStrobe[16] Inst_LE_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A11
+ VPWR VGND sg13g2_dlhq_1
X_2441_ FrameData[10] FrameStrobe[18] Inst_LA_LUT4c_frame_config_dffesr.c_reset_value
+ VPWR VGND sg13g2_dlhq_1
X_2372_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame0_bit29.Q _0334_ _0969_ _0968_ sg13g2_a21oi_1
X_1323_ VPWR _1158_ _1157_ VGND sg13g2_inv_1
X_1254_ _1093_ Inst_LUT4AB_ConfigMem.Inst_frame4_bit9.Q _1092_ VPWR VGND sg13g2_nand2b_1
X_1185_ VPWR _1026_ W2MID[4] VGND sg13g2_inv_1
XFILLER_24_216 VPWR VGND sg13g2_fill_1
X_2639_ FrameData[16] FrameStrobe[12] Inst_LUT4AB_ConfigMem.Inst_frame12_bit16.Q VPWR
+ VGND sg13g2_dlhq_1
X_2708_ FrameData[21] FrameStrobe[10] Inst_LUT4AB_switch_matrix.DEBUG_select_LB_EN[0]
+ VPWR VGND sg13g2_dlhq_1
X_1872_ _0530_ _0531_ Inst_LG_LUT4c_frame_config_dffesr.c_I0mux _0532_ VPWR VGND sg13g2_mux2_1
X_1941_ _0599_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit18.Q D VPWR VGND sg13g2_nand2b_1
X_2990_ FrameData[15] FrameStrobe[1] Inst_LUT4AB_ConfigMem.Inst_frame1_bit15.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_36_0 VPWR VGND sg13g2_fill_2
X_2286_ Inst_LUT4AB_ConfigMem.Inst_frame13_bit31.Q N1END[1] E1END[1] S1END[1] D Inst_LUT4AB_ConfigMem.Inst_frame12_bit0.Q
+ _0916_ VPWR VGND sg13g2_mux4_1
X_1306_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit6.Q A B C E Inst_LUT4AB_ConfigMem.Inst_frame2_bit7.Q
+ _1142_ VPWR VGND sg13g2_mux4_1
X_2424_ FrameData[25] FrameStrobe[19] Inst_LA_LUT4c_frame_config_dffesr.inst_cus_mux161_buf.A1
+ VPWR VGND sg13g2_dlhq_1
X_2355_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit11.Q E Inst_LUT4AB_switch_matrix.E2BEG3
+ _0453_ _0129_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit10.Q Inst_LUT4AB_switch_matrix.S1BEG0
+ VPWR VGND sg13g2_mux4_1
X_1237_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit8.Q _1076_ _1077_ VPWR VGND sg13g2_nor2_1
XFILLER_52_399 VPWR VGND sg13g2_fill_2
XFILLER_38_116 VPWR VGND sg13g2_fill_1
X_2140_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit27.Q _0781_ _0785_ _0784_ sg13g2_a21oi_1
XFILLER_15_5 VPWR VGND sg13g2_fill_2
XFILLER_34_322 VPWR VGND sg13g2_fill_2
X_2071_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame1_bit23.Q _0720_ _0722_ _0721_ sg13g2_a21oi_1
X_1924_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q _0580_ _0583_ _0582_ sg13g2_a21oi_1
X_1855_ Inst_LUT4AB_switch_matrix.JN2BEG6 _0509_ _0515_ _0507_ _0501_ VPWR VGND sg13g2_a22oi_1
X_2973_ FrameData[30] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit30.Q VPWR
+ VGND sg13g2_dlhq_1
XFILLER_39_18 VPWR VGND sg13g2_fill_1
X_1786_ Inst_LUT4AB_ConfigMem.Inst_frame7_bit8.Q W2MID[0] _0449_ VPWR VGND sg13g2_nor2_1
X_2269_ VGND VPWR W1END[2] Inst_LUT4AB_ConfigMem.Inst_frame12_bit6.Q _0901_ Inst_LUT4AB_ConfigMem.Inst_frame12_bit7.Q
+ sg13g2_a21oi_1
X_2338_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame13_bit2.Q _1084_ _0961_ _0960_ sg13g2_a21oi_1
X_2407_ Inst_LD_LUT4c_frame_config_dffesr.c_reset_value _0688_ _0999_ _1000_ VPWR
+ VGND sg13g2_mux2_1
XFILLER_29_40 VPWR VGND sg13g2_fill_1
X_1640_ VPWR _0309_ _0308_ VGND sg13g2_inv_1
X_1571_ _0241_ VPWR _0242_ VGND Inst_LUT4AB_ConfigMem.Inst_frame9_bit10.Q _0236_ sg13g2_o21ai_1
XANTENNA_4 VPWR VGND EE4END[4] sg13g2_antennanp
X_3241_ Inst_LUT4AB_switch_matrix.S4BEG2 S4BEG[14] VPWR VGND sg13g2_buf_1
X_2123_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit27.Q _0767_ _0769_ _0768_ sg13g2_a21oi_1
X_3172_ N2MID[5] N2BEGb[5] VPWR VGND sg13g2_buf_1
XFILLER_26_108 VPWR VGND sg13g2_fill_2
X_2054_ _0706_ Inst_LUT4AB_ConfigMem.Inst_frame2_bit22.Q W1END[2] VPWR VGND sg13g2_nand2b_1
X_1838_ E F Inst_LUT4AB_ConfigMem.Inst_frame4_bit18.Q _0499_ VPWR VGND sg13g2_mux2_1
X_1907_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit18.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame3_bit19.Q
+ _0566_ VPWR VGND sg13g2_mux4_1
X_2956_ FrameData[13] FrameStrobe[2] Inst_LUT4AB_ConfigMem.Inst_frame2_bit13.Q VPWR
+ VGND sg13g2_dlhq_1
X_2887_ FrameData[8] FrameStrobe[4] Inst_LUT4AB_ConfigMem.Inst_frame4_bit8.Q VPWR
+ VGND sg13g2_dlhq_1
X_1769_ Inst_LUT4AB_ConfigMem.Inst_frame1_bit10.Q A B C D Inst_LUT4AB_ConfigMem.Inst_frame1_bit11.Q
+ _0433_ VPWR VGND sg13g2_mux4_1
XFILLER_15_64 VPWR VGND sg13g2_fill_2
XFILLER_31_133 VPWR VGND sg13g2_fill_1
XFILLER_31_111 VPWR VGND sg13g2_fill_1
XFILLER_16_196 VPWR VGND sg13g2_fill_2
X_2741_ FrameData[22] FrameStrobe[9] Inst_LUT4AB_ConfigMem.Inst_frame9_bit22.Q VPWR
+ VGND sg13g2_dlhq_1
X_2672_ FrameData[17] FrameStrobe[11] Inst_LUT4AB_ConfigMem.Inst_frame11_bit17.Q VPWR
+ VGND sg13g2_dlhq_1
X_2810_ FrameData[27] FrameStrobe[7] Inst_LUT4AB_ConfigMem.Inst_frame7_bit27.Q VPWR
+ VGND sg13g2_dlhq_1
X_1623_ _0293_ Inst_LUT4AB_ConfigMem.Inst_frame3_bit16.Q _0292_ VPWR VGND sg13g2_nand2b_1
X_1554_ S1END[2] S2END[6] Inst_LUT4AB_ConfigMem.Inst_frame4_bit14.Q _0226_ VPWR VGND
+ sg13g2_mux2_1
X_3224_ S2MID[5] S2BEGb[5] VPWR VGND sg13g2_buf_1
X_1485_ VGND VPWR Inst_LUT4AB_ConfigMem.Inst_frame2_bit3.Q _0158_ _0159_ _1037_ sg13g2_a21oi_1
.ends

